magic
tech sky130B
magscale 1 2
timestamp 1687809653
<< locali >>
rect -1900 660 -432 698
rect -1900 644 -520 660
rect -1900 -544 -1846 644
rect -540 -544 -520 644
rect -1900 -560 -520 -544
rect -460 -560 -432 660
rect -1900 -592 -432 -560
<< viali >>
rect -520 -560 -460 660
<< metal1 >>
rect -1732 398 -1300 1506
rect -304 1486 22 1506
rect -304 1446 60 1486
rect -304 1354 22 1446
rect 1650 1354 2352 1506
rect -540 660 -432 698
rect -1084 380 -652 532
rect -1084 320 -900 380
rect -840 320 -652 380
rect -1734 190 -1302 236
rect -1734 130 -1406 190
rect -1346 130 -1302 190
rect -1084 166 -652 320
rect -1734 -130 -1302 130
rect -1084 -212 -652 -60
rect -1084 -272 -800 -212
rect -740 -272 -652 -212
rect -1734 -1716 -1302 -356
rect -1084 -426 -652 -272
rect -1734 -1776 -1372 -1716
rect -1312 -1776 -1302 -1716
rect -1734 -1906 -1302 -1776
rect -540 -560 -520 660
rect -460 -560 -432 660
rect -304 -400 -152 1354
rect 0 656 10 716
rect 70 656 80 716
rect 2200 600 2352 1354
rect 1172 410 1182 470
rect 1242 410 1252 470
rect 20 20 60 60
rect 1650 0 1954 152
rect -304 -552 0 -400
rect -540 -1754 -432 -560
rect 1802 -754 1954 0
rect 2200 -240 2240 -200
rect 3380 -240 3420 -200
rect 1802 -906 2214 -754
rect 1172 -1116 1182 -1056
rect 1242 -1116 1252 -1056
rect 0 -1250 10 -1190
rect 70 -1250 80 -1190
rect 1802 -1754 1954 -906
rect -540 -1906 0 -1754
rect 1650 -1906 1954 -1754
<< via1 >>
rect -900 320 -840 380
rect -1406 130 -1346 190
rect -800 -272 -740 -212
rect -1372 -1776 -1312 -1716
rect 10 656 70 716
rect 1182 410 1242 470
rect 1182 -1116 1242 -1056
rect 10 -1250 70 -1190
<< metal2 >>
rect -910 1306 870 1386
rect -910 380 -830 1306
rect -910 320 -900 380
rect -840 320 -830 380
rect -910 310 -830 320
rect 0 716 80 726
rect 0 656 10 716
rect 70 656 80 716
rect -1420 194 -60 204
rect -1420 190 -134 194
rect -1420 130 -1406 190
rect -1346 130 -134 190
rect -1420 126 -134 130
rect -68 126 -60 194
rect -1420 116 -60 126
rect -810 -212 -730 -202
rect -810 -272 -800 -212
rect -740 -272 -730 -212
rect -810 -516 -730 -272
rect -810 -526 -60 -516
rect -810 -594 -134 -526
rect -68 -594 -60 -526
rect -810 -604 -60 -594
rect 0 -1190 80 656
rect 1170 474 1434 484
rect 1170 470 1366 474
rect 1170 410 1182 470
rect 1242 410 1366 470
rect 1170 406 1366 410
rect 1170 396 1434 406
rect 1800 474 3780 484
rect 1800 406 1806 474
rect 1874 406 3780 474
rect 1800 396 3780 406
rect 140 194 1710 204
rect 140 126 146 194
rect 212 126 1710 194
rect 140 116 1710 126
rect 140 -526 1580 -516
rect 140 -594 146 -526
rect 214 -594 1580 -526
rect 140 -604 1580 -594
rect 3070 -1042 3150 -786
rect 1170 -1052 1252 -1042
rect 1170 -1120 1178 -1052
rect 1246 -1120 1252 -1052
rect 1170 -1130 1252 -1120
rect 1800 -1052 3150 -1042
rect 1800 -1120 1806 -1052
rect 1874 -1120 3150 -1052
rect 1800 -1130 3150 -1120
rect 0 -1250 10 -1190
rect 70 -1250 80 -1190
rect 0 -1260 80 -1250
rect -1382 -1716 870 -1706
rect -1382 -1776 -1372 -1716
rect -1312 -1776 870 -1716
rect -1382 -1786 870 -1776
<< via2 >>
rect -134 126 -68 194
rect -134 -594 -68 -526
rect 1366 406 1434 474
rect 1806 406 1874 474
rect 146 126 212 194
rect 146 -594 214 -526
rect 1178 -1056 1246 -1052
rect 1178 -1116 1182 -1056
rect 1182 -1116 1242 -1056
rect 1242 -1116 1246 -1056
rect 1178 -1120 1246 -1116
rect 1806 -1120 1874 -1052
<< metal3 >>
rect 1356 474 1884 480
rect 1356 406 1366 474
rect 1434 406 1806 474
rect 1874 406 1884 474
rect 1356 400 1884 406
rect -146 194 226 204
rect -146 126 -134 194
rect -68 126 146 194
rect 212 126 226 194
rect -146 116 226 126
rect -146 -526 226 -516
rect -146 -594 -134 -526
rect -68 -594 146 -526
rect 214 -594 226 -526
rect -146 -604 226 -594
rect 1160 -1052 1884 -1046
rect 1160 -1120 1178 -1052
rect 1246 -1120 1806 -1052
rect 1874 -1120 1884 -1052
rect 1160 -1126 1884 -1120
use sw  X1
timestamp 1687764782
transform 1 0 0 0 1 786
box 0 -786 1720 720
use sw  X2
timestamp 1687764782
transform 1 0 0 0 1 -1120
box 0 -786 1720 720
use sw  X3
timestamp 1687764782
transform 1 0 2200 0 1 -120
box 0 -786 1720 720
use sky130_fd_pr__res_high_po_0p35_2NY7PZ  XR1
timestamp 1687795939
transform 0 -1 -1193 1 0 497
box -201 -707 201 707
use sky130_fd_pr__res_high_po_0p35_2NY7PZ  XR2
timestamp 1687795939
transform 0 -1 -1193 1 0 201
box -201 -707 201 707
use sky130_fd_pr__res_high_po_0p35_2NY7PZ  XR3
timestamp 1687795939
transform 0 -1 -1193 1 0 -95
box -201 -707 201 707
use sky130_fd_pr__res_high_po_0p35_2NY7PZ  XR4
timestamp 1687795939
transform 0 -1 -1193 1 0 -391
box -201 -707 201 707
<< labels >>
flabel metal1 0 666 40 706 0 FreeSans 256 0 0 0 d0
port 4 nsew
flabel metal1 20 1446 60 1486 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 20 20 60 60 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 2200 -240 2240 -200 0 FreeSans 256 0 0 0 d1
port 5 nsew
flabel metal1 3380 -240 3420 -200 0 FreeSans 256 0 0 0 vout
port 6 nsew
flabel metal1 -1638 1396 -1598 1436 0 FreeSans 256 0 0 0 vrefh
port 2 nsew
flabel metal1 -1540 -1840 -1500 -1800 0 FreeSans 256 0 0 0 vrefl
port 3 nsew
<< end >>
