magic
tech sky130B
magscale 1 2
timestamp 1687357769
<< metal1 >>
rect -702 972 -502 1172
rect 640 930 720 940
rect 640 870 650 930
rect 710 870 720 930
rect 26 578 66 860
rect 102 618 240 820
rect 0 500 92 576
rect -200 300 92 500
rect 0 268 92 300
rect 154 450 240 618
rect 412 578 452 860
rect 640 820 720 870
rect 488 808 588 820
rect 488 630 510 808
rect 570 630 588 808
rect 488 618 588 630
rect 640 618 762 820
rect 800 578 840 860
rect 874 618 1148 820
rect 386 450 478 538
rect 772 450 864 538
rect 154 350 864 450
rect 26 74 66 222
rect 154 190 240 350
rect 386 222 478 350
rect 772 222 864 350
rect 102 106 240 190
rect 280 -20 340 190
rect 410 74 450 222
rect 488 178 588 190
rect 488 118 510 178
rect 570 118 588 178
rect 488 106 588 118
rect 798 74 838 222
rect 960 190 1060 618
rect 1184 578 1224 860
rect 1260 618 1442 820
rect 1158 430 1250 538
rect 1158 370 1174 430
rect 1234 370 1250 430
rect 1158 222 1250 370
rect 1872 300 2072 500
rect 874 106 1146 190
rect 1184 74 1224 222
rect 1260 178 1400 190
rect 1260 118 1328 178
rect 1388 118 1400 178
rect 1260 106 1400 118
rect -200 -234 0 -34
rect -750 -944 -550 -744
rect -788 -1224 -588 -1024
<< via1 >>
rect 650 870 710 930
rect 510 630 570 808
rect 510 118 570 178
rect 1174 370 1234 430
rect 1328 118 1388 178
<< metal2 >>
rect 640 930 1388 940
rect 640 870 650 930
rect 710 870 1388 930
rect 640 860 1388 870
rect 500 808 600 818
rect 500 630 510 808
rect 570 630 600 808
rect 500 440 600 630
rect 500 430 1240 440
rect 500 370 1174 430
rect 1234 370 1240 430
rect 500 360 1240 370
rect 500 178 600 360
rect 500 118 510 178
rect 570 118 600 178
rect 500 108 600 118
rect 1328 178 1388 860
rect 1328 108 1388 118
use sky130_fd_pr__pfet_01v8_XPYSY6  sky130_fd_pr__pfet_01v8_XPYSY6_0
timestamp 1687352469
transform 1 0 46 0 1 719
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_XHX9Y6  XM2
timestamp 1687352469
transform 1 0 432 0 1 719
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_XHX9Y6  XM3
timestamp 1687352469
transform 1 0 818 0 1 719
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_XPYSY6  XM4
timestamp 1687352469
transform 1 0 1204 0 1 719
box -246 -319 246 319
use sky130_fd_pr__nfet_01v8_ZFH27D  XM5
timestamp 1687352469
transform 1 0 46 0 1 148
box -246 -252 246 252
use sky130_fd_pr__nfet_01v8_HEL24J  XM6
timestamp 1687352469
transform 1 0 432 0 1 148
box -246 -252 246 252
use sky130_fd_pr__nfet_01v8_HEL24J  XM7
timestamp 1687352469
transform 1 0 818 0 1 148
box -246 -252 246 252
use sky130_fd_pr__nfet_01v8_ZFH27D  XM8
timestamp 1687352469
transform 1 0 1204 0 1 148
box -246 -252 246 252
<< labels >>
flabel metal1 -750 -944 -550 -744 0 FreeSans 256 0 0 0 vin1
port 3 nsew
flabel metal1 -788 -1224 -588 -1024 0 FreeSans 256 0 0 0 vin2
port 4 nsew
flabel metal1 -200 -234 0 -34 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 -702 972 -502 1172 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 -200 300 0 500 0 FreeSans 256 0 0 0 din
port 2 nsew
flabel metal1 1872 300 2072 500 0 FreeSans 256 0 0 0 vout
port 5 nsew
<< end >>
