magic
tech sky130B
timestamp 1688377021
<< metal1 >>
rect 540 7280 640 7380
rect 1100 7370 1140 7410
rect 1350 7380 1390 7420
rect 1350 6994 1390 7034
rect 2450 6541 2490 6581
rect 2600 5568 2640 5608
rect 2600 3682 2640 3722
rect 2703 3687 2708 3717
rect 2738 3687 2743 3717
rect 3680 3715 3720 3720
rect 3680 3685 3685 3715
rect 3715 3685 3720 3715
rect 3186 3600 3191 3630
rect 3221 3600 3226 3630
rect 3186 3513 3191 3543
rect 3221 3513 3226 3543
rect 3390 2110 3575 2186
rect 3499 300 3575 2110
rect 3390 224 3575 300
rect 483 -200 699 0
rect 1080 -200 1156 2
rect 2450 -377 2526 199
rect 2600 -130 2640 -90
rect 3185 -130 3225 -90
rect 2450 -453 2600 -377
rect 3185 -3720 3190 -3690
rect 3220 -3720 3225 -3690
rect 3680 -3905 3720 3685
rect 2703 -3937 2708 -3907
rect 2738 -3937 2743 -3907
rect 3565 -3910 3720 -3905
rect 3565 -3940 3570 -3910
rect 3600 -3940 3720 -3910
rect 3565 -3945 3720 -3940
rect 540 -7580 640 -7480
<< via1 >>
rect 2708 3687 2738 3717
rect 3685 3685 3715 3715
rect 3191 3600 3221 3630
rect 3191 3513 3221 3543
rect 3190 -3720 3220 -3690
rect 2708 -3937 2738 -3907
rect 3570 -3940 3600 -3910
<< metal2 >>
rect 2700 3719 2893 3724
rect 2700 3717 2850 3719
rect 2700 3687 2708 3717
rect 2738 3687 2850 3717
rect 2700 3685 2850 3687
rect 2884 3685 2893 3719
rect 2700 3680 2893 3685
rect 3500 3719 3720 3724
rect 3534 3715 3720 3719
rect 3534 3685 3685 3715
rect 3715 3685 3720 3715
rect 3500 3679 3720 3685
rect 3186 3631 3290 3636
rect 3186 3630 3252 3631
rect 3186 3600 3191 3630
rect 3221 3600 3252 3630
rect 3186 3599 3252 3600
rect 3284 3599 3290 3631
rect 3186 3594 3290 3599
rect 3581 3631 3621 3636
rect 3581 3599 3585 3631
rect 3617 3599 3621 3631
rect 3186 3543 3226 3548
rect 3186 3513 3191 3543
rect 3221 3513 3226 3543
rect 3186 3508 3226 3513
rect 2295 1545 2335 1551
rect 2295 1511 2298 1545
rect 2332 1511 2335 1545
rect 590 323 1390 363
rect 590 -400 630 323
rect 2295 285 2335 1511
rect 2295 251 2298 285
rect 2332 251 2335 285
rect 2295 246 2335 251
rect 2274 -200 2350 0
rect 2295 -356 2335 -350
rect 2295 -390 2298 -356
rect 2332 -390 2335 -356
rect 590 -440 1390 -400
rect 1350 -630 1390 -440
rect 2295 -1635 2335 -390
rect 2450 -1043 2490 823
rect 3581 240 3621 3599
rect 3390 200 3621 240
rect 3455 -393 3620 -353
rect 2295 -1669 2298 -1635
rect 2332 -1669 2335 -1635
rect 2295 -1674 2335 -1669
rect 3185 -3689 3289 -3684
rect 3185 -3690 3251 -3689
rect 3185 -3720 3190 -3690
rect 3220 -3720 3251 -3690
rect 3185 -3721 3251 -3720
rect 3283 -3721 3289 -3689
rect 3185 -3726 3289 -3721
rect 3581 -3689 3620 -393
rect 3581 -3721 3584 -3689
rect 3616 -3721 3620 -3689
rect 3581 -3726 3620 -3721
rect 2700 -3905 2893 -3900
rect 2700 -3907 2850 -3905
rect 2700 -3937 2708 -3907
rect 2738 -3937 2850 -3907
rect 2700 -3939 2850 -3937
rect 2884 -3939 2893 -3905
rect 2700 -3944 2893 -3939
rect 3494 -3905 3605 -3900
rect 3494 -3939 3500 -3905
rect 3534 -3910 3605 -3905
rect 3534 -3939 3570 -3910
rect 3494 -3940 3570 -3939
rect 3600 -3940 3605 -3910
rect 3494 -3945 3605 -3940
<< via2 >>
rect 2850 3685 2884 3719
rect 3500 3685 3534 3719
rect 3252 3599 3284 3631
rect 3585 3599 3617 3631
rect 2298 1511 2332 1545
rect 2298 251 2332 285
rect 2298 -390 2332 -356
rect 2298 -1669 2332 -1635
rect 3251 -3721 3283 -3689
rect 3584 -3721 3616 -3689
rect 2850 -3939 2884 -3905
rect 3500 -3939 3534 -3905
<< metal3 >>
rect 2840 3719 3540 3724
rect 2840 3685 2850 3719
rect 2884 3685 3500 3719
rect 3534 3685 3540 3719
rect 2840 3679 3540 3685
rect 3245 3631 3625 3636
rect 3245 3599 3252 3631
rect 3284 3599 3585 3631
rect 3617 3599 3625 3631
rect 3245 3594 3625 3599
rect 2293 1545 2337 1754
rect 2293 1511 2298 1545
rect 2332 1511 2337 1545
rect 2293 1506 2337 1511
rect 2293 285 2337 290
rect 2293 251 2298 285
rect 2332 251 2337 285
rect 2293 -356 2337 251
rect 2293 -390 2298 -356
rect 2332 -390 2337 -356
rect 2293 -395 2337 -390
rect 2293 -1635 2337 -1630
rect 2293 -1669 2298 -1635
rect 2332 -1669 2337 -1635
rect 2293 -2014 2337 -1669
rect 3245 -3689 3625 -3684
rect 3245 -3721 3251 -3689
rect 3283 -3721 3584 -3689
rect 3616 -3721 3625 -3689
rect 3245 -3726 3625 -3721
rect 2840 -3905 3540 -3900
rect 2840 -3939 2850 -3905
rect 2884 -3939 3500 -3905
rect 3534 -3939 3540 -3905
rect 2840 -3945 3540 -3939
use 4bit_dac  X1
timestamp 1688377021
transform 1 0 -200 0 1 3512
box 600 -3512 3720 3912
use 4bit_dac  X2
timestamp 1688377021
transform 1 0 -200 0 1 -4112
box 600 -3512 3720 3912
use sw  X3
timestamp 1687966408
transform 1 0 2600 0 1 -60
box 0 -393 860 360
<< labels >>
flabel metal1 540 7280 640 7380 0 FreeSans 128 0 0 0 vrefh
port 2 nsew
flabel metal1 540 -7580 640 -7480 0 FreeSans 128 0 0 0 vrefl
port 3 nsew
flabel metal1 1350 7380 1390 7420 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 1100 7370 1140 7410 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 1350 6994 1390 7034 0 FreeSans 128 0 0 0 d0
port 4 nsew
flabel metal1 2450 6541 2490 6581 0 FreeSans 128 0 0 0 d1
port 5 nsew
flabel metal1 2600 5568 2640 5608 0 FreeSans 128 0 0 0 d2
port 6 nsew
flabel metal1 2600 3682 2640 3722 0 FreeSans 128 0 0 0 d3
port 7 nsew
flabel metal1 2600 -130 2640 -90 0 FreeSans 128 0 0 0 d4
port 8 nsew
flabel metal1 3185 -130 3225 -90 0 FreeSans 128 0 0 0 vout
port 9 nsew
<< end >>
