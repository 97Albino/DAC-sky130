* NGSPICE file created from 8bit_dac.ext - technology: sky130B

.subckt x8bit_dac vrefh vrefl d0 d1 d2 d3 d4 d5 d6 d7 vout vss vdd
X0 X1.X2.X1.X2.X3.vin2 a_19722_10916# X1.X2.X1.X3.vin2 vdd.t1362 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 X1.X1.X1.X2.X1.X2.X1.vin2 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin1 vdd.t360 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X3 X2.X2.X1.X2.X1.X1.X3.vin2 a_46116_15634# X2.X2.X1.X2.X1.X2.vrefh vss.t288 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X4 X2.X2.X1.X3.vin1 a_49002_18540# X2.X2.X3.vin1 vss.t757 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X5 vdd.t128 a_11072_4110# a_10686_4110# vdd.t127 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X6 a_46502_9916# a_46116_9916# vdd.t125 vdd.t124 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X7 X2.X1.X1.X1.X1.X2.X3.vin1 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin2 vss.t1425 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X8 vss.t684 a_52492_18358# a_52106_18358# vss.t683 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X9 X1.X2.X2.X2.X1.X1.X3.vin2 a_23512_20264# X1.X2.X2.X2.X1.X1.vout vss.t672 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X10 a_35312_892# a_34926_892# vdd.t1430 vdd.t1429 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 a_2582_13728# a_2196_13728# vss.t755 vss.t754 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X12 a_16836_25164# d0.t0 vss.t634 vss.t633 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X13 vdd.t283 a_8872_16452# a_8486_16452# vdd.t282 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 a_33676_12822# d1.t0 vss.t788 vss.t787 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X15 X1.X1.X2.X1.X2.X1.X1.vin2 a_11072_11734# X1.X1.X2.X1.X2.X1.X3.vin1 vss.t1431 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X16 X2.X2.X1.X1.X1.X2.X3.vin1 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin1 vdd.t957 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X17 a_46502_4198# a_46116_4198# vdd.t832 vdd.t831 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X19 X2.X2.X2.X1.X1.X2.X3.vin1 a_54606_7922# X2.X2.X2.X1.X1.X2.X1.vin2 vdd.t1447 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X20 X2.X1.X1.X1.X2.X2.X3.vin2 a_34062_20446# X2.X1.X1.X1.X2.X2.vout vdd.t1258 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 X2.X2.X2.X2.X1.X2.X1.vin1 a_54992_23170# X2.X2.X2.X2.X1.X2.X3.vin1 vdd.t1370 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X22 X2.X1.X2.X2.X1.X1.vout a_37766_20264# X2.X1.X2.X2.X1.X1.X3.vin2 vdd.t1412 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X23 a_16836_4198# d0.t1 vss.t636 vss.t635 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X24 X1.X2.X2.X1.X1.X1.vout a_23126_5016# X1.X2.X2.X1.X1.X1.X3.vin1 vss.t1291 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X25 X2.X2.X1.X2.X3.vin1 a_49002_10916# X2.X2.X1.X3.vin2 vss.t1426 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X26 X1.X1.X1.X2.X1.X1.X3.vin2 a_4782_16634# X1.X1.X1.X2.X1.X1.vout vdd.t1366 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X27 X1.X1.X2.X1.X1.X1.X1.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 vss.t242 sky130_fd_pr__res_high_po_0p35 l=1.09
X28 vss.t1369 d0.t2 a_54992_13640# vss.t1368 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X29 vdd.t887 a_23212_6962# a_22826_6962# vdd.t886 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 a_46502_15634# a_46116_15634# vss.t287 vss.t286 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X31 vss.t1371 d0.t3 a_25712_17452# vss.t1370 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X32 X1.X1.X2.X3.vin2 a_8186_25982# X1.X1.X2.X2.X3.vin1 vss.t1397 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X33 a_17222_19446# a_16836_19446# vss.t1536 vss.t1535 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X34 X2.X1.X1.X1.X2.X1.vout a_34362_22312# X2.X1.X1.X1.X3.vin2 vss.t812 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X35 X1.X2.X1.X1.X1.X2.X3.vin2 a_19422_28070# X1.X2.X1.X1.X1.X2.vout vdd.t658 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X36 vdd.t1341 d0.t4 a_11072_17452# vdd.t1340 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X37 X2.X1.X1.X2.X2.X2.X1.vin2 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin1 vdd.t441 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X38 X1.X1.X1.X1.X1.X1.X3.vin2 a_2196_30882# X1.X1.X1.X1.X1.X1.X2.vin1 vdd.t1087 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X39 X1.X2.X2.X2.X1.X2.X1.vin2 a_25712_23170# X1.X2.X2.X2.X1.X2.X3.vin1 vss.t902 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X40 a_19422_31882# a_19036_31882# vdd.t1081 vdd.t1080 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X41 X2.X2.X2.X2.X2.X1.vout a_52492_29834# X2.X2.X2.X2.X3.vin2 vdd.t118 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X42 X2.X2.vrefh X2.X2.X1.X1.X1.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X43 X2.X2.X1.X1.X2.X2.vout a_49002_22312# X2.X2.X1.X1.X3.vin2 vdd.t1106 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X44 a_46502_28976# a_46116_28976# vdd.t956 vdd.t955 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X45 vdd.t845 d1.t1 a_38152_27888# vdd.t844 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X46 a_4782_31882# a_4396_31882# vss.t251 vss.t250 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X47 vdd.t1343 d0.t5 a_25712_9828# vdd.t1342 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X48 X1.X1.X1.X2.X1.X2.X2.vin1 a_2582_11822# X1.X1.X1.X2.X1.X2.X3.vin2 vss.t300 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X49 vss.t898 a_25712_28888# a_25326_28888# vss.t897 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X50 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X51 X1.X2.X1.X2.vrefh a_17222_19446# X1.X2.X1.X1.X2.X2.X3.vin2 vdd.t1108 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X52 a_2582_32788# a_2196_32788# vdd.t1084 vdd.t1083 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X53 X2.X2.X2.X2.X2.X2.X3.vin1 a_52792_31700# X2.X2.X2.X2.X2.X2.vout vdd.t877 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X54 X1.X2.X1.X1.X2.X2.vout a_19036_20446# X1.X2.X1.X1.X2.X2.X3.vin1 vdd.t640 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X55 X2.X1.X2.X2.X1.X2.X3.vin1 a_39966_23170# X2.X1.X2.X2.X1.X2.X1.vin2 vdd.t114 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X56 X2.X2.X2.X2.X2.X2.X3.vin2 a_54606_32700# vrefl.t1 vdd.t1423 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X57 X2.X2.X2.X2.X2.X2.X3.vin1 a_54606_30794# X2.X2.X2.X2.X2.X2.X1.vin1 vss.t971 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X58 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X59 a_5082_18540# a_4696_18540# vdd.t1418 vdd.t1417 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X60 X1.X1.X1.X1.X3.vin1 a_4696_29936# X1.X1.X1.X1.X1.X1.vout vdd.t653 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X61 vdd.t1345 d0.t6 a_54992_21264# vdd.t1344 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X62 vdd.t1347 d0.t7 a_25712_25076# vdd.t1346 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X63 a_4782_5198# a_4396_5198# vss.t974 vss.t973 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X64 vdd.t1155 d3.t0 a_23212_10734# vdd.t1154 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X65 X1.X1.X1.X1.X2.X1.X1.vin2 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin1 vdd.t960 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X66 vss.t1442 a_40352_15546# a_39966_15546# vss.t1441 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X67 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X68 X2.X1.X1.X1.X2.X1.vout a_33676_24258# X2.X1.X1.X1.X2.X1.X3.vin1 vdd.t330 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X69 a_5646_892# d5.t0 vss.t36 vss.t35 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X70 a_4396_20446# d1.t2 vdd.t847 vdd.t846 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X71 X2.X1.X1.X3.vin1 a_33976_26164# X2.X1.X1.X1.X3.vin1 vdd.t1517 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X72 X2.X1.X2.X2.X3.vin2 a_37466_29834# X2.X1.X2.X2.X2.X2.vout vdd.t660 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X73 a_5082_10916# a_4696_10916# vdd.t1365 vdd.t1364 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X74 X2.X1.X2.X2.X1.X1.X1.vin1 a_40352_19358# X2.X1.X2.X2.X1.X1.X3.vin1 vdd.t421 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X75 a_17222_6104# a_16836_6104# vss.t372 vss.t371 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X76 X1.X2.X1.X1.X2.X1.X1.vin1 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin1 vss.t1133 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X77 X2.X1.X1.X2.X2.X1.vout a_34362_7064# X2.X1.X1.X2.X3.vin2 vss.t339 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X78 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X79 vrefl.t2 a_54992_32700# X2.X2.X2.X2.X2.X2.X3.vin2 vss.t1462 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X80 X2.X1.X2.X2.X2.X2.vout a_37766_31700# X2.X1.X2.X2.X2.X2.X3.vin2 vdd.t1411 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X81 vdd.t252 a_23512_8828# a_23126_8828# vdd.t251 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X82 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X83 X1.X1.X2.X1.X1.X1.X3.vin1 a_8872_5016# X1.X1.X2.X1.X1.X1.vout vdd.t288 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X84 X1.X1.X1.X2.X1.X2.X3.vin1 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin1 vdd.t727 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X85 X2.X1.X1.X2.X2.X2.X3.vin2 a_34062_5198# X2.X1.X1.X2.X2.X2.vout vdd.t1367 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X86 a_31862_19446# a_31476_19446# vss.t2 vss.t1 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X87 X1.X1.X2.X2.X2.X1.vout a_8486_27888# X1.X1.X2.X2.X2.X1.X3.vin2 vdd.t49 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X88 X2.X2.X2.X1.X1.X1.X3.vin1 a_52792_5016# X2.X2.X2.X1.X1.X1.vout vdd.t1224 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X89 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X90 X2.X2.X2.vrefh.t2 a_46502_4198# X2.X2.X1.X2.X2.X2.X3.vin2 vdd.t1123 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X91 vdd.t410 a_54992_7922# a_54606_7922# vdd.t409 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X92 vss.t763 a_11072_6016# a_10686_6016# vss.t762 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X93 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X94 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X95 a_34062_31882# a_33676_31882# vdd.t715 vdd.t714 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X96 X1.X2.X1.X1.X3.vin1 a_19336_29936# X1.X2.X1.X1.X1.X1.vout vdd.t764 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X97 vss.t1373 d0.t8 a_11072_26982# vss.t1372 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X98 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X99 X1.X1.X2.X2.X2.X2.X1.vin1 a_11072_30794# X1.X1.X2.X2.X2.X2.X3.vin1 vdd.t509 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X100 X2.X1.X1.X2.X2.vrefh a_31862_11822# X2.X1.X1.X2.X1.X2.X3.vin2 vdd.t1026 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X101 X1.X1.X2.X1.X2.X1.X3.vin1 a_10686_11734# X1.X1.X2.X1.X2.X1.X1.vin1 vss.t983 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X102 X2.X2.X2.X1.X2.X2.X3.vin1 a_54606_15546# X2.X2.X2.X1.X2.X2.X1.vin2 vdd.t65 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X103 X1.X2.X2.X2.X1.X1.X3.vin1 a_25326_19358# X1.X2.X2.X2.X1.X1.X1.vin2 vdd.t536 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X104 vss.t548 a_25712_19358# a_25326_19358# vss.t547 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X105 a_4782_28070# a_4396_28070# vdd.t782 vdd.t781 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X106 vss.t402 a_52792_16452# a_52406_16452# vss.t401 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X107 X2.X1.X2.X2.X2.X2.X3.vin2 a_39966_32700# X2.X1.X2.X2.X2.X2.X2.vin1 vss.t277 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X108 a_48316_28070# d1.t3 vss.t873 vss.t872 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X109 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X110 vdd.t1349 d0.t9 a_54992_32700# vdd.t1348 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X111 X1.X3.vin2 a_20286_892# X1.X2.X3.vin1.t1 vdd.t709 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X112 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X113 a_46116_30882# d0.t10 vdd.t1351 vdd.t1350 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X114 vss.t1375 d0.t11 a_54992_30794# vss.t1374 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X115 a_49002_18540# a_48616_18540# vss.t640 vss.t639 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X116 X2.X1.X1.X1.X3.vin2 a_33976_22312# X2.X1.X1.X1.X2.X2.vout vss.t1539 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X117 a_17222_23258# a_16836_23258# vdd.t757 vdd.t756 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X118 a_16836_19446# d0.t12 vss.t1377 vss.t1376 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X119 X1.X2.X1.X2.X2.X1.X3.vin2 a_16836_8010# X1.X2.X1.X2.X2.X1.X2.vin1 vdd.t546 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X120 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X121 a_19036_31882# d1.t4 vdd.t849 vdd.t848 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X122 X2.X1.X1.X2.X1.X1.X1.vin1 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin1 vss.t146 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X123 X2.X2.X2.X1.X2.X2.X2.vin1 a_54992_17452# X2.X2.X2.X1.X2.X2.X3.vin2 vdd.t160 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X124 X1.X2.X1.X2.X1.X2.X3.vin2 a_16836_11822# X1.X2.X1.X2.X1.X2.X2.vin1 vdd.t401 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X125 X1.X1.X1.X3.vin1 a_4696_26164# X1.X1.X1.X1.X3.vin2 vss.t1415 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X126 vss.t1152 d4.t0 a_37852_18358# vss.t1151 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X127 a_48316_20446# d1.t5 vss.t875 vss.t874 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X128 X2.X1.X2.X2.X2.X2.vrefh a_40352_28888# X2.X1.X2.X2.X2.X1.X3.vin2 vss.t748 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X129 X1.X2.X2.X2.X2.X1.vout a_23126_27888# X1.X2.X2.X2.X2.X1.X3.vin2 vdd.t1112 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X130 vdd.t233 a_52792_24076# a_52406_24076# vdd.t232 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X131 X1.X1.X1.X2.X1.X2.X3.vin2 a_2196_11822# X1.X1.X1.X2.X2.vrefh vss.t158 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X132 a_19422_12822# a_19036_12822# vss.t774 vss.t773 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X133 a_49002_10916# a_48616_10916# vss.t1449 vss.t1448 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X134 vss.t654 d2.t0 a_8572_6962# vss.t653 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X135 vss.t1379 d0.t13 a_54992_4110# vss.t1378 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X136 vdd.t448 a_37852_6962# a_37466_6962# vdd.t447 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X137 a_2582_6104# a_2196_6104# vss.t1523 vss.t1522 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X138 vss.t877 d1.t6 a_8872_31700# vss.t876 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X139 vss.t656 d2.t1 a_52492_6962# vss.t655 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X140 a_2196_11822# d0.t14 vdd.t1353 vdd.t1352 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X141 X1.X1.X1.X1.X2.X1.X3.vin1 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin1 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X142 X1.X2.X2.X2.vrefh a_25712_17452# X1.X2.X2.X1.X2.X2.X3.vin2 vss.t987 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X143 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X144 X2.X2.X1.X2.X2.X1.X3.vin1 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin2 vss.t135 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X145 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X146 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X147 a_19722_7064# a_19336_7064# vss.t1060 vss.t1059 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X148 X1.X1.X2.X2.X1.X2.vout a_8572_22210# X1.X1.X2.X2.X3.vin1 vss.t1457 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X149 X1.X2.X1.X2.X1.X1.X3.vin1 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin2 vss.t225 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X150 X2.X2.X2.X2.X2.X2.vout a_52492_29834# X2.X2.X2.X2.X3.vin2 vss.t128 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X151 a_2196_6104# d0.t15 vdd.t1355 vdd.t1354 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X152 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X2.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X153 X2.X1.X2.X1.X2.X2.X3.vin2 a_39966_17452# X2.X1.X2.X2.vrefh vdd.t308 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X154 a_49002_22312# a_48616_22312# vdd.t135 vdd.t134 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X155 X1.X1.X1.X2.X2.X1.X3.vin2 a_4782_9010# X1.X1.X1.X2.X2.X1.vout vdd.t742 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X156 X1.X1.X2.X1.X1.X2.X3.vin1 a_10686_7922# X1.X1.X2.X1.X1.X2.X1.vin2 vdd.t336 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X157 vdd.t732 a_54992_26982# a_54606_26982# vdd.t731 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X158 a_31476_21352# d0.t16 vss.t1381 vss.t1380 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X159 X1.X2.X2.X2.X2.X1.X3.vin2 a_25326_28888# X1.X2.X2.X2.X2.X1.X2.vin1 vss.t899 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X160 vdd.t1357 d0.t17 a_54992_15546# vdd.t1356 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X161 vss.t1144 a_54992_25076# a_54606_25076# vss.t1143 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X162 a_46116_13728# d0.t18 vdd.t1359 vdd.t1358 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X163 vdd.t1361 d0.t19 a_25712_19358# vdd.t1360 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X164 vdd.t457 d0.t20 a_40352_28888# vdd.t456 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X165 vss.t141 a_23212_22210# a_22826_22210# vss.t140 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X166 X2.X1.X2.X1.X3.vin2 a_37852_10734# X2.X1.X2.X3.vin1 vss.t1269 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X167 a_19336_7064# d2.t2 vdd.t628 vdd.t627 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X168 X1.X2.X1.X1.X2.X2.X3.vin2 a_19422_20446# X1.X2.X1.X1.X2.X2.vout vdd.t1062 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X169 X1.X2.X2.X2.X1.X2.X2.vin1 a_25712_25076# X1.X2.X2.X2.X1.X2.X3.vin2 vdd.t1450 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X170 a_2196_17540# d0.t21 vss.t467 vss.t466 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X171 X2.X1.X2.X1.X1.X2.X3.vin1 a_39966_7922# X2.X1.X2.X1.X1.X2.X1.vin2 vdd.t951 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X172 X1.X2.X1.X3.vin1 a_19336_26164# X1.X2.X1.X1.X3.vin2 vss.t100 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X173 a_31862_23258# a_31476_23258# vdd.t678 vdd.t677 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X174 X2.X2.X1.X1.X1.X2.X3.vin1 a_48702_28070# X2.X2.X1.X1.X1.X2.vout vss.t745 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X175 X2.X2.X2.X1.X1.X2.X1.vin2 a_54992_7922# X2.X2.X2.X1.X1.X2.X3.vin1 vss.t422 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X176 X2.X2.X2.X2.X1.X1.vout a_52492_22210# X2.X2.X2.X2.X3.vin1 vdd.t843 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X177 X1.X1.X3.vin2.t3 a_8186_18358# X1.X1.X2.X3.vin1 vss.t1067 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X178 X2.X2.X1.X1.X1.X2.vrefh a_46502_30882# X2.X2.X1.X1.X1.X1.X3.vin2 vdd.t916 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X179 X1.X2.X1.X1.X2.X2.X2.vin1 a_17222_19446# X1.X2.X1.X1.X2.X2.X3.vin2 vss.t1134 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X180 X1.X1.X2.X2.X2.X2.X3.vin1 a_10686_30794# X1.X1.X2.X2.X2.X2.X1.vin2 vdd.t1182 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X181 X2.X1.X1.X1.X1.X2.X1.vin1 a_31862_28976# X2.X1.X1.X1.X1.X2.X3.vin1 vss.t491 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X182 X2.X1.X2.X2.X3.vin2 a_37466_29834# X2.X1.X2.X2.X2.X1.vout vss.t688 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X183 X2.X2.X2.X2.X2.X1.X1.vin2 a_54992_26982# X2.X2.X2.X2.X2.X1.X3.vin1 vss.t760 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X184 X2.X1.X2.X2.X1.X1.X1.vin2 a_40352_19358# X2.X1.X2.X2.X1.X1.X3.vin1 vss.t433 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X185 X1.X1.X1.X1.X3.vin1 a_4696_29936# X1.X1.X1.X1.X1.X2.vout vss.t681 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X186 vdd.t669 a_38152_8828# a_37766_8828# vdd.t668 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X187 X1.X1.X2.X2.X1.X2.X1.vin2 a_11072_23170# X1.X1.X2.X2.X1.X2.X3.vin1 vss.t766 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X188 a_33676_24258# d1.t7 vss.t879 vss.t878 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X189 X1.X2.X1.X2.X2.X2.X1.vin2 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin1 vdd.t728 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X190 X1.X1.X1.X2.X2.X1.X3.vin2 a_2196_8010# X1.X1.X1.X2.X2.X1.X2.vin1 vdd.t1162 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X191 a_34062_12822# a_33676_12822# vss.t1421 vss.t1420 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X192 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X193 vdd.t851 d1.t8 a_8872_16452# vdd.t850 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X194 a_48316_16634# d1.t9 vdd.t853 vdd.t852 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X195 vdd.t855 d1.t10 a_23512_27888# vdd.t854 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X196 X2.X2.X1.X1.X2.X2.X3.vin1 a_48702_20446# X2.X2.X1.X1.X2.X2.vout vss.t1249 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X197 X1.X2.X2.X2.X1.X2.vout a_23212_22210# X1.X2.X2.X2.X3.vin1 vss.t139 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X198 a_13696_892# d6.t0 vdd.t985 vdd.t984 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X199 X1.X2.X1.X2.X2.X2.vout a_19036_5198# X1.X2.X1.X2.X2.X2.X3.vin2 vss.t691 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X200 X2.X2.X2.X1.X2.X1.vout a_52492_14586# X2.X2.X2.X1.X3.vin2 vdd.t370 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X201 a_16836_23258# d0.t22 vdd.t459 vdd.t458 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X202 X2.X1.X2.X2.X3.vin1 a_37466_22210# X2.X1.X2.X2.X1.X2.vout vdd.t607 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X203 a_4396_5198# d1.t11 vdd.t937 vdd.t936 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X204 X1.X1.X1.X2.X1.X2.vout a_4396_12822# X1.X1.X1.X2.X1.X2.X3.vin1 vdd.t610 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X205 vss.t103 a_54992_9828# a_54606_9828# vss.t102 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X206 X1.X1.X2.X2.X3.vin2 a_8572_25982# X1.X1.X2.X3.vin2 vss.t152 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X207 a_46116_11822# d0.t23 vss.t469 vss.t468 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X208 X3.vin1.t3 a_28482_892# vout.t3 vss.t1271 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X209 vss.t86 a_25712_13640# a_25326_13640# vss.t85 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X210 X2.X2.X1.X2.vrefh X2.X2.X1.X1.X2.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X211 X1.X2.X1.X1.X1.X2.X3.vin1 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin2 vss.t312 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X212 vdd.t1146 a_11072_13640# a_10686_13640# vdd.t1145 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X213 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X214 X2.X1.X2.X2.X2.X1.X3.vin1 a_39966_26982# X2.X1.X2.X2.X2.X1.X1.vin1 vss.t495 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X215 X1.X2.X2.X2.X1.X1.X3.vin1 a_25326_19358# X1.X2.X2.X2.X1.X1.X1.vin1 vss.t550 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X216 a_31476_32788# d0.t24 vss.t471 vss.t470 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X217 X2.X1.X2.X2.X1.X2.X3.vin2 a_38152_24076# X2.X1.X2.X2.X1.X2.vout vss.t331 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X218 a_5082_7064# a_4696_7064# vss.t1274 vss.t1273 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X219 a_19036_12822# d1.t12 vss.t947 vss.t946 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X220 X2.X1.X2.X1.X1.X2.vout a_37852_6962# X2.X1.X2.X1.X3.vin1 vss.t458 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X221 X2.X2.X2.X1.X2.X2.vout a_52406_16452# X2.X2.X2.X1.X2.X2.X3.vin1 vss.t403 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X222 a_31476_17540# d0.t25 vdd.t461 vdd.t460 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X223 X1.X1.X1.X1.X2.X1.X2.vin1 a_2582_23258# X1.X1.X1.X1.X2.X1.X3.vin2 vss.t1168 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X224 a_46116_25164# d0.t26 vdd.t463 vdd.t462 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X225 vss.t1411 a_23212_25982# a_22826_25982# vss.t1410 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X226 vss.t473 d0.t27 a_25712_28888# vss.t472 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X227 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X228 X2.X2.X1.X2.X1.X2.X1.vin2 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin1 vdd.t1202 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X229 X1.X1.X1.X1.X1.X2.vout a_5082_29936# X1.X1.X1.X1.X3.vin1 vdd.t260 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X230 a_2196_28976# d0.t28 vss.t475 vss.t474 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X231 a_31476_8010# d0.t29 vss.t477 vss.t476 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X232 X1.X2.X1.X1.X3.vin1 a_19336_29936# X1.X2.X1.X1.X1.X2.vout vss.t794 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X233 vss.t949 d1.t13 a_38152_5016# vss.t948 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X234 vss.t479 d0.t30 a_40352_4110# vss.t478 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X235 X2.X1.X2.X1.X3.vin2 a_37466_14586# X2.X1.X2.X1.X2.X2.vout vdd.t1256 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X236 vdd.t326 a_25712_21264# a_25326_21264# vdd.t325 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X237 a_4696_7064# d2.t3 vdd.t630 vdd.t629 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X238 X2.X1.X1.X1.X2.X1.X3.vin2 a_34062_24258# X2.X1.X1.X1.X2.X1.vout vdd.t23 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X239 a_34062_9010# a_33676_9010# vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X240 a_31476_9916# d0.t31 vdd.t465 vdd.t464 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X241 a_4782_20446# a_4396_20446# vdd.t1402 vdd.t1401 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X242 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X243 X2.X1.X1.X2.X2.X1.X3.vin1 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin2 vss.t710 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X244 X2.X2.X2.X2.X1.X2.vout a_52406_24076# X2.X2.X2.X2.X1.X2.X3.vin2 vdd.t1131 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X245 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X246 X2.X1.X2.X2.X2.X1.vout a_37852_29834# X2.X1.X2.X2.X3.vin2 vdd.t1505 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X247 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X248 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X249 vdd.t720 a_40352_28888# a_39966_28888# vdd.t719 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X250 X1.X2.X2.X2.X3.vin2 a_23212_25982# X1.X2.X2.X3.vin2 vss.t1409 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X251 X2.X1.X1.X1.X1.X1.X3.vin2 a_31476_30882# X2.X1.X1.X1.X1.X2.vrefh vss.t410 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X252 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X253 X2.X2.X1.X2.X1.X1.X3.vin2 a_48702_16634# X2.X2.X1.X2.X1.X1.vout vdd.t1156 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X254 X2.X2.X1.X1.X1.X2.vout a_48316_28070# X2.X2.X1.X1.X1.X2.X3.vin2 vss.t1124 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X255 a_49566_892# d5.t1 vss.t38 vss.t37 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X256 X2.X2.X1.X1.X1.X1.X3.vin2 a_46116_30882# X2.X2.X1.X1.X1.X1.X2.vin1 vdd.t618 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X257 a_17222_4198# a_16836_4198# vdd.t1520 vdd.t1519 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X258 X1.X1.X2.X2.X2.X1.X3.vin1 a_8872_27888# X1.X1.X2.X2.X2.X1.vout vdd.t359 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X259 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X260 X1.X2.X2.X1.X1.X2.X3.vin1 a_25326_7922# X1.X2.X2.X1.X1.X2.X1.vin2 vdd.t143 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X261 X1.X2.X1.X1.X2.X2.vrefh a_17222_23258# X1.X2.X1.X1.X2.X1.X3.vin2 vdd.t758 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X262 a_31476_15634# d0.t32 vss.t481 vss.t480 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X263 a_34362_18540# a_33976_18540# vss.t805 vss.t804 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X264 X1.X2.X1.X1.X2.X1.vout a_19036_24258# X1.X2.X1.X1.X2.X1.X3.vin1 vdd.t139 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X265 vdd.t467 d0.t33 a_54992_6016# vdd.t466 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X266 X2.X1.X2.X1.X1.X2.X1.vin2 a_40352_7922# X2.X1.X2.X1.X1.X2.X3.vin1 vss.t1261 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X267 X2.X2.X1.X2.X1.X2.X2.vin1 a_46502_11822# X2.X2.X1.X2.X1.X2.X3.vin2 vss.t828 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X268 X2.X2.X2.X2.X2.X1.X3.vin1 a_54606_26982# X2.X2.X2.X2.X2.X1.X1.vin2 vdd.t747 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X269 X2.X2.X2.X2.X1.X2.X3.vin2 a_52792_24076# X2.X2.X2.X2.X1.X2.vout vss.t239 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X270 X1.X1.X2.X2.X1.X2.X3.vin1 a_10686_23170# X1.X1.X2.X2.X1.X2.X1.vin1 vss.t541 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X271 X2.X2.X2.X2.X1.X2.X3.vin2 a_54606_25076# X2.X2.X2.X2.X1.X2.X2.vin1 vss.t1145 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X272 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X273 X1.X2.X2.X2.X1.X1.X1.vin1 a_25712_19358# X1.X2.X2.X2.X1.X1.X3.vin1 vdd.t534 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X274 X2.X2.X1.X1.X2.X2.vout a_48316_20446# X2.X2.X1.X1.X2.X2.X3.vin2 vss.t1402 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X275 vss.t483 d0.t34 a_25712_19358# vss.t482 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X276 X2.X2.X1.X1.X3.vin1 a_48616_29936# X2.X2.X1.X1.X1.X1.vout vdd.t334 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X277 a_31476_28976# d0.t35 vdd.t469 vdd.t468 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X278 vdd.t1177 a_23512_27888# a_23126_27888# vdd.t1176 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X279 X1.X2.X2.X2.X3.vin1 a_22826_22210# X1.X2.X2.X2.X1.X1.vout vss.t343 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X280 a_17222_21352# a_16836_21352# vss.t1012 vss.t1011 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X281 X1.X2.X1.X2.X2.X2.X3.vin1 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin2 vss.t370 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X282 a_14082_892# a_13696_892# vss.t1141 vss.t1140 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X283 vss.t951 d1.t14 a_52792_16452# vss.t950 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X284 a_4396_24258# d1.t15 vdd.t939 vdd.t938 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X285 X2.X2.X1.X1.X2.X1.X1.vin2 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin1 vdd.t236 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X286 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X287 a_34362_10916# a_33976_10916# vss.t751 vss.t750 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X288 a_48702_28070# a_48316_28070# vss.t1123 vss.t1122 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X289 a_4696_26164# d3.t1 vdd.t576 vdd.t575 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X290 a_46502_30882# a_46116_30882# vdd.t617 vdd.t616 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X291 vdd.t1065 a_25712_32700# a_25326_32700# vdd.t1064 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X292 X2.X1.X2.X1.X2.X2.vrefh a_40352_13640# X2.X1.X2.X1.X2.X1.X3.vin2 vss.t1257 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X293 vss.t536 a_25712_30794# a_25326_30794# vss.t535 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X294 vss.t658 d2.t4 a_8572_14586# vss.t657 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X295 X1.X1.X2.X2.vrefh a_11072_17452# X1.X1.X2.X1.X2.X2.X3.vin2 vss.t1533 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X296 a_19336_18540# d4.t1 vss.t1154 vss.t1153 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X297 vss.t306 a_52792_27888# a_52406_27888# vss.t305 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X298 vss.t953 d1.t16 a_8872_8828# vss.t952 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X299 X2.X1.X2.X2.X1.X2.vout a_37766_24076# X2.X1.X2.X2.X1.X2.X3.vin1 vss.t1306 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X300 X2.X2.X2.X1.X1.X2.X2.vin1 a_54992_9828# X2.X2.X2.X1.X1.X2.X3.vin2 vdd.t85 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X301 vss.t955 d1.t17 a_52792_8828# vss.t954 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X302 a_34362_22312# a_33976_22312# vdd.t1529 vdd.t1528 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X303 X1.X1.X1.X1.X2.X1.X3.vin2 a_2196_23258# X1.X1.X1.X1.X2.X2.vrefh vss.t364 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X304 X1.X2.X2.X2.X2.X1.X3.vin1 a_23512_27888# X1.X2.X2.X2.X2.X1.vout vdd.t1175 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X305 X1.X1.X1.X1.X3.vin1 a_5082_26164# X1.X1.X1.X3.vin1 vss.t722 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X306 a_48702_20446# a_48316_20446# vss.t1401 vss.t1400 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X307 vdd.t941 d1.t18 a_52792_24076# vdd.t940 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X308 a_19422_24258# a_19036_24258# vss.t149 vss.t148 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X309 vss.t1408 a_11072_21264# a_10686_21264# vss.t1407 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X310 X1.X2.X2.X1.X1.X1.X1.vin2 a_25712_4110# X1.X2.X2.X1.X1.X1.X3.vin1 vss.t733 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X311 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X312 X2.X2.X1.X2.X1.X2.X3.vin1 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin1 vdd.t291 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X313 X2.X2.X1.X2.X2.X1.vout a_48316_9010# X2.X2.X1.X2.X2.X1.X3.vin2 vss.t275 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X314 vss.t526 a_38152_16452# a_37766_16452# vss.t525 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X315 X2.X1.X1.X1.X1.X2.X3.vin2 a_31476_27070# X2.X1.X1.X1.X1.X2.X2.vin1 vdd.t583 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X316 X1.X2.X2.X1.X1.X2.vout a_23212_6962# X1.X2.X2.X1.X3.vin1 vss.t905 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X317 a_19336_10916# d3.t2 vss.t586 vss.t585 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X318 X2.X1.X2.X2.X1.X1.X2.vin1 a_40352_21264# X2.X1.X2.X2.X1.X1.X3.vin2 vdd.t346 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X319 a_2582_11822# a_2196_11822# vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X320 X1.X1.X2.X2.X1.X2.X2.vin1 a_11072_25076# X1.X1.X2.X2.X1.X2.X3.vin2 vdd.t530 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X321 a_16836_9916# d0.t36 vss.t485 vss.t484 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X322 X2.X2.X2.X1.X1.X2.X3.vin2 a_54606_9828# X2.X2.X2.X1.X1.X2.X2.vin1 vss.t1048 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X323 X1.X2.X2.X1.X2.X1.X3.vin2 a_25326_13640# X1.X2.X2.X1.X2.X1.X2.vin1 vss.t314 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X324 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X325 vss.t487 d0.t37 a_40352_11734# vss.t486 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X326 X2.X1.X1.X2.X1.X1.vout a_33676_16634# X2.X1.X1.X2.X1.X1.X3.vin2 vss.t661 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X327 a_2582_4198# a_2196_4198# vdd.t1198 vdd.t1197 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X328 a_31862_21352# a_31476_21352# vss.t1164 vss.t1163 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X329 X1.X2.X2.X3.vin2 a_22826_25982# X1.X2.X2.X2.X3.vin1 vss.t285 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X330 vdd.t196 d0.t38 a_54992_26982# vdd.t195 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X331 a_19336_22312# d2.t5 vdd.t766 vdd.t765 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X332 X1.X2.X2.X2.X2.X2.vrefh a_25712_28888# X1.X2.X2.X2.X2.X1.X3.vin2 vss.t896 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X333 vss.t202 d0.t39 a_54992_25076# vss.t201 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X334 vdd.t323 a_38152_24076# a_37766_24076# vdd.t322 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X335 a_46116_8010# d0.t40 vss.t204 vss.t203 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X336 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X337 a_17222_32788# a_16836_32788# vss.t1469 vss.t1468 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X338 vdd.t919 a_54992_11734# a_54606_11734# vdd.t918 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X339 a_46502_13728# a_46116_13728# vdd.t290 vdd.t289 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X340 X2.X2.X1.X2.X1.X1.vout a_48316_16634# X2.X2.X1.X2.X1.X1.X3.vin1 vdd.t801 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X341 a_4696_22312# d2.t6 vss.t796 vss.t795 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X342 vdd.t932 a_25712_7922# a_25326_7922# vdd.t931 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X343 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X2.vrefh vss.t242 sky130_fd_pr__res_high_po_0p35 l=1.09
X344 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X345 vdd.t1093 a_25712_15546# a_25326_15546# vdd.t1092 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X346 a_17222_17540# a_16836_17540# vdd.t219 vdd.t218 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X347 vss.t798 d2.t7 a_23212_22210# vss.t797 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X348 a_2582_17540# a_2196_17540# vss.t1209 vss.t1208 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X349 X1.X2.X2.X2.X1.X1.X3.vin2 a_25326_21264# X1.X2.X2.X2.X1.X2.vrefh vdd.t70 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X350 a_48702_9010# a_48316_9010# vdd.t267 vdd.t266 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X351 X1.X1.X1.X2.X3.vin1 a_4696_14688# X1.X1.X1.X2.X1.X2.vout vss.t271 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X352 X1.X1.X1.X2.X2.X2.X3.vin1 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin2 vss.t1521 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X353 X1.X1.X2.X1.X1.X1.vout a_8486_5016# X1.X1.X2.X1.X1.X1.X3.vin1 vss.t512 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X354 X1.X1.X2.X3.vin2 a_8572_18358# X1.X1.X3.vin2.t0 vss.t419 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X355 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X356 a_33976_18540# d4.t2 vss.t1156 vss.t1155 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X357 X2.X2.X1.X3.vin1 a_48616_26164# X2.X2.X1.X1.X3.vin2 vss.t416 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X358 X2.X2.X1.X2.X1.X2.X3.vin2 a_46116_11822# X2.X2.X1.X2.X2.vrefh vss.t1305 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X359 vdd.t578 d3.t3 a_8572_25982# vdd.t577 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X360 a_17222_9916# a_16836_9916# vdd.t626 vdd.t625 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X361 X2.X1.X2.X2.X2.X2.vout a_37852_29834# X2.X1.X2.X2.X3.vin2 vss.t1515 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X362 X1.X1.X1.X1.X1.X1.vout a_5082_29936# X1.X1.X1.X1.X3.vin1 vss.t268 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X363 vdd.t198 d0.t41 a_40352_6016# vdd.t197 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X364 a_34062_24258# a_33676_24258# vss.t338 vss.t337 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X365 a_16836_21352# d0.t42 vss.t206 vss.t205 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X366 vdd.t515 a_8872_12640# a_8486_12640# vdd.t514 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X367 vss.t556 a_23212_18358# a_22826_18358# vss.t555 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X368 a_48702_16634# a_48316_16634# vdd.t800 vdd.t799 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X369 X2.X2.X1.X1.X2.X1.X3.vin1 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin1 vdd.t923 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X370 a_33976_10916# d3.t4 vss.t588 vss.t587 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X371 X2.X2.X2.X1.X1.X1.X3.vin1 a_54606_4110# X2.X2.X2.X1.X1.X1.X1.vin2 vdd.t893 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X372 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X373 X2.X2.X2.X3.vin1 a_52492_18358# X2.X2.X3.vin2 vdd.t656 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X374 X2.X1.X2.X2.X2.X2.X2.vin1 a_40352_32700# X2.X1.X2.X2.X2.X2.X3.vin2 vdd.t506 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X375 X2.X1.X2.X2.X2.X2.X1.vin2 a_40352_30794# X2.X1.X2.X2.X2.X2.X3.vin1 vss.t407 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X376 vss.t909 a_8572_14586# a_8186_14586# vss.t908 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X377 X1.X1.X2.X1.X2.X2.X3.vin2 a_10686_17452# X1.X1.X2.X1.X2.X2.X2.vin1 vss.t1270 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X378 X2.X1.X2.X2.X1.X1.vout a_37852_22210# X2.X1.X2.X2.X3.vin1 vdd.t109 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X379 vss.t208 d0.t43 a_54992_9828# vss.t207 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X380 X1.X1.X1.X2.X1.X2.X3.vin2 a_4782_12822# X1.X1.X1.X2.X1.X2.vout vdd.t253 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X381 a_46116_23258# d0.t44 vss.t210 vss.t209 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X382 vss.t212 d0.t45 a_25712_4110# vss.t211 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X383 a_46502_11822# a_46116_11822# vss.t1304 vss.t1303 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X384 vss.t214 d0.t46 a_25712_13640# vss.t213 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X385 X1.X2.X1.X1.X2.X1.X3.vin2 a_19422_24258# X1.X2.X1.X1.X2.X1.vout vdd.t66 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X386 a_17222_15634# a_16836_15634# vss.t1297 vss.t1296 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X387 vdd.t200 d0.t47 a_11072_13640# vdd.t199 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X388 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X389 a_33976_22312# d2.t8 vdd.t768 vdd.t767 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X390 X1.X2.X1.X2.X3.vin1 a_19336_14688# X1.X2.X1.X2.X1.X2.vout vss.t811 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X391 a_48616_29936# d2.t9 vdd.t770 vdd.t769 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X392 X1.X2.X1.X1.X3.vin2 a_19722_26164# X1.X2.X1.X3.vin1 vdd.t1089 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X393 X1.X2.X2.X2.X1.X1.X1.vin2 a_25712_19358# X1.X2.X2.X2.X1.X1.X3.vin1 vss.t546 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X394 a_31862_32788# a_31476_32788# vss.t791 vss.t790 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X395 a_19036_24258# d1.t19 vss.t957 vss.t956 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X396 X1.X2.X2.X3.vin2 a_23212_18358# X1.X2.X3.vin2.t0 vss.t554 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X397 X1.X2.vrefh X1.X2.X1.X1.X1.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X398 a_31862_17540# a_31476_17540# vdd.t1281 vdd.t1280 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X399 a_46502_25164# a_46116_25164# vdd.t922 vdd.t921 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X400 vss.t590 d3.t5 a_23212_25982# vss.t589 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X401 a_17222_28976# a_16836_28976# vdd.t304 vdd.t303 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X402 X2.X1.X2.X1.X1.X2.X2.vin1 a_40352_9828# X2.X1.X2.X1.X1.X2.X3.vin2 vdd.t472 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X403 a_2582_28976# a_2196_28976# vss.t347 vss.t346 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X404 X1.X1.X2.X2.X1.X2.X3.vin2 a_10686_25076# X1.X1.X2.X2.X2.vrefh vdd.t1120 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X405 X2.X1.X3.vin2.t0 a_37466_18358# X2.X1.X2.X3.vin2 vdd.t411 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X406 X1.X2.X2.X2.X2.X2.X3.vin2 a_25326_32700# X2.vrefh vdd.t1066 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X407 X2.X1.X1.X2.X2.X1.vout a_33676_9010# X2.X1.X1.X2.X2.X1.X3.vin2 vss.t30 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X408 X1.X2.X2.X2.X2.X2.X3.vin1 a_25326_30794# X1.X2.X2.X2.X2.X2.X1.vin1 vss.t1055 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X409 X1.X2.X1.X2.X2.X1.X3.vin2 a_19422_9010# X1.X2.X1.X2.X2.X1.vout vdd.t523 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X410 X2.X1.X2.X1.X2.X1.vout a_37852_14586# X2.X1.X2.X1.X3.vin2 vdd.t367 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X411 vdd.t202 d0.t48 a_25712_21264# vdd.t201 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X412 vdd.t204 d0.t49 a_40352_30794# vdd.t203 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X413 X2.X2.X2.X2.X2.X1.vout a_52406_27888# X2.X2.X2.X2.X2.X1.X3.vin1 vss.t939 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X414 X2.X2.X1.X1.X3.vin1 a_48616_29936# X2.X2.X1.X1.X1.X2.vout vss.t342 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X415 vss.t1453 a_40352_11734# a_39966_11734# vss.t1452 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X416 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X417 a_31862_9916# a_31476_9916# vdd.t682 vdd.t681 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X418 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X419 vss.t584 a_11072_15546# a_10686_15546# vss.t583 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X420 X2.X2.X1.X2.X2.X1.X3.vin2 a_48702_9010# X2.X2.X1.X2.X2.X1.vout vdd.t1203 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X421 a_16836_32788# d0.t50 vss.t216 vss.t215 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X422 X2.X1.X2.X1.X2.X2.X1.vin1 a_40352_15546# X2.X1.X2.X1.X2.X2.X3.vin1 vdd.t1426 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X423 a_16836_17540# d0.t51 vdd.t206 vdd.t205 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X424 X1.X1.X2.X2.X1.X1.X1.vin1 a_11072_19358# X1.X1.X2.X2.X1.X1.X3.vin1 vdd.t163 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X425 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X426 X1.X2.X1.X1.X2.X2.X1.vin1 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin1 vss.t1013 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X427 X2.X1.X1.X1.X1.X1.X2.vin1 a_31862_30882# X2.X1.X1.X1.X1.X1.X3.vin2 vss.t154 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X428 X1.X2.X2.X1.X1.X1.X2.vin1 a_25712_6016# X1.X2.X2.X1.X1.X1.X3.vin2 vdd.t225 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X429 a_31862_15634# a_31476_15634# vss.t1187 vss.t1186 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X430 vdd.t142 a_8572_25982# a_8186_25982# vdd.t141 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X431 X1.X2.X1.X1.X2.X1.vout a_19722_22312# X1.X2.X1.X1.X3.vin2 vss.t1223 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X432 X2.X1.X2.X1.X1.X1.X3.vin1 a_38152_5016# X2.X1.X2.X1.X1.X1.vout vdd.t698 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X433 a_16836_9916# d0.t52 vdd.t208 vdd.t207 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X434 vdd.t349 a_54992_4110# a_54606_4110# vdd.t348 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X435 X2.X2.X1.X1.X2.X1.X2.vin1 a_46502_23258# X2.X2.X1.X1.X2.X1.X3.vin2 vss.t627 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X436 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X437 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X438 a_31476_4198# d0.t53 vss.t218 vss.t217 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X439 X2.X1.X1.X2.X1.X2.vout a_34362_14688# X2.X1.X1.X2.X3.vin1 vdd.t671 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X440 X2.X1.X1.X1.X2.X2.X3.vin2 a_31476_19446# X2.X1.X1.X1.X2.X2.X2.vin1 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X441 X2.X2.X2.X1.X2.X1.X3.vin1 a_54606_11734# X2.X2.X2.X1.X2.X1.X1.vin2 vdd.t920 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X442 X2.X2.X1.X1.X1.X2.vout a_49002_29936# X2.X2.X1.X1.X3.vin1 vdd.t1027 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X443 a_31862_28976# a_31476_28976# vdd.t1409 vdd.t1408 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X444 X2.X2.X1.X2.X2.X1.X3.vin2 a_46116_8010# X2.X2.X1.X2.X2.X1.X2.vin1 vdd.t1137 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X445 X1.X2.X2.X1.X2.X2.X3.vin1 a_25326_15546# X1.X2.X2.X1.X2.X2.X1.vin2 vdd.t1094 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X446 X3.vin2.t3 a_28482_892# vout.t2 vdd.t1243 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X447 a_4782_24258# a_4396_24258# vdd.t689 vdd.t688 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X448 X1.X2.X1.X1.X1.X1.X3.vin2 a_16836_30882# X1.X2.X1.X1.X1.X2.vrefh vss.t264 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X449 X1.X1.X1.X2.X2.X2.X1.vin2 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin1 vdd.t1514 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X450 X2.X2.X2.X1.X1.X1.X3.vin2 a_54606_6016# X2.X2.X2.X1.X1.X1.X2.vin1 vss.t1063 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X451 vss.t694 a_52792_12640# a_52406_12640# vss.t693 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X452 vdd.t210 d0.t54 a_11072_7922# vdd.t209 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X453 vss.t280 a_8872_20264# a_8486_20264# vss.t279 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X454 a_5082_26164# a_4696_26164# vdd.t1399 vdd.t1398 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X455 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X456 vdd.t212 d0.t55 a_25712_32700# vdd.t211 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X457 a_48616_26164# d3.t6 vss.t592 vss.t591 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X458 vss.t610 d0.t56 a_25712_30794# vss.t609 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X459 X2.X2.X2.X1.X1.X1.X1.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X460 a_16836_15634# d0.t57 vss.t612 vss.t611 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X461 a_19722_18540# a_19336_18540# vss.t1229 vss.t1228 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X462 a_2196_30882# d0.t58 vss.t614 vss.t613 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X463 vss.t959 d1.t20 a_52792_27888# vss.t958 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X464 X1.X2.X1.X2.X2.X2.X3.vin2 a_16836_4198# X1.X2.X1.X2.X2.X2.X2.vin1 vdd.t1518 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X465 X2.X1.X1.X1.X2.X1.X3.vin1 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin2 vss.t1237 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X466 X1.X2.X2.X1.X1.X2.X3.vin2 a_23512_8828# X1.X2.X2.X1.X1.X2.vout vss.t260 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X467 X2.X2.X2.X1.X2.X1.X2.vin1 a_54992_13640# X2.X2.X2.X1.X2.X1.X3.vin2 vdd.t789 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X468 X1.X2.X3.vin2.t1 a_22826_18358# X1.X2.X2.X3.vin1 vss.t557 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X469 vss.t1260 a_40352_7922# a_39966_7922# vss.t1259 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X470 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X471 a_16836_28976# d0.t59 vdd.t588 vdd.t587 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X472 vdd.t1219 a_52792_20264# a_52406_20264# vdd.t1218 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X473 vss.t616 d0.t60 a_11072_21264# vss.t615 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X474 X1.X2.X1.X1.X1.X1.X1.vin1 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin1 vss.t662 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X475 a_19036_9010# d1.t21 vss.t961 vss.t960 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X476 X1.X1.X2.X2.X2.X2.vrefh a_11072_28888# X1.X1.X2.X2.X2.X1.X3.vin2 vss.t325 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X477 vss.t963 d1.t22 a_38152_16452# vss.t962 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X478 X1.X2.X1.X2.X1.X1.X1.vin2 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin1 vdd.t413 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X479 X2.X1.X1.X1.X2.vrefh a_31862_27070# X2.X1.X1.X1.X1.X2.X3.vin2 vdd.t424 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X480 a_20672_892# a_20286_892# vss.t737 vss.t736 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X481 a_19722_10916# a_19336_10916# vss.t721 vss.t720 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X482 X2.X2.X2.X1.X3.vin1 a_52106_6962# X2.X2.X2.X1.X1.X2.vout vdd.t1121 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X483 X2.X1.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X484 vdd.t395 a_40352_30794# a_39966_30794# vdd.t394 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X485 X1.X2.X2.X1.X2.X2.vrefh a_25712_13640# X1.X2.X2.X1.X2.X1.X3.vin2 vss.t84 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X486 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X487 X1.X3.vin2 a_14082_892# X3.vin1.t0 vdd.t237 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X488 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X489 vss.t618 d0.t61 a_40352_23170# vss.t617 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X490 vss.t1137 a_38152_27888# a_37766_27888# vss.t1136 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X491 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X492 X2.X1.X1.X2.X1.X1.X3.vin1 a_34062_16634# X2.X1.X1.X2.X1.X1.vout vss.t313 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X493 X1.X2.X1.X2.X2.X1.X1.vin2 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin1 vdd.t235 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X494 X2.X1.X2.X1.X2.X1.X3.vin2 a_39966_13640# X2.X1.X2.X1.X2.X2.vrefh vdd.t1090 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X495 X1.X1.X1.X2.X2.X2.X3.vin2 a_4782_5198# X1.X1.X1.X2.X2.X2.vout vdd.t285 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X496 a_19722_22312# a_19336_22312# vdd.t586 vdd.t585 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X497 X1.X1.X2.X1.X1.X1.X3.vin1 a_10686_4110# X1.X1.X2.X1.X1.X1.X1.vin2 vdd.t122 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X498 X1.X1.X2.X2.X1.X1.X3.vin1 a_10686_19358# X1.X1.X2.X2.X1.X1.X1.vin2 vdd.t1238 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X499 vdd.t943 d1.t23 a_38152_24076# vdd.t942 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X500 vdd.t1369 a_54992_23170# a_54606_23170# vdd.t1368 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X501 vdd.t184 a_25712_26982# a_25326_26982# vdd.t183 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X502 vdd.t590 d0.t62 a_25712_6016# vdd.t589 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X503 vdd.t592 d0.t63 a_54992_11734# vdd.t591 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X504 a_5082_22312# a_4696_22312# vss.t309 vss.t308 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X505 X1.X1.X2.X1.X1.X2.X1.vin2 a_11072_7922# X1.X1.X2.X1.X1.X2.X3.vin1 vss.t937 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X506 vss.t1466 a_25712_25076# a_25326_25076# vss.t1465 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X507 vdd.t594 d0.t64 a_25712_15546# vdd.t593 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X508 X1.X2.X1.X1.X1.X2.X3.vin2 a_16836_27070# X1.X2.X1.X1.X1.X2.X2.vin1 vdd.t190 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X509 a_33676_28070# d1.t24 vss.t965 vss.t964 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X510 X1.X2.X2.X2.X1.X1.X2.vin1 a_25712_21264# X1.X2.X2.X2.X1.X1.X3.vin2 vdd.t324 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X511 a_31476_30882# d0.t65 vdd.t596 vdd.t595 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X512 a_48616_29936# d2.t10 vss.t800 vss.t799 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X513 X2.X1.X2.X1.X1.X1.X3.vin1 a_39966_4110# X2.X1.X2.X1.X1.X1.X1.vin2 vdd.t230 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X514 X1.X1.X1.X2.X1.X1.vout a_5082_14688# X1.X1.X1.X2.X3.vin1 vss.t1128 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X515 X1.X1.X1.X1.X2.X2.X1.vin2 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin1 vdd.t1023 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X516 X2.X2.X1.X1.X2.X1.X3.vin2 a_46116_23258# X2.X2.X1.X1.X2.X2.vrefh vss.t228 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X517 X2.X2.X1.X1.X3.vin1 a_49002_26164# X2.X2.X1.X3.vin1 vss.t1258 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X518 X2.X1.X1.X2.X2.X1.X2.vin1 a_31862_8010# X2.X1.X1.X2.X2.X1.X3.vin2 vss.t641 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X519 X2.X2.X1.X2.X2.X2.vout a_48316_5198# X2.X2.X1.X2.X2.X2.X3.vin2 vss.t678 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X520 X2.X1.X1.X2.X3.vin1 a_33976_14688# X2.X1.X1.X2.X1.X1.vout vdd.t1206 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X521 vss.t1096 a_54992_6016# a_54606_6016# vss.t1095 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X522 X1.X2.X1.X2.X1.X1.X2.vin1 a_17222_15634# X1.X2.X1.X2.X1.X1.X3.vin2 vss.t1298 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X523 X1.X1.X2.X1.X2.X2.vout a_8486_16452# X1.X1.X2.X1.X2.X2.X3.vin1 vss.t982 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X524 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X525 a_2196_27070# d0.t66 vdd.t598 vdd.t597 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X526 X1.X2.X1.X2.X1.X1.vout a_19036_16634# X1.X2.X1.X2.X1.X1.X3.vin2 vss.t97 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X527 vdd.t580 d3.t7 a_8572_10734# vdd.t579 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X528 X1.X1.X1.X1.X1.X1.vout a_4396_31882# X1.X1.X1.X1.X1.X1.X3.vin2 vss.t249 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X529 X1.X1.X1.X2.X2.X2.vout a_5082_7064# X1.X1.X1.X2.X3.vin2 vdd.t1247 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X530 X2.X2.X2.X1.X1.X2.vout a_52406_8828# X2.X2.X2.X1.X1.X2.X3.vin2 vdd.t309 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X531 vss.t1158 d4.t3 a_23212_18358# vss.t1157 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X532 a_33676_20446# d1.t25 vss.t967 vss.t966 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X533 a_31862_6104# a_31476_6104# vdd.t476 vdd.t475 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X534 X1.X1.X1.X2.X2.X2.X3.vin2 a_2196_4198# X1.X1.X1.X2.X2.X2.X2.vin1 vdd.t1196 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X535 vdd.t966 d1.t26 a_8872_12640# vdd.t965 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X536 X1.X1.X2.X2.X1.X1.X1.vin2 a_11072_19358# X1.X1.X2.X2.X1.X1.X3.vin1 vss.t173 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X537 vdd.t876 a_52792_31700# a_52406_31700# vdd.t875 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X538 a_48316_12822# d1.t27 vdd.t968 vdd.t967 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X539 X1.X1.X3.vin1.t3 a_4696_18540# X1.X1.X1.X3.vin1 vdd.t1416 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X540 X1.X2.X1.X1.X1.X2.X1.vin2 a_17222_28976# X1.X2.X1.X1.X1.X2.X3.vin1 vdd.t353 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X541 vdd.t1274 a_23512_5016# a_23126_5016# vdd.t1273 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X542 X2.X1.X1.X2.X2.X1.X3.vin2 a_31476_8010# X2.X1.X1.X2.X2.X1.X2.vin1 vdd.t686 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X543 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X544 vss.t990 d1.t28 a_23512_8828# vss.t989 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X545 a_4396_16634# d1.t29 vss.t992 vss.t991 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X546 X1.X1.X1.X1.X1.X2.X2.vin1 a_2582_27070# X1.X1.X1.X1.X1.X2.X3.vin2 vss.t430 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X547 a_46116_4198# d0.t67 vss.t620 vss.t619 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X548 X1.X1.X2.X2.X1.X2.vout a_8486_24076# X1.X1.X2.X2.X1.X2.X3.vin2 vdd.t641 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X549 a_46502_23258# a_46116_23258# vss.t227 vss.t226 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X550 vss.t1294 a_25712_9828# a_25326_9828# vss.t1293 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X551 X1.X1.X1.X3.vin2 a_4696_10916# X1.X1.X1.X2.X3.vin1 vdd.t1363 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X552 a_49002_29936# a_48616_29936# vdd.t333 vdd.t332 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X553 a_34926_892# d5.t2 vss.t40 vss.t39 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X554 X1.X2.X1.X2.vrefh X1.X2.X1.X1.X2.X2.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X555 X2.X2.X2.X3.vin1 a_52106_10734# X2.X2.X2.X1.X3.vin1 vss.t1459 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X556 X1.X1.X2.X2.X2.X1.X3.vin2 a_10686_28888# X1.X1.X2.X2.X2.X1.X2.vin1 vss.t1299 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X557 vss.t1461 a_54992_32700# a_54606_32700# vss.t1460 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X558 X2.X2.X2.X1.X2.X1.vout a_52406_12640# X2.X2.X2.X1.X2.X1.X3.vin1 vss.t711 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X559 a_31476_13728# d0.t68 vdd.t600 vdd.t599 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X560 X2.X2.X1.X2.X3.vin1 a_48616_14688# X2.X2.X1.X2.X1.X2.vout vss.t284 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X561 X2.X2.X2.X2.X1.X2.vrefh a_54992_21264# X2.X2.X2.X2.X1.X1.X3.vin2 vss.t665 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X562 X1.X2.X2.X1.X2.X2.vout a_23126_16452# X1.X2.X2.X1.X2.X2.X3.vin1 vss.t646 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X563 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X564 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X565 X2.X1.X2.X3.vin1 a_37852_18358# X2.X1.X3.vin2 vdd.t416 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X566 a_34362_7064# a_33976_7064# vss.t779 vss.t778 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X567 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X568 X1.X2.X2.X2.X2.X2.X2.vin1 a_25712_32700# X1.X2.X2.X2.X2.X2.X3.vin2 vdd.t1063 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X569 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X570 X1.X2.X2.X2.X2.X2.X1.vin2 a_25712_30794# X1.X2.X2.X2.X2.X2.X3.vin1 vss.t534 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X571 X2.X1.X1.X1.X2.X2.X3.vin2 a_31476_19446# X2.X1.X1.X2.vrefh vss.t0 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X572 vss.t1213 a_40352_23170# a_39966_23170# vss.t1212 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X573 X1.X2.X3.vin1.t3 a_19336_18540# X1.X2.X1.X3.vin1 vdd.t1201 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X574 X2.X2.X1.X1.X1.X1.vout a_49002_29936# X2.X2.X1.X1.X3.vin1 vss.t1057 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X575 X2.X1.X1.X1.X1.X1.vout a_33676_31882# X2.X1.X1.X1.X1.X1.X3.vin1 vdd.t713 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X576 vss.t622 d0.t69 a_11072_15546# vss.t621 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X577 a_34062_5198# a_33676_5198# vdd.t1171 vdd.t1170 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X578 X3.vin1 a_13696_892# X1.X3.vin2 vss.t1139 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X579 a_19422_9010# a_19036_9010# vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X580 X2.X2.X2.X2.X1.X1.vout a_52406_20264# X2.X2.X2.X2.X1.X1.X3.vin2 vdd.t1220 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X581 X2.X1.X2.X2.X2.X1.X1.vin1 a_40352_26982# X2.X1.X2.X2.X2.X1.X3.vin1 vdd.t623 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X582 X1.X1.X2.X1.X1.X1.X3.vin2 a_10686_6016# X1.X1.X2.X1.X1.X1.X2.vin1 vss.t552 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X583 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X584 X1.X1.X1.X1.X1.X2.vout a_4396_28070# X1.X1.X1.X1.X1.X2.X3.vin1 vdd.t780 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X585 X2.X1.X2.X2.X2.vrefh a_40352_25076# X2.X1.X2.X2.X1.X2.X3.vin2 vss.t729 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X586 X1.X2.X2.X2.X1.X2.vout a_23126_24076# X1.X2.X2.X2.X1.X2.X3.vin2 vdd.t1442 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X587 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X588 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X1.X2.X2.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X589 a_33676_16634# d1.t30 vdd.t970 vdd.t969 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X590 vdd.t317 a_11072_28888# a_10686_28888# vdd.t316 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X591 X2.X1.X2.X2.X1.X1.X3.vin2 a_39966_21264# X2.X1.X2.X2.X1.X1.X2.vin1 vss.t197 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X592 X1.X2.X1.X3.vin2 a_19336_10916# X1.X2.X1.X2.X3.vin1 vdd.t693 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X593 X2.X2.X1.X2.X1.X2.X3.vin2 a_48702_12822# X2.X2.X1.X2.X1.X2.vout vdd.t1282 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X594 vdd.t295 a_8872_8828# a_8486_8828# vdd.t294 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X595 vss.t624 d0.t70 a_40352_17452# vss.t623 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X596 vdd.t471 a_40352_9828# a_39966_9828# vdd.t470 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X597 X2.X1.X2.X1.X1.X1.X3.vin2 a_39966_6016# X2.X1.X2.X1.X1.X1.X2.vin1 vss.t1206 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X598 X1.X1.X1.X1.X2.X2.X3.vin1 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin1 vdd.t259 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X599 vdd.t954 a_52792_8828# a_52406_8828# vdd.t953 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X600 X2.X2.X1.X2.X2.X2.X3.vin1 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin2 vss.t61 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X601 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X602 X1.X2.X2.X1.X1.X1.X3.vin1 a_25326_4110# X1.X2.X2.X1.X1.X1.X1.vin2 vdd.t1088 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X603 a_31476_11822# d0.t71 vss.t626 vss.t625 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X604 vdd.t159 a_54992_17452# a_54606_17452# vdd.t158 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X605 vdd.t741 a_8572_10734# a_8186_10734# vdd.t740 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X606 X2.X1.X1.X2.vrefh a_31862_19446# X2.X1.X1.X1.X2.X2.X3.vin2 vdd.t429 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X607 a_16836_8010# d0.t72 vdd.t602 vdd.t601 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X608 X1.X1.X2.X2.X1.X1.X3.vin1 a_10686_19358# X1.X1.X2.X2.X1.X1.X1.vin1 vss.t1266 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X609 X2.X2.X2.X2.X1.X2.X3.vin1 a_54606_23170# X2.X2.X2.X2.X1.X2.X1.vin2 vdd.t86 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X610 X1.X2.X2.X2.X2.X1.X3.vin1 a_25326_26982# X1.X2.X2.X2.X2.X1.X1.vin2 vdd.t979 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X611 X2.X1.X1.X2.X2.X2.vout a_33676_5198# X2.X1.X1.X2.X2.X2.X3.vin2 vss.t1199 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X612 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X613 X2.X1.X2.X2.X2.X2.X3.vin2 a_38152_31700# X2.X1.X2.X2.X2.X2.vout vss.t515 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X614 X1.X2.X2.X2.X1.X2.X3.vin2 a_25326_25076# X1.X2.X2.X2.X1.X2.X2.vin1 vss.t771 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X615 X1.X2.X2.X1.X2.X2.X1.vin1 a_25712_15546# X1.X2.X2.X1.X2.X2.X3.vin1 vdd.t1091 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X616 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X617 a_31476_25164# d0.t73 vdd.t604 vdd.t603 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X618 vss.t594 d3.t8 a_52492_10734# vss.t593 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X619 vdd.t1305 d0.t74 a_40352_25076# vdd.t1304 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X620 vss.t994 d1.t31 a_52792_12640# vss.t993 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X621 X1.X1.X1.X2.X1.X2.vrefh a_2582_15634# X1.X1.X1.X2.X1.X1.X3.vin2 vdd.t1019 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X622 vss.t996 d1.t32 a_23512_16452# vss.t995 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X623 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X624 vss.t998 d1.t33 a_8872_20264# vss.t997 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X625 X1.X1.X1.X1.X1.X2.X3.vin2 a_2196_27070# X1.X1.X1.X1.X2.vrefh vss.t1052 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X626 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X627 X2.X2.X3.vin1.t2 a_49952_892# X2.X3.vin2 vss.t776 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X628 a_19422_28070# a_19036_28070# vss.t945 vss.t944 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X629 X1.X1.X2.X1.X1.X2.vout a_8572_6962# X1.X1.X2.X1.X3.vin1 vss.t675 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X630 X2.X2.X2.X1.X1.X1.X1.vin2 a_54992_4110# X2.X2.X2.X1.X1.X1.X3.vin1 vss.t357 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X631 a_49002_26164# a_48616_26164# vss.t415 vss.t414 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X632 X2.X1.X2.X1.X3.vin1 a_37466_6962# X2.X1.X2.X1.X1.X2.vout vdd.t145 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X633 X1.X3.vin1 a_5646_892# X1.X1.X3.vin1.t2 vdd.t912 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X634 a_17222_30882# a_16836_30882# vdd.t256 vdd.t255 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X635 X2.X1.X2.X1.X2.vrefh a_40352_9828# X2.X1.X2.X1.X1.X2.X3.vin2 vss.t490 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X636 X1.X1.X2.X1.X1.X2.X2.vin1 a_11072_9828# X1.X1.X2.X1.X1.X2.X3.vin2 vdd.t352 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X637 X2.X2.X2.X2.X3.vin2 a_52106_29834# X2.X2.X2.X2.X2.X2.vout vdd.t516 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X638 X2.X2.X2.X1.X1.X2.vout a_52492_6962# X2.X2.X2.X1.X3.vin1 vss.t1218 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X639 X1.X1.X2.X1.X2.X2.vrefh a_11072_13640# X1.X1.X2.X1.X2.X1.X3.vin2 vss.t1176 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X640 a_2582_30882# a_2196_30882# vss.t1113 vss.t1112 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X641 X2.X3.vin2 a_49566_892# X2.X2.X3.vin1.t3 vdd.t1153 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X642 X2.X1.X1.X1.X2.X1.X1.vin1 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin1 vss.t832 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X643 a_2196_8010# d0.t75 vss.t1333 vss.t1332 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X644 a_46502_6104# a_46116_6104# vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X645 vss.t1000 d1.t34 a_8872_5016# vss.t999 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X646 X1.X2.X1.X1.X2.X2.X3.vin2 a_16836_19446# X1.X2.X1.X1.X2.X2.X2.vin1 vdd.t1526 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X647 X2.X2.X2.X2.X2.X2.vout a_52406_31700# X2.X2.X2.X2.X2.X2.X3.vin2 vdd.t606 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X648 vdd.t697 a_38152_5016# a_37766_5016# vdd.t696 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X649 X1.X2.X1.X2.X1.X1.X3.vin1 a_19422_16634# X1.X2.X1.X2.X1.X1.vout vss.t80 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X650 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X651 vss.t1002 d1.t35 a_52792_5016# vss.t1001 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X652 vdd.t972 d1.t36 a_52792_20264# vdd.t971 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X653 vss.t1268 a_37852_10734# a_37466_10734# vss.t1267 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X654 a_19422_20446# a_19036_20446# vss.t668 vss.t667 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X655 vdd.t974 d1.t37 a_23512_24076# vdd.t973 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X656 a_4782_9010# a_4396_9010# vdd.t1236 vdd.t1235 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X657 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X658 vss.t235 a_38152_12640# a_37766_12640# vss.t234 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X659 X2.X1.X1.X1.X2.X1.X3.vin2 a_31476_23258# X2.X1.X1.X1.X2.X1.X2.vin1 vdd.t676 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X660 a_2196_19446# d0.t76 vdd.t1307 vdd.t1306 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X661 X1.X1.X2.X2.X1.X1.X2.vin1 a_11072_21264# X1.X1.X2.X2.X1.X1.X3.vin2 vdd.t1392 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X662 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X663 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X664 X1.X2.X2.X1.X1.X2.X3.vin2 a_25326_9828# X1.X2.X2.X1.X1.X2.X2.vin1 vss.t1104 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X665 X2.X1.X2.X1.X2.X2.X3.vin1 a_38152_16452# X2.X1.X2.X1.X2.X2.vout vdd.t512 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X666 vss.t1004 d1.t38 a_38152_27888# vss.t1003 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X667 vss.t759 a_54992_26982# a_54606_26982# vss.t758 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X668 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X669 X1.X1.X1.X2.X1.X2.X1.vin1 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin1 vss.t368 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X670 X1.X2.X1.X1.X2.X1.X3.vin1 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin2 vss.t838 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X671 X2.X2.X2.X1.X2.X2.X1.vin2 a_54992_15546# X2.X2.X2.X1.X2.X2.X3.vin1 vss.t321 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X672 X1.X2.X1.X2.X2.X1.X2.vin1 a_17222_8010# X1.X2.X1.X2.X2.X1.X3.vin2 vss.t440 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X673 X2.X1.X1.X2.X1.X2.vout a_33676_12822# X2.X1.X1.X2.X1.X2.X3.vin2 vss.t1419 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X674 X2.X2.X2.X2.X2.X2.X3.vin2 a_52792_31700# X2.X2.X2.X2.X2.X2.vout vss.t895 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X675 X2.X2.X2.X2.X2.X2.X3.vin2 a_54606_32700# X2.X2.X2.X2.X2.X2.X2.vin1 vss.t1439 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X676 a_48616_14688# d2.t11 vss.t802 vss.t801 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X677 vdd.t1309 d0.t77 a_54992_23170# vdd.t1308 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X678 vdd.t1311 d0.t78 a_25712_26982# vdd.t1310 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X679 vdd.t1168 a_38152_20264# a_37766_20264# vdd.t1167 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X680 a_46116_21352# d0.t79 vdd.t1313 vdd.t1312 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X681 vss.t1335 d0.t80 a_25712_25076# vss.t1334 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X682 vdd.t705 a_25712_4110# a_25326_4110# vdd.t704 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X683 X2.X1.X2.X1.X1.X2.vout a_37766_8828# X2.X1.X2.X1.X1.X2.X3.vin2 vdd.t670 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X684 X2.X2.X1.X2.X1.X2.vout a_48316_12822# X2.X2.X1.X2.X1.X2.X3.vin1 vdd.t1212 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X685 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X2.vin1 vss.t257 sky130_fd_pr__res_high_po_0p35 l=1.09
X686 a_17222_13728# a_16836_13728# vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X687 vss.t1127 a_40352_17452# a_39966_17452# vss.t1126 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X688 vdd.t1254 a_25712_11734# a_25326_11734# vdd.t1253 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X689 a_34062_28070# a_33676_28070# vss.t1244 vss.t1243 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X690 a_2196_25164# d0.t81 vss.t1337 vss.t1336 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X691 a_31862_30882# a_31476_30882# vdd.t398 vdd.t397 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X692 a_49002_29936# a_48616_29936# vss.t341 vss.t340 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X693 a_48702_5198# a_48316_5198# vdd.t650 vdd.t649 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X694 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X695 a_19036_5198# d1.t39 vss.t1006 vss.t1005 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X696 X1.X2.X2.X1.X1.X1.X3.vin2 a_25326_6016# X1.X2.X2.X1.X1.X1.X2.vin1 vss.t1254 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X697 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X698 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X699 X1.X1.X2.X1.X2.X2.X3.vin2 a_8872_16452# X1.X1.X2.X1.X2.X2.vout vss.t291 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X700 vdd.t772 d2.t12 a_52492_29834# vdd.t771 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X701 X2.X1.X1.X2.X2.X2.X3.vin1 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin2 vss.t494 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X702 a_2582_27070# a_2196_27070# vdd.t1022 vdd.t1021 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X703 X2.X1.X2.X1.X2.X2.X3.vin1 a_39966_15546# X2.X1.X2.X1.X2.X2.X1.vin1 vss.t1443 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X704 X1.X1.X1.X1.X1.X1.X3.vin1 a_4782_31882# X1.X1.X1.X1.X1.X1.vout vss.t434 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X705 X2.X1.X2.X2.X2.X2.vout a_37766_31700# X2.X1.X2.X2.X2.X2.X3.vin1 vss.t1427 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X706 a_34362_29936# a_33976_29936# vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X707 vss.t1100 a_52492_10734# a_52106_10734# vss.t1099 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X708 a_34062_20446# a_33676_20446# vss.t1222 vss.t1221 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X709 a_46116_27070# d0.t82 vss.t1339 vss.t1338 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X710 X1.X1.X1.X1.X1.X1.X1.vin2 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin1 vdd.t829 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X711 vdd.t976 d1.t40 a_52792_31700# vdd.t975 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X712 vdd.t701 a_40352_25076# a_39966_25076# vdd.t700 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X713 a_48702_12822# a_48316_12822# vdd.t1211 vdd.t1210 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X714 X1.X1.X1.X2.X1.X1.X3.vin2 a_2196_15634# X1.X1.X1.X2.X1.X1.X2.vin1 vdd.t1077 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X715 X1.X1.X1.X3.vin2 a_5082_18540# X1.X1.X3.vin1.t0 vdd.t659 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X716 a_19422_16634# a_19036_16634# vdd.t79 vdd.t78 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X717 vss.t328 a_23512_16452# a_23126_16452# vss.t327 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X718 X1.X1.X2.X2.X2.X1.vout a_8486_27888# X1.X1.X2.X2.X2.X1.X3.vin1 vss.t62 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X719 X2.X2.X1.X2.X2.X2.X1.vin2 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin1 vdd.t695 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X720 vss.t936 a_11072_7922# a_10686_7922# vss.t935 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X721 a_4782_16634# a_4396_16634# vss.t1290 vss.t1289 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X722 a_19036_28070# d1.t41 vss.t1031 vss.t1030 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X723 a_34926_892# d5.t3 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X724 X1.X1.X2.X2.X2.X2.X2.vin1 a_11072_32700# X1.X1.X2.X2.X2.X2.X3.vin2 vdd.t342 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X725 a_16836_30882# d0.t83 vdd.t1315 vdd.t1314 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X726 a_49002_7064# a_48616_7064# vdd.t1510 vdd.t1509 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X727 X2.X2.X2.X1.X2.X2.X3.vin1 a_52792_16452# X2.X2.X2.X1.X2.X2.vout vdd.t390 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X728 X1.X1.X2.X2.X2.X2.X1.vin2 a_11072_30794# X1.X1.X2.X2.X2.X2.X3.vin1 vss.t523 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X729 X2.X2.X2.X1.X2.X2.X3.vin2 a_54606_17452# X2.X2.X2.X2.vrefh vdd.t268 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X730 X1.X1.X2.X2.X1.X2.X3.vin1 a_8872_24076# X1.X1.X2.X2.X1.X2.vout vdd.t1250 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X731 X1.X1.X2.X1.X2.X1.X3.vin2 a_10686_13640# X1.X1.X2.X1.X2.X1.X2.vin1 vss.t1177 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X732 X1.X1.X1.X1.X2.X2.vout a_4396_20446# X1.X1.X1.X1.X2.X2.X3.vin1 vdd.t1400 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X733 X2.X1.X2.X1.X1.X1.X1.vin2 a_40352_4110# X2.X1.X2.X1.X1.X1.X3.vin1 vss.t1066 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X734 vss.t1341 d0.t84 a_25712_9828# vss.t1340 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X735 vdd.t1504 a_37852_29834# a_37466_29834# vdd.t1503 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X736 a_17222_11822# a_16836_11822# vss.t413 vss.t412 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X737 X1.X1.X1.X2.X3.vin2 a_5082_10916# X1.X1.X1.X3.vin2 vdd.t964 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X738 vdd.t1317 d0.t85 a_40352_19358# vdd.t1316 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X739 a_19336_29936# d2.t13 vdd.t774 vdd.t773 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X740 vdd.t249 a_23512_24076# a_23126_24076# vdd.t248 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X741 a_31476_9916# d0.t86 vss.t1343 vss.t1342 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X742 a_19036_20446# d1.t42 vss.t1033 vss.t1032 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X743 vss.t1345 d0.t87 a_54992_32700# vss.t1344 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X744 vdd.t501 a_38152_31700# a_37766_31700# vdd.t500 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X745 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X746 X2.X2.X1.X2.X1.X1.vout a_49002_14688# X2.X2.X1.X2.X3.vin1 vss.t32 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X747 a_31862_13728# a_31476_13728# vdd.t194 vdd.t193 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X748 X1.X2.X2.X1.X2.X2.X3.vin2 a_23512_16452# X1.X2.X2.X1.X2.X2.vout vss.t326 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X749 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X750 a_17222_25164# a_16836_25164# vdd.t808 vdd.t807 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X751 X2.X1.X1.X2.X2.X2.X2.vin1 a_31862_4198# X2.X1.X1.X2.X2.X2.X3.vin2 vss.t322 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X752 X2.X2.X1.X1.X2.X2.X1.vin2 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin1 vdd.t361 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X753 a_4696_14688# d2.t14 vdd.t776 vdd.t775 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X754 X1.X1.X2.X2.X1.X1.X3.vin2 a_10686_21264# X1.X1.X2.X2.X1.X2.vrefh vdd.t535 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X755 X2.X1.X1.X1.X2.X2.X2.vin1 a_31862_19446# X2.X1.X1.X1.X2.X2.X3.vin2 vss.t441 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X756 vdd.t358 a_8872_27888# a_8486_27888# vdd.t357 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X757 X1.X2.X1.X2.X2.X2.X3.vin2 a_19422_5198# X1.X2.X1.X2.X2.X2.vout vdd.t1191 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X758 X2.X1.X2.X1.X2.X2.vout a_37766_16452# X2.X1.X2.X1.X2.X2.X3.vin2 vdd.t1165 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X759 X2.X2.X2.X2.X3.vin2 a_52106_29834# X2.X2.X2.X2.X2.X1.vout vss.t530 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X760 X2.X1.X1.X1.X1.X1.X3.vin2 a_34062_31882# X2.X1.X1.X1.X1.X1.vout vdd.t716 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X761 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X762 X1.X1.X1.X2.X1.X2.X3.vin1 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin2 vss.t753 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X763 X1.X2.X2.X2.X2.X1.vout a_23126_27888# X1.X2.X2.X2.X2.X1.X3.vin1 vss.t1138 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X764 vss.t238 a_52792_24076# a_52406_24076# vss.t237 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X765 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X766 vss.t1430 a_11072_11734# a_10686_11734# vss.t1429 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X767 X2.X2.X3.vin1.t0 a_48616_18540# X2.X2.X1.X3.vin1 vdd.t614 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X768 X2.X2.X2.X1.X1.X1.X2.vin1 a_54992_6016# X2.X2.X2.X1.X1.X1.X3.vin2 vdd.t1070 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X769 X1.X1.X1.X1.X1.X2.X3.vin2 a_4782_28070# X1.X1.X1.X1.X1.X2.vout vdd.t1438 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X770 X1.X2.X2.X2.X1.X2.X3.vin1 a_23512_24076# X1.X2.X2.X2.X1.X2.vout vdd.t247 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X771 X2.X2.X1.X2.X2.X2.X3.vin2 a_48702_5198# X2.X2.X1.X2.X2.X2.vout vdd.t1061 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X772 X2.X1.X2.X1.X2.X1.X1.vin1 a_40352_11734# X2.X1.X2.X1.X2.X1.X3.vin1 vdd.t1437 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X773 a_34062_16634# a_33676_16634# vdd.t633 vdd.t632 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X774 X2.X2.X1.X1.X1.X2.X2.vin1 a_46502_27070# X2.X2.X1.X1.X1.X2.X3.vin2 vss.t404 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X775 a_16836_13728# d0.t88 vdd.t1319 vdd.t1318 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X776 X1.X1.X2.X1.X2.X2.X1.vin1 a_11072_15546# X1.X1.X2.X1.X2.X2.X3.vin1 vdd.t574 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X777 vdd.t1321 d0.t89 a_11072_28888# vdd.t1320 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X778 vss.t231 a_25712_6016# a_25326_6016# vss.t230 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X779 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X780 X2.X2.X2.X2.X3.vin1 a_52106_22210# X2.X2.X2.X2.X1.X2.vout vdd.t226 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X781 a_35312_892# a_34926_892# vss.t1446 vss.t1445 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X782 a_16836_6104# d0.t90 vss.t1347 vss.t1346 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X783 X1.X2.X2.X1.X1.X2.vout a_23126_8828# X1.X2.X2.X1.X1.X2.X3.vin2 vdd.t874 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X784 X1.X2.X1.X1.X2.X2.X3.vin2 a_16836_19446# X1.X2.X1.X2.vrefh vss.t1534 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X785 X2.X2.X1.X3.vin2 a_48616_10916# X2.X2.X1.X2.X3.vin1 vdd.t1433 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X786 X2.X1.X1.X2.X3.vin2 a_33976_7064# X2.X1.X1.X2.X2.X2.vout vss.t777 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X787 X1.X2.X1.X2.X2.X2.vout a_19722_7064# X1.X2.X1.X2.X3.vin2 vdd.t1031 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X788 X1.X2.X1.X1.X1.X2.vrefh a_17222_30882# X1.X2.X1.X1.X1.X1.X3.vin2 vdd.t1143 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X789 X2.X2.X2.X2.X2.X1.X3.vin1 a_54606_26982# X2.X2.X2.X2.X2.X1.X1.vin1 vss.t775 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X790 a_31476_23258# d0.t91 vss.t1349 vss.t1348 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X791 a_34362_26164# a_33976_26164# vss.t1527 vss.t1526 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X792 X1.X2.X1.X1.X1.X1.vout a_19036_31882# X1.X2.X1.X1.X1.X1.X3.vin1 vdd.t1079 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X793 vdd.t117 a_52492_29834# a_52106_29834# vdd.t116 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X794 a_31862_11822# a_31476_11822# vss.t970 vss.t969 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X795 vdd.t372 d0.t92 a_54992_17452# vdd.t371 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X796 a_46116_15634# d0.t93 vdd.t374 vdd.t373 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X797 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X798 vss.t380 d0.t94 a_40352_28888# vss.t379 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X799 X2.X3.vin1 a_34926_892# X2.X1.X3.vin1.t3 vdd.t1428 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X800 a_33976_29936# d2.t15 vdd.t165 vdd.t164 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X801 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X802 X1.X2.X2.X2.X2.X1.X1.vin1 a_25712_26982# X1.X2.X2.X2.X2.X1.X3.vin1 vdd.t182 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X803 a_2196_19446# d0.t95 vss.t382 vss.t381 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X804 X1.X1.X1.X1.X1.X1.X3.vin1 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin1 vdd.t1082 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X805 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.X1.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X806 X1.X2.X2.X2.X2.vrefh a_25712_25076# X1.X2.X2.X2.X1.X2.X3.vin2 vss.t1464 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X807 X2.X2.X1.X2.X2.X2.vout a_49002_7064# X2.X2.X1.X2.X3.vin2 vdd.t310 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X808 X1.X2.X1.X2.X2.X1.vout a_19036_9010# X1.X2.X1.X2.X2.X1.X3.vin1 vdd.t176 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X809 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X810 X2.X2.X1.X2.X2.X2.X3.vin2 a_46116_4198# X2.X2.X1.X2.X2.X2.X2.vin1 vdd.t830 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X811 X1.X1.X2.X1.X1.X2.X3.vin2 a_8872_8828# X1.X1.X2.X1.X1.X2.vout vss.t303 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X812 a_31862_25164# a_31476_25164# vdd.t1209 vdd.t1208 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X813 X1.X2.X2.X1.X2.X1.X3.vin1 a_25326_11734# X1.X2.X2.X1.X2.X1.X1.vin2 vdd.t1255 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X814 a_19036_16634# d1.t43 vdd.t1007 vdd.t1006 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X815 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X816 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X817 a_4396_31882# d1.t44 vdd.t1009 vdd.t1008 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X818 X2.X2.X2.X1.X3.vin2 a_52106_14586# X2.X2.X2.X1.X2.X2.vout vdd.t132 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X819 X2.X2.X2.X1.X1.X2.X3.vin2 a_52792_8828# X2.X2.X2.X1.X1.X2.vout vss.t978 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X820 vdd.t376 d0.t96 a_11072_4110# vdd.t375 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X821 X1.X1.X2.X2.X2.X2.X3.vin2 a_10686_32700# X1.X2.vrefh vdd.t1071 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X822 X1.X1.X2.X2.X2.X2.X3.vin1 a_10686_30794# X1.X1.X2.X2.X2.X2.X1.vin1 vss.t1210 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X823 vss.t175 d2.t16 a_8572_22210# vss.t174 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X824 vss.t177 d2.t17 a_52492_29834# vss.t176 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X825 a_19336_26164# d3.t9 vss.t596 vss.t595 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X826 a_16836_11822# d0.t97 vss.t384 vss.t383 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X827 vdd.t420 a_40352_19358# a_39966_19358# vdd.t419 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X828 vss.t1035 d1.t45 a_23512_27888# vss.t1034 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X829 X1.X1.X1.X2.X2.X1.vout a_4396_9010# X1.X1.X1.X2.X2.X1.X3.vin2 vss.t1264 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X830 X2.X1.X1.X1.X2.X2.X3.vin1 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin2 vss.t1162 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X831 X1.X2.X2.X1.X1.X1.X3.vin2 a_23512_5016# X1.X2.X2.X1.X1.X1.vout vss.t1302 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X832 a_42976_892# d6.t1 vss.t1015 vss.t1014 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X833 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X834 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X835 vss.t598 d3.t10 a_37852_10734# vss.t597 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X836 a_16836_25164# d0.t98 vdd.t378 vdd.t377 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X837 X2.X2.X2.X1.X2.X2.vout a_52492_14586# X2.X2.X2.X1.X3.vin2 vss.t378 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X838 X2.X2.X1.X1.X2.X2.X3.vin1 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin1 vdd.t215 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X839 vdd.t167 d2.t18 a_23212_6962# vdd.t166 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X840 vss.t1037 d1.t46 a_38152_12640# vss.t1036 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X841 X1.X2.X1.X2.X1.X2.X1.vin2 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin1 vdd.t155 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X842 X2.X1.X1.X1.X2.X2.vrefh a_31862_23258# X2.X1.X1.X1.X2.X1.X3.vin2 vdd.t679 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X843 a_46116_13728# d0.t99 vss.t386 vss.t385 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X844 a_2582_19446# a_2196_19446# vdd.t805 vdd.t804 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X845 vdd.t169 d2.t19 a_52492_22210# vdd.t168 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X846 a_34362_29936# a_33976_29936# vss.t193 vss.t192 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X847 vdd.t508 a_11072_30794# a_10686_30794# vdd.t507 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X848 X1.X2.X2.X1.X2.vrefh a_25712_9828# X1.X2.X2.X1.X1.X2.X3.vin2 vss.t1292 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X849 vss.t674 a_8572_6962# a_8186_6962# vss.t673 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X850 vss.t1514 a_37852_29834# a_37466_29834# vss.t1513 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X851 vss.t388 d0.t100 a_54992_26982# vss.t387 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X852 a_46116_9916# d0.t101 vss.t390 vss.t389 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X853 vss.t392 d0.t102 a_40352_19358# vss.t391 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X854 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X855 X2.X1.X1.X1.X2.X1.vout a_33676_24258# X2.X1.X1.X1.X2.X1.X3.vin2 vss.t336 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X856 vdd.t351 a_11072_9828# a_10686_9828# vdd.t350 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X857 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X858 vss.t1217 a_52492_6962# a_52106_6962# vss.t1216 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X859 X2.X1.X1.X2.X1.X2.X3.vin1 a_34062_12822# X2.X1.X1.X2.X1.X2.vout vss.t253 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X860 X1.X2.X1.X2.X1.X2.vout a_19722_14688# X1.X2.X1.X2.X3.vin1 vdd.t1024 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X861 X2.X2.X1.X2.X1.X2.vrefh a_46502_15634# X2.X2.X1.X2.X1.X1.X3.vin2 vdd.t245 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X862 a_6032_892# a_5646_892# vss.t922 vss.t921 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X863 a_49002_14688# a_48616_14688# vss.t283 vss.t282 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X864 X1.X1.X2.X1.X2.X2.X3.vin1 a_10686_15546# X1.X1.X2.X1.X2.X2.X1.vin2 vdd.t156 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X865 X2.X2.X1.X1.X1.X2.X3.vin2 a_46116_27070# X2.X2.X1.X1.X2.vrefh vss.t1171 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X866 vdd.t1011 d1.t47 a_38152_20264# vdd.t1010 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X867 a_46502_21352# a_46116_21352# vdd.t214 vdd.t213 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X868 X2.X1.X2.X1.X1.X1.X2.vin1 a_40352_6016# X2.X1.X2.X1.X1.X1.X3.vin2 vdd.t151 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X869 X2.X1.X2.X1.X3.vin2 a_37466_14586# X2.X1.X2.X1.X2.X1.vout vss.t1284 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X870 vdd.t884 a_25712_23170# a_25326_23170# vdd.t883 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X871 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X872 vdd.t380 d0.t103 a_25712_11734# vdd.t379 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X873 X2.X2.X2.X2.X2.X1.X2.vin1 a_54992_28888# X2.X2.X2.X2.X2.X1.X3.vin2 vdd.t1040 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X874 a_2196_4198# d0.t104 vss.t394 vss.t393 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X875 a_2582_25164# a_2196_25164# vss.t75 vss.t74 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X876 vdd.t171 d2.t20 a_52492_14586# vdd.t170 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X877 X1.X2.X1.X1.X2.X1.X3.vin2 a_16836_23258# X1.X2.X1.X1.X2.X1.X2.vin1 vdd.t755 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X878 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X879 vdd.t108 a_37852_22210# a_37466_22210# vdd.t107 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X880 a_48316_31882# d1.t48 vss.t1039 vss.t1038 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X881 vss.t600 d3.t11 a_8572_25982# vss.t599 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X882 a_33976_26164# d3.t12 vss.t602 vss.t601 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X883 a_19336_29936# d2.t21 vss.t179 vss.t178 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X884 X2.X2.X2.X2.X1.X2.vout a_52406_24076# X2.X2.X2.X2.X1.X2.X3.vin1 vss.t1161 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X885 a_46116_32788# d0.t105 vdd.t382 vdd.t381 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X886 X1.X1.X2.X3.vin1 a_8186_10734# X1.X1.X2.X1.X3.vin1 vss.t1148 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X887 a_48616_18540# d4.t4 vdd.t1126 vdd.t1125 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X888 vss.t747 a_40352_28888# a_39966_28888# vss.t746 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X889 X1.X2.X1.X2.X3.vin2 a_19336_7064# X1.X2.X1.X2.X2.X2.vout vss.t1058 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X890 X1.X1.X2.X1.X2.X1.vout a_8486_12640# X1.X1.X2.X1.X2.X1.X3.vin1 vss.t125 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X891 X2.X1.X1.X1.X1.X1.X3.vin1 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin2 vss.t789 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X892 X1.X2.X1.X2.X1.X2.X2.vin1 a_17222_11822# X1.X2.X1.X2.X1.X2.X3.vin2 vss.t561 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X893 a_2196_23258# d0.t106 vdd.t384 vdd.t383 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X894 X1.X2.X1.X2.X1.X2.vout a_19036_12822# X1.X2.X1.X2.X1.X2.X3.vin2 vss.t772 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X895 X2.X1.X1.X2.X1.X1.X3.vin1 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin1 vdd.t1279 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X896 a_46502_27070# a_46116_27070# vss.t1170 vss.t1169 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X897 a_17222_6104# a_16836_6104# vdd.t364 vdd.t363 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X898 X1.X1.X2.X2.X2.X1.X3.vin2 a_8872_27888# X1.X1.X2.X2.X2.X1.vout vss.t367 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X899 X1.X2.X1.X1.X2.X1.X1.vin2 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin1 vdd.t1107 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X900 X2.X1.X1.X2.X2.X2.vout a_34362_7064# X2.X1.X1.X2.X3.vin2 vdd.t331 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X901 X2.X1.X2.X2.X2.X1.X3.vin2 a_39966_28888# X2.X1.X2.X2.X2.X2.vrefh vdd.t63 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X902 X2.X2.X2.X2.X3.vin1 a_52492_25982# X2.X2.X2.X3.vin2 vdd.t674 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X903 X2.X1.X1.X2.X2.X2.X3.vin2 a_31476_4198# X2.X1.X1.X2.X2.X2.X2.vin1 vdd.t121 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X904 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X905 vdd.t386 d0.t107 a_54992_7922# vdd.t385 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X906 vss.t396 d0.t108 a_11072_6016# vss.t395 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X907 a_48616_10916# d3.t13 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X908 vdd.t366 a_37852_14586# a_37466_14586# vdd.t365 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X909 X1.X2.X1.X2.X2.X2.X2.vin1 a_17222_4198# X1.X2.X1.X2.X2.X2.X3.vin2 vss.t94 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X910 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X1.X2.X1.X1.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X911 a_4396_12822# d1.t49 vss.t1041 vss.t1040 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X912 vss.t1043 d1.t50 a_23512_5016# vss.t1042 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X913 X2.X2.X1.X2.X1.X2.X1.vin1 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin1 vss.t1230 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X914 vss.t1456 a_8572_22210# a_8186_22210# vss.t1455 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X915 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X916 X2.X1.X1.X2.X2.X1.X3.vin1 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin1 vdd.t680 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X917 X1.X1.X1.X1.X2.X2.X3.vin2 a_4782_20446# X1.X1.X1.X1.X2.X2.vout vdd.t1454 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X918 vss.t127 a_52492_29834# a_52106_29834# vss.t126 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X919 X1.X1.X2.X2.X1.X1.vout a_8486_20264# X1.X1.X2.X2.X1.X1.X3.vin2 vdd.t273 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X920 a_33676_9010# d1.t51 vss.t1045 vss.t1044 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X921 vss.t1205 a_23512_27888# a_23126_27888# vss.t1204 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X922 a_17222_23258# a_16836_23258# vss.t785 vss.t784 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X923 X1.X2.X1.X1.X1.X1.X3.vin2 a_19422_31882# X1.X2.X1.X1.X1.X1.vout vdd.t284 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X924 vdd.t173 d2.t22 a_37852_29834# vdd.t172 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X925 a_19722_29936# a_19336_29936# vdd.t763 vdd.t762 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X926 vdd.t1013 d1.t52 a_38152_31700# vdd.t1012 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X927 vss.t1091 a_25712_32700# a_25326_32700# vss.t1090 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X928 X1.X2.X2.X1.X2.X1.vout a_23126_12640# X1.X2.X2.X1.X2.X1.X3.vin1 vss.t1516 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X929 a_5082_14688# a_4696_14688# vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X930 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X931 vdd.t842 a_52492_22210# a_52106_22210# vdd.t841 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X932 X2.X1.X2.X3.vin2 a_37466_25982# X2.X1.X2.X2.X3.vin2 vdd.t1067 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X933 vdd.t1015 d1.t53 a_8872_27888# vdd.t1014 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X934 a_33976_29936# d2.t23 vss.t181 vss.t180 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X935 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X936 X2.X1.X1.X2.X1.X1.X3.vin2 a_31476_15634# X2.X1.X1.X2.X1.X2.vrefh vss.t1185 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X937 X2.X1.X1.X3.vin1 a_34362_18540# X2.X1.X3.vin1 vss.t938 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X938 a_48316_28070# d1.t54 vdd.t1017 vdd.t1016 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X939 X2.X2.X1.X1.X1.X1.X3.vin1 a_48702_31882# X2.X2.X1.X1.X1.X1.vout vss.t435 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X940 vss.t432 a_40352_19358# a_39966_19358# vss.t431 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X941 X1.X2.X2.X2.X2.X1.X3.vin2 a_23512_27888# X1.X2.X2.X2.X2.X1.vout vss.t1203 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X942 vss.t1047 d1.t55 a_52792_24076# vss.t1046 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X943 vss.t765 a_11072_23170# a_10686_23170# vss.t764 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X944 X2.X2.X1.X1.X1.X1.X1.vin2 a_46502_32788# X2.X2.X1.X1.X1.X1.X3.vin1 vdd.t1213 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X945 vss.t398 d0.t109 a_11072_11734# vss.t397 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X946 X2.X2.X1.X2.X1.X1.X3.vin2 a_46116_15634# X2.X2.X1.X2.X1.X1.X2.vin1 vdd.t280 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X947 X2.X2.X1.X3.vin2 a_49002_18540# X2.X2.X3.vin1.t1 vdd.t729 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X948 a_19422_5198# a_19036_5198# vdd.t663 vdd.t662 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X949 X2.X1.X1.X1.X1.X2.X3.vin1 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin1 vdd.t1407 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X950 vdd.t175 d2.t24 a_37852_6962# vdd.t174 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X951 vss.t1065 a_40352_4110# a_39966_4110# vss.t1064 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X952 X2.X1.X2.X2.X1.X2.X1.vin1 a_40352_23170# X2.X1.X2.X2.X1.X2.X3.vin1 vdd.t1185 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X953 X1.X1.X2.X2.X2.X1.X1.vin1 a_11072_26982# X1.X1.X2.X2.X2.X1.X3.vin1 vdd.t915 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X954 X1.X1.X1.X1.X2.X1.vout a_4396_24258# X1.X1.X1.X1.X2.X1.X3.vin1 vdd.t687 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X955 X1.X2.X2.X2.X1.X1.vout a_23126_20264# X1.X2.X2.X2.X1.X1.X3.vin2 vdd.t22 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X956 X1.X1.X1.X2.X2.X1.X2.vin1 a_2582_8010# X1.X1.X1.X2.X2.X1.X3.vin2 vss.t429 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X957 X1.X1.X2.X2.X2.vrefh a_11072_25076# X1.X1.X2.X2.X1.X2.X3.vin2 vss.t544 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X958 X2.X1.X1.X2.X3.vin1 a_34362_10916# X2.X1.X1.X3.vin2 vss.t752 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X959 a_33676_12822# d1.t56 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X960 X1.X1.X1.X3.vin1 a_4696_26164# X1.X1.X1.X1.X3.vin1 vdd.t1397 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X961 vdd.t369 a_52492_14586# a_52106_14586# vdd.t368 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X962 X1.X1.X2.X2.X3.vin2 a_8186_29834# X1.X1.X2.X2.X2.X2.vout vdd.t1396 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X963 a_28482_892# a_28096_892# vdd.t551 vdd.t550 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X964 vss.t1072 d0.t110 a_40352_13640# vss.t1071 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X965 vss.t151 a_8572_25982# a_8186_25982# vss.t150 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X966 a_2582_6104# a_2196_6104# vdd.t1513 vdd.t1512 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X967 X2.X2.X1.X2.X3.vin2 a_49002_10916# X2.X2.X1.X3.vin2 vdd.t1410 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X968 X1.X1.X2.X2.X2.X2.vout a_8486_31700# X1.X1.X2.X2.X2.X2.X3.vin2 vdd.t619 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X969 a_31862_23258# a_31476_23258# vss.t706 vss.t705 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X970 vss.t330 a_38152_24076# a_37766_24076# vss.t329 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X971 a_46502_15634# a_46116_15634# vdd.t279 vdd.t278 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X972 vdd.t788 a_54992_13640# a_54606_13640# vdd.t787 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X973 X2.X1.X1.X1.X2.X2.vout a_34362_22312# X2.X1.X1.X1.X3.vin2 vdd.t786 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X974 vdd.t963 a_25712_17452# a_25326_17452# vdd.t962 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X975 a_19722_7064# a_19336_7064# vdd.t1030 vdd.t1029 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X976 a_2582_19446# a_2196_19446# vss.t835 vss.t834 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X977 a_16836_4198# d0.t111 vdd.t1042 vdd.t1041 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X978 X2.X2.X3.vin2 a_52106_18358# X2.X2.X2.X3.vin2 vdd.t657 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X979 X1.X2.X2.X2.X1.X2.X3.vin1 a_25326_23170# X1.X2.X2.X2.X1.X2.X1.vin2 vdd.t1285 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X980 X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X981 X1.X2.X2.X1.X2.X1.X1.vin1 a_25712_11734# X1.X2.X2.X1.X2.X1.X3.vin1 vdd.t1252 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X982 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X983 X1.X1.X2.X1.X1.X1.X1.vin2 a_11072_4110# X1.X1.X2.X1.X1.X1.X3.vin1 vss.t138 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X984 a_4782_31882# a_4396_31882# vdd.t244 vdd.t243 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X985 vdd.t1044 d0.t112 a_40352_21264# vdd.t1043 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X986 X1.X1.X1.X2.X2.vrefh a_2582_11822# X1.X1.X1.X2.X1.X2.X3.vin2 vdd.t292 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X987 X2.X2.X1.X2.X1.X2.X3.vin1 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin2 vss.t299 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X988 vss.t44 d1.t57 a_23512_12640# vss.t43 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X989 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X990 vdd.t35 d1.t58 a_38152_8828# vdd.t34 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X991 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X992 vdd.t1046 d0.t113 a_40352_7922# vdd.t1045 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X993 X1.X2.X1.X3.vin1 a_19336_26164# X1.X2.X1.X1.X3.vin1 vdd.t82 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X994 a_19722_26164# a_19336_26164# vss.t99 vss.t98 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X995 a_16836_23258# d0.t114 vss.t1074 vss.t1073 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X996 X2.X2.X1.X1.X1.X2.X3.vin2 a_48702_28070# X2.X2.X1.X1.X1.X2.vout vdd.t717 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X997 X1.X1.X2.X1.X2.vrefh a_11072_9828# X1.X1.X2.X1.X1.X2.X3.vin2 vss.t360 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X998 X2.X1.X1.X1.X2.X2.X1.vin1 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin1 vss.t637 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X999 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1000 X2.X1.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1001 a_14082_892# a_13696_892# vdd.t1115 vdd.t1114 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1002 X1.X2.X1.X2.X1.X2.X3.vin1 a_19422_12822# X1.X2.X1.X2.X1.X2.vout vss.t703 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1003 X1.X1.X1.X1.X3.vin2 a_4696_22312# X1.X1.X1.X1.X2.X2.vout vss.t307 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1004 X2.X2.X2.X1.X1.X1.vout a_52406_5016# X2.X2.X2.X1.X1.X1.X3.vin2 vdd.t1142 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1005 X2.X2.vrefh a_40352_32700# X2.X1.X2.X2.X2.X2.X3.vin2 vss.t520 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1006 X2.X1.X2.X1.X1.X1.X1.vin1 X2.X1.X2.vrefh.t1 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1007 X1.X2.X2.X2.X2.X2.vout a_23126_31700# X1.X2.X2.X2.X2.X2.X3.vin2 vdd.t1149 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1008 a_34362_14688# a_33976_14688# vss.t1234 vss.t1233 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1009 a_4782_5198# a_4396_5198# vdd.t950 vdd.t949 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1010 X1.X1.X1.X2.X1.X1.X1.vin1 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin1 vss.t1312 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1011 vdd.t37 d1.t59 a_23512_20264# vdd.t36 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1012 a_46502_13728# a_46116_13728# vss.t298 vss.t297 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1013 a_48316_9010# d1.t60 vss.t46 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1014 vss.t1160 d4.t5 a_8572_18358# vss.t1159 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1015 X2.X1.X3.vin1 a_33976_18540# X2.X1.X1.X3.vin2 vss.t803 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1016 X2.X2.X1.X1.X1.X1.vout a_48316_31882# X2.X2.X1.X1.X1.X1.X3.vin2 vss.t540 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1017 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1018 vdd.t1048 d0.t115 a_11072_30794# vdd.t1047 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1019 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1020 X2.X2.X1.X1.X1.X1.X3.vin1 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin1 vdd.t181 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1021 X2.X1.X2.X1.X2.X1.X3.vin1 a_38152_12640# X2.X1.X2.X1.X2.X1.vout vdd.t229 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1022 vss.t64 d2.t25 a_37852_29834# vss.t63 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1023 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1024 X1.X2.X2.X1.X3.vin1 a_22826_6962# X1.X2.X2.X1.X1.X1.vout vss.t839 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1025 X2.X1.X1.X1.X2.X1.X3.vin1 a_34062_24258# X2.X1.X1.X1.X2.X1.vout vss.t34 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1026 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1027 X2.X2.X2.X1.X2.X1.X1.vin2 a_54992_11734# X2.X2.X2.X1.X2.X1.X3.vin1 vss.t929 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1028 X1.X2.X1.X1.X2.X2.X3.vin1 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin2 vss.t1010 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1029 vss.t190 a_25712_26982# a_25326_26982# vss.t189 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1030 X2.X3.vin2 a_43362_892# X3.vin2.t1 vdd.t1150 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1031 a_31862_8010# a_31476_8010# vss.t714 vss.t713 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1032 X1.X1.X2.X2.X2.X1.X3.vin1 a_10686_26982# X1.X1.X2.X2.X2.X1.X1.vin2 vdd.t977 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1033 X1.X1.X2.X2.X1.X2.X3.vin2 a_10686_25076# X1.X1.X2.X2.X1.X2.X2.vin1 vss.t1146 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1034 X1.X2.X2.X2.X2.X2.X3.vin2 a_25326_32700# X1.X2.X2.X2.X2.X2.X2.vin1 vss.t1092 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1035 X2.X1.X1.X3.vin2 a_33976_10916# X2.X1.X1.X2.X3.vin2 vss.t749 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1036 a_19336_14688# d2.t26 vss.t66 vss.t65 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1037 X2.X1.X2.X1.X2.X2.vout a_37852_14586# X2.X1.X2.X1.X3.vin2 vss.t375 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1038 vdd.t1128 d4.t6 a_52492_18358# vdd.t1127 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1039 vdd.t1050 d0.t116 a_25712_23170# vdd.t1049 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1040 vdd.t1052 d0.t117 a_40352_32700# vdd.t1051 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1041 a_5082_7064# a_4696_7064# vdd.t1246 vdd.t1245 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1042 vss.t1076 d0.t118 a_40352_30794# vss.t1075 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1043 vss.t1256 a_40352_13640# a_39966_13640# vss.t1255 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1044 X1.X1.X1.X2.X2.X2.vout a_4396_5198# X1.X1.X1.X2.X2.X2.X3.vin2 vss.t972 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1045 X2.X1.X1.X2.X2.X1.X1.vin1 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin1 vss.t240 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1046 vss.t1532 a_11072_17452# a_10686_17452# vss.t1531 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1047 a_2196_21352# d0.t119 vss.t1078 vss.t1077 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1048 vdd.t51 d2.t27 a_37852_22210# vdd.t50 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1049 a_48702_31882# a_48316_31882# vss.t539 vss.t538 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1050 a_43362_892# a_42976_892# vss.t1202 vss.t1201 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1051 X1.X2.X1.X1.X3.vin2 a_19336_22312# X1.X2.X1.X1.X2.X2.vout vss.t608 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1052 a_31476_8010# d0.t120 vdd.t1054 vdd.t1053 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1053 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1054 a_19722_29936# a_19336_29936# vss.t793 vss.t792 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1055 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1056 a_46502_32788# a_46116_32788# vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1057 a_49952_892# a_49566_892# vss.t1183 vss.t1182 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1058 X1.X1.X2.X1.X3.vin2 a_8572_10734# X1.X1.X2.X3.vin1 vss.t769 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1059 X2.X1.X2.X1.X2.X2.X2.vin1 a_40352_17452# X2.X1.X2.X1.X2.X2.X3.vin2 vdd.t1101 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1060 a_49002_18540# a_48616_18540# vdd.t613 vdd.t612 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1061 X2.X1.X1.X1.X3.vin2 a_33976_22312# X2.X1.X1.X1.X2.X1.vout vdd.t1527 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1062 X1.X2.X1.X1.X2.X1.X2.vin1 a_17222_23258# X1.X2.X1.X1.X2.X1.X3.vin2 vss.t786 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1063 X2.X1.X1.X1.X1.X1.X1.vin1 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin1 vss.t335 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1064 X1.X2.X1.X1.X2.X1.vout a_19036_24258# X1.X2.X1.X1.X2.X1.X3.vin2 vss.t147 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1065 X1.X1.X2.X1.X2.X1.X3.vin2 a_8872_12640# X1.X1.X2.X1.X2.X1.vout vss.t529 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1066 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1067 a_2582_23258# a_2196_23258# vdd.t356 vdd.t355 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1068 X2.X1.X2.X1.X2.X1.X3.vin1 a_39966_11734# X2.X1.X2.X1.X2.X1.X1.vin1 vss.t1253 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1069 X2.X1.X1.X2.X1.X1.X1.vin2 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin1 vdd.t136 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1070 X1.X1.X2.X1.X3.vin1 a_8186_6962# X1.X1.X2.X1.X1.X2.vout vdd.t1251 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1071 vss.t664 a_54992_21264# a_54606_21264# vss.t663 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1072 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1073 a_48316_20446# d1.t61 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1074 vdd.t345 a_40352_21264# a_39966_21264# vdd.t344 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1075 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1076 vss.t454 a_23212_10734# a_22826_10734# vss.t453 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1077 X1.X1.X1.X2.X1.X2.X3.vin2 a_2196_11822# X1.X1.X1.X2.X1.X2.X2.vin1 vdd.t146 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1078 vdd.t41 d1.t62 a_23512_31700# vdd.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1079 X1.X1.X1.X1.X1.X2.X1.vin1 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin1 vss.t562 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1080 vdd.t529 a_11072_25076# a_10686_25076# vdd.t528 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1081 vdd.t415 a_37852_18358# a_37466_18358# vdd.t414 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1082 X1.X2.X2.X1.X1.X2.X1.vin1 a_25712_7922# X1.X2.X2.X1.X1.X2.X3.vin1 vdd.t930 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1083 X2.X3.vin1 a_34926_892# X2.X1.X3.vin2.t4 vss.t1444 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1084 X1.X1.X2.X2.X3.vin2 a_8186_29834# X1.X1.X2.X2.X2.X1.vout vss.t1412 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1085 vss.t533 a_23512_12640# a_23126_12640# vss.t532 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1086 a_19422_12822# a_19036_12822# vdd.t746 vdd.t745 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1087 a_49002_10916# a_48616_10916# vdd.t1432 vdd.t1431 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1088 vdd.t53 d2.t28 a_37852_14586# vdd.t52 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1089 a_4396_24258# d1.t63 vss.t48 vss.t47 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1090 vdd.t287 a_8872_5016# a_8486_5016# vdd.t286 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1091 vdd.t150 a_40352_6016# a_39966_6016# vdd.t149 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1092 a_4782_12822# a_4396_12822# vss.t632 vss.t631 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1093 X2.X2.X2.X1.X3.vin1 a_52492_10734# X2.X2.X2.X3.vin1 vdd.t1074 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1094 vdd.t1223 a_52792_5016# a_52406_5016# vdd.t1222 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1095 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1096 X2.X2.X2.X1.X2.X1.X3.vin1 a_52792_12640# X2.X2.X2.X1.X2.X1.vout vdd.t666 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1097 X2.X2.X1.X1.X1.X2.vout a_48316_28070# X2.X2.X1.X1.X1.X2.X3.vin1 vdd.t1098 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1098 X2.X1.X1.X2.X2.X1.X1.vin2 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin1 vdd.t234 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1099 X1.X1.X2.X1.X1.X2.X3.vin2 a_10686_9828# X1.X1.X2.X1.X1.X2.X2.vin1 vss.t222 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1100 X2.X2.X2.X1.X2.X1.X3.vin2 a_54606_13640# X2.X2.X2.X1.X2.X2.vrefh vdd.t1283 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1101 X1.X1.X2.X2.X1.X1.X3.vin1 a_8872_20264# X1.X1.X2.X2.X1.X1.vout vdd.t272 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1102 X1.X2.X2.X1.X2.X2.X3.vin2 a_25326_17452# X1.X2.X2.X2.vrefh vdd.t978 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1103 X1.X2.X1.X1.X1.X1.X3.vin1 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin2 vss.t1467 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1104 X2.X2.X2.X1.X1.X2.X3.vin1 a_54606_7922# X2.X2.X2.X1.X1.X2.X1.vin1 vss.t1463 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1105 vdd.t1056 d0.t121 a_40352_15546# vdd.t1055 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1106 X1.X2.X1.X2.X1.X1.X3.vin1 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin1 vdd.t217 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1107 X1.X1.X2.X2.X3.vin1 a_8186_22210# X1.X1.X2.X2.X1.X2.vout vdd.t307 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1108 a_33976_14688# d2.t29 vss.t68 vss.t67 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1109 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1110 X1.X2.X2.X1.X3.vin2 a_23212_10734# X1.X2.X2.X3.vin1 vss.t452 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1111 X1.X1.X1.X2.X1.X1.X3.vin1 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin2 vss.t1207 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1112 vdd.t644 a_23512_20264# a_23126_20264# vdd.t643 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1113 a_31476_21352# d0.t122 vdd.t1058 vdd.t1057 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1114 X2.X2.X2.vrefh.t0 X2.X2.X1.X2.X2.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1115 vss.t1080 d0.t123 a_25712_32700# vss.t1079 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1116 X1.X2.X2.X1.X2.X1.X3.vin2 a_23512_12640# X1.X2.X2.X1.X2.X1.vout vss.t531 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1117 vss.t904 a_23212_6962# a_22826_6962# vss.t903 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1118 X2.X1.X2.X2.X3.vin1 a_37852_25982# X2.X1.X2.X3.vin2 vdd.t712 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1119 X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X2.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1120 vss.t418 a_8572_18358# a_8186_18358# vss.t417 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1121 a_2196_32788# d0.t124 vss.t1082 vss.t1081 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1122 X1.X2.X1.X2.X2.X2.X3.vin1 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin1 vdd.t362 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1123 X2.X1.X2.X3.vin1 a_37466_10734# X2.X1.X2.X1.X3.vin2 vdd.t455 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1124 X2.X1.X1.X2.X1.X1.X2.vin1 a_31862_15634# X2.X1.X1.X2.X1.X1.X3.vin2 vss.t399 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1125 a_2196_17540# d0.t125 vdd.t1060 vdd.t1059 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1126 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1127 a_48702_28070# a_48316_28070# vdd.t1097 vdd.t1096 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1128 X1.X2.X1.X2.X2.X1.X3.vin1 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin1 vdd.t624 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1129 X2.X1.X2.X1.X2.X1.vout a_37766_12640# X2.X1.X2.X1.X2.X1.X3.vin2 vdd.t72 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1130 X1.X1.X2.X1.X1.X1.X2.vin1 a_11072_6016# X1.X1.X2.X1.X1.X1.X3.vin2 vdd.t735 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1131 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1132 X1.X1.X2.X1.X1.X2.vout a_8486_8828# X1.X1.X2.X1.X1.X2.X3.vin2 vdd.t539 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1133 X2.X2.X2.X2.X2.X2.X1.vin1 a_54992_30794# X2.X2.X2.X2.X2.X2.X3.vin1 vdd.t113 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1134 X2.X1.X2.X2.X2.X1.X1.vin2 a_40352_26982# X2.X1.X2.X2.X2.X1.X3.vin1 vss.t649 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1135 vss.t1084 d0.t126 a_11072_23170# vss.t1083 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1136 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1137 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1138 X1.X1.X2.X1.X3.vin2 a_8186_14586# X1.X1.X2.X1.X2.X2.vout vdd.t531 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1139 X2.X1.X1.X1.X1.X2.X1.vin2 a_31862_28976# X2.X1.X1.X1.X1.X2.X3.vin1 vdd.t473 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1140 X2.X1.X2.X2.X1.X1.X3.vin2 a_38152_20264# X2.X1.X2.X2.X1.X1.vout vss.t1196 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1141 a_31476_27070# d0.t127 vss.t1086 vss.t1085 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1142 X1.X1.X1.X1.X2.X1.X3.vin2 a_4782_24258# X1.X1.X1.X1.X2.X1.vout vdd.t702 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1143 X1.X2.X2.X2.X1.X1.X3.vin1 a_23512_20264# X1.X2.X2.X2.X1.X1.vout vdd.t642 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1144 vdd.t655 a_52492_18358# a_52106_18358# vdd.t654 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1145 vdd.t505 a_40352_32700# a_39966_32700# vdd.t504 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1146 a_2196_9916# d0.t128 vdd.t1323 vdd.t1322 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1147 a_34062_12822# a_33676_12822# vdd.t1405 vdd.t1404 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1148 vss.t406 a_40352_30794# a_39966_30794# vss.t405 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1149 X1.X1.X1.X1.X3.vin2 a_5082_26164# X1.X1.X1.X3.vin1 vdd.t694 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1150 a_33676_5198# d1.t64 vss.t50 vss.t49 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1151 X1.X1.X2.X1.X2.X1.X1.vin1 a_11072_11734# X1.X1.X2.X1.X2.X1.X3.vin1 vdd.t1415 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1152 X2.X2.X2.X2.X2.X2.X2.vin1 vrefl.t0 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1153 X2.X2.X1.X1.X2.X2.X3.vin2 a_48702_20446# X2.X2.X1.X1.X2.X2.vout vdd.t1221 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1154 X1.X1.X2.X2.X2.X1.vout a_8572_29834# X1.X1.X2.X2.X3.vin2 vdd.t106 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1155 X2.X2.X1.X2.X2.X1.vout a_48316_9010# X2.X2.X1.X2.X2.X1.X3.vin1 vdd.t265 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1156 X1.X2.X1.X2.X1.X1.X3.vin2 a_16836_15634# X1.X2.X1.X2.X1.X2.vrefh vss.t1295 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1157 X1.X1.X2.X2.X2.X2.X3.vin1 a_8872_31700# X1.X1.X2.X2.X2.X2.vout vdd.t754 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1158 a_46502_8010# a_46116_8010# vss.t1167 vss.t1166 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1159 X2.X1.X2.X2.X2.X2.X3.vin1 a_39966_30794# X2.X1.X2.X2.X2.X2.X1.vin2 vdd.t440 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1160 X1.X2.X2.X2.X2.X1.X3.vin1 a_25326_26982# X1.X2.X2.X2.X2.X1.X1.vin1 vss.t1009 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1161 vss.t52 d1.t65 a_38152_24076# vss.t51 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1162 vdd.t1325 d0.t129 a_54992_13640# vdd.t1324 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1163 vdd.t1327 d0.t130 a_25712_7922# vdd.t1326 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1164 vdd.t451 a_23212_29834# a_22826_29834# vdd.t450 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1165 a_5646_892# d5.t4 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1166 a_46116_11822# d0.t131 vdd.t1329 vdd.t1328 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1167 vdd.t1331 d0.t132 a_25712_17452# vdd.t1330 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1168 X1.X2.X1.X1.X1.X2.X3.vin1 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin1 vdd.t302 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1169 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1170 X1.X2.X2.X2.X1.X2.X1.vin1 a_25712_23170# X1.X2.X2.X2.X1.X2.X3.vin1 vdd.t882 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1171 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1172 a_2196_15634# d0.t133 vss.t1351 vss.t1350 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1173 vdd.t1421 a_23512_31700# a_23126_31700# vdd.t1420 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1174 X1.X1.X1.X1.X1.X2.X3.vin1 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin2 vss.t345 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1175 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1176 X1.X2.X1.X2.X2.X2.vout a_19036_5198# X1.X2.X1.X2.X2.X2.X3.vin1 vdd.t661 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1177 X1.X1.X2.X1.X1.X1.X3.vin2 a_8872_5016# X1.X1.X2.X1.X1.X1.vout vss.t296 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1178 a_19036_12822# d1.t66 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1179 X2.X1.X2.X1.X1.X1.vout a_37766_5016# X2.X1.X2.X1.X1.X1.X3.vin2 vdd.t1148 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1180 X1.X2.X2.X1.X1.X1.X1.vin1 X1.X2.X2.vrefh.t0 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1181 a_46116_8010# d0.t134 vdd.t1333 vdd.t1332 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1182 X2.X2.X2.X1.X1.X1.X3.vin2 a_52792_5016# X2.X2.X2.X1.X1.X1.vout vss.t1252 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1183 X2.X1.X2.X1.X1.X2.X3.vin2 a_38152_8828# X2.X1.X2.X1.X1.X2.vout vss.t697 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1184 vss.t421 a_54992_7922# a_54606_7922# vss.t420 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1185 a_2196_28976# d0.t135 vdd.t1335 vdd.t1334 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1186 a_2196_9916# d0.t136 vss.t1353 vss.t1352 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1187 X1.X3.vin1 a_5646_892# X1.X1.X3.vin2.t2 vss.t920 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1188 vout.t1 a_28096_892# X3.vin1.t1 vdd.t549 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1189 X1.X1.X1.X2.X2.X2.X3.vin1 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin1 vdd.t1511 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1190 X1.X1.X1.X2.X2.X2.X2.vin1 a_2582_4198# X1.X1.X1.X2.X2.X2.X3.vin2 vss.t718 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1191 vss.t320 a_54992_15546# a_54606_15546# vss.t319 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1192 a_46116_17540# d0.t137 vss.t1355 vss.t1354 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1193 vss.t894 a_52792_31700# a_52406_31700# vss.t893 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1194 X1.X2.X2.X2.X2.X1.vout a_23212_29834# X1.X2.X2.X2.X3.vin2 vdd.t449 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1195 vdd.t1425 a_40352_15546# a_39966_15546# vdd.t1424 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1196 vdd.t162 a_11072_19358# a_10686_19358# vdd.t161 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1197 X2.X2.X2.X2.X1.X1.X3.vin2 a_52792_20264# X2.X2.X2.X2.X1.X1.vout vss.t1247 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1198 X2.X2.X1.X3.vin1 a_48616_26164# X2.X2.X1.X1.X3.vin1 vdd.t404 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1199 X2.X2.X2.X2.X1.X1.X3.vin2 a_54606_21264# X2.X2.X2.X2.X1.X1.X2.vin1 vss.t120 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1200 X1.X2.X1.X1.X2.X1.X3.vin1 a_19422_24258# X1.X2.X1.X1.X2.X1.vout vss.t82 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1201 X1.X1.X1.X1.X2.X1.vout a_5082_22312# X1.X1.X1.X1.X3.vin2 vss.t516 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1202 X1.X2.X2.X3.vin1 a_22826_10734# X1.X2.X2.X1.X3.vin1 vss.t910 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1203 X1.X2.X2.X2.X2.X2.X3.vin1 a_23512_31700# X1.X2.X2.X2.X2.X2.vout vdd.t1419 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1204 X2.X1.X1.X1.X1.X2.vout a_33676_28070# X2.X1.X1.X1.X1.X2.X3.vin2 vss.t1242 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1205 X1.X1.X2.X2.X1.X2.vout a_8486_24076# X1.X1.X2.X2.X1.X2.X3.vin1 vss.t669 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1206 a_28096_892# d7.t0 vss.t1215 vss.t1214 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1207 X2.X1.X1.X1.X1.X1.X3.vin2 a_31476_30882# X2.X1.X1.X1.X1.X1.X2.vin1 vdd.t396 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1208 vss.t137 a_11072_4110# a_10686_4110# vss.t136 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1209 X1.X2.X1.X2.X2.X1.X1.vin1 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin1 vss.t241 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1210 vss.t290 a_8872_16452# a_8486_16452# vss.t289 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1211 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1212 a_31476_15634# d0.t138 vdd.t1337 vdd.t1336 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1213 a_34362_18540# a_33976_18540# vdd.t779 vdd.t778 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1214 X2.X2.X2.X2.X1.X2.X1.vin2 a_54992_23170# X2.X2.X2.X2.X1.X2.X3.vin1 vss.t1390 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1215 vss.t1357 d0.t139 a_25712_26982# vss.t1356 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1216 X2.X1.X1.X1.X2.X2.vout a_33676_20446# X2.X1.X1.X1.X2.X2.X3.vin2 vss.t1220 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1217 X2.X1.X2.X2.X1.X1.vout a_37766_20264# X2.X1.X2.X2.X1.X1.X3.vin1 vss.t1428 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1218 vss.t457 a_37852_6962# a_37466_6962# vss.t456 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1219 X1.X1.X1.X2.X3.vin2 a_4696_7064# X1.X1.X1.X2.X2.X2.vout vss.t1272 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1220 X2.X2.X1.X2.X2.vrefh a_46502_11822# X2.X2.X1.X2.X1.X2.X3.vin2 vdd.t798 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1221 a_31476_6104# d0.t140 vss.t1359 vss.t1358 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1222 X2.X1.X1.X2.X2.X1.X3.vin1 a_34062_9010# X2.X1.X1.X2.X2.X1.vout vss.t31 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1223 X2.vrefh a_25712_32700# X1.X2.X2.X2.X2.X2.X3.vin2 vss.t1089 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1224 X1.X1.X2.X1.X2.X1.X3.vin1 a_10686_11734# X1.X1.X2.X1.X2.X1.X1.vin2 vdd.t959 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1225 a_19722_14688# a_19336_14688# vss.t810 vss.t809 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1226 X2.X2.X1.X2.X2.X1.X2.vin1 a_46502_8010# X2.X2.X1.X2.X2.X1.X3.vin2 vss.t1150 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1227 X2.X2.X1.X1.X2.X2.vout a_48316_20446# X2.X2.X1.X1.X2.X2.X3.vin1 vdd.t1386 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1228 X1.X1.X1.X2.X1.X1.vout a_4396_16634# X1.X1.X1.X2.X1.X1.X3.vin2 vss.t1288 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1229 a_17222_21352# a_16836_21352# vdd.t982 vdd.t981 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1230 X2.X2.X2.X1.X1.X2.X3.vin2 a_54606_9828# X2.X2.X2.X1.X2.vrefh vdd.t1018 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1231 vss.t1361 d0.t141 a_11072_17452# vss.t1360 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1232 a_2582_21352# a_2196_21352# vss.t267 vss.t266 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1233 vdd.t389 a_52792_16452# a_52406_16452# vdd.t388 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1234 vdd.t1249 a_8872_24076# a_8486_24076# vdd.t1248 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1235 a_34362_10916# a_33976_10916# vdd.t723 vdd.t722 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1236 X2.X1.X1.X2.X2.X1.vout a_33676_9010# X2.X1.X1.X2.X2.X1.X3.vin1 vdd.t17 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1237 X1.X1.X2.X1.X1.X2.X3.vin1 a_10686_7922# X1.X1.X2.X1.X1.X2.X1.vin1 vss.t344 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1238 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1239 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1240 X2.X2.X1.X1.X3.vin2 a_48616_22312# X2.X2.X1.X1.X2.X2.vout vss.t145 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1241 X1.X2.X2.X2.X1.X2.vout a_23126_24076# X1.X2.X2.X2.X1.X2.X3.vin1 vss.t1458 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1242 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1243 a_46116_28976# d0.t142 vss.t1363 vss.t1362 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1244 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1245 X2.X1.X2.X2.X1.X2.X3.vin1 a_39966_23170# X2.X1.X2.X2.X1.X2.X1.vin1 vss.t124 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1246 a_19336_18540# d4.t7 vdd.t1130 vdd.t1129 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1247 X2.X2.X1.X2.X1.X1.X1.vin1 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin1 vss.t1399 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1248 vss.t324 a_11072_28888# a_10686_28888# vss.t323 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1249 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1250 a_48316_5198# d1.t67 vss.t54 vss.t53 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1251 a_4696_18540# d4.t8 vss.t1392 vss.t1391 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1252 X2.X1.X1.X2.X1.X2.X3.vin1 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin1 vdd.t192 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1253 vss.t1365 d0.t143 a_54992_21264# vss.t1364 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1254 X2.X1.X2.X1.X1.X2.X3.vin1 a_39966_7922# X2.X1.X2.X1.X1.X2.X1.vin1 vss.t975 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1255 a_17222_27070# a_16836_27070# vss.t196 vss.t195 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1256 vss.t106 d3.t14 a_23212_10734# vss.t105 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1257 a_48702_20446# a_48316_20446# vdd.t1385 vdd.t1384 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1258 vdd.t1372 d4.t9 a_37852_18358# vdd.t1371 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1259 vdd.t1339 d0.t144 a_11072_25076# vdd.t1338 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1260 X1.X1.X2.X2.X2.X2.vout a_8572_29834# X1.X1.X2.X2.X3.vin2 vss.t116 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1261 a_4782_24258# a_4396_24258# vss.t717 vss.t716 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1262 X2.X1.X2.vrefh.t2 X2.X1.X1.X2.X2.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1263 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1264 a_31476_13728# d0.t145 vss.t1367 vss.t1366 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1265 vdd.t553 d0.t146 a_54992_4110# vdd.t552 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1266 X1.X2.X2.X1.X1.X1.vout a_23126_5016# X1.X2.X2.X1.X1.X1.X3.vin2 vdd.t1263 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1267 X1.X1.X2.X1.X1.X1.X1.vin1 X1.X1.X2.vrefh.t2 vss.t242 sky130_fd_pr__res_high_po_0p35 l=1.09
X1268 a_31862_4198# a_31476_4198# vss.t131 vss.t130 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1269 a_19336_10916# d3.t15 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1270 a_4696_10916# d3.t16 vss.t108 vss.t107 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1271 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1272 X1.X2.X2.X2.X3.vin2 a_22826_29834# X1.X2.X2.X2.X2.X2.vout vdd.t343 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1273 X1.X2.X2.X1.X2.X2.X2.vin1 a_25712_17452# X1.X2.X2.X1.X2.X2.X3.vin2 vdd.t961 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1274 vss.t461 a_23212_29834# a_22826_29834# vss.t460 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1275 vdd.t555 d0.t147 a_40352_26982# vdd.t554 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1276 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1277 vss.t567 d0.t148 a_40352_25076# vss.t566 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1278 vss.t259 a_23512_8828# a_23126_8828# vss.t258 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1279 X1.X1.X2.X2.X1.X1.vout a_8572_22210# X1.X1.X2.X2.X3.vin1 vdd.t1441 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1280 X2.X1.X1.X2.X1.X1.vout a_33676_16634# X2.X1.X1.X2.X1.X1.X3.vin1 vdd.t631 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1281 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X1.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1282 a_31862_21352# a_31476_21352# vdd.t1134 vdd.t1133 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1283 a_4696_22312# d2.t30 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1284 a_2582_32788# a_2196_32788# vss.t1110 vss.t1109 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1285 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1286 vdd.t131 a_23212_22210# a_22826_22210# vdd.t130 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1287 X2.X1.X2.X1.X3.vin1 a_37852_10734# X2.X1.X2.X3.vin1 vdd.t1241 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1288 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1289 a_33676_31882# d1.t68 vss.t56 vss.t55 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1290 a_2582_17540# a_2196_17540# vdd.t1181 vdd.t1180 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1291 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1292 X2.X1.X1.X2.X1.X2.X3.vin2 a_31476_11822# X2.X1.X1.X2.X2.vrefh vss.t968 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1293 X2.X2.X2.X1.X2.X2.X3.vin1 a_54606_15546# X2.X2.X2.X1.X2.X2.X1.vin1 vss.t81 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1294 X2.X2.X2.X2.X2.X2.vout a_52406_31700# X2.X2.X2.X2.X2.X2.X3.vin1 vss.t628 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1295 a_48316_24258# d1.t69 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1296 a_31476_32788# d0.t149 vdd.t557 vdd.t556 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1297 X1.X2.X2.X2.X2.X2.vout a_23212_29834# X1.X2.X2.X2.X3.vin2 vss.t459 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1298 a_33976_18540# d4.t10 vdd.t1374 vdd.t1373 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1299 a_48616_26164# d3.t17 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1300 X1.X1.X3.vin2 a_8186_18358# X1.X1.X2.X3.vin2 vdd.t1037 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1301 a_33976_7064# d2.t31 vss.t70 vss.t69 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1302 vss.t172 a_11072_19358# a_10686_19358# vss.t171 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1303 X2.X2.X1.X1.X1.X2.X1.vin1 a_46502_28976# X2.X2.X1.X1.X1.X2.X3.vin1 vss.t1287 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1304 vss.t58 d1.t70 a_23512_24076# vss.t57 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1305 X2.X2.X1.X2.X1.X2.X3.vin2 a_46116_11822# X2.X2.X1.X2.X1.X2.X2.vin1 vdd.t1277 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1306 X1.X1.X2.X1.X2.X1.vout a_8572_14586# X1.X1.X2.X1.X3.vin2 vdd.t891 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1307 vdd.t84 a_54992_9828# a_54606_9828# vdd.t83 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1308 X2.X1.X1.X1.X2.X1.X3.vin1 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin1 vdd.t1207 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1309 a_31862_27070# a_31476_27070# vss.t605 vss.t604 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1310 a_2582_9916# a_2196_9916# vdd.t1389 vdd.t1388 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1311 a_16836_21352# d0.t150 vdd.t559 vdd.t558 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1312 X1.X1.X2.X2.X1.X2.X1.vin1 a_11072_23170# X1.X1.X2.X2.X1.X2.X3.vin1 vdd.t738 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1313 a_19036_9010# d1.t71 vdd.t989 vdd.t988 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1314 a_33976_10916# d3.t18 vdd.t94 vdd.t93 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1315 vdd.t240 a_23212_14586# a_22826_14586# vdd.t239 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1316 X1.X2.X2.X2.X1.X1.vout a_23212_22210# X1.X2.X2.X2.X3.vin1 vdd.t129 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1317 vss.t569 d0.t151 a_40352_9828# vss.t568 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1318 X2.X2.X2.X2.vrefh a_54992_17452# X2.X2.X2.X1.X2.X2.X3.vin2 vss.t170 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1319 X1.X1.X1.X1.X1.X1.X2.vin1 a_2582_30882# X1.X1.X1.X1.X1.X1.X3.vin2 vss.t1192 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1320 X1.X2.X2.X2.X2.X2.X1.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1321 X1.X2.X2.X2.X2.X1.X1.vin2 a_25712_26982# X1.X2.X2.X2.X2.X1.X3.vin1 vss.t188 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1322 a_46116_6104# d0.t152 vss.t571 vss.t570 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1323 X2.X2.X1.X2.X1.X1.X3.vin1 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin2 vss.t439 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1324 vdd.t57 d2.t32 a_23212_29834# vdd.t56 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1325 vdd.t734 a_11072_6016# a_10686_6016# vdd.t733 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1326 a_46502_11822# a_46116_11822# vdd.t1276 vdd.t1275 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1327 vdd.t69 a_25712_13640# a_25326_13640# vdd.t68 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1328 a_17222_15634# a_16836_15634# vdd.t1269 vdd.t1268 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1329 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1330 a_2582_15634# a_2196_15634# vss.t1103 vss.t1102 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1331 a_16836_27070# d0.t153 vss.t573 vss.t572 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1332 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1333 a_4396_9010# d1.t72 vss.t1019 vss.t1018 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1334 X2.X2.X2.X1.X2.X2.vout a_52406_16452# X2.X2.X2.X1.X2.X2.X3.vin2 vdd.t391 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1335 X2.X2.X2.X2.X1.X2.X2.vin1 a_54992_25076# X2.X2.X2.X2.X1.X2.X3.vin2 vdd.t1118 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1336 X1.X2.X2.X1.X2.X1.vout a_23212_14586# X1.X2.X2.X1.X3.vin2 vdd.t238 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1337 X1.X2.X2.X1.X1.X2.X3.vin1 a_25326_7922# X1.X2.X2.X1.X1.X2.X1.vin1 vss.t153 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1338 vss.t575 d0.t154 a_54992_6016# vss.t574 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1339 a_2582_28976# a_2196_28976# vdd.t339 vdd.t338 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1340 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1341 X2.X1.X2.X1.X2.X2.X3.vin2 a_39966_17452# X2.X1.X2.X1.X2.X2.X2.vin1 vss.t316 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1342 X1.X2.X1.X3.vin1 a_19722_18540# X1.X2.X3.vin1 vss.t272 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1343 a_48616_22312# d2.t33 vss.t72 vss.t71 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1344 a_33676_28070# d1.t73 vdd.t991 vdd.t990 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1345 X1.X2.X2.vrefh.t2 X1.X2.X1.X2.X2.X2.X2.vin1 vss.t257 sky130_fd_pr__res_high_po_0p35 l=1.09
X1346 vdd.t561 d0.t155 a_40352_4110# vdd.t560 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1347 vss.t577 d0.t156 a_54992_15546# vss.t576 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1348 vdd.t622 a_40352_26982# a_39966_26982# vdd.t621 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1349 a_46502_17540# a_46116_17540# vss.t438 vss.t437 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1350 X2.X2.X1.X1.X2.X1.X3.vin2 a_48702_24258# X2.X2.X1.X1.X2.X1.vout vdd.t445 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1351 vss.t1021 d1.t74 a_52792_31700# vss.t1020 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1352 vss.t728 a_40352_25076# a_39966_25076# vss.t727 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1353 X2.X2.X1.X1.X3.vin2 a_49002_26164# X2.X2.X1.X3.vin1 vdd.t1230 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1354 vdd.t563 d0.t157 a_11072_19358# vdd.t562 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1355 X2.X1.X1.X2.X2.X2.vrefh a_31862_8010# X2.X1.X1.X2.X2.X1.X3.vin2 vdd.t615 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1356 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1357 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1358 X1.X1.X2.X1.X1.X2.X3.vin2 a_10686_9828# X1.X1.X2.X1.X2.vrefh vdd.t216 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1359 X2.X2.X2.X2.X1.X2.vout a_52492_22210# X2.X2.X2.X2.X3.vin1 vss.t871 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1360 vdd.t1039 a_54992_28888# a_54606_28888# vdd.t1038 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1361 a_46502_4198# a_46116_4198# vss.t856 vss.t855 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1362 X1.X2.X1.X2.X3.vin1 a_19722_10916# X1.X2.X1.X3.vin2 vss.t1382 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1363 X1.X2.vrefh a_11072_32700# X1.X1.X2.X2.X2.X2.X3.vin2 vss.t350 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1364 X2.X1.X1.X1.X1.X2.X3.vin1 a_34062_28070# X2.X1.X1.X1.X1.X2.vout vss.t934 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1365 X1.X1.X2.X2.X1.X2.X3.vin2 a_8872_24076# X1.X1.X2.X2.X1.X2.vout vss.t1278 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1366 X1.X2.X1.X1.X2.X2.X1.vin2 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin1 vdd.t983 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1367 X2.X1.X1.X1.X1.X2.vrefh a_31862_30882# X2.X1.X1.X1.X1.X1.X3.vin2 vdd.t144 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1368 X2.X1.X2.X2.X1.X2.X3.vin2 a_39966_25076# X2.X1.X2.X2.X2.vrefh vdd.t537 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1369 vdd.t59 d2.t34 a_8572_6962# vdd.t58 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1370 a_17222_13728# a_16836_13728# vss.t164 vss.t163 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1371 vdd.t834 d2.t35 a_52492_6962# vdd.t833 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1372 X2.X1.X2.X1.X1.X2.X3.vin2 a_39966_9828# X2.X1.X2.X1.X2.vrefh vdd.t1032 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1373 vss.t696 a_38152_8828# a_37766_8828# vss.t695 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1374 X1.X2.X2.X2.X3.vin2 a_22826_29834# X1.X2.X2.X2.X2.X1.vout vss.t351 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1375 vss.t1023 d1.t75 a_8872_16452# vss.t1022 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1376 X1.X1.X1.X1.X2.vrefh a_2582_27070# X1.X1.X1.X1.X1.X2.X3.vin2 vdd.t418 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1377 X1.X3.vin2 a_20286_892# X1.X2.X3.vin2.t2 vss.t735 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1378 vss.t256 a_23512_24076# a_23126_24076# vss.t255 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1379 a_31862_15634# a_31476_15634# vdd.t1159 vdd.t1158 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1380 vss.t514 a_38152_31700# a_37766_31700# vss.t513 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1381 X2.X2.X1.X1.X1.X1.X1.vin2 X2.X2.X1.X1.X1.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1382 X2.X2.X1.X1.X1.X2.X3.vin1 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin2 vss.t981 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1383 X1.X2.X1.X1.X2.X2.vout a_19722_22312# X1.X2.X1.X1.X3.vin2 vdd.t1195 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1384 X2.X1.X1.X1.X1.X2.vout a_34362_29936# X2.X1.X1.X1.X3.vin1 vdd.t1237 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1385 X2.X1.X1.X1.X2.X2.X3.vin1 a_34062_20446# X2.X1.X1.X1.X2.X2.vout vss.t1286 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1386 X1.X3.vin1 a_14082_892# X3.vin1 vss.t244 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1387 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1388 X1.X1.X2.X2.X1.X2.X3.vin1 a_10686_23170# X1.X1.X2.X2.X1.X2.X1.vin2 vdd.t527 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1389 a_17222_8010# a_16836_8010# vss.t560 vss.t559 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1390 vss.t366 a_8872_27888# a_8486_27888# vss.t365 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1391 X1.X2.X1.X1.X1.X2.X2.vin1 a_17222_27070# X1.X2.X1.X1.X1.X2.X3.vin2 vss.t1517 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1392 X2.X1.X2.X2.X3.vin1 a_37466_22210# X2.X1.X2.X2.X1.X1.vout vss.t629 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1393 X1.X1.X1.X2.X1.X1.X3.vin1 a_4782_16634# X1.X1.X1.X2.X1.X1.vout vss.t1386 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1394 X1.X2.X1.X1.X1.X2.vout a_19036_28070# X1.X2.X1.X1.X1.X2.X3.vin2 vss.t943 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1395 X1.X2.X2.X2.X3.vin1 a_22826_22210# X1.X2.X2.X2.X1.X2.vout vdd.t335 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1396 X1.X2.X1.X1.X1.X1.X3.vin2 a_16836_30882# X1.X2.X1.X1.X1.X1.X2.vin1 vdd.t254 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1397 vss.t489 a_40352_9828# a_39966_9828# vss.t488 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1398 vdd.t993 d1.t76 a_52792_16452# vdd.t992 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1399 a_20286_892# d5.t5 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1400 vdd.t995 d1.t77 a_8872_24076# vdd.t994 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1401 vss.t1175 a_11072_13640# a_10686_13640# vss.t1174 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1402 X1.X1.X1.X1.X1.X1.X3.vin2 a_2196_30882# X1.X1.X1.X1.X1.X2.vrefh vss.t1111 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1403 a_48616_7064# d2.t36 vss.t858 vss.t857 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1404 a_34362_7064# a_33976_7064# vdd.t751 vdd.t750 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1405 a_19422_31882# a_19036_31882# vss.t1107 vss.t1106 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1406 a_31476_4198# d0.t158 vdd.t565 vdd.t564 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1407 X2.X2.X2.X1.X1.X2.X1.vin1 a_54992_7922# X2.X2.X2.X1.X1.X2.X3.vin1 vdd.t408 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1408 X2.X2.X1.X1.X2.X1.vout a_49002_22312# X2.X2.X1.X1.X3.vin2 vss.t1132 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1409 a_46502_28976# a_46116_28976# vss.t980 vss.t979 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1410 X1.X2.X2.X2.X1.X2.X3.vin2 a_23512_24076# X1.X2.X2.X2.X1.X2.vout vss.t254 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1411 X2.X1.X2.X1.X2.X1.X2.vin1 a_40352_13640# X2.X1.X2.X1.X2.X1.X3.vin2 vdd.t1229 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1412 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1413 a_4396_28070# d1.t78 vss.t1025 vss.t1024 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1414 a_28482_892# a_28096_892# vss.t565 vss.t564 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1415 a_17222_32788# a_16836_32788# vdd.t1453 vdd.t1452 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1416 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1417 a_16836_15634# d0.t159 vdd.t567 vdd.t566 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1418 X1.X1.X2.X1.X2.X2.X2.vin1 a_11072_17452# X1.X1.X2.X1.X2.X2.X3.vin2 vdd.t1523 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1419 vss.t942 a_25712_7922# a_25326_7922# vss.t941 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1420 a_19722_18540# a_19336_18540# vdd.t1200 vdd.t1199 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1421 a_49566_892# d5.t6 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1422 a_2196_30882# d0.t160 vdd.t569 vdd.t568 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1423 vss.t579 d0.t161 a_11072_28888# vss.t578 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1424 X1.X2.X1.X1.X2.X2.vout a_19036_20446# X1.X2.X1.X1.X2.X2.X3.vin2 vss.t666 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1425 a_5082_18540# a_4696_18540# vss.t1434 vss.t1433 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1426 vdd.t997 d1.t79 a_8872_8828# vdd.t996 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1427 X2.X1.X1.X2.X1.X2.X1.vin2 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin1 vdd.t503 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1428 X2.X2.X2.X2.X3.vin2 a_52492_25982# X2.X2.X2.X3.vin2 vss.t702 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1429 X2.X1.X2.X2.X2.X1.X3.vin1 a_38152_27888# X2.X1.X2.X2.X2.X1.vout vdd.t1111 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1430 vdd.t999 d1.t80 a_52792_8828# vdd.t998 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1431 X1.X1.X1.X2.X3.vin1 a_4696_14688# X1.X1.X1.X2.X1.X1.vout vdd.t261 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1432 vss.t334 a_25712_21264# a_25326_21264# vss.t333 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1433 X1.X2.X2.X1.X3.vin2 a_22826_14586# X1.X2.X2.X1.X2.X2.vout vdd.t241 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1434 X1.X2.X1.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1435 vdd.t1391 a_11072_21264# a_10686_21264# vdd.t1390 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1436 X1.X2.X2.X1.X1.X1.X1.vin1 a_25712_4110# X1.X2.X2.X1.X1.X1.X3.vin1 vdd.t703 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1437 a_31862_13728# a_31476_13728# vss.t200 vss.t199 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1438 vdd.t511 a_38152_16452# a_37766_16452# vdd.t510 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1439 a_4396_20446# d1.t81 vss.t1027 vss.t1026 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1440 a_19722_10916# a_19336_10916# vdd.t692 vdd.t691 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1441 X2.X1.X1.X2.X2.X2.X3.vin1 a_34062_5198# X2.X1.X1.X2.X2.X2.vout vss.t1387 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1442 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1443 a_5082_10916# a_4696_10916# vss.t1385 vss.t1384 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1444 X2.X2.X1.X1.X2.X1.vout a_48316_24258# X2.X2.X1.X1.X2.X1.X3.vin1 vdd.t75 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1445 vss.t581 d0.t162 a_40352_6016# vss.t580 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1446 X2.X2.X1.X2.X2.X2.X2.vin1 a_46502_4198# X2.X2.X1.X2.X2.X2.X3.vin2 vss.t1149 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1447 vss.t860 d2.t37 a_23212_29834# vss.t859 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1448 X2.X2.X1.X2.X2.X2.X3.vin1 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin1 vdd.t46 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1449 X1.X2.X2.X1.X2.X1.X3.vin2 a_25326_13640# X1.X2.X2.X1.X2.X2.vrefh vdd.t306 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1450 X2.X2.X2.X1.X3.vin2 a_52106_14586# X2.X2.X2.X1.X2.X1.vout vss.t142 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1451 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1452 vdd.t571 d0.t163 a_40352_11734# vdd.t570 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1453 X2.X1.X1.X2.X1.X1.X3.vin2 a_34062_16634# X2.X1.X1.X2.X1.X1.vout vdd.t305 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1454 X2.X2.X2.X2.X1.X1.X1.vin1 a_54992_19358# X2.X2.X2.X2.X1.X1.X3.vin1 vdd.t1105 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1455 X1.X2.X1.X2.X1.X2.X3.vin1 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin1 vdd.t152 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1456 X1.X1.X2.X2.X2.X2.X3.vin2 a_10686_32700# X1.X1.X2.X2.X2.X2.X2.vin1 vss.t1097 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1457 X2.X1.X2.X3.vin2 a_37466_25982# X2.X1.X2.X2.X3.vin1 vss.t1093 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1458 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1459 X2.X1.X2.X1.X1.X1.vout a_37852_6962# X2.X1.X2.X1.X3.vin1 vdd.t446 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1460 X1.X1.X3.vin2.t1 a_6032_892# X1.X3.vin1 vdd.t706 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1461 a_5082_22312# a_4696_22312# vdd.t301 vdd.t300 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1462 X2.X2.X3.vin2.t2 a_49952_892# X2.X3.vin2 vdd.t748 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1463 a_16836_13728# d0.t164 vss.t497 vss.t496 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1464 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1465 a_2582_8010# a_2196_8010# vss.t1190 vss.t1189 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1466 vdd.t836 d2.t38 a_23212_22210# vdd.t835 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1467 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1468 a_34062_31882# a_33676_31882# vss.t743 vss.t742 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1469 X2.X1.X1.X1.X2.X1.X3.vin2 a_31476_23258# X2.X1.X1.X1.X2.X2.vrefh vss.t704 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1470 X2.X1.X1.X1.X3.vin1 a_34362_26164# X2.X1.X1.X3.vin1 vss.t1438 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1471 vdd.t1001 d1.t82 a_38152_5016# vdd.t1000 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1472 X2.X1.X1.X2.X1.X2.X2.vin1 a_31862_11822# X2.X1.X1.X2.X1.X2.X3.vin2 vss.t1056 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1473 a_2196_13728# d0.t165 vdd.t479 vdd.t478 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1474 X1.X2.X1.X2.X3.vin1 a_19336_14688# X1.X2.X1.X2.X1.X1.vout vdd.t785 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1475 X1.X1.X1.X1.X1.X2.X3.vin2 a_2196_27070# X1.X1.X1.X1.X1.X2.X2.vin1 vdd.t1020 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1476 a_48702_24258# a_48316_24258# vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1477 a_31862_32788# a_31476_32788# vdd.t761 vdd.t760 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1478 a_19422_28070# a_19036_28070# vdd.t935 vdd.t934 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1479 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1480 a_49002_26164# a_48616_26164# vdd.t403 vdd.t402 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1481 X1.X1.X2.X3.vin1 a_8572_18358# X1.X1.X3.vin2 vdd.t407 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1482 X2.X1.X1.X1.X3.vin1 a_33976_29936# X2.X1.X1.X1.X1.X1.vout vdd.t185 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1483 X1.X2.X2.X1.X1.X2.X3.vin2 a_25326_9828# X1.X2.X2.X1.X2.vrefh vdd.t1078 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1484 vss.t499 d0.t166 a_11072_19358# vss.t498 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1485 X1.X1.X1.X2.X2.X1.X1.vin1 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin1 vss.t88 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1486 X1.X1.X2.X2.X2.X1.X1.vin2 a_11072_26982# X1.X1.X2.X2.X2.X1.X3.vin1 vss.t925 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1487 X1.X2.X1.X2.X1.X2.vrefh a_17222_15634# X1.X2.X1.X2.X1.X1.X3.vin2 vdd.t1270 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1488 X2.X2.X2.X2.X2.X1.X3.vin1 a_52792_27888# X2.X2.X2.X2.X2.X1.vout vdd.t298 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1489 X2.X1.X1.X1.X2.X1.X1.vin2 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin1 vdd.t802 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1490 a_2196_8010# d0.t167 vdd.t481 vdd.t480 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1491 X1.X2.X1.X2.X1.X1.vout a_19036_16634# X1.X2.X1.X2.X1.X1.X3.vin1 vdd.t77 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1492 X2.X1.X2.X2.X1.X1.X3.vin1 a_39966_19358# X2.X1.X2.X2.X1.X1.X1.vin2 vdd.t810 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1493 X2.X2.X2.X2.X2.X1.X3.vin2 a_54606_28888# X2.X2.X2.X2.X2.X2.vrefh vdd.t103 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1494 X2.X2.X1.X2.X3.vin2 a_48616_7064# X2.X2.X1.X2.X2.X2.vout vss.t1520 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1495 X1.X1.X1.X1.X1.X1.vout a_4396_31882# X1.X1.X1.X1.X1.X1.X3.vin1 vdd.t242 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1496 a_46116_30882# d0.t168 vss.t501 vss.t500 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1497 a_33676_20446# d1.t83 vdd.t1003 vdd.t1002 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1498 vdd.t542 a_23212_18358# a_22826_18358# vdd.t541 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1499 vdd.t341 a_11072_32700# a_10686_32700# vdd.t340 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1500 vss.t522 a_11072_30794# a_10686_30794# vss.t521 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1501 vdd.t838 d2.t39 a_23212_14586# vdd.t837 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1502 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1503 X2.X2.X1.X2.X2.X2.vout a_48316_5198# X2.X2.X1.X2.X2.X2.X3.vin1 vdd.t648 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1504 a_19036_31882# d1.t84 vss.t1029 vss.t1028 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1505 a_4396_16634# d1.t85 vdd.t1005 vdd.t1004 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1506 X1.X2.X1.X2.X1.X2.X3.vin2 a_16836_11822# X1.X2.X1.X2.X2.vrefh vss.t411 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1507 a_16836_32788# d0.t169 vdd.t483 vdd.t482 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1508 X1.X1.X2.X1.X2.X2.X3.vin2 a_10686_17452# X1.X1.X2.X2.vrefh vdd.t1242 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1509 vdd.t485 d0.t170 a_25712_4110# vdd.t484 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1510 X2.X1.X2.X1.X1.X2.X1.vin1 a_40352_7922# X2.X1.X2.X1.X1.X2.X3.vin1 vdd.t1233 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1511 vdd.t487 d0.t171 a_25712_13640# vdd.t486 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1512 X2.X2.X2.X2.X2.X2.vrefh a_54992_28888# X2.X2.X2.X2.X2.X1.X3.vin2 vss.t1070 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1513 X2.X1.X2.X2.X2.X1.vout a_37766_27888# X2.X1.X2.X2.X2.X1.X3.vin2 vdd.t888 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1514 X2.X1.X2.X2.X1.X2.vrefh a_40352_21264# X2.X1.X2.X2.X1.X1.X3.vin2 vss.t354 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1515 X1.X2.X1.X1.X2.X1.X3.vin1 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin1 vdd.t806 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1516 X2.X2.X2.X3.vin2 a_52106_25982# X2.X2.X2.X2.X3.vin2 vdd.t1163 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1517 vss.t862 d2.t40 a_52492_14586# vss.t861 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1518 X1.X2.X1.X2.X2.X2.vrefh a_17222_8010# X1.X2.X1.X2.X2.X1.X3.vin2 vdd.t428 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1519 a_2196_11822# d0.t172 vss.t503 vss.t502 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1520 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1521 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1522 X1.X2.X2.X3.vin1 a_23212_18358# X1.X2.X3.vin2 vdd.t540 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1523 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X2.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1524 X1.X2.X2.X1.X1.X2.vrefh a_25712_6016# X1.X2.X2.X1.X1.X1.X3.vin2 vss.t229 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1525 a_46116_4198# d0.t173 vdd.t489 vdd.t488 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1526 X1.X1.X1.X2.vrefh a_2582_19446# X1.X1.X1.X1.X2.X2.X3.vin2 vdd.t1257 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1527 X1.X2.X1.X1.X1.X2.X3.vin1 a_19422_28070# X1.X2.X1.X1.X1.X2.vout vss.t686 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1528 vrefh.t0 X1.X1.X1.X1.X1.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1529 X2.X1.X1.X2.X2.X2.X1.vin1 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin1 vss.t451 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1530 X2.X1.X2.X1.X1.X1.X3.vin2 a_38152_5016# X2.X1.X2.X1.X1.X1.vout vss.t726 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1531 X2.X1.X1.X1.X1.X1.vout a_34362_29936# X2.X1.X1.X1.X3.vin1 vss.t1265 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1532 X1.X2.X1.X2.X1.X2.X1.vin1 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin1 vss.t165 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1533 a_2196_25164# d0.t174 vdd.t491 vdd.t490 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1534 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1535 a_49002_22312# a_48616_22312# vss.t144 vss.t143 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1536 a_34062_28070# a_33676_28070# vdd.t1216 vdd.t1215 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1537 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1538 vss.t928 a_54992_11734# a_54606_11734# vss.t927 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1539 vdd.t1436 a_40352_11734# a_39966_11734# vdd.t1435 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1540 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X1.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1541 vss.t1119 a_25712_15546# a_25326_15546# vss.t1118 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1542 vdd.t573 a_11072_15546# a_10686_15546# vdd.t572 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1543 X2.X1.X1.X2.X2.X2.X3.vin1 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin1 vdd.t474 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1544 vss.t505 d0.t175 a_11072_7922# vss.t504 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1545 X1.X2.X1.X1.X2.X2.X3.vin1 a_19422_20446# X1.X2.X1.X1.X2.X2.vout vss.t1088 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1546 X2.X1.X2.X2.X2.X1.X3.vin2 a_39966_28888# X2.X1.X2.X2.X2.X1.X2.vin1 vss.t78 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1547 X1.X2.X2.X2.X1.X1.X3.vin2 a_25326_21264# X1.X2.X2.X2.X1.X1.X2.vin1 vss.t87 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1548 vss.t374 a_37852_14586# a_37466_14586# vss.t373 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1549 vdd.t493 d0.t176 a_54992_28888# vdd.t492 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1550 X1.X1.X1.X1.X2.X1.X1.vin1 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin1 vss.t984 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1551 a_46116_27070# d0.t177 vdd.t495 vdd.t494 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1552 a_43362_892# a_42976_892# vdd.t1174 vdd.t1173 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1553 X2.X2.X1.X1.X1.X1.X2.vin1 a_46502_30882# X2.X2.X1.X1.X1.X1.X3.vin2 vss.t926 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1554 vdd.t1266 a_25712_9828# a_25326_9828# vdd.t1265 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1555 X2.X1.X1.X3.vin1 a_33976_26164# X2.X1.X1.X1.X3.vin2 vss.t1525 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1556 X1.X2.X2.X1.X1.X1.vout a_23212_6962# X1.X2.X2.X1.X3.vin1 vdd.t885 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1557 a_19036_28070# d1.t86 vdd.t857 vdd.t856 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1558 a_4396_5198# d1.t87 vss.t881 vss.t880 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1559 a_31862_9916# a_31476_9916# vss.t709 vss.t708 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1560 vss.t528 a_8872_12640# a_8486_12640# vss.t527 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1561 X1.X1.X2.X2.X2.X1.X3.vin1 a_10686_26982# X1.X1.X2.X2.X2.X1.X1.vin1 vss.t1007 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1562 a_48316_16634# d1.t88 vss.t883 vss.t882 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1563 X1.X2.X1.X1.X1.X1.X1.vin2 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin1 vdd.t634 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1564 vss.t885 d1.t89 a_38152_31700# vss.t884 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1565 a_31476_11822# d0.t178 vdd.t497 vdd.t496 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1566 X2.X2.X2.X2.X1.X1.X1.vin2 a_54992_19358# X2.X2.X2.X2.X1.X1.X3.vin1 vss.t1131 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1567 X2.X2.X2.X1.X1.X1.X3.vin1 a_54606_4110# X2.X2.X2.X1.X1.X1.X1.vin1 vss.t911 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1568 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1569 X2.X2.X2.X3.vin2 a_52492_18358# X2.X2.X3.vin2.t0 vss.t682 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1570 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1571 X2.X2.X2.X1.X3.vin1 a_52106_6962# X2.X2.X2.X1.X1.X1.vout vss.t1147 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1572 vss.t887 d1.t90 a_8872_27888# vss.t886 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1573 vdd.t96 d3.t19 a_52492_25982# vdd.t95 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1574 X2.X1.X2.X2.X1.X2.vout a_37852_22210# X2.X1.X2.X2.X3.vin1 vss.t119 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1575 X1.X1.X1.X2.X1.X2.vout a_4396_12822# X1.X1.X1.X2.X1.X2.X3.vin2 vss.t630 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1576 vdd.t665 a_52792_12640# a_52406_12640# vdd.t664 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1577 vss.t507 d0.t179 a_11072_13640# vss.t506 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1578 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1579 vdd.t271 a_8872_20264# a_8486_20264# vdd.t270 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1580 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1581 X1.X1.X2.X1.X1.X1.vout a_8486_5016# X1.X1.X2.X1.X1.X1.X3.vin2 vdd.t498 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1582 X2.X1.X1.X2.X2.X2.vout a_33676_5198# X2.X1.X1.X2.X2.X2.X3.vin1 vdd.t1169 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1583 a_4782_28070# a_4396_28070# vss.t808 vss.t807 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1584 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1585 a_31476_17540# d0.t180 vss.t509 vss.t508 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1586 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1587 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1588 vss.t511 d0.t181 a_25712_6016# vss.t510 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1589 a_2582_30882# a_2196_30882# vdd.t1086 vdd.t1085 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1590 vss.t377 a_52492_14586# a_52106_14586# vss.t376 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1591 X2.X1.X2.X2.X1.X1.X3.vin1 a_39966_19358# X2.X1.X2.X2.X1.X1.X1.vin1 vss.t840 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1592 X2.X1.X3.vin2.t1 a_37466_18358# X2.X1.X2.X3.vin1 vss.t423 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1593 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1594 X1.X2.X2.X1.X1.X2.X3.vin1 a_23512_8828# X1.X2.X2.X1.X1.X2.vout vdd.t250 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1595 X1.X2.X1.X2.X1.X1.X3.vin2 a_19422_16634# X1.X2.X1.X2.X1.X1.vout vdd.t64 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1596 X1.X2.X3.vin2 a_22826_18358# X1.X2.X2.X3.vin2 vdd.t543 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1597 X1.X2.X3.vin1.t2 a_20672_892# X1.X3.vin2 vss.t1121 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1598 X1.X1.X1.X2.X1.X2.vout a_5082_14688# X1.X1.X1.X2.X3.vin1 vdd.t1102 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1599 X1.X1.X1.X1.X2.X2.X3.vin2 a_2196_19446# X1.X1.X1.X1.X2.X2.X2.vin1 vdd.t803 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1600 vss.t1315 d0.t182 a_25712_21264# vss.t1314 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1601 vdd.t711 a_37852_25982# a_37466_25982# vdd.t710 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1602 a_19422_20446# a_19036_20446# vdd.t639 vdd.t638 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1603 vdd.t1287 d0.t183 a_11072_21264# vdd.t1286 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1604 X1.X2.X1.X2.X2.X1.X3.vin2 a_16836_8010# X1.X2.X1.X2.X2.X2.vrefh vss.t558 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1605 X1.X1.X2.X2.X2.X2.vout a_8486_31700# X1.X1.X2.X2.X2.X2.X3.vin1 vss.t645 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1606 X2.X1.X1.X1.X3.vin1 a_33976_29936# X2.X1.X1.X1.X1.X2.vout vss.t191 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1607 X2.X2.X1.X1.X2.vrefh a_46502_27070# X2.X2.X1.X1.X1.X2.X3.vin2 vdd.t392 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1608 vdd.t859 d1.t91 a_38152_16452# vdd.t858 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1609 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1610 a_4782_20446# a_4396_20446# vss.t1418 vss.t1417 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1611 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1612 X2.X1.X3.vin2.t3 a_35312_892# X2.X3.vin1 vdd.t1382 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1613 vdd.t112 a_54992_30794# a_54606_30794# vdd.t111 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1614 a_17222_4198# a_16836_4198# vss.t1530 vss.t1529 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1615 a_16836_6104# d0.t184 vdd.t1289 vdd.t1288 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1616 X2.X1.X2.X1.X2.X2.X1.vin2 a_40352_15546# X2.X1.X2.X1.X2.X2.X3.vin1 vss.t1440 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1617 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1618 X2.X1.X1.X2.X3.vin2 a_33976_7064# X2.X1.X1.X2.X2.X1.vout vdd.t749 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1619 X1.X2.X2.X1.X2.X1.X2.vin1 a_25712_13640# X1.X2.X2.X1.X2.X1.X3.vin2 vdd.t67 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1620 a_34362_26164# a_33976_26164# vdd.t1516 vdd.t1515 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1621 vdd.t1291 d0.t185 a_40352_23170# vdd.t1290 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1622 vss.t1301 a_23512_5016# a_23126_5016# vss.t1300 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1623 X2.X2.X1.X2.X1.X1.X3.vin1 a_48702_16634# X2.X2.X1.X2.X1.X1.vout vss.t1184 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1624 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1625 X2.X1.X1.X2.X1.X2.vout a_33676_12822# X2.X1.X1.X2.X1.X2.X3.vin1 vdd.t1403 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1626 X2.X1.X2.X2.X3.vin2 a_37852_25982# X2.X1.X2.X3.vin2 vss.t740 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1627 X1.X1.X1.X1.X2.X1.X3.vin1 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin2 vss.t73 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1628 X2.X2.X1.X1.X1.X1.X3.vin2 a_46116_30882# X2.X2.X1.X1.X1.X2.vrefh vss.t644 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1629 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1630 vss.t356 a_54992_4110# a_54606_4110# vss.t355 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1631 a_2196_6104# d0.t186 vss.t1317 vss.t1316 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1632 X1.X1.X1.X2.X2.X1.X3.vin1 a_4782_9010# X1.X1.X1.X2.X2.X1.vout vss.t770 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1633 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1634 X2.X1.X1.X1.X2.X1.X2.vin1 a_31862_23258# X2.X1.X1.X1.X2.X1.X3.vin2 vss.t707 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1635 vdd.t753 a_8872_31700# a_8486_31700# vdd.t752 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1636 a_2582_13728# a_2196_13728# vdd.t726 vdd.t725 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1637 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1638 X2.X2.X2.X1.X2.X1.X3.vin1 a_54606_11734# X2.X2.X2.X1.X2.X1.X1.vin1 vss.t930 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1639 X1.X2.X2.X1.X2.X2.X3.vin1 a_25326_15546# X1.X2.X2.X1.X2.X2.X1.vin1 vss.t1120 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1640 a_31476_28976# d0.t187 vss.t1319 vss.t1318 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1641 X1.X2.X2.X2.X2.X2.vout a_23126_31700# X1.X2.X2.X2.X2.X2.X3.vin1 vss.t1179 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1642 X2.X2.X1.X2.X3.vin1 a_48616_14688# X2.X2.X1.X2.X1.X1.vout vdd.t276 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1643 X1.X1.X1.X1.X2.X2.X2.vin1 a_2582_19446# X1.X1.X1.X1.X2.X2.X3.vin2 vss.t1285 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1644 a_19336_26164# d3.t20 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1645 a_19336_7064# d2.t41 vss.t864 vss.t863 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1646 X1.X1.X2.X1.X2.X2.vout a_8486_16452# X1.X1.X2.X1.X2.X2.X3.vin2 vdd.t958 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1647 X1.X1.X1.X1.X1.X1.X3.vin2 a_4782_31882# X1.X1.X1.X1.X1.X1.vout vdd.t422 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1648 vdd.t673 a_52492_25982# a_52106_25982# vdd.t672 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1649 X1.X1.X1.X2.X2.X1.vout a_4396_9010# X1.X1.X1.X2.X2.X1.X3.vin1 vdd.t1234 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1650 a_46502_30882# a_46116_30882# vss.t643 vss.t642 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1651 a_34062_20446# a_33676_20446# vdd.t1194 vdd.t1193 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1652 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1653 vdd.t1376 d4.t11 a_23212_18358# vdd.t1375 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1654 vdd.t1293 d0.t188 a_11072_32700# vdd.t1292 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1655 vss.t1321 d0.t189 a_11072_30794# vss.t1320 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1656 a_19036_5198# d1.t92 vdd.t861 vdd.t860 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1657 a_46502_9916# a_46116_9916# vss.t134 vss.t133 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1658 vdd.t1295 d0.t190 a_11072_9828# vdd.t1294 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1659 a_4782_16634# a_4396_16634# vdd.t1262 vdd.t1261 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1660 X2.X2.X2.X1.X2.X2.vrefh a_54992_13640# X2.X2.X2.X1.X2.X1.X3.vin2 vss.t815 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1661 X1.X2.X1.X1.X2.X1.X3.vin2 a_16836_23258# X1.X2.X1.X1.X2.X2.vrefh vss.t783 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1662 vdd.t863 d1.t93 a_23512_8828# vdd.t862 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1663 X1.X1.X1.X2.X2.X1.X3.vin2 a_2196_8010# X1.X1.X1.X2.X2.X2.vrefh vss.t1188 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1664 X1.X2.X1.X2.X2.X2.X1.vin1 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin1 vss.t756 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1665 a_34362_22312# a_33976_22312# vss.t1538 vss.t1537 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1666 vss.t1246 a_52792_20264# a_52406_20264# vss.t1245 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1667 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1668 a_46116_19446# d0.t191 vdd.t1297 vdd.t1296 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1669 a_28096_892# d7.t1 vdd.t1187 vdd.t1186 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1670 a_2582_4198# a_2196_4198# vss.t1226 vss.t1225 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1671 vss.t1323 d0.t192 a_40352_32700# vss.t1322 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1672 a_17222_11822# a_16836_11822# vdd.t400 vdd.t399 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1673 X2.X1.X1.X2.X1.X1.vout a_34362_14688# X2.X1.X1.X2.X3.vin1 vss.t699 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1674 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 vss.t242 sky130_fd_pr__res_high_po_0p35 l=1.09
X1675 a_2196_23258# d0.t193 vss.t1325 vss.t1324 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1676 a_2582_11822# a_2196_11822# vss.t157 vss.t156 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1677 X2.X2.X2.X3.vin1 a_52106_10734# X2.X2.X2.X1.X3.vin2 vdd.t1443 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1678 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1679 a_19036_20446# d1.t94 vdd.t865 vdd.t864 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1680 X1.X1.X1.X2.vrefh X1.X1.X1.X1.X2.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1681 X2.X2.X1.X1.X1.X2.X3.vin2 a_46116_27070# X2.X2.X1.X1.X1.X2.X2.vin1 vdd.t1141 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1682 X2.X2.X2.X1.X2.X1.vout a_52406_12640# X2.X2.X2.X1.X2.X1.X3.vin2 vdd.t683 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1683 a_4696_29936# d2.t42 vdd.t840 vdd.t839 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1684 X2.X2.X2.X2.X1.X1.X2.vin1 a_54992_21264# X2.X2.X2.X2.X1.X1.X3.vin2 vdd.t637 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1685 X2.X2.X2.X1.X1.X1.X3.vin2 a_54606_6016# X2.X2.X2.X1.X1.X2.vrefh vdd.t1033 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1686 X1.X2.X2.X1.X2.X2.vout a_23126_16452# X1.X2.X2.X1.X2.X2.X3.vin2 vdd.t620 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1687 a_2582_25164# a_2196_25164# vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1688 X2.X2.X2.X1.X1.X1.X1.vin1 X2.X2.X2.vrefh.t3 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1689 X2.X1.X2.X1.X2.X1.X3.vin2 a_39966_13640# X2.X1.X2.X1.X2.X1.X2.vin1 vss.t1116 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1690 X1.X1.X2.X1.X1.X1.X3.vin1 a_10686_4110# X1.X1.X2.X1.X1.X1.X1.vin1 vss.t132 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1691 a_33676_24258# d1.t95 vdd.t867 vdd.t866 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1692 a_19336_22312# d2.t43 vss.t866 vss.t865 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1693 vss.t1389 a_54992_23170# a_54606_23170# vss.t1388 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1694 a_46116_25164# d0.t194 vss.t1327 vss.t1326 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1695 a_33976_26164# d3.t21 vdd.t100 vdd.t99 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1696 X1.X2.X3.vin2.t3 a_20672_892# X1.X3.vin2 vdd.t1095 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1697 vss.t1329 d0.t195 a_54992_11734# vss.t1328 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1698 X2.X2.X1.X2.X1.X1.vout a_48316_16634# X2.X2.X1.X2.X1.X1.X3.vin2 vss.t831 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1699 vss.t1331 d0.t196 a_25712_15546# vss.t1330 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1700 vdd.t1184 a_40352_23170# a_39966_23170# vdd.t1183 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1701 vdd.t914 a_11072_26982# a_10686_26982# vdd.t913 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1702 a_17222_17540# a_16836_17540# vss.t224 vss.t223 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1703 vss.t889 d1.t96 a_23512_31700# vss.t888 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1704 vss.t543 a_11072_25076# a_10686_25076# vss.t542 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1705 vdd.t1299 d0.t197 a_11072_15546# vdd.t1298 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1706 X2.X1.X2.vrefh.t3 a_31862_4198# X2.X1.X1.X2.X2.X2.X3.vin2 vdd.t314 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1707 X1.X2.X1.X2.X3.vin2 a_19336_7064# X1.X2.X1.X2.X2.X1.vout vdd.t1028 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1708 vss.t868 d2.t44 a_37852_14586# vss.t867 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1709 X1.X2.X2.X2.X1.X2.vrefh a_25712_21264# X1.X2.X2.X2.X1.X1.X3.vin2 vss.t332 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1710 vdd.t1232 a_40352_7922# a_39966_7922# vdd.t1231 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1711 X2.X1.X2.X1.X1.X1.X3.vin1 a_39966_4110# X2.X1.X2.X1.X1.X1.X1.vin1 vss.t236 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1712 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1713 a_46502_27070# a_46116_27070# vdd.t1140 vdd.t1139 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1714 a_4696_7064# d2.t45 vss.t817 vss.t816 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1715 X2.X1.X2.X1.X3.vin1 a_37466_6962# X2.X1.X2.X1.X1.X1.vout vss.t155 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1716 vdd.t880 a_25712_28888# a_25326_28888# vdd.t879 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1717 a_34062_9010# a_33676_9010# vss.t29 vss.t28 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1718 X2.X1.X2.X2.X1.X1.X3.vin2 a_39966_21264# X2.X1.X2.X2.X1.X2.vrefh vdd.t191 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1719 X2.X2.X2.X2.X2.X2.X3.vin1 a_54606_30794# X2.X2.X2.X2.X2.X2.X1.vin2 vdd.t947 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1720 vss.t110 d3.t22 a_8572_10734# vss.t109 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1721 vdd.t1301 d0.t198 a_40352_17452# vdd.t1300 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1722 vss.t725 a_38152_5016# a_37766_5016# vss.t724 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1723 X2.X2.X2.X1.X1.X2.vout a_52406_8828# X2.X2.X2.X1.X1.X2.X3.vin1 vss.t317 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1724 vss.t891 d1.t97 a_8872_12640# vss.t890 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1725 X1.X1.X1.X1.X2.X2.vrefh a_2582_23258# X1.X1.X1.X1.X2.X1.X3.vin2 vdd.t1138 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1726 a_48702_16634# a_48316_16634# vss.t830 vss.t829 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1727 X1.X1.X1.X1.X2.X2.X3.vin2 a_2196_19446# X1.X1.X1.X2.vrefh vss.t833 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1728 a_31862_11822# a_31476_11822# vdd.t946 vdd.t945 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1729 X2.X2.X1.X2.X2.X1.X1.vin1 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin1 vss.t1422 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1730 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1731 a_33676_9010# d1.t98 vdd.t869 vdd.t868 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1732 X2.X2.X1.X2.vrefh a_46502_19446# X2.X2.X1.X1.X2.X2.X3.vin2 vdd.t1434 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1733 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1734 X1.X1.X1.X1.X2.X1.vout a_4396_24258# X1.X1.X1.X1.X2.X1.X3.vin2 vss.t715 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1735 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1736 X1.X1.X2.X1.X1.X2.X1.vin1 a_11072_7922# X1.X1.X2.X1.X1.X2.X3.vin1 vdd.t927 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1737 X1.X1.X1.X2.X1.X2.X3.vin1 a_4782_12822# X1.X1.X1.X2.X1.X2.vout vss.t261 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1738 X1.X2.X2.X2.X2.X2.X2.vin1 X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1739 vdd.t102 d3.t23 a_52492_10734# vdd.t101 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1740 X2.X2.X2.X2.X2.X2.X2.vin1 a_54992_32700# X2.X2.X2.X2.X2.X2.X3.vin2 vdd.t1446 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1741 X2.X2.X2.X2.X2.X2.X1.vin2 a_54992_30794# X2.X2.X2.X2.X2.X2.X3.vin1 vss.t123 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1742 X3.vin2.t2 a_42976_892# X2.X3.vin1 vdd.t1172 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1743 vdd.t871 d1.t99 a_52792_12640# vdd.t870 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1744 vss.t359 a_11072_9828# a_10686_9828# vss.t358 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1745 vdd.t873 d1.t100 a_23512_16452# vdd.t872 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1746 vdd.t812 d1.t101 a_8872_20264# vdd.t811 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1747 a_33976_22312# d2.t46 vss.t819 vss.t818 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1748 X1.X1.X2.X1.X3.vin2 a_8186_14586# X1.X1.X2.X1.X2.X1.vout vss.t545 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1749 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1750 X2.X2.X2.X1.X1.X1.X1.vin1 a_54992_4110# X2.X2.X2.X1.X1.X1.X3.vin1 vdd.t347 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1751 a_48616_14688# d2.t47 vdd.t791 vdd.t790 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1752 a_31862_17540# a_31476_17540# vss.t1309 vss.t1308 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1753 vss.t519 a_40352_32700# a_39966_32700# vss.t518 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1754 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1755 a_17222_28976# a_16836_28976# vss.t311 vss.t310 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1756 X2.X2.X1.X1.X2.X1.X1.vin1 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin1 vss.t243 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1757 vdd.t1069 a_54992_6016# a_54606_6016# vdd.t1068 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1758 a_16836_11822# d0.t199 vdd.t1303 vdd.t1302 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1759 X1.X1.X2.X1.X2.X1.X2.vin1 a_11072_13640# X1.X1.X2.X1.X2.X1.X3.vin2 vdd.t1144 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1760 X2.X1.X1.X2.X3.vin1 a_33976_14688# X2.X1.X1.X2.X1.X2.vout vss.t1232 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1761 a_4696_26164# d3.t24 vss.t112 vss.t111 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1762 X2.X1.X2.X3.vin2 a_37852_18358# X2.X1.X3.vin2.t2 vss.t428 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1763 X2.X1.X1.X1.X2.X2.X3.vin1 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin1 vdd.t1132 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1764 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1765 X2.vrefh X2.X1.X1.X1.X1.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1766 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1767 vdd.t1456 d3.t25 a_37852_25982# vdd.t1455 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1768 X1.X1.X2.X2.X2.X2.X3.vin2 a_8872_31700# X1.X1.X2.X2.X2.X2.vout vss.t782 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1769 X1.X1.X1.X2.X2.X2.vrefh a_2582_8010# X1.X1.X1.X2.X2.X1.X3.vin2 vdd.t417 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1770 vdd.t1240 a_37852_10734# a_37466_10734# vdd.t1239 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1771 X2.X1.X2.X2.X2.X2.X3.vin2 a_39966_32700# X2.X2.vrefh vdd.t269 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1772 X2.X1.X2.X2.X2.X2.X3.vin1 a_39966_30794# X2.X1.X2.X2.X2.X2.X1.vin1 vss.t450 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1773 vdd.t228 a_38152_12640# a_37766_12640# vdd.t227 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1774 vdd.t4 d0.t200 a_54992_30794# vdd.t3 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1775 vss.t4 d0.t201 a_40352_26982# vss.t3 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1776 X2.X2.X2.X2.X1.X1.vout a_52406_20264# X2.X2.X2.X2.X1.X1.X3.vin1 vss.t1248 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1777 X2.X2.X2.X2.X2.X2.X2.vin1 X2.X2.X2.X2.X2.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1778 a_13696_892# d6.t2 vss.t1017 vss.t1016 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1779 a_16836_17540# d0.t202 vss.t6 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1780 vss.t1437 a_23512_31700# a_23126_31700# vss.t1436 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1781 X1.X2.X1.X1.X1.X2.vout a_19722_29936# X1.X2.X1.X1.X3.vin1 vdd.t412 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1782 X2.X1.X1.X1.X1.X2.X3.vin2 a_31476_27070# X2.X1.X1.X1.X2.vrefh vss.t603 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1783 vss.t302 a_8872_8828# a_8486_8828# vss.t301 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1784 X2.X2.X2.X1.X2.X2.X1.vin1 a_54992_15546# X2.X2.X2.X1.X2.X2.X3.vin1 vdd.t313 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1785 X2.X1.X1.X2.X1.X2.X3.vin2 a_34062_12822# X2.X1.X1.X2.X1.X2.vout vdd.t246 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1786 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1787 X2.X1.X2.X2.X2.X1.X2.vin1 a_40352_28888# X2.X1.X2.X2.X2.X1.X3.vin2 vdd.t718 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1788 vss.t977 a_52792_8828# a_52406_8828# vss.t976 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1789 vdd.t793 d2.t48 a_8572_29834# vdd.t792 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1790 X1.X2.X2.X1.X1.X1.X3.vin1 a_25326_4110# X1.X2.X2.X1.X1.X1.X1.vin1 vss.t1114 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1791 vss.t169 a_54992_17452# a_54606_17452# vss.t168 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1792 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1793 a_46116_19446# d0.t203 vss.t8 vss.t7 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1794 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1795 vss.t768 a_8572_10734# a_8186_10734# vss.t767 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1796 vdd.t1100 a_40352_17452# a_39966_17452# vdd.t1099 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1797 vdd.t814 d1.t102 a_8872_31700# vdd.t813 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1798 X2.X2.X2.X2.X1.X2.X3.vin1 a_54606_23170# X2.X2.X2.X2.X1.X2.X1.vin1 vss.t104 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1799 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1800 a_48316_31882# d1.t103 vdd.t816 vdd.t815 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1801 X1.X1.X1.X1.X2.X1.X3.vin2 a_2196_23258# X1.X1.X1.X1.X2.X1.X2.vin1 vdd.t354 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1802 X1.X2.X2.X1.X2.X2.X1.vin2 a_25712_15546# X1.X2.X2.X1.X2.X2.X3.vin1 vss.t1117 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1803 a_31862_28976# a_31476_28976# vss.t1424 vss.t1423 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1804 a_19422_24258# a_19036_24258# vdd.t138 vdd.t137 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1805 X1.X2.X2.X2.X2.X2.X3.vin2 a_23512_31700# X1.X2.X2.X2.X2.X2.vout vss.t1435 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1806 X1.X1.X2.X3.vin2 a_8186_25982# X1.X1.X2.X2.X3.vin2 vdd.t1381 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1807 X1.X2.X1.X2.X2.X2.X3.vin2 a_16836_4198# X1.X2.X2.vrefh.t3 vss.t1528 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1808 X2.X2.X1.X2.X1.X2.vout a_49002_14688# X2.X2.X1.X2.X3.vin1 vdd.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1809 a_4696_29936# d2.t49 vss.t821 vss.t820 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1810 a_19722_26164# a_19336_26164# vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1811 X2.X2.X1.X1.X2.X2.X3.vin2 a_46116_19446# X2.X2.X1.X1.X2.X2.X2.vin1 vdd.t454 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1812 X1.X1.X2.X1.X2.X2.X3.vin1 a_8872_16452# X1.X1.X2.X1.X2.X2.vout vdd.t281 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1813 X1.X2.X1.X2.X2.vrefh a_17222_11822# X1.X2.X1.X2.X1.X2.X3.vin2 vdd.t547 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1814 a_2196_4198# d0.t204 vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1815 a_48702_9010# a_48316_9010# vss.t274 vss.t273 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1816 X1.X2.X1.X2.X1.X2.vout a_19036_12822# X1.X2.X1.X2.X1.X2.X3.vin1 vdd.t744 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1817 X2.X1.X2.X1.X2.X2.X3.vin1 a_39966_15546# X2.X1.X2.X1.X2.X2.X1.vin2 vdd.t1427 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1818 X1.X1.X2.X1.X1.X1.X3.vin2 a_10686_6016# X1.X1.X2.X1.X1.X2.vrefh vdd.t538 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1819 X1.X2.X2.X2.X2.X1.X3.vin2 a_25326_28888# X1.X2.X2.X2.X2.X2.vrefh vdd.t881 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1820 vdd.t1117 a_54992_25076# a_54606_25076# vdd.t1116 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1821 vdd.t1073 a_52492_10734# a_52106_10734# vdd.t1072 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1822 vdd.t320 a_23512_16452# a_23126_16452# vdd.t319 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1823 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1824 X2.X1.X2.X1.X1.X1.X3.vin2 a_39966_6016# X2.X1.X2.X1.X1.X2.vrefh vdd.t1178 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1825 a_4396_12822# d1.t104 vdd.t818 vdd.t817 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1826 a_48316_9010# d1.t105 vdd.t820 vdd.t819 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1827 X2.X2.X2.X1.X1.X2.vrefh a_54992_6016# X2.X2.X2.X1.X1.X1.X3.vin2 vss.t1094 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1828 vss.t842 d1.t106 a_52792_20264# vss.t841 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1829 a_16836_28976# d0.t205 vss.t10 vss.t9 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1830 X2.X2.X1.X1.X2.X1.X3.vin1 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin2 vss.t933 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1831 X1.X1.X2.X1.X2.X1.X3.vin2 a_10686_13640# X1.X1.X2.X1.X2.X2.vrefh vdd.t1147 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1832 a_46502_19446# a_46116_19446# vdd.t453 vdd.t452 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1833 X2.X1.X2.X1.X1.X1.X1.vin1 a_40352_4110# X2.X1.X2.X1.X1.X1.X3.vin1 vdd.t1036 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1834 X1.X2.X1.X2.X1.X1.X1.vin1 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin1 vss.t425 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1835 X1.X1.X1.X2.X2.X2.X3.vin1 a_4782_5198# X1.X1.X1.X2.X2.X2.vout vss.t293 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1836 a_2582_23258# a_2196_23258# vss.t363 vss.t362 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1837 vss.t1277 a_8872_24076# a_8486_24076# vss.t1276 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1838 X1.X2.X2.vrefh.t1 a_17222_4198# X1.X2.X1.X2.X2.X2.X3.vin2 vdd.t76 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1839 X1.X1.X2.X2.X1.X2.vrefh a_11072_21264# X1.X1.X2.X2.X1.X1.X3.vin2 vss.t1406 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1840 a_31862_8010# a_31476_8010# vdd.t685 vdd.t684 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1841 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1842 X2.X1.X2.X1.X2.X2.X3.vin2 a_38152_16452# X2.X1.X2.X1.X2.X2.vout vss.t524 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1843 a_5082_29936# a_4696_29936# vdd.t652 vdd.t651 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1844 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1845 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1846 X1.X2.X2.X1.X2.X2.X3.vin1 a_23512_16452# X1.X2.X2.X1.X2.X2.vout vdd.t318 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1847 vss.t648 a_40352_26982# a_39966_26982# vss.t647 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1848 X2.X1.X3.vin1.t2 a_35312_892# X2.X3.vin1 vss.t1398 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1849 X1.X2.X1.X1.X3.vin1 a_19722_26164# X1.X2.X1.X3.vin1 vss.t1115 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1850 X2.X2.X1.X1.X2.X2.X2.vin1 a_46502_19446# X2.X2.X1.X1.X2.X2.X3.vin2 vss.t1450 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1851 a_34062_24258# a_33676_24258# vdd.t329 vdd.t328 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1852 X1.X1.X2.X1.X1.X1.vout a_8572_6962# X1.X1.X2.X1.X3.vin1 vdd.t647 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1853 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1854 X2.X1.X1.X2.X1.X1.X3.vin2 a_31476_15634# X2.X1.X1.X2.X1.X1.X2.vin1 vdd.t1157 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1855 a_19722_22312# a_19336_22312# vss.t607 vss.t606 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1856 X2.X1.X1.X3.vin2 a_34362_18540# X2.X1.X3.vin1.t1 vdd.t928 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1857 vss.t12 d0.t206 a_54992_23170# vss.t11 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1858 X2.X2.X1.X1.X1.X1.X3.vin2 a_48702_31882# X2.X2.X1.X1.X1.X1.vout vdd.t423 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1859 a_46502_25164# a_46116_25164# vss.t932 vss.t931 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1860 vss.t1195 a_38152_20264# a_37766_20264# vss.t1194 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1861 X2.X2.X2.X1.X1.X1.vout a_52492_6962# X2.X2.X2.X1.X3.vin1 vdd.t1190 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1862 vdd.t8 d0.t207 a_11072_26982# vdd.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1863 vss.t732 a_25712_4110# a_25326_4110# vss.t731 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1864 X2.X1.X2.X1.X1.X2.vout a_37766_8828# X2.X1.X2.X1.X1.X2.X3.vin1 vss.t698 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1865 vss.t1282 a_25712_11734# a_25326_11734# vss.t1281 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1866 vss.t14 d0.t208 a_11072_25076# vss.t13 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1867 vdd.t822 d1.t107 a_8872_5016# vdd.t821 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1868 vdd.t1414 a_11072_11734# a_10686_11734# vdd.t1413 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1869 X1.X2.X1.X2.X2.X1.X3.vin1 a_19422_9010# X1.X2.X1.X2.X2.X1.vout vss.t537 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1870 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1871 vdd.t105 a_8572_29834# a_8186_29834# vdd.t104 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1872 X2.X1.X2.X2.X1.X2.X3.vin1 a_38152_24076# X2.X1.X2.X2.X1.X2.vout vdd.t321 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1873 X1.X1.X1.X2.X2.X2.X3.vin2 a_2196_4198# X1.X1.X2.vrefh.t3 vss.t1224 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1874 a_31476_30882# d0.t209 vss.t16 vss.t15 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1875 vdd.t824 d1.t108 a_52792_5016# vdd.t823 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1876 X1.X1.X1.X1.X2.X2.X1.vin1 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin1 vss.t1053 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1877 vdd.t10 d0.t210 a_25712_28888# vdd.t9 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1878 a_46116_23258# d0.t211 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1879 X2.X1.X1.X2.X3.vin2 a_34362_10916# X2.X1.X1.X3.vin2 vdd.t724 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1880 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1881 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X1882 X2.X2.X1.X2.X2.X1.X3.vin1 a_48702_9010# X2.X2.X1.X2.X2.X1.vout vss.t1231 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1883 a_19036_24258# d1.t109 vdd.t826 vdd.t825 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1884 X1.X1.X1.X2.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1885 a_17222_9916# a_16836_9916# vss.t652 vss.t651 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1886 a_48316_12822# d1.t110 vss.t844 vss.t843 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1887 X1.X1.X3.vin1 a_4696_18540# X1.X1.X1.X3.vin2 vss.t1432 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1888 X1.X2.X1.X1.X1.X2.X1.vin1 a_17222_28976# X1.X2.X1.X1.X1.X2.X3.vin1 vss.t361 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1889 vss.t823 d2.t50 a_23212_6962# vss.t822 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1890 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X1891 vss.t825 d2.t51 a_8572_29834# vss.t824 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1892 X2.X2.X2.X1.X2.X2.X3.vin2 a_52792_16452# X2.X2.X2.X1.X2.X2.vout vss.t400 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1893 X2.X2.X2.X1.X2.X2.X3.vin2 a_54606_17452# X2.X2.X2.X1.X2.X2.X2.vin1 vss.t276 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1894 X1.X1.X1.X1.X2.X1.X3.vin1 a_4782_24258# X1.X1.X1.X1.X2.X1.vout vss.t730 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1895 X2.X1.X1.X2.X1.X2.X3.vin1 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin2 vss.t198 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1896 X1.X1.X2.X1.X1.X2.X3.vin1 a_8872_8828# X1.X1.X2.X1.X1.X2.vout vdd.t293 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1897 X2.X2.X2.X1.X1.X2.X3.vin1 a_52792_8828# X2.X2.X2.X1.X1.X2.vout vdd.t952 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1898 X1.X2.X1.X1.X1.X1.vout a_19722_29936# X1.X2.X1.X1.X3.vin1 vss.t424 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1899 vss.t18 d0.t212 a_11072_9828# vss.t17 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1900 X1.X1.X1.X3.vin2 a_4696_10916# X1.X1.X1.X2.X3.vin2 vss.t1383 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1901 X1.X1.X2.X1.X2.X2.vout a_8572_14586# X1.X1.X2.X1.X3.vin2 vss.t907 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1902 X2.X2.X1.X2.X2.X1.X3.vin2 a_46116_8010# X2.X2.X1.X2.X2.X2.vrefh vss.t1165 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1903 a_49002_14688# a_48616_14688# vdd.t275 vdd.t274 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1904 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1905 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X1906 X1.X2.X1.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1907 X1.X2.X2.X1.X1.X1.X3.vin2 a_25326_6016# X1.X2.X2.X1.X1.X2.vrefh vdd.t1226 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1908 X3.vin2 a_42976_892# X2.X3.vin2 vss.t1200 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1909 vdd.t1104 a_54992_19358# a_54606_19358# vdd.t1103 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1910 vdd.t795 d2.t52 a_8572_22210# vdd.t794 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1911 X1.X1.X1.X2.X2.X2.X1.vin1 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin1 vss.t1524 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1912 a_34062_5198# a_33676_5198# vss.t1198 vss.t1197 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1913 X2.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X2.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1914 X2.X1.X2.X1.X1.X2.vrefh a_40352_6016# X2.X1.X2.X1.X1.X1.X3.vin2 vss.t161 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1915 a_5082_26164# a_4696_26164# vss.t1414 vss.t1413 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1916 X2.X2.X2.X2.X1.X2.X3.vin1 a_52792_24076# X2.X2.X2.X2.X1.X2.vout vdd.t231 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1917 X2.X1.X1.X1.X2.X2.X1.vin2 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin1 vdd.t611 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1918 X2.X2.X2.X2.X1.X2.X3.vin2 a_54606_25076# X2.X2.X2.X2.X2.vrefh vdd.t1119 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1919 X1.X1.X2.X2.X1.X1.X3.vin2 a_10686_21264# X1.X1.X2.X2.X1.X1.X2.vin1 vss.t549 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1920 vss.t247 a_23212_14586# a_22826_14586# vss.t246 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1921 X1.X2.X1.X2.X1.X2.X3.vin2 a_19422_12822# X1.X2.X1.X2.X1.X2.vout vdd.t675 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1922 X1.X1.X1.X1.X3.vin2 a_4696_22312# X1.X1.X1.X1.X2.X1.vout vdd.t299 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1923 X2.X1.X2.X1.X2.X2.vout a_37766_16452# X2.X1.X2.X1.X2.X2.X3.vin1 vss.t1193 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1924 X1.X1.X1.X1.X1.X1.X1.vin1 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin1 vss.t853 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1925 a_31476_27070# d0.t213 vdd.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1926 X1.X2.X3.vin1 a_19336_18540# X1.X2.X1.X3.vin2 vss.t1227 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1927 vdd.t1458 d3.t26 a_37852_10734# vdd.t1457 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1928 X2.X1.X1.X1.X1.X1.vout a_33676_31882# X2.X1.X1.X1.X1.X1.X3.vin2 vss.t741 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1929 X1.X1.X1.X2.X1.X1.X1.vin2 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin1 vdd.t1284 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1930 X2.X2.X1.X1.X2.X2.vrefh a_46502_23258# X2.X2.X1.X1.X2.X1.X3.vin2 vdd.t605 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1931 X2.X2.X1.X1.X2.X2.X3.vin2 a_46116_19446# X2.X2.X1.X2.vrefh vss.t464 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1932 a_6032_892# a_5646_892# vdd.t911 vdd.t910 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1933 vdd.t828 d1.t111 a_38152_12640# vdd.t827 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1934 vdd.t926 a_11072_7922# a_10686_7922# vdd.t925 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1935 X2.X1.X1.X1.X1.X1.X3.vin1 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin1 vdd.t759 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1936 X2.X1.X3.vin1.t0 a_33976_18540# X2.X1.X1.X3.vin1 vdd.t777 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1937 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X1938 X2.X2.X1.X1.X1.X1.vout a_48316_31882# X2.X2.X1.X1.X1.X1.X3.vin1 vdd.t526 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1939 vdd.t522 a_25712_30794# a_25326_30794# vdd.t521 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1940 X1.X1.X3.vin1.t1 a_6032_892# X1.X3.vin1 vss.t734 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1941 X2.X1.X2.X1.X2.X1.X1.vin2 a_40352_11734# X2.X1.X2.X1.X2.X1.X3.vin1 vss.t1451 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1942 vdd.t797 d2.t53 a_8572_14586# vdd.t796 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1943 a_33676_16634# d1.t112 vss.t846 vss.t845 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1944 X1.X1.X2.X1.X2.X2.X1.vin2 a_11072_15546# X1.X1.X2.X1.X2.X2.X3.vin1 vss.t582 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1945 vdd.t297 a_52792_27888# a_52406_27888# vdd.t296 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1946 X2.X1.X1.X1.X1.X2.X2.vin1 a_31862_27070# X2.X1.X1.X1.X1.X2.X3.vin2 vss.t436 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1947 a_46502_8010# a_46116_8010# vdd.t1136 vdd.t1135 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1948 X2.X2.X2.X2.X3.vin1 a_52106_22210# X2.X2.X2.X2.X1.X1.vout vss.t232 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1949 X2.X2.X2.X2.X2.X1.X1.vin1 a_54992_26982# X2.X2.X2.X2.X2.X1.X3.vin1 vdd.t730 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1950 X1.X2.X1.X3.vin2 a_19336_10916# X1.X2.X1.X2.X3.vin2 vss.t719 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1951 X2.X2.X1.X2.X1.X2.X3.vin1 a_48702_12822# X2.X2.X1.X2.X1.X2.vout vss.t1310 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1952 X2.X2.X2.X2.X2.vrefh a_54992_25076# X2.X2.X2.X2.X1.X2.X3.vin2 vss.t1142 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1953 X2.X1.X2.X2.X1.X2.vout a_37766_24076# X2.X1.X2.X2.X1.X2.X3.vin2 vdd.t1278 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1954 X1.X1.X1.X2.X2.X1.X1.vin2 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin1 vdd.t71 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1955 X1.X2.X2.X1.X2.X2.vout a_23212_14586# X1.X2.X2.X1.X3.vin2 vss.t245 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1956 X1.X2.X1.X1.X2.X2.X3.vin1 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin1 vdd.t980 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1957 vss.t20 d0.t214 a_54992_7922# vss.t19 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1958 X1.X2.X2.X1.X1.X2.vout a_23126_8828# X1.X2.X2.X1.X1.X2.X3.vin1 vss.t892 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1959 X1.X2.X2.X2.X2.X2.X1.vin1 X1.X2.X2.X2.X2.X2.vrefh vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1960 a_2582_9916# a_2196_9916# vss.t1405 vss.t1404 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1961 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X1962 X1.X1.X1.X1.X2.X2.X3.vin1 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin2 vss.t265 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1963 X2.X1.X1.X3.vin2 a_33976_10916# X2.X1.X1.X2.X3.vin1 vdd.t721 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1964 vss.t22 d0.t215 a_54992_17452# vss.t21 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1965 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1966 a_46502_19446# a_46116_19446# vss.t463 vss.t462 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1967 a_4696_14688# d2.t54 vss.t827 vss.t826 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1968 a_2196_21352# d0.t216 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1969 X1.X2.X1.X1.X3.vin2 a_19336_22312# X1.X2.X1.X1.X2.X1.vout vdd.t584 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1970 a_48702_31882# a_48316_31882# vdd.t525 vdd.t524 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1971 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1972 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X1973 X1.X1.X2.X2.X3.vin1 a_8572_25982# X1.X1.X2.X3.vin2 vdd.t140 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1974 X1.X2.X2.X1.X2.X1.X3.vin1 a_25326_11734# X1.X2.X2.X1.X2.X1.X1.vin1 vss.t1283 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1975 X3.vin1.t2 a_13696_892# X1.X3.vin1 vdd.t1113 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1976 a_5082_29936# a_4696_29936# vss.t680 vss.t679 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1977 vss.t1069 a_54992_28888# a_54606_28888# vss.t1068 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1978 X1.X1.X2.X3.vin1 a_8186_10734# X1.X1.X2.X1.X3.vin2 vdd.t1122 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1979 X1.X1.X1.X2.X1.X1.X2.vin1 a_2582_15634# X1.X1.X1.X2.X1.X1.X3.vin2 vss.t1049 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1980 X1.X2.X1.X1.X1.X2.X3.vin2 a_16836_27070# X1.X2.X1.X1.X2.vrefh vss.t194 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1981 a_20286_892# d5.t7 vss.t42 vss.t41 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1982 X2.X1.X2.X2.X2.X1.X3.vin1 a_39966_26982# X2.X1.X2.X2.X2.X1.X1.vin2 vdd.t477 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1983 vss.t24 d0.t217 a_11072_4110# vss.t23 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1984 X1.X1.X2.X1.X2.X1.vout a_8486_12640# X1.X1.X2.X1.X2.X1.X3.vin2 vdd.t115 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1985 vss.t115 a_8572_29834# a_8186_29834# vss.t114 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1986 X2.X1.X2.X2.X1.X2.X3.vin2 a_39966_25076# X2.X1.X2.X2.X1.X2.X2.vin1 vss.t551 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1987 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X1988 X1.X1.X1.X2.X2.X2.vout a_4396_5198# X1.X1.X1.X2.X2.X2.X3.vin1 vdd.t948 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1989 X1.X2.X2.X2.X2.X1.X2.vin1 a_25712_28888# X1.X2.X2.X2.X2.X1.X3.vin2 vdd.t878 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1990 vdd.t1482 d0.t218 a_54992_25076# vdd.t1481 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1991 vdd.t1395 a_23212_25982# a_22826_25982# vdd.t1394 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1992 a_17222_30882# a_16836_30882# vss.t263 vss.t262 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1993 vdd.t224 a_25712_6016# a_25326_6016# vdd.t223 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1994 X1.X1.X1.X1.X1.X2.X1.vin2 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin1 vdd.t548 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1995 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X1996 X2.X1.X1.X1.X1.X2.vout a_33676_28070# X2.X1.X1.X1.X1.X2.X3.vin1 vdd.t1214 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1997 a_2196_27070# d0.t219 vss.t1498 vss.t1497 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1998 X2.X2.X2.X1.X2.vrefh a_54992_9828# X2.X2.X2.X1.X1.X2.X3.vin2 vss.t101 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1999 a_4782_12822# a_4396_12822# vdd.t609 vdd.t608 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2000 vss.t443 d2.t55 a_37852_6962# vss.t442 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2001 X1.X1.X1.X2.X2.X1.vout a_5082_7064# X1.X1.X1.X2.X3.vin2 vss.t1275 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2002 a_31862_6104# a_31476_6104# vss.t493 vss.t492 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2003 vdd.t1440 a_8572_22210# a_8186_22210# vdd.t1439 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2004 X2.X2.X2.X3.vin2 a_52106_25982# X2.X2.X2.X2.X3.vin1 vss.t1191 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2005 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X2.vrefh vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X2006 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X2007 X2.X1.X1.X2.X2.X1.X3.vin2 a_31476_8010# X2.X1.X1.X2.X2.X2.vrefh vss.t712 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2008 X1.X1.X1.X2.X2.X2.vrefh X1.X1.X1.X2.X2.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X2009 vss.t445 d2.t56 a_52492_22210# vss.t444 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2010 X1.X1.X1.X1.X1.X1.X3.vin1 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin2 vss.t1108 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2011 X2.X2.X1.X1.X1.X1.X1.vin2 X2.X2.X1.X1.X1.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X2012 X1.X2.X2.X2.X3.vin1 a_23212_25982# X1.X2.X2.X3.vin2 vdd.t1393 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2013 vss.t848 d1.t113 a_8872_24076# vss.t847 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2014 X1.X1.X1.X2.X3.vin2 a_4696_7064# X1.X1.X1.X2.X2.X1.vout vdd.t1244 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2015 a_31476_6104# d0.t220 vdd.t1484 vdd.t1483 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2016 X1.X1.X1.X2.X1.X1.X3.vin1 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin1 vdd.t1179 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2017 X2.X1.X1.X2.X2.X1.X3.vin2 a_34062_9010# X2.X1.X1.X2.X2.X1.vout vdd.t20 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2018 X2.X2.X1.X1.X2.X1.X3.vin2 a_46116_23258# X2.X2.X1.X1.X2.X1.X2.vin1 vdd.t222 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2019 X2.X2.X1.X2.X2.X2.vrefh a_46502_8010# X2.X2.X1.X2.X2.X1.X3.vin2 vdd.t1124 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2020 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X2021 X1.X2.X2.X1.X2.X1.vout a_23126_12640# X1.X2.X2.X1.X2.X1.X3.vin2 vdd.t1506 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2022 X2.X1.X2.X2.X2.X2.X1.vin1 a_40352_30794# X2.X1.X2.X2.X2.X2.X3.vin1 vdd.t393 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2023 a_48702_5198# a_48316_5198# vss.t677 vss.t676 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2024 X2.X1.X2.X1.X1.X2.X3.vin2 a_39966_9828# X2.X1.X2.X1.X1.X2.X2.vin1 vss.t1062 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2025 vdd.t890 a_8572_14586# a_8186_14586# vdd.t889 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2026 X2.X1.X1.X2.X1.X2.vrefh a_31862_15634# X2.X1.X1.X2.X1.X1.X3.vin2 vdd.t387 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2027 X1.X1.X2.X1.X2.X2.X3.vin1 a_10686_15546# X1.X1.X2.X1.X2.X2.X1.vin1 vss.t166 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2028 X2.X2.X2.X2.X1.X1.X3.vin1 a_54606_19358# X2.X2.X2.X2.X1.X1.X1.vin2 vdd.t157 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2029 vss.t850 d1.t114 a_38152_20264# vss.t849 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2030 vss.t1130 a_54992_19358# a_54606_19358# vss.t1129 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2031 X2.X1.X2.X2.X2.X1.X3.vin2 a_38152_27888# X2.X1.X2.X2.X2.X1.vout vss.t1135 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2032 a_46116_21352# d0.t221 vss.t1500 vss.t1499 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2033 vss.t901 a_25712_23170# a_25326_23170# vss.t900 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2034 X1.X1.X1.X2.X2.X1.X3.vin1 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin1 vdd.t1387 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2035 X2.X2.X1.X2.X1.X2.vout a_48316_12822# X2.X2.X1.X2.X1.X2.X3.vin2 vss.t1240 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2036 vss.t1502 d0.t222 a_25712_11734# vss.t1501 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2037 X1.X2.X2.X1.X3.vin2 a_22826_14586# X1.X2.X2.X1.X2.X1.vout vss.t248 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2038 vdd.t737 a_11072_23170# a_10686_23170# vdd.t736 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2039 vdd.t1486 d0.t223 a_11072_11734# vdd.t1485 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2040 vss.t118 a_37852_22210# a_37466_22210# vss.t117 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2041 X1.X2.X2.X1.X1.X1.X3.vin1 a_23512_5016# X1.X2.X2.X1.X1.X1.vout vdd.t1272 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2042 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X2043 vdd.t1035 a_40352_4110# a_39966_4110# vdd.t1034 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2044 a_31862_30882# a_31476_30882# vss.t409 vss.t408 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2045 a_46502_23258# a_46116_23258# vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2046 vss.t1504 d0.t224 a_40352_7922# vss.t1503 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2047 a_17222_27070# a_16836_27070# vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2048 a_19422_9010# a_19036_9010# vss.t184 vss.t183 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2049 X1.X2.X2.X2.X2.X2.X3.vin1 a_25326_30794# X1.X2.X2.X2.X2.X2.X1.vin2 vdd.t1025 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2050 vdd.t1488 d0.t225 a_40352_13640# vdd.t1487 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2051 X1.X1.X1.X1.X1.X2.vout a_4396_28070# X1.X1.X1.X1.X1.X2.X3.vin2 vss.t806 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2052 X1.X2.X1.X2.X1.X1.X3.vin2 a_16836_15634# X1.X2.X1.X2.X1.X1.X2.vin1 vdd.t1267 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2053 X2.X2.X2.X2.X2.X1.vout a_52406_27888# X2.X2.X2.X2.X2.X1.X3.vin2 vdd.t929 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2054 X2.X2.X2.X1.X1.X1.vout a_52406_5016# X2.X2.X2.X1.X1.X1.X3.vin1 vss.t1172 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2055 a_48316_24258# d1.t115 vss.t852 vss.t851 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2056 a_34362_14688# a_33976_14688# vdd.t1205 vdd.t1204 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2057 vdd.t646 a_8572_6962# a_8186_6962# vdd.t645 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2058 a_48702_12822# a_48316_12822# vss.t1239 vss.t1238 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2059 X1.X1.X1.X2.X1.X1.X3.vin2 a_2196_15634# X1.X1.X1.X2.X1.X2.vrefh vss.t1101 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2060 X1.X1.X1.X3.vin1 a_5082_18540# X1.X1.X3.vin1 vss.t687 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2061 a_31476_19446# d0.t226 vdd.t1490 vdd.t1489 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2062 a_19422_16634# a_19036_16634# vss.t96 vss.t95 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2063 vss.t1472 d3.t27 a_52492_25982# vss.t1471 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2064 a_33676_5198# d1.t116 vdd.t895 vdd.t894 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2065 X2.X1.X2.X1.X1.X1.X1.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X2066 X1.X2.X1.X2.X1.X1.vout a_19722_14688# X1.X2.X1.X2.X3.vin1 vss.t1054 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2067 vdd.t1189 a_52492_6962# a_52106_6962# vdd.t1188 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2068 a_16836_30882# d0.t227 vss.t1506 vss.t1505 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2069 X2.X1.X1.X2.X1.X2.X1.vin1 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin1 vss.t517 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2070 a_2196_15634# d0.t228 vdd.t1492 vdd.t1491 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2071 X1.X1.X1.X1.X1.X2.X3.vin1 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin1 vdd.t337 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2072 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X2073 X1.X1.X2.X2.X1.X1.vout a_8486_20264# X1.X1.X2.X2.X1.X1.X3.vin1 vss.t281 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2074 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X2075 X1.X1.X1.X1.X2.X2.vout a_4396_20446# X1.X1.X1.X1.X2.X2.X3.vin2 vss.t1416 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2076 X1.X1.X2.X1.X1.X1.X1.vin1 a_11072_4110# X1.X1.X2.X1.X1.X1.X3.vin1 vdd.t126 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2077 X1.X1.X1.X2.X3.vin1 a_5082_10916# X1.X1.X1.X3.vin2 vss.t988 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2078 vdd.t1494 d0.t229 a_54992_9828# vdd.t1493 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2079 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X2.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X2080 a_16836_8010# d0.t230 vss.t1508 vss.t1507 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2081 vdd.t897 d1.t117 a_23512_12640# vdd.t896 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2082 X1.X2.X1.X2.X2.X2.X3.vin1 a_19422_5198# X1.X2.X1.X2.X2.X2.vout vss.t1219 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2083 X2.X2.X2.X2.X2.X1.X3.vin2 a_52792_27888# X2.X2.X2.X2.X2.X1.vout vss.t304 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2084 X2.X2.X2.X2.X2.X1.X3.vin2 a_54606_28888# X2.X2.X2.X2.X2.X1.X2.vin1 vss.t113 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2085 a_31476_25164# d0.t231 vss.t1510 vss.t1509 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2086 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X1.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X2087 a_46116_32788# d0.t232 vss.t1512 vss.t1511 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2088 a_19336_14688# d2.t57 vdd.t431 vdd.t430 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2089 vdd.t1496 d0.t233 a_54992_19358# vdd.t1495 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2090 a_46116_17540# d0.t234 vdd.t1498 vdd.t1497 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2091 X2.X2.X1.X1.X2.X2.X1.vin1 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin1 vss.t369 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2092 vss.t870 a_52492_22210# a_52106_22210# vss.t869 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2093 vss.t349 a_11072_32700# a_10686_32700# vss.t348 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2094 vss.t739 a_37852_25982# a_37466_25982# vss.t738 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2095 a_33976_7064# d2.t58 vdd.t433 vdd.t432 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2096 X1.X2.X1.X2.X2.X1.X3.vin1 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin2 vss.t650 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2097 vss.t447 d2.t59 a_23212_14586# vss.t446 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2098 X1.X2.X2.X3.vin2 a_22826_25982# X1.X2.X2.X2.X3.vin2 vdd.t277 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2099 X2.X2.X1.X2.X2.X2.X3.vin1 a_48702_5198# X2.X2.X1.X2.X2.X2.vout vss.t1087 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2100 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X2101 X1.X1.X1.X1.X2.X2.vout a_5082_22312# X1.X1.X1.X1.X3.vin2 vdd.t502 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2102 a_31862_27070# a_31476_27070# vdd.t582 vdd.t581 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2103 X1.X2.X1.X2.X1.X2.X3.vin1 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin2 vss.t162 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2104 X2.X1.X1.X1.X1.X1.X3.vin1 a_34062_31882# X2.X1.X1.X1.X1.X1.vout vss.t744 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2105 X1.X1.X2.vrefh.t1 a_2582_4198# X1.X1.X1.X2.X2.X2.X3.vin2 vdd.t690 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2106 a_46502_6104# a_46116_6104# vss.t60 vss.t59 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2107 vdd.t1500 d0.t235 a_11072_6016# vdd.t1499 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2108 X2.X1.X1.X1.X1.X1.X1.vin2 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin1 vdd.t327 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2109 a_46116_9916# d0.t236 vdd.t1502 vdd.t1501 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2110 X2.X2.X3.vin1 a_48616_18540# X2.X2.X1.X3.vin2 vss.t638 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2111 vdd.t899 d1.t118 a_23512_5016# vdd.t898 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2112 vdd.t1378 d4.t12 a_8572_18358# vdd.t1377 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2113 X2.X1.X2.X2.X1.X2.X1.vin2 a_40352_23170# X2.X1.X2.X2.X1.X2.X3.vin1 vss.t1211 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2114 vdd.t1464 d0.t237 a_25712_30794# vdd.t1463 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2115 X2.X1.X2.X2.X2.X1.vout a_37766_27888# X2.X1.X2.X2.X2.X1.X3.vin1 vss.t906 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2116 X1.X1.X2.X1.X3.vin1 a_8186_6962# X1.X1.X2.X1.X1.X1.vout vss.t1279 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2117 X1.X2.X2.X2.X1.X1.vout a_23126_20264# X1.X2.X2.X2.X1.X1.X3.vin1 vss.t33 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2118 a_4782_9010# a_4396_9010# vss.t1263 vss.t1262 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2119 a_2196_13728# d0.t238 vss.t1478 vss.t1477 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2120 a_34062_16634# a_33676_16634# vss.t660 vss.t659 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2121 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X2.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X2122 vdd.t901 d1.t119 a_52792_27888# vdd.t900 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2123 X2.X2.X1.X1.X2.X1.X3.vin1 a_48702_24258# X2.X2.X1.X1.X2.X1.vout vss.t455 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2124 a_46116_6104# d0.t239 vdd.t1466 vdd.t1465 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2125 X2.X3.vin2 a_49566_892# X2.X2.X3.vin2.t3 vss.t1181 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2126 X1.X2.X2.X1.X1.X2.X1.vin2 a_25712_7922# X1.X2.X2.X1.X1.X2.X3.vin1 vss.t940 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2127 vss.t295 a_8872_5016# a_8486_5016# vss.t294 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2128 X2.X1.X1.X1.X2.X2.vout a_33676_20446# X2.X1.X1.X1.X2.X2.X3.vin1 vdd.t1192 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2129 X2.X2.X2.X1.X2.X1.X1.vin1 a_54992_11734# X2.X2.X2.X1.X2.X1.X3.vin1 vdd.t917 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2130 vss.t160 a_40352_6016# a_39966_6016# vss.t159 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2131 X2.X2.X1.X2.X2.X2.X3.vin2 a_46116_4198# X2.X2.X2.vrefh.t1 vss.t854 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2132 X2.X2.X1.X3.vin2 a_48616_10916# X2.X2.X1.X2.X3.vin2 vss.t1447 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2133 vss.t1251 a_52792_5016# a_52406_5016# vss.t1250 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2134 X1.X1.X2.X2.X2.X1.X2.vin1 a_11072_28888# X1.X1.X2.X2.X2.X1.X3.vin2 vdd.t315 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2135 a_16836_27070# d0.t240 vdd.t1468 vdd.t1467 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2136 X2.X3.vin1 a_43362_892# X3.vin2 vss.t1180 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2137 X1.X2.X1.X1.X1.X1.X2.vin1 a_17222_30882# X1.X2.X1.X1.X1.X1.X3.vin2 vss.t1173 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2138 X1.X2.X1.X1.X1.X1.vout a_19036_31882# X1.X2.X1.X1.X1.X1.X3.vin2 vss.t1105 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2139 a_4396_9010# d1.t120 vdd.t903 vdd.t902 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2140 vss.t814 a_54992_13640# a_54606_13640# vss.t813 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2141 a_5082_14688# a_4696_14688# vss.t270 vss.t269 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2142 X1.X1.X1.X2.X1.X1.vout a_4396_16634# X1.X1.X1.X2.X1.X1.X3.vin1 vdd.t1260 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2143 a_46116_15634# d0.t241 vss.t1480 vss.t1479 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2144 vss.t986 a_25712_17452# a_25326_17452# vss.t985 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2145 vdd.t1228 a_40352_13640# a_39966_13640# vdd.t1227 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2146 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X2.vrefh vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X2147 X1.X2.X1.X1.X1.X1.X3.vin1 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin1 vdd.t1451 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2148 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X1.X2.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X2149 a_2582_21352# a_2196_21352# vdd.t258 vdd.t257 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2150 vdd.t1522 a_11072_17452# a_10686_17452# vdd.t1521 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2151 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X2152 X2.X2.X2.X2.X1.X1.X3.vin1 a_54606_19358# X2.X2.X2.X2.X1.X1.X1.vin1 vss.t167 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2153 X1.X2.X2.X2.X1.X2.X3.vin1 a_25326_23170# X1.X2.X2.X2.X1.X2.X1.vin1 vss.t1313 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2154 a_33976_14688# d2.t60 vdd.t435 vdd.t434 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2155 X2.X2.X3.vin2.t1 a_52106_18358# X2.X2.X2.X3.vin1 vss.t685 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2156 X1.X2.X2.X1.X2.X1.X1.vin2 a_25712_11734# X1.X2.X2.X1.X2.X1.X3.vin1 vss.t1280 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2157 a_19036_16634# d1.t121 vss.t913 vss.t912 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2158 X2.X2.X1.X1.X3.vin2 a_48616_22312# X2.X2.X1.X1.X2.X1.vout vdd.t133 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2159 vss.t1482 d0.t242 a_54992_28888# vss.t1481 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2160 vdd.t1110 a_38152_27888# a_37766_27888# vdd.t1109 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2161 vss.t701 a_52492_25982# a_52106_25982# vss.t700 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2162 X1.X1.X2.X1.X3.vin1 a_8572_10734# X1.X1.X2.X3.vin1 vdd.t739 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2163 a_4396_31882# d1.t122 vss.t915 vss.t914 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2164 a_46116_28976# d0.t243 vdd.t1470 vdd.t1469 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2165 vss.t1484 d0.t244 a_40352_21264# vss.t1483 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2166 X2.X2.X1.X1.X1.X1.X1.vin1 a_46502_32788# X2.X2.X1.X1.X1.X1.X3.vin1 vss.t1241 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2167 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X2168 X1.X1.X2.X1.X2.X1.X3.vin1 a_8872_12640# X1.X1.X2.X1.X2.X1.vout vdd.t513 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2169 X2.X2.X1.X2.X1.X1.X1.vin2 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin1 vdd.t1383 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2170 a_2196_32788# d0.t245 vdd.t1472 vdd.t1471 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2171 X2.X1.X2.X1.X2.X1.X3.vin1 a_39966_11734# X2.X1.X2.X1.X2.X1.X1.vin2 vdd.t1225 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2172 a_4696_18540# d4.t13 vdd.t1380 vdd.t1379 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2173 vdd.t1460 d3.t28 a_23212_25982# vdd.t1459 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2174 vss.t917 d1.t123 a_38152_8828# vss.t916 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2175 vdd.t636 a_54992_21264# a_54606_21264# vdd.t635 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2176 vdd.t1449 a_25712_25076# a_25326_25076# vdd.t1448 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2177 X1.X1.X2.X1.X1.X2.vrefh a_11072_6016# X1.X1.X2.X1.X1.X1.X3.vin2 vss.t761 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2178 X1.X1.X1.X2.X2.X1.X3.vin1 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin2 vss.t1403 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2179 vdd.t444 a_23212_10734# a_22826_10734# vdd.t443 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2180 X2.X1.X1.X1.X1.X2.X3.vin2 a_34062_28070# X2.X1.X1.X1.X1.X2.vout vdd.t924 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2181 a_2582_27070# a_2196_27070# vss.t1051 vss.t1050 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2182 vdd.t519 a_23512_12640# a_23126_12640# vdd.t518 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2183 a_48316_5198# d1.t124 vdd.t905 vdd.t904 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2184 X2.X2.X1.X2.X2.X1.X1.vin2 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin1 vdd.t1406 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2185 vdd.t1474 d0.t246 a_40352_9828# vdd.t1473 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2186 a_4696_10916# d3.t29 vdd.t1462 vdd.t1461 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2187 X2.X2.X1.X1.X2.X2.X3.vin1 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin2 vss.t221 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2188 vss.t919 d1.t125 a_23512_20264# vss.t918 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2189 X2.X2.X1.X2.X2.X2.X1.vin1 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin1 vss.t723 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2190 a_17222_19446# a_16836_19446# vdd.t1525 vdd.t1524 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2191 a_20672_892# a_20286_892# vdd.t708 vdd.t707 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2192 a_49002_7064# a_48616_7064# vss.t1519 vss.t1518 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2193 a_31862_4198# a_31476_4198# vdd.t120 vdd.t119 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2194 X1.X2.X2.X1.X3.vin1 a_23212_10734# X1.X2.X2.X3.vin1 vdd.t442 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2195 a_17222_8010# a_16836_8010# vdd.t545 vdd.t544 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2196 X2.X1.X2.X1.X2.X1.X3.vin2 a_38152_12640# X2.X1.X2.X1.X2.X1.vout vss.t233 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2197 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X2.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X2198 X1.X2.X1.X1.X2.vrefh a_17222_27070# X1.X2.X1.X1.X1.X2.X3.vin2 vdd.t1507 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2199 a_31476_19446# d0.t247 vss.t1486 vss.t1485 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2200 X1.X2.X2.X1.X2.X1.X3.vin1 a_23512_12640# X1.X2.X2.X1.X2.X1.vout vdd.t517 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2201 X1.X2.X1.X1.X1.X2.vout a_19036_28070# X1.X2.X1.X1.X1.X2.X3.vin1 vdd.t933 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2202 vss.t1488 d0.t248 a_25712_7922# vss.t1487 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2203 a_49952_892# a_49566_892# vdd.t1152 vdd.t1151 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2204 vdd.t406 a_8572_18358# a_8186_18358# vdd.t405 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2205 X2.X2.X1.X2.X1.X1.X2.vin1 a_46502_15634# X2.X2.X1.X2.X1.X1.X3.vin2 vss.t252 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2206 a_33676_31882# d1.t126 vdd.t907 vdd.t906 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2207 vss.t924 a_11072_26982# a_10686_26982# vss.t923 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2208 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X2.vrefh vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X2209 a_48616_7064# d2.t61 vdd.t437 vdd.t436 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2210 X2.X1.X1.X2.X1.X2.X3.vin2 a_31476_11822# X2.X1.X1.X2.X1.X2.X2.vin1 vdd.t944 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2211 vss.t1490 d0.t249 a_54992_19358# vss.t1489 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2212 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X2213 a_46502_21352# a_46116_21352# vss.t220 vss.t219 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2214 vss.t1492 d0.t250 a_25712_23170# vss.t1491 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2215 X2.X2.X1.X1.X2.X1.vout a_48316_24258# X2.X2.X1.X1.X2.X1.X3.vin2 vss.t93 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2216 vss.t1394 d4.t14 a_52492_18358# vss.t1393 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2217 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X2.X1.vin1 vss.t77 sky130_fd_pr__res_high_po_0p35 l=1.09
X2218 a_17222_25164# a_16836_25164# vss.t837 vss.t836 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2219 X2.X1.X2.X1.X1.X1.vout a_37766_5016# X2.X1.X2.X1.X1.X1.X3.vin1 vss.t1178 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2220 vdd.t1476 d0.t251 a_11072_23170# vdd.t1475 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2221 a_4396_28070# d1.t127 vdd.t909 vdd.t908 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2222 X2.X2.X1.X1.X1.X2.X1.vin2 a_46502_28976# X2.X2.X1.X1.X1.X2.X3.vin1 vdd.t1259 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2223 vss.t449 d2.t62 a_37852_22210# vss.t448 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2224 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X2225 X1.X1.X2.X2.X2.X1.X3.vin2 a_10686_28888# X1.X1.X2.X2.X2.X2.vrefh vdd.t1271 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2226 X1.X2.X2.X1.X1.X1.X1.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 vss.t27 sky130_fd_pr__res_high_po_0p35 l=1.09
X2227 X2.X1.X2.X2.X1.X1.X3.vin1 a_38152_20264# X2.X1.X2.X2.X1.X1.vout vdd.t1166 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2228 vdd.t1445 a_54992_32700# a_54606_32700# vdd.t1444 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2229 vss.t122 a_54992_30794# a_54606_30794# vss.t121 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2230 X2.X1.X2.X2.vrefh a_40352_17452# X2.X1.X2.X1.X2.X2.X3.vin2 vss.t1125 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2231 a_48616_18540# d4.t15 vss.t1396 vss.t1395 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2232 X2.X1.X1.X2.X2.X2.X3.vin2 a_31476_4198# X2.X1.X2.vrefh.t0 vss.t129 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2233 X1.X2.X2.X2.X2.X2.X1.vin1 a_25712_30794# X1.X2.X2.X2.X2.X2.X3.vin1 vdd.t520 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2234 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 vss.t83 sky130_fd_pr__res_high_po_0p35 l=1.09
X2235 X1.X1.X1.X1.X1.X2.X3.vin1 a_4782_28070# X1.X1.X1.X1.X1.X2.vout vss.t1454 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2236 X2.X1.X1.X2.X1.X1.X3.vin1 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin2 vss.t1307 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2237 a_42976_892# d6.t3 vdd.t987 vdd.t986 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2238 X1.X1.X1.X1.X1.X2.vrefh a_2582_30882# X1.X1.X1.X1.X1.X1.X3.vin2 vdd.t1164 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2239 a_48702_24258# a_48316_24258# vss.t92 vss.t91 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2240 X1.X1.X2.vrefh.t0 X1.X1.X1.X2.X2.X2.X2.vin1 vss.t26 sky130_fd_pr__res_high_po_0p35 l=1.09
X2241 vss.t353 a_40352_21264# a_39966_21264# vss.t352 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2242 a_31862_19446# a_31476_19446# vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2243 X2.X2.X1.X1.X1.X1.X3.vin1 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin2 vss.t187 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2244 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 vss.t90 sky130_fd_pr__res_high_po_0p35 l=1.09
X2245 vss.t427 a_37852_18358# a_37466_18358# vss.t426 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2246 X1.X2.X2.X1.X3.vin1 a_22826_6962# X1.X2.X2.X1.X1.X2.vout vdd.t809 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2247 X2.X2.X1.X2.X1.X1.X3.vin1 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin1 vdd.t427 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2248 a_48616_10916# d3.t30 vss.t1474 vss.t1473 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2249 X2.X2.X2.X1.X3.vin2 a_52492_10734# X2.X2.X2.X3.vin1 vss.t1098 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2250 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 vss.t79 sky130_fd_pr__res_high_po_0p35 l=1.09
X2251 X2.X1.X2.X2.X1.X2.X2.vin1 a_40352_25076# X2.X1.X2.X2.X1.X2.X3.vin2 vdd.t699 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2252 vss.t781 a_8872_31700# a_8486_31700# vss.t780 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2253 X1.X2.X1.X2.X2.X1.vout a_19722_7064# X1.X2.X1.X2.X3.vin2 vss.t1061 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2254 X2.X2.X2.X1.X2.X1.X3.vin2 a_52792_12640# X2.X2.X2.X1.X2.X1.vout vss.t692 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2255 a_2582_15634# a_2196_15634# vdd.t1076 vdd.t1075 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2256 X2.X2.X2.X1.X2.X1.X3.vin2 a_54606_13640# X2.X2.X2.X1.X2.X1.X2.vin1 vss.t1311 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2257 X1.X1.X1.X1.X2.X2.X3.vin1 a_4782_20446# X1.X1.X1.X1.X2.X2.vout vss.t1470 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2258 X1.X1.X2.X2.X1.X1.X3.vin2 a_8872_20264# X1.X1.X2.X2.X1.X1.vout vss.t278 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2259 X1.X2.X2.X1.X2.X2.X3.vin2 a_25326_17452# X1.X2.X2.X1.X2.X2.X2.vin1 vss.t1008 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2260 X1.X2.X2.X1.X1.X2.X2.vin1 a_25712_9828# X1.X2.X2.X1.X1.X2.X3.vin2 vdd.t1264 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2261 X1.X2.X1.X1.X1.X1.X3.vin1 a_19422_31882# X1.X2.X1.X1.X1.X1.vout vss.t292 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2262 vss.t1494 d0.t252 a_40352_15546# vss.t1493 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2263 X2.X1.X2.X1.X1.X2.X3.vin1 a_38152_8828# X2.X1.X2.X1.X1.X2.vout vdd.t667 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2264 X2.X2.X1.X2.X2.X1.X3.vin1 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin1 vdd.t123 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2265 X1.X1.X2.X2.X3.vin1 a_8186_22210# X1.X1.X2.X2.X1.X1.vout vss.t315 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2266 a_2582_8010# a_2196_8010# vdd.t1161 vdd.t1160 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2267 X2.X2.X1.X2.X2.X1.vout a_49002_7064# X2.X2.X1.X2.X3.vin2 vss.t318 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2268 X1.X2.X1.X2.X2.X1.vout a_19036_9010# X1.X2.X1.X2.X2.X1.X3.vin2 vss.t182 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2269 a_48616_22312# d2.t63 vdd.t439 vdd.t438 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2270 X1.X2.X1.X3.vin2 a_19722_18540# X1.X2.X3.vin1.t0 vdd.t264 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2271 X2.X1.X1.X1.X3.vin2 a_34362_26164# X2.X1.X1.X3.vin1 vdd.t1422 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2272 a_31862_25164# a_31476_25164# vss.t1236 vss.t1235 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2273 vss.t671 a_23512_20264# a_23126_20264# vss.t670 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2274 a_46502_32788# a_46116_32788# vss.t186 vss.t185 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2275 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin1 vss.t76 sky130_fd_pr__res_high_po_0p35 l=1.09
X2276 a_19722_14688# a_19336_14688# vdd.t784 vdd.t783 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2277 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin1 vss.t25 sky130_fd_pr__res_high_po_0p35 l=1.09
X2278 a_16836_19446# d0.t253 vdd.t1478 vdd.t1477 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2279 vdd.t312 a_54992_15546# a_54606_15546# vdd.t311 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2280 a_46502_17540# a_46116_17540# vdd.t426 vdd.t425 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2281 vss.t1496 d0.t254 a_11072_32700# vss.t1495 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2282 vss.t1476 d3.t31 a_37852_25982# vss.t1475 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2283 vdd.t533 a_25712_19358# a_25326_19358# vdd.t532 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2284 a_19422_5198# a_19036_5198# vss.t690 vss.t689 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2285 X2.X2.X2.X2.X1.X1.X3.vin1 a_52792_20264# X2.X2.X2.X2.X1.X1.vout vdd.t1217 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2286 X2.X1.X2.X3.vin1 a_37466_10734# X2.X1.X2.X1.X3.vin1 vss.t465 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2287 X2.X2.X2.X2.X1.X1.X3.vin2 a_54606_21264# X2.X2.X2.X2.X1.X2.vrefh vdd.t110 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2288 vout.t0 a_28096_892# X3.vin2.t0 vss.t563 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2289 X2.X1.X2.X2.X2.X2.X3.vin1 a_38152_31700# X2.X1.X2.X2.X2.X2.vout vdd.t499 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2290 X1.X2.X2.X2.X1.X2.X3.vin2 a_25326_25076# X1.X2.X2.X2.X2.vrefh vdd.t743 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2291 X1.X2.X2.X3.vin1 a_22826_10734# X1.X2.X2.X1.X3.vin2 vdd.t892 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2292 X2.X2.X1.X2.X3.vin2 a_48616_7064# X2.X2.X1.X2.X2.X1.vout vdd.t1508 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2293 X2.X1.X2.X1.X2.X1.vout a_37766_12640# X2.X1.X2.X1.X2.X1.X3.vin1 vss.t89 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2294 X1.X1.X2.X1.X1.X2.vout a_8486_8828# X1.X1.X2.X1.X1.X2.X3.vin1 vss.t553 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2295 a_31476_23258# d0.t255 vdd.t1480 vdd.t1479 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
R0 vdd.n130 vdd.n129 1560
R1 vdd.n117 vdd.n109 1560
R2 vdd.n176 vdd.n175 1560
R3 vdd.n163 vdd.n155 1560
R4 vdd.n273 vdd.n272 1560
R5 vdd.n260 vdd.n252 1560
R6 vdd.n319 vdd.n318 1560
R7 vdd.n306 vdd.n298 1560
R8 vdd.n365 vdd.n364 1560
R9 vdd.n352 vdd.n344 1560
R10 vdd.n411 vdd.n410 1560
R11 vdd.n398 vdd.n390 1560
R12 vdd.n508 vdd.n507 1560
R13 vdd.n495 vdd.n487 1560
R14 vdd.n554 vdd.n553 1560
R15 vdd.n541 vdd.n533 1560
R16 vdd.n6701 vdd.n6700 1560
R17 vdd.n6716 vdd.n6715 1560
R18 vdd.n6747 vdd.n6746 1560
R19 vdd.n6762 vdd.n6761 1560
R20 vdd.n6845 vdd.n6844 1560
R21 vdd.n6860 vdd.n6859 1560
R22 vdd.n6891 vdd.n6890 1560
R23 vdd.n6906 vdd.n6905 1560
R24 vdd.n6937 vdd.n6936 1560
R25 vdd.n6952 vdd.n6951 1560
R26 vdd.n6983 vdd.n6982 1560
R27 vdd.n6998 vdd.n6997 1560
R28 vdd.n7081 vdd.n7080 1560
R29 vdd.n7096 vdd.n7095 1560
R30 vdd.n8539 vdd.n8538 1560
R31 vdd.n8554 vdd.n8553 1560
R32 vdd.n7146 vdd.n7145 1560
R33 vdd.n7133 vdd.n7125 1560
R34 vdd.n7192 vdd.n7191 1560
R35 vdd.n7179 vdd.n7171 1560
R36 vdd.n7289 vdd.n7288 1560
R37 vdd.n7276 vdd.n7268 1560
R38 vdd.n7335 vdd.n7334 1560
R39 vdd.n7322 vdd.n7314 1560
R40 vdd.n7381 vdd.n7380 1560
R41 vdd.n7368 vdd.n7360 1560
R42 vdd.n7427 vdd.n7426 1560
R43 vdd.n7414 vdd.n7406 1560
R44 vdd.n7524 vdd.n7523 1560
R45 vdd.n7511 vdd.n7503 1560
R46 vdd.n6673 vdd.n6672 1560
R47 vdd.n6660 vdd.n6652 1560
R48 vdd.n7568 vdd.n7567 1560
R49 vdd.n7555 vdd.n7547 1560
R50 vdd.n7613 vdd.n7612 1560
R51 vdd.n7600 vdd.n7592 1560
R52 vdd.n7663 vdd.n7662 1560
R53 vdd.n7650 vdd.n7642 1560
R54 vdd.n7709 vdd.n7708 1560
R55 vdd.n7696 vdd.n7688 1560
R56 vdd.n7757 vdd.n7756 1560
R57 vdd.n7744 vdd.n7736 1560
R58 vdd.n7469 vdd.n7468 1560
R59 vdd.n7481 vdd.n7440 1560
R60 vdd.n7804 vdd.n7803 1560
R61 vdd.n7791 vdd.n7783 1560
R62 vdd.n7849 vdd.n7848 1560
R63 vdd.n7836 vdd.n7828 1560
R64 vdd.n7895 vdd.n7894 1560
R65 vdd.n7882 vdd.n7874 1560
R66 vdd.n7946 vdd.n7945 1560
R67 vdd.n7933 vdd.n7925 1560
R68 vdd.n7992 vdd.n7991 1560
R69 vdd.n7979 vdd.n7971 1560
R70 vdd.n8040 vdd.n8039 1560
R71 vdd.n8027 vdd.n8019 1560
R72 vdd.n8086 vdd.n8085 1560
R73 vdd.n8073 vdd.n8065 1560
R74 vdd.n8131 vdd.n8130 1560
R75 vdd.n8118 vdd.n8110 1560
R76 vdd.n8181 vdd.n8180 1560
R77 vdd.n8168 vdd.n8160 1560
R78 vdd.n8227 vdd.n8226 1560
R79 vdd.n8214 vdd.n8206 1560
R80 vdd.n8275 vdd.n8274 1560
R81 vdd.n8262 vdd.n8254 1560
R82 vdd.n7234 vdd.n7233 1560
R83 vdd.n7246 vdd.n7205 1560
R84 vdd.n8322 vdd.n8321 1560
R85 vdd.n8309 vdd.n8301 1560
R86 vdd.n8367 vdd.n8366 1560
R87 vdd.n8354 vdd.n8346 1560
R88 vdd.n8417 vdd.n8416 1560
R89 vdd.n8404 vdd.n8396 1560
R90 vdd.n8463 vdd.n8462 1560
R91 vdd.n8450 vdd.n8442 1560
R92 vdd.n8511 vdd.n8510 1560
R93 vdd.n8498 vdd.n8490 1560
R94 vdd.n8632 vdd.n8631 1560
R95 vdd.n8647 vdd.n8646 1560
R96 vdd.n8586 vdd.n8585 1560
R97 vdd.n8601 vdd.n8600 1560
R98 vdd.n8679 vdd.n8678 1560
R99 vdd.n8694 vdd.n8693 1560
R100 vdd.n8727 vdd.n8726 1560
R101 vdd.n8742 vdd.n8741 1560
R102 vdd.n8773 vdd.n8772 1560
R103 vdd.n8788 vdd.n8787 1560
R104 vdd.n7035 vdd.n7029 1560
R105 vdd.n7053 vdd.n7014 1560
R106 vdd.n8915 vdd.n8914 1560
R107 vdd.n8930 vdd.n8929 1560
R108 vdd.n8868 vdd.n8867 1560
R109 vdd.n8883 vdd.n8882 1560
R110 vdd.n8822 vdd.n8821 1560
R111 vdd.n8837 vdd.n8836 1560
R112 vdd.n8962 vdd.n8961 1560
R113 vdd.n8977 vdd.n8976 1560
R114 vdd.n9010 vdd.n9009 1560
R115 vdd.n9025 vdd.n9024 1560
R116 vdd.n9056 vdd.n9055 1560
R117 vdd.n9071 vdd.n9070 1560
R118 vdd.n9150 vdd.n9149 1560
R119 vdd.n9165 vdd.n9164 1560
R120 vdd.n9104 vdd.n9103 1560
R121 vdd.n9119 vdd.n9118 1560
R122 vdd.n9197 vdd.n9196 1560
R123 vdd.n9212 vdd.n9211 1560
R124 vdd.n9245 vdd.n9244 1560
R125 vdd.n9260 vdd.n9259 1560
R126 vdd.n9291 vdd.n9290 1560
R127 vdd.n9306 vdd.n9305 1560
R128 vdd.n6799 vdd.n6793 1560
R129 vdd.n6817 vdd.n6778 1560
R130 vdd.n9386 vdd.n9385 1560
R131 vdd.n9401 vdd.n9400 1560
R132 vdd.n9340 vdd.n9339 1560
R133 vdd.n9355 vdd.n9354 1560
R134 vdd.n9433 vdd.n9432 1560
R135 vdd.n9448 vdd.n9447 1560
R136 vdd.n9481 vdd.n9480 1560
R137 vdd.n9496 vdd.n9495 1560
R138 vdd.n9527 vdd.n9526 1560
R139 vdd.n9542 vdd.n9541 1560
R140 vdd.n3687 vdd.n3686 1560
R141 vdd.n3702 vdd.n3701 1560
R142 vdd.n3733 vdd.n3732 1560
R143 vdd.n3748 vdd.n3747 1560
R144 vdd.n3831 vdd.n3830 1560
R145 vdd.n3846 vdd.n3845 1560
R146 vdd.n3877 vdd.n3876 1560
R147 vdd.n3892 vdd.n3891 1560
R148 vdd.n3923 vdd.n3922 1560
R149 vdd.n3938 vdd.n3937 1560
R150 vdd.n3969 vdd.n3968 1560
R151 vdd.n3984 vdd.n3983 1560
R152 vdd.n4067 vdd.n4066 1560
R153 vdd.n4082 vdd.n4081 1560
R154 vdd.n5525 vdd.n5524 1560
R155 vdd.n5540 vdd.n5539 1560
R156 vdd.n4132 vdd.n4131 1560
R157 vdd.n4119 vdd.n4111 1560
R158 vdd.n4178 vdd.n4177 1560
R159 vdd.n4165 vdd.n4157 1560
R160 vdd.n4275 vdd.n4274 1560
R161 vdd.n4262 vdd.n4254 1560
R162 vdd.n4321 vdd.n4320 1560
R163 vdd.n4308 vdd.n4300 1560
R164 vdd.n4367 vdd.n4366 1560
R165 vdd.n4354 vdd.n4346 1560
R166 vdd.n4413 vdd.n4412 1560
R167 vdd.n4400 vdd.n4392 1560
R168 vdd.n4510 vdd.n4509 1560
R169 vdd.n4497 vdd.n4489 1560
R170 vdd.n3659 vdd.n3658 1560
R171 vdd.n3646 vdd.n3638 1560
R172 vdd.n4554 vdd.n4553 1560
R173 vdd.n4541 vdd.n4533 1560
R174 vdd.n4599 vdd.n4598 1560
R175 vdd.n4586 vdd.n4578 1560
R176 vdd.n4649 vdd.n4648 1560
R177 vdd.n4636 vdd.n4628 1560
R178 vdd.n4695 vdd.n4694 1560
R179 vdd.n4682 vdd.n4674 1560
R180 vdd.n4743 vdd.n4742 1560
R181 vdd.n4730 vdd.n4722 1560
R182 vdd.n4455 vdd.n4454 1560
R183 vdd.n4467 vdd.n4426 1560
R184 vdd.n4790 vdd.n4789 1560
R185 vdd.n4777 vdd.n4769 1560
R186 vdd.n4835 vdd.n4834 1560
R187 vdd.n4822 vdd.n4814 1560
R188 vdd.n4881 vdd.n4880 1560
R189 vdd.n4868 vdd.n4860 1560
R190 vdd.n4932 vdd.n4931 1560
R191 vdd.n4919 vdd.n4911 1560
R192 vdd.n4978 vdd.n4977 1560
R193 vdd.n4965 vdd.n4957 1560
R194 vdd.n5026 vdd.n5025 1560
R195 vdd.n5013 vdd.n5005 1560
R196 vdd.n5072 vdd.n5071 1560
R197 vdd.n5059 vdd.n5051 1560
R198 vdd.n5117 vdd.n5116 1560
R199 vdd.n5104 vdd.n5096 1560
R200 vdd.n5167 vdd.n5166 1560
R201 vdd.n5154 vdd.n5146 1560
R202 vdd.n5213 vdd.n5212 1560
R203 vdd.n5200 vdd.n5192 1560
R204 vdd.n5261 vdd.n5260 1560
R205 vdd.n5248 vdd.n5240 1560
R206 vdd.n4220 vdd.n4219 1560
R207 vdd.n4232 vdd.n4191 1560
R208 vdd.n5308 vdd.n5307 1560
R209 vdd.n5295 vdd.n5287 1560
R210 vdd.n5353 vdd.n5352 1560
R211 vdd.n5340 vdd.n5332 1560
R212 vdd.n5403 vdd.n5402 1560
R213 vdd.n5390 vdd.n5382 1560
R214 vdd.n5449 vdd.n5448 1560
R215 vdd.n5436 vdd.n5428 1560
R216 vdd.n5497 vdd.n5496 1560
R217 vdd.n5484 vdd.n5476 1560
R218 vdd.n5618 vdd.n5617 1560
R219 vdd.n5633 vdd.n5632 1560
R220 vdd.n5572 vdd.n5571 1560
R221 vdd.n5587 vdd.n5586 1560
R222 vdd.n5665 vdd.n5664 1560
R223 vdd.n5680 vdd.n5679 1560
R224 vdd.n5713 vdd.n5712 1560
R225 vdd.n5728 vdd.n5727 1560
R226 vdd.n5759 vdd.n5758 1560
R227 vdd.n5774 vdd.n5773 1560
R228 vdd.n4021 vdd.n4015 1560
R229 vdd.n4039 vdd.n4000 1560
R230 vdd.n5901 vdd.n5900 1560
R231 vdd.n5916 vdd.n5915 1560
R232 vdd.n5854 vdd.n5853 1560
R233 vdd.n5869 vdd.n5868 1560
R234 vdd.n5808 vdd.n5807 1560
R235 vdd.n5823 vdd.n5822 1560
R236 vdd.n5948 vdd.n5947 1560
R237 vdd.n5963 vdd.n5962 1560
R238 vdd.n5996 vdd.n5995 1560
R239 vdd.n6011 vdd.n6010 1560
R240 vdd.n6042 vdd.n6041 1560
R241 vdd.n6057 vdd.n6056 1560
R242 vdd.n6136 vdd.n6135 1560
R243 vdd.n6151 vdd.n6150 1560
R244 vdd.n6090 vdd.n6089 1560
R245 vdd.n6105 vdd.n6104 1560
R246 vdd.n6183 vdd.n6182 1560
R247 vdd.n6198 vdd.n6197 1560
R248 vdd.n6231 vdd.n6230 1560
R249 vdd.n6246 vdd.n6245 1560
R250 vdd.n6277 vdd.n6276 1560
R251 vdd.n6292 vdd.n6291 1560
R252 vdd.n3785 vdd.n3779 1560
R253 vdd.n3803 vdd.n3764 1560
R254 vdd.n6372 vdd.n6371 1560
R255 vdd.n6387 vdd.n6386 1560
R256 vdd.n6326 vdd.n6325 1560
R257 vdd.n6341 vdd.n6340 1560
R258 vdd.n6419 vdd.n6418 1560
R259 vdd.n6434 vdd.n6433 1560
R260 vdd.n6467 vdd.n6466 1560
R261 vdd.n6482 vdd.n6481 1560
R262 vdd.n6513 vdd.n6512 1560
R263 vdd.n6528 vdd.n6527 1560
R264 vdd.n673 vdd.n672 1560
R265 vdd.n688 vdd.n687 1560
R266 vdd.n719 vdd.n718 1560
R267 vdd.n734 vdd.n733 1560
R268 vdd.n817 vdd.n816 1560
R269 vdd.n832 vdd.n831 1560
R270 vdd.n863 vdd.n862 1560
R271 vdd.n878 vdd.n877 1560
R272 vdd.n909 vdd.n908 1560
R273 vdd.n924 vdd.n923 1560
R274 vdd.n955 vdd.n954 1560
R275 vdd.n970 vdd.n969 1560
R276 vdd.n1053 vdd.n1052 1560
R277 vdd.n1068 vdd.n1067 1560
R278 vdd.n2511 vdd.n2510 1560
R279 vdd.n2526 vdd.n2525 1560
R280 vdd.n1118 vdd.n1117 1560
R281 vdd.n1105 vdd.n1097 1560
R282 vdd.n1164 vdd.n1163 1560
R283 vdd.n1151 vdd.n1143 1560
R284 vdd.n1261 vdd.n1260 1560
R285 vdd.n1248 vdd.n1240 1560
R286 vdd.n1307 vdd.n1306 1560
R287 vdd.n1294 vdd.n1286 1560
R288 vdd.n1353 vdd.n1352 1560
R289 vdd.n1340 vdd.n1332 1560
R290 vdd.n1399 vdd.n1398 1560
R291 vdd.n1386 vdd.n1378 1560
R292 vdd.n1496 vdd.n1495 1560
R293 vdd.n1483 vdd.n1475 1560
R294 vdd.n645 vdd.n644 1560
R295 vdd.n632 vdd.n624 1560
R296 vdd.n1540 vdd.n1539 1560
R297 vdd.n1527 vdd.n1519 1560
R298 vdd.n1585 vdd.n1584 1560
R299 vdd.n1572 vdd.n1564 1560
R300 vdd.n1635 vdd.n1634 1560
R301 vdd.n1622 vdd.n1614 1560
R302 vdd.n1681 vdd.n1680 1560
R303 vdd.n1668 vdd.n1660 1560
R304 vdd.n1729 vdd.n1728 1560
R305 vdd.n1716 vdd.n1708 1560
R306 vdd.n1441 vdd.n1440 1560
R307 vdd.n1453 vdd.n1412 1560
R308 vdd.n1776 vdd.n1775 1560
R309 vdd.n1763 vdd.n1755 1560
R310 vdd.n1821 vdd.n1820 1560
R311 vdd.n1808 vdd.n1800 1560
R312 vdd.n1867 vdd.n1866 1560
R313 vdd.n1854 vdd.n1846 1560
R314 vdd.n1918 vdd.n1917 1560
R315 vdd.n1905 vdd.n1897 1560
R316 vdd.n1964 vdd.n1963 1560
R317 vdd.n1951 vdd.n1943 1560
R318 vdd.n2012 vdd.n2011 1560
R319 vdd.n1999 vdd.n1991 1560
R320 vdd.n2058 vdd.n2057 1560
R321 vdd.n2045 vdd.n2037 1560
R322 vdd.n2103 vdd.n2102 1560
R323 vdd.n2090 vdd.n2082 1560
R324 vdd.n2153 vdd.n2152 1560
R325 vdd.n2140 vdd.n2132 1560
R326 vdd.n2199 vdd.n2198 1560
R327 vdd.n2186 vdd.n2178 1560
R328 vdd.n2247 vdd.n2246 1560
R329 vdd.n2234 vdd.n2226 1560
R330 vdd.n1206 vdd.n1205 1560
R331 vdd.n1218 vdd.n1177 1560
R332 vdd.n2294 vdd.n2293 1560
R333 vdd.n2281 vdd.n2273 1560
R334 vdd.n2339 vdd.n2338 1560
R335 vdd.n2326 vdd.n2318 1560
R336 vdd.n2389 vdd.n2388 1560
R337 vdd.n2376 vdd.n2368 1560
R338 vdd.n2435 vdd.n2434 1560
R339 vdd.n2422 vdd.n2414 1560
R340 vdd.n2483 vdd.n2482 1560
R341 vdd.n2470 vdd.n2462 1560
R342 vdd.n2604 vdd.n2603 1560
R343 vdd.n2619 vdd.n2618 1560
R344 vdd.n2558 vdd.n2557 1560
R345 vdd.n2573 vdd.n2572 1560
R346 vdd.n2651 vdd.n2650 1560
R347 vdd.n2666 vdd.n2665 1560
R348 vdd.n2699 vdd.n2698 1560
R349 vdd.n2714 vdd.n2713 1560
R350 vdd.n2745 vdd.n2744 1560
R351 vdd.n2760 vdd.n2759 1560
R352 vdd.n1007 vdd.n1001 1560
R353 vdd.n1025 vdd.n986 1560
R354 vdd.n2887 vdd.n2886 1560
R355 vdd.n2902 vdd.n2901 1560
R356 vdd.n2840 vdd.n2839 1560
R357 vdd.n2855 vdd.n2854 1560
R358 vdd.n2794 vdd.n2793 1560
R359 vdd.n2809 vdd.n2808 1560
R360 vdd.n2934 vdd.n2933 1560
R361 vdd.n2949 vdd.n2948 1560
R362 vdd.n2982 vdd.n2981 1560
R363 vdd.n2997 vdd.n2996 1560
R364 vdd.n3028 vdd.n3027 1560
R365 vdd.n3043 vdd.n3042 1560
R366 vdd.n3122 vdd.n3121 1560
R367 vdd.n3137 vdd.n3136 1560
R368 vdd.n3076 vdd.n3075 1560
R369 vdd.n3091 vdd.n3090 1560
R370 vdd.n3169 vdd.n3168 1560
R371 vdd.n3184 vdd.n3183 1560
R372 vdd.n3217 vdd.n3216 1560
R373 vdd.n3232 vdd.n3231 1560
R374 vdd.n3263 vdd.n3262 1560
R375 vdd.n3278 vdd.n3277 1560
R376 vdd.n771 vdd.n765 1560
R377 vdd.n789 vdd.n750 1560
R378 vdd.n3358 vdd.n3357 1560
R379 vdd.n3373 vdd.n3372 1560
R380 vdd.n3312 vdd.n3311 1560
R381 vdd.n3327 vdd.n3326 1560
R382 vdd.n3405 vdd.n3404 1560
R383 vdd.n3420 vdd.n3419 1560
R384 vdd.n3453 vdd.n3452 1560
R385 vdd.n3468 vdd.n3467 1560
R386 vdd.n3499 vdd.n3498 1560
R387 vdd.n3514 vdd.n3513 1560
R388 vdd.n581 vdd.n580 1560
R389 vdd.n596 vdd.n595 1560
R390 vdd.n3594 vdd.n3593 1560
R391 vdd.n3609 vdd.n3608 1560
R392 vdd.n3548 vdd.n3547 1560
R393 vdd.n3563 vdd.n3562 1560
R394 vdd.n6608 vdd.n6607 1560
R395 vdd.n6623 vdd.n6622 1560
R396 vdd.n6562 vdd.n6561 1560
R397 vdd.n6577 vdd.n6576 1560
R398 vdd.n9622 vdd.n9621 1560
R399 vdd.n9637 vdd.n9636 1560
R400 vdd.n9576 vdd.n9575 1560
R401 vdd.n9591 vdd.n9590 1560
R402 vdd.n9668 vdd.n9667 1560
R403 vdd.n9683 vdd.n9682 1560
R404 vdd.n9714 vdd.n9713 1560
R405 vdd.n9729 vdd.n9728 1560
R406 vdd.n9812 vdd.n9811 1560
R407 vdd.n9827 vdd.n9826 1560
R408 vdd.n9858 vdd.n9857 1560
R409 vdd.n9873 vdd.n9872 1560
R410 vdd.n9904 vdd.n9903 1560
R411 vdd.n9919 vdd.n9918 1560
R412 vdd.n9950 vdd.n9949 1560
R413 vdd.n9965 vdd.n9964 1560
R414 vdd.n10048 vdd.n10047 1560
R415 vdd.n10063 vdd.n10062 1560
R416 vdd.n64 vdd.n63 1560
R417 vdd.n79 vdd.n78 1560
R418 vdd.n18 vdd.n17 1560
R419 vdd.n33 vdd.n32 1560
R420 vdd.n10094 vdd.n10093 1560
R421 vdd.n10109 vdd.n10108 1560
R422 vdd.n10142 vdd.n10141 1560
R423 vdd.n10157 vdd.n10156 1560
R424 vdd.n10188 vdd.n10187 1560
R425 vdd.n10203 vdd.n10202 1560
R426 vdd.n10002 vdd.n9996 1560
R427 vdd.n10020 vdd.n9981 1560
R428 vdd.n10330 vdd.n10329 1560
R429 vdd.n10345 vdd.n10344 1560
R430 vdd.n10283 vdd.n10282 1560
R431 vdd.n10298 vdd.n10297 1560
R432 vdd.n10237 vdd.n10236 1560
R433 vdd.n10252 vdd.n10251 1560
R434 vdd.n10377 vdd.n10376 1560
R435 vdd.n10392 vdd.n10391 1560
R436 vdd.n10425 vdd.n10424 1560
R437 vdd.n10440 vdd.n10439 1560
R438 vdd.n10471 vdd.n10470 1560
R439 vdd.n10486 vdd.n10485 1560
R440 vdd.n10565 vdd.n10564 1560
R441 vdd.n10580 vdd.n10579 1560
R442 vdd.n10519 vdd.n10518 1560
R443 vdd.n10534 vdd.n10533 1560
R444 vdd.n10612 vdd.n10611 1560
R445 vdd.n10627 vdd.n10626 1560
R446 vdd.n10660 vdd.n10659 1560
R447 vdd.n10675 vdd.n10674 1560
R448 vdd.n10706 vdd.n10705 1560
R449 vdd.n10721 vdd.n10720 1560
R450 vdd.n9766 vdd.n9760 1560
R451 vdd.n9784 vdd.n9745 1560
R452 vdd.n10801 vdd.n10800 1560
R453 vdd.n10816 vdd.n10815 1560
R454 vdd.n10755 vdd.n10754 1560
R455 vdd.n10770 vdd.n10769 1560
R456 vdd.n10848 vdd.n10847 1560
R457 vdd.n10863 vdd.n10862 1560
R458 vdd.n10896 vdd.n10895 1560
R459 vdd.n10911 vdd.n10910 1560
R460 vdd.n10942 vdd.n10941 1560
R461 vdd.n10957 vdd.n10956 1560
R462 vdd.n11008 vdd.n11007 1560
R463 vdd.n10995 vdd.n10987 1560
R464 vdd.n11053 vdd.n11052 1560
R465 vdd.n11040 vdd.n11032 1560
R466 vdd.n11103 vdd.n11102 1560
R467 vdd.n11090 vdd.n11082 1560
R468 vdd.n11149 vdd.n11148 1560
R469 vdd.n11136 vdd.n11128 1560
R470 vdd.n11197 vdd.n11196 1560
R471 vdd.n11184 vdd.n11176 1560
R472 vdd.n453 vdd.n452 1560
R473 vdd.n465 vdd.n424 1560
R474 vdd.n11244 vdd.n11243 1560
R475 vdd.n11231 vdd.n11223 1560
R476 vdd.n11289 vdd.n11288 1560
R477 vdd.n11276 vdd.n11268 1560
R478 vdd.n11335 vdd.n11334 1560
R479 vdd.n11322 vdd.n11314 1560
R480 vdd.n11386 vdd.n11385 1560
R481 vdd.n11373 vdd.n11365 1560
R482 vdd.n11432 vdd.n11431 1560
R483 vdd.n11419 vdd.n11411 1560
R484 vdd.n11480 vdd.n11479 1560
R485 vdd.n11467 vdd.n11459 1560
R486 vdd.n11526 vdd.n11525 1560
R487 vdd.n11513 vdd.n11505 1560
R488 vdd.n11571 vdd.n11570 1560
R489 vdd.n11558 vdd.n11550 1560
R490 vdd.n11621 vdd.n11620 1560
R491 vdd.n11608 vdd.n11600 1560
R492 vdd.n11667 vdd.n11666 1560
R493 vdd.n11654 vdd.n11646 1560
R494 vdd.n11715 vdd.n11714 1560
R495 vdd.n11702 vdd.n11694 1560
R496 vdd.n218 vdd.n217 1560
R497 vdd.n230 vdd.n189 1560
R498 vdd.n11762 vdd.n11761 1560
R499 vdd.n11749 vdd.n11741 1560
R500 vdd.n11807 vdd.n11806 1560
R501 vdd.n11794 vdd.n11786 1560
R502 vdd.n11857 vdd.n11856 1560
R503 vdd.n11844 vdd.n11836 1560
R504 vdd.n11903 vdd.n11902 1560
R505 vdd.n11890 vdd.n11882 1560
R506 vdd.n11951 vdd.n11950 1560
R507 vdd.n11938 vdd.n11930 1560
R508 vdd.n127 vdd.n99 878.823
R509 vdd.n134 vdd.n99 878.823
R510 vdd.n106 vdd.n102 878.823
R511 vdd.n106 vdd.n98 878.823
R512 vdd.n108 vdd.n104 878.823
R513 vdd.n118 vdd.n108 878.823
R514 vdd.n173 vdd.n145 878.823
R515 vdd.n180 vdd.n145 878.823
R516 vdd.n152 vdd.n148 878.823
R517 vdd.n152 vdd.n144 878.823
R518 vdd.n154 vdd.n150 878.823
R519 vdd.n164 vdd.n154 878.823
R520 vdd.n270 vdd.n242 878.823
R521 vdd.n277 vdd.n242 878.823
R522 vdd.n249 vdd.n245 878.823
R523 vdd.n249 vdd.n241 878.823
R524 vdd.n251 vdd.n247 878.823
R525 vdd.n261 vdd.n251 878.823
R526 vdd.n316 vdd.n288 878.823
R527 vdd.n323 vdd.n288 878.823
R528 vdd.n295 vdd.n291 878.823
R529 vdd.n295 vdd.n287 878.823
R530 vdd.n297 vdd.n293 878.823
R531 vdd.n307 vdd.n297 878.823
R532 vdd.n362 vdd.n334 878.823
R533 vdd.n369 vdd.n334 878.823
R534 vdd.n341 vdd.n337 878.823
R535 vdd.n341 vdd.n333 878.823
R536 vdd.n343 vdd.n339 878.823
R537 vdd.n353 vdd.n343 878.823
R538 vdd.n408 vdd.n380 878.823
R539 vdd.n415 vdd.n380 878.823
R540 vdd.n387 vdd.n383 878.823
R541 vdd.n387 vdd.n379 878.823
R542 vdd.n389 vdd.n385 878.823
R543 vdd.n399 vdd.n389 878.823
R544 vdd.n505 vdd.n477 878.823
R545 vdd.n512 vdd.n477 878.823
R546 vdd.n484 vdd.n480 878.823
R547 vdd.n484 vdd.n476 878.823
R548 vdd.n486 vdd.n482 878.823
R549 vdd.n496 vdd.n486 878.823
R550 vdd.n551 vdd.n523 878.823
R551 vdd.n558 vdd.n523 878.823
R552 vdd.n530 vdd.n526 878.823
R553 vdd.n530 vdd.n522 878.823
R554 vdd.n532 vdd.n528 878.823
R555 vdd.n542 vdd.n532 878.823
R556 vdd.n6694 vdd.n6686 878.823
R557 vdd.n6695 vdd.n6694 878.823
R558 vdd.n6707 vdd.n6697 878.823
R559 vdd.n6697 vdd.n6693 878.823
R560 vdd.n6721 vdd.n6687 878.823
R561 vdd.n6721 vdd.n6720 878.823
R562 vdd.n6740 vdd.n6732 878.823
R563 vdd.n6741 vdd.n6740 878.823
R564 vdd.n6753 vdd.n6743 878.823
R565 vdd.n6743 vdd.n6739 878.823
R566 vdd.n6767 vdd.n6733 878.823
R567 vdd.n6767 vdd.n6766 878.823
R568 vdd.n6838 vdd.n6830 878.823
R569 vdd.n6839 vdd.n6838 878.823
R570 vdd.n6851 vdd.n6841 878.823
R571 vdd.n6841 vdd.n6837 878.823
R572 vdd.n6865 vdd.n6831 878.823
R573 vdd.n6865 vdd.n6864 878.823
R574 vdd.n6884 vdd.n6876 878.823
R575 vdd.n6885 vdd.n6884 878.823
R576 vdd.n6897 vdd.n6887 878.823
R577 vdd.n6887 vdd.n6883 878.823
R578 vdd.n6911 vdd.n6877 878.823
R579 vdd.n6911 vdd.n6910 878.823
R580 vdd.n6930 vdd.n6922 878.823
R581 vdd.n6931 vdd.n6930 878.823
R582 vdd.n6943 vdd.n6933 878.823
R583 vdd.n6933 vdd.n6929 878.823
R584 vdd.n6957 vdd.n6923 878.823
R585 vdd.n6957 vdd.n6956 878.823
R586 vdd.n6976 vdd.n6968 878.823
R587 vdd.n6977 vdd.n6976 878.823
R588 vdd.n6989 vdd.n6979 878.823
R589 vdd.n6979 vdd.n6975 878.823
R590 vdd.n7003 vdd.n6969 878.823
R591 vdd.n7003 vdd.n7002 878.823
R592 vdd.n7074 vdd.n7066 878.823
R593 vdd.n7075 vdd.n7074 878.823
R594 vdd.n7087 vdd.n7077 878.823
R595 vdd.n7077 vdd.n7073 878.823
R596 vdd.n7101 vdd.n7067 878.823
R597 vdd.n7101 vdd.n7100 878.823
R598 vdd.n8532 vdd.n8524 878.823
R599 vdd.n8533 vdd.n8532 878.823
R600 vdd.n8545 vdd.n8535 878.823
R601 vdd.n8535 vdd.n8531 878.823
R602 vdd.n8559 vdd.n8525 878.823
R603 vdd.n8559 vdd.n8558 878.823
R604 vdd.n7143 vdd.n7115 878.823
R605 vdd.n7150 vdd.n7115 878.823
R606 vdd.n7122 vdd.n7118 878.823
R607 vdd.n7122 vdd.n7114 878.823
R608 vdd.n7124 vdd.n7120 878.823
R609 vdd.n7134 vdd.n7124 878.823
R610 vdd.n7189 vdd.n7161 878.823
R611 vdd.n7196 vdd.n7161 878.823
R612 vdd.n7168 vdd.n7164 878.823
R613 vdd.n7168 vdd.n7160 878.823
R614 vdd.n7170 vdd.n7166 878.823
R615 vdd.n7180 vdd.n7170 878.823
R616 vdd.n7286 vdd.n7258 878.823
R617 vdd.n7293 vdd.n7258 878.823
R618 vdd.n7265 vdd.n7261 878.823
R619 vdd.n7265 vdd.n7257 878.823
R620 vdd.n7267 vdd.n7263 878.823
R621 vdd.n7277 vdd.n7267 878.823
R622 vdd.n7332 vdd.n7304 878.823
R623 vdd.n7339 vdd.n7304 878.823
R624 vdd.n7311 vdd.n7307 878.823
R625 vdd.n7311 vdd.n7303 878.823
R626 vdd.n7313 vdd.n7309 878.823
R627 vdd.n7323 vdd.n7313 878.823
R628 vdd.n7378 vdd.n7350 878.823
R629 vdd.n7385 vdd.n7350 878.823
R630 vdd.n7357 vdd.n7353 878.823
R631 vdd.n7357 vdd.n7349 878.823
R632 vdd.n7359 vdd.n7355 878.823
R633 vdd.n7369 vdd.n7359 878.823
R634 vdd.n7424 vdd.n7396 878.823
R635 vdd.n7431 vdd.n7396 878.823
R636 vdd.n7403 vdd.n7399 878.823
R637 vdd.n7403 vdd.n7395 878.823
R638 vdd.n7405 vdd.n7401 878.823
R639 vdd.n7415 vdd.n7405 878.823
R640 vdd.n7521 vdd.n7493 878.823
R641 vdd.n7528 vdd.n7493 878.823
R642 vdd.n7500 vdd.n7496 878.823
R643 vdd.n7500 vdd.n7492 878.823
R644 vdd.n7502 vdd.n7498 878.823
R645 vdd.n7512 vdd.n7502 878.823
R646 vdd.n6670 vdd.n6642 878.823
R647 vdd.n6677 vdd.n6642 878.823
R648 vdd.n6649 vdd.n6645 878.823
R649 vdd.n6649 vdd.n6641 878.823
R650 vdd.n6651 vdd.n6647 878.823
R651 vdd.n6661 vdd.n6651 878.823
R652 vdd.n7565 vdd.n7537 878.823
R653 vdd.n7572 vdd.n7537 878.823
R654 vdd.n7544 vdd.n7540 878.823
R655 vdd.n7544 vdd.n7536 878.823
R656 vdd.n7546 vdd.n7542 878.823
R657 vdd.n7556 vdd.n7546 878.823
R658 vdd.n7610 vdd.n7582 878.823
R659 vdd.n7617 vdd.n7582 878.823
R660 vdd.n7589 vdd.n7585 878.823
R661 vdd.n7589 vdd.n7581 878.823
R662 vdd.n7591 vdd.n7587 878.823
R663 vdd.n7601 vdd.n7591 878.823
R664 vdd.n7660 vdd.n7632 878.823
R665 vdd.n7667 vdd.n7632 878.823
R666 vdd.n7639 vdd.n7635 878.823
R667 vdd.n7639 vdd.n7631 878.823
R668 vdd.n7641 vdd.n7637 878.823
R669 vdd.n7651 vdd.n7641 878.823
R670 vdd.n7706 vdd.n7678 878.823
R671 vdd.n7713 vdd.n7678 878.823
R672 vdd.n7685 vdd.n7681 878.823
R673 vdd.n7685 vdd.n7677 878.823
R674 vdd.n7687 vdd.n7683 878.823
R675 vdd.n7697 vdd.n7687 878.823
R676 vdd.n7754 vdd.n7726 878.823
R677 vdd.n7761 vdd.n7726 878.823
R678 vdd.n7733 vdd.n7729 878.823
R679 vdd.n7733 vdd.n7725 878.823
R680 vdd.n7735 vdd.n7731 878.823
R681 vdd.n7745 vdd.n7735 878.823
R682 vdd.n7466 vdd.n7447 878.823
R683 vdd.n7473 vdd.n7447 878.823
R684 vdd.n7452 vdd.n7451 878.823
R685 vdd.n7451 vdd.n7443 878.823
R686 vdd.n7458 vdd.n7441 878.823
R687 vdd.n7480 vdd.n7441 878.823
R688 vdd.n7801 vdd.n7773 878.823
R689 vdd.n7808 vdd.n7773 878.823
R690 vdd.n7780 vdd.n7776 878.823
R691 vdd.n7780 vdd.n7772 878.823
R692 vdd.n7782 vdd.n7778 878.823
R693 vdd.n7792 vdd.n7782 878.823
R694 vdd.n7846 vdd.n7818 878.823
R695 vdd.n7853 vdd.n7818 878.823
R696 vdd.n7825 vdd.n7821 878.823
R697 vdd.n7825 vdd.n7817 878.823
R698 vdd.n7827 vdd.n7823 878.823
R699 vdd.n7837 vdd.n7827 878.823
R700 vdd.n7892 vdd.n7864 878.823
R701 vdd.n7899 vdd.n7864 878.823
R702 vdd.n7871 vdd.n7867 878.823
R703 vdd.n7871 vdd.n7863 878.823
R704 vdd.n7873 vdd.n7869 878.823
R705 vdd.n7883 vdd.n7873 878.823
R706 vdd.n7943 vdd.n7915 878.823
R707 vdd.n7950 vdd.n7915 878.823
R708 vdd.n7922 vdd.n7918 878.823
R709 vdd.n7922 vdd.n7914 878.823
R710 vdd.n7924 vdd.n7920 878.823
R711 vdd.n7934 vdd.n7924 878.823
R712 vdd.n7989 vdd.n7961 878.823
R713 vdd.n7996 vdd.n7961 878.823
R714 vdd.n7968 vdd.n7964 878.823
R715 vdd.n7968 vdd.n7960 878.823
R716 vdd.n7970 vdd.n7966 878.823
R717 vdd.n7980 vdd.n7970 878.823
R718 vdd.n8037 vdd.n8009 878.823
R719 vdd.n8044 vdd.n8009 878.823
R720 vdd.n8016 vdd.n8012 878.823
R721 vdd.n8016 vdd.n8008 878.823
R722 vdd.n8018 vdd.n8014 878.823
R723 vdd.n8028 vdd.n8018 878.823
R724 vdd.n8083 vdd.n8055 878.823
R725 vdd.n8090 vdd.n8055 878.823
R726 vdd.n8062 vdd.n8058 878.823
R727 vdd.n8062 vdd.n8054 878.823
R728 vdd.n8064 vdd.n8060 878.823
R729 vdd.n8074 vdd.n8064 878.823
R730 vdd.n8128 vdd.n8100 878.823
R731 vdd.n8135 vdd.n8100 878.823
R732 vdd.n8107 vdd.n8103 878.823
R733 vdd.n8107 vdd.n8099 878.823
R734 vdd.n8109 vdd.n8105 878.823
R735 vdd.n8119 vdd.n8109 878.823
R736 vdd.n8178 vdd.n8150 878.823
R737 vdd.n8185 vdd.n8150 878.823
R738 vdd.n8157 vdd.n8153 878.823
R739 vdd.n8157 vdd.n8149 878.823
R740 vdd.n8159 vdd.n8155 878.823
R741 vdd.n8169 vdd.n8159 878.823
R742 vdd.n8224 vdd.n8196 878.823
R743 vdd.n8231 vdd.n8196 878.823
R744 vdd.n8203 vdd.n8199 878.823
R745 vdd.n8203 vdd.n8195 878.823
R746 vdd.n8205 vdd.n8201 878.823
R747 vdd.n8215 vdd.n8205 878.823
R748 vdd.n8272 vdd.n8244 878.823
R749 vdd.n8279 vdd.n8244 878.823
R750 vdd.n8251 vdd.n8247 878.823
R751 vdd.n8251 vdd.n8243 878.823
R752 vdd.n8253 vdd.n8249 878.823
R753 vdd.n8263 vdd.n8253 878.823
R754 vdd.n7231 vdd.n7212 878.823
R755 vdd.n7238 vdd.n7212 878.823
R756 vdd.n7217 vdd.n7216 878.823
R757 vdd.n7216 vdd.n7208 878.823
R758 vdd.n7223 vdd.n7206 878.823
R759 vdd.n7245 vdd.n7206 878.823
R760 vdd.n8319 vdd.n8291 878.823
R761 vdd.n8326 vdd.n8291 878.823
R762 vdd.n8298 vdd.n8294 878.823
R763 vdd.n8298 vdd.n8290 878.823
R764 vdd.n8300 vdd.n8296 878.823
R765 vdd.n8310 vdd.n8300 878.823
R766 vdd.n8364 vdd.n8336 878.823
R767 vdd.n8371 vdd.n8336 878.823
R768 vdd.n8343 vdd.n8339 878.823
R769 vdd.n8343 vdd.n8335 878.823
R770 vdd.n8345 vdd.n8341 878.823
R771 vdd.n8355 vdd.n8345 878.823
R772 vdd.n8414 vdd.n8386 878.823
R773 vdd.n8421 vdd.n8386 878.823
R774 vdd.n8393 vdd.n8389 878.823
R775 vdd.n8393 vdd.n8385 878.823
R776 vdd.n8395 vdd.n8391 878.823
R777 vdd.n8405 vdd.n8395 878.823
R778 vdd.n8460 vdd.n8432 878.823
R779 vdd.n8467 vdd.n8432 878.823
R780 vdd.n8439 vdd.n8435 878.823
R781 vdd.n8439 vdd.n8431 878.823
R782 vdd.n8441 vdd.n8437 878.823
R783 vdd.n8451 vdd.n8441 878.823
R784 vdd.n8508 vdd.n8480 878.823
R785 vdd.n8515 vdd.n8480 878.823
R786 vdd.n8487 vdd.n8483 878.823
R787 vdd.n8487 vdd.n8479 878.823
R788 vdd.n8489 vdd.n8485 878.823
R789 vdd.n8499 vdd.n8489 878.823
R790 vdd.n8625 vdd.n8617 878.823
R791 vdd.n8626 vdd.n8625 878.823
R792 vdd.n8638 vdd.n8628 878.823
R793 vdd.n8628 vdd.n8624 878.823
R794 vdd.n8652 vdd.n8618 878.823
R795 vdd.n8652 vdd.n8651 878.823
R796 vdd.n8579 vdd.n8571 878.823
R797 vdd.n8580 vdd.n8579 878.823
R798 vdd.n8592 vdd.n8582 878.823
R799 vdd.n8582 vdd.n8578 878.823
R800 vdd.n8606 vdd.n8572 878.823
R801 vdd.n8606 vdd.n8605 878.823
R802 vdd.n8672 vdd.n8664 878.823
R803 vdd.n8673 vdd.n8672 878.823
R804 vdd.n8685 vdd.n8675 878.823
R805 vdd.n8675 vdd.n8671 878.823
R806 vdd.n8699 vdd.n8665 878.823
R807 vdd.n8699 vdd.n8698 878.823
R808 vdd.n8720 vdd.n8712 878.823
R809 vdd.n8721 vdd.n8720 878.823
R810 vdd.n8733 vdd.n8723 878.823
R811 vdd.n8723 vdd.n8719 878.823
R812 vdd.n8747 vdd.n8713 878.823
R813 vdd.n8747 vdd.n8746 878.823
R814 vdd.n8766 vdd.n8758 878.823
R815 vdd.n8767 vdd.n8766 878.823
R816 vdd.n8779 vdd.n8769 878.823
R817 vdd.n8769 vdd.n8765 878.823
R818 vdd.n8793 vdd.n8759 878.823
R819 vdd.n8793 vdd.n8792 878.823
R820 vdd.n7025 vdd.n7022 878.823
R821 vdd.n7026 vdd.n7025 878.823
R822 vdd.n7030 vdd.n7021 878.823
R823 vdd.n7031 vdd.n7030 878.823
R824 vdd.n7052 vdd.n7051 878.823
R825 vdd.n7051 vdd.n7016 878.823
R826 vdd.n8908 vdd.n8900 878.823
R827 vdd.n8909 vdd.n8908 878.823
R828 vdd.n8921 vdd.n8911 878.823
R829 vdd.n8911 vdd.n8907 878.823
R830 vdd.n8935 vdd.n8901 878.823
R831 vdd.n8935 vdd.n8934 878.823
R832 vdd.n8861 vdd.n8853 878.823
R833 vdd.n8862 vdd.n8861 878.823
R834 vdd.n8874 vdd.n8864 878.823
R835 vdd.n8864 vdd.n8860 878.823
R836 vdd.n8888 vdd.n8854 878.823
R837 vdd.n8888 vdd.n8887 878.823
R838 vdd.n8815 vdd.n8807 878.823
R839 vdd.n8816 vdd.n8815 878.823
R840 vdd.n8828 vdd.n8818 878.823
R841 vdd.n8818 vdd.n8814 878.823
R842 vdd.n8842 vdd.n8808 878.823
R843 vdd.n8842 vdd.n8841 878.823
R844 vdd.n8955 vdd.n8947 878.823
R845 vdd.n8956 vdd.n8955 878.823
R846 vdd.n8968 vdd.n8958 878.823
R847 vdd.n8958 vdd.n8954 878.823
R848 vdd.n8982 vdd.n8948 878.823
R849 vdd.n8982 vdd.n8981 878.823
R850 vdd.n9003 vdd.n8995 878.823
R851 vdd.n9004 vdd.n9003 878.823
R852 vdd.n9016 vdd.n9006 878.823
R853 vdd.n9006 vdd.n9002 878.823
R854 vdd.n9030 vdd.n8996 878.823
R855 vdd.n9030 vdd.n9029 878.823
R856 vdd.n9049 vdd.n9041 878.823
R857 vdd.n9050 vdd.n9049 878.823
R858 vdd.n9062 vdd.n9052 878.823
R859 vdd.n9052 vdd.n9048 878.823
R860 vdd.n9076 vdd.n9042 878.823
R861 vdd.n9076 vdd.n9075 878.823
R862 vdd.n9143 vdd.n9135 878.823
R863 vdd.n9144 vdd.n9143 878.823
R864 vdd.n9156 vdd.n9146 878.823
R865 vdd.n9146 vdd.n9142 878.823
R866 vdd.n9170 vdd.n9136 878.823
R867 vdd.n9170 vdd.n9169 878.823
R868 vdd.n9097 vdd.n9089 878.823
R869 vdd.n9098 vdd.n9097 878.823
R870 vdd.n9110 vdd.n9100 878.823
R871 vdd.n9100 vdd.n9096 878.823
R872 vdd.n9124 vdd.n9090 878.823
R873 vdd.n9124 vdd.n9123 878.823
R874 vdd.n9190 vdd.n9182 878.823
R875 vdd.n9191 vdd.n9190 878.823
R876 vdd.n9203 vdd.n9193 878.823
R877 vdd.n9193 vdd.n9189 878.823
R878 vdd.n9217 vdd.n9183 878.823
R879 vdd.n9217 vdd.n9216 878.823
R880 vdd.n9238 vdd.n9230 878.823
R881 vdd.n9239 vdd.n9238 878.823
R882 vdd.n9251 vdd.n9241 878.823
R883 vdd.n9241 vdd.n9237 878.823
R884 vdd.n9265 vdd.n9231 878.823
R885 vdd.n9265 vdd.n9264 878.823
R886 vdd.n9284 vdd.n9276 878.823
R887 vdd.n9285 vdd.n9284 878.823
R888 vdd.n9297 vdd.n9287 878.823
R889 vdd.n9287 vdd.n9283 878.823
R890 vdd.n9311 vdd.n9277 878.823
R891 vdd.n9311 vdd.n9310 878.823
R892 vdd.n6789 vdd.n6786 878.823
R893 vdd.n6790 vdd.n6789 878.823
R894 vdd.n6794 vdd.n6785 878.823
R895 vdd.n6795 vdd.n6794 878.823
R896 vdd.n6816 vdd.n6815 878.823
R897 vdd.n6815 vdd.n6780 878.823
R898 vdd.n9379 vdd.n9371 878.823
R899 vdd.n9380 vdd.n9379 878.823
R900 vdd.n9392 vdd.n9382 878.823
R901 vdd.n9382 vdd.n9378 878.823
R902 vdd.n9406 vdd.n9372 878.823
R903 vdd.n9406 vdd.n9405 878.823
R904 vdd.n9333 vdd.n9325 878.823
R905 vdd.n9334 vdd.n9333 878.823
R906 vdd.n9346 vdd.n9336 878.823
R907 vdd.n9336 vdd.n9332 878.823
R908 vdd.n9360 vdd.n9326 878.823
R909 vdd.n9360 vdd.n9359 878.823
R910 vdd.n9426 vdd.n9418 878.823
R911 vdd.n9427 vdd.n9426 878.823
R912 vdd.n9439 vdd.n9429 878.823
R913 vdd.n9429 vdd.n9425 878.823
R914 vdd.n9453 vdd.n9419 878.823
R915 vdd.n9453 vdd.n9452 878.823
R916 vdd.n9474 vdd.n9466 878.823
R917 vdd.n9475 vdd.n9474 878.823
R918 vdd.n9487 vdd.n9477 878.823
R919 vdd.n9477 vdd.n9473 878.823
R920 vdd.n9501 vdd.n9467 878.823
R921 vdd.n9501 vdd.n9500 878.823
R922 vdd.n9520 vdd.n9512 878.823
R923 vdd.n9521 vdd.n9520 878.823
R924 vdd.n9533 vdd.n9523 878.823
R925 vdd.n9523 vdd.n9519 878.823
R926 vdd.n9547 vdd.n9513 878.823
R927 vdd.n9547 vdd.n9546 878.823
R928 vdd.n3680 vdd.n3672 878.823
R929 vdd.n3681 vdd.n3680 878.823
R930 vdd.n3693 vdd.n3683 878.823
R931 vdd.n3683 vdd.n3679 878.823
R932 vdd.n3707 vdd.n3673 878.823
R933 vdd.n3707 vdd.n3706 878.823
R934 vdd.n3726 vdd.n3718 878.823
R935 vdd.n3727 vdd.n3726 878.823
R936 vdd.n3739 vdd.n3729 878.823
R937 vdd.n3729 vdd.n3725 878.823
R938 vdd.n3753 vdd.n3719 878.823
R939 vdd.n3753 vdd.n3752 878.823
R940 vdd.n3824 vdd.n3816 878.823
R941 vdd.n3825 vdd.n3824 878.823
R942 vdd.n3837 vdd.n3827 878.823
R943 vdd.n3827 vdd.n3823 878.823
R944 vdd.n3851 vdd.n3817 878.823
R945 vdd.n3851 vdd.n3850 878.823
R946 vdd.n3870 vdd.n3862 878.823
R947 vdd.n3871 vdd.n3870 878.823
R948 vdd.n3883 vdd.n3873 878.823
R949 vdd.n3873 vdd.n3869 878.823
R950 vdd.n3897 vdd.n3863 878.823
R951 vdd.n3897 vdd.n3896 878.823
R952 vdd.n3916 vdd.n3908 878.823
R953 vdd.n3917 vdd.n3916 878.823
R954 vdd.n3929 vdd.n3919 878.823
R955 vdd.n3919 vdd.n3915 878.823
R956 vdd.n3943 vdd.n3909 878.823
R957 vdd.n3943 vdd.n3942 878.823
R958 vdd.n3962 vdd.n3954 878.823
R959 vdd.n3963 vdd.n3962 878.823
R960 vdd.n3975 vdd.n3965 878.823
R961 vdd.n3965 vdd.n3961 878.823
R962 vdd.n3989 vdd.n3955 878.823
R963 vdd.n3989 vdd.n3988 878.823
R964 vdd.n4060 vdd.n4052 878.823
R965 vdd.n4061 vdd.n4060 878.823
R966 vdd.n4073 vdd.n4063 878.823
R967 vdd.n4063 vdd.n4059 878.823
R968 vdd.n4087 vdd.n4053 878.823
R969 vdd.n4087 vdd.n4086 878.823
R970 vdd.n5518 vdd.n5510 878.823
R971 vdd.n5519 vdd.n5518 878.823
R972 vdd.n5531 vdd.n5521 878.823
R973 vdd.n5521 vdd.n5517 878.823
R974 vdd.n5545 vdd.n5511 878.823
R975 vdd.n5545 vdd.n5544 878.823
R976 vdd.n4129 vdd.n4101 878.823
R977 vdd.n4136 vdd.n4101 878.823
R978 vdd.n4108 vdd.n4104 878.823
R979 vdd.n4108 vdd.n4100 878.823
R980 vdd.n4110 vdd.n4106 878.823
R981 vdd.n4120 vdd.n4110 878.823
R982 vdd.n4175 vdd.n4147 878.823
R983 vdd.n4182 vdd.n4147 878.823
R984 vdd.n4154 vdd.n4150 878.823
R985 vdd.n4154 vdd.n4146 878.823
R986 vdd.n4156 vdd.n4152 878.823
R987 vdd.n4166 vdd.n4156 878.823
R988 vdd.n4272 vdd.n4244 878.823
R989 vdd.n4279 vdd.n4244 878.823
R990 vdd.n4251 vdd.n4247 878.823
R991 vdd.n4251 vdd.n4243 878.823
R992 vdd.n4253 vdd.n4249 878.823
R993 vdd.n4263 vdd.n4253 878.823
R994 vdd.n4318 vdd.n4290 878.823
R995 vdd.n4325 vdd.n4290 878.823
R996 vdd.n4297 vdd.n4293 878.823
R997 vdd.n4297 vdd.n4289 878.823
R998 vdd.n4299 vdd.n4295 878.823
R999 vdd.n4309 vdd.n4299 878.823
R1000 vdd.n4364 vdd.n4336 878.823
R1001 vdd.n4371 vdd.n4336 878.823
R1002 vdd.n4343 vdd.n4339 878.823
R1003 vdd.n4343 vdd.n4335 878.823
R1004 vdd.n4345 vdd.n4341 878.823
R1005 vdd.n4355 vdd.n4345 878.823
R1006 vdd.n4410 vdd.n4382 878.823
R1007 vdd.n4417 vdd.n4382 878.823
R1008 vdd.n4389 vdd.n4385 878.823
R1009 vdd.n4389 vdd.n4381 878.823
R1010 vdd.n4391 vdd.n4387 878.823
R1011 vdd.n4401 vdd.n4391 878.823
R1012 vdd.n4507 vdd.n4479 878.823
R1013 vdd.n4514 vdd.n4479 878.823
R1014 vdd.n4486 vdd.n4482 878.823
R1015 vdd.n4486 vdd.n4478 878.823
R1016 vdd.n4488 vdd.n4484 878.823
R1017 vdd.n4498 vdd.n4488 878.823
R1018 vdd.n3656 vdd.n3628 878.823
R1019 vdd.n3663 vdd.n3628 878.823
R1020 vdd.n3635 vdd.n3631 878.823
R1021 vdd.n3635 vdd.n3627 878.823
R1022 vdd.n3637 vdd.n3633 878.823
R1023 vdd.n3647 vdd.n3637 878.823
R1024 vdd.n4551 vdd.n4523 878.823
R1025 vdd.n4558 vdd.n4523 878.823
R1026 vdd.n4530 vdd.n4526 878.823
R1027 vdd.n4530 vdd.n4522 878.823
R1028 vdd.n4532 vdd.n4528 878.823
R1029 vdd.n4542 vdd.n4532 878.823
R1030 vdd.n4596 vdd.n4568 878.823
R1031 vdd.n4603 vdd.n4568 878.823
R1032 vdd.n4575 vdd.n4571 878.823
R1033 vdd.n4575 vdd.n4567 878.823
R1034 vdd.n4577 vdd.n4573 878.823
R1035 vdd.n4587 vdd.n4577 878.823
R1036 vdd.n4646 vdd.n4618 878.823
R1037 vdd.n4653 vdd.n4618 878.823
R1038 vdd.n4625 vdd.n4621 878.823
R1039 vdd.n4625 vdd.n4617 878.823
R1040 vdd.n4627 vdd.n4623 878.823
R1041 vdd.n4637 vdd.n4627 878.823
R1042 vdd.n4692 vdd.n4664 878.823
R1043 vdd.n4699 vdd.n4664 878.823
R1044 vdd.n4671 vdd.n4667 878.823
R1045 vdd.n4671 vdd.n4663 878.823
R1046 vdd.n4673 vdd.n4669 878.823
R1047 vdd.n4683 vdd.n4673 878.823
R1048 vdd.n4740 vdd.n4712 878.823
R1049 vdd.n4747 vdd.n4712 878.823
R1050 vdd.n4719 vdd.n4715 878.823
R1051 vdd.n4719 vdd.n4711 878.823
R1052 vdd.n4721 vdd.n4717 878.823
R1053 vdd.n4731 vdd.n4721 878.823
R1054 vdd.n4452 vdd.n4433 878.823
R1055 vdd.n4459 vdd.n4433 878.823
R1056 vdd.n4438 vdd.n4437 878.823
R1057 vdd.n4437 vdd.n4429 878.823
R1058 vdd.n4444 vdd.n4427 878.823
R1059 vdd.n4466 vdd.n4427 878.823
R1060 vdd.n4787 vdd.n4759 878.823
R1061 vdd.n4794 vdd.n4759 878.823
R1062 vdd.n4766 vdd.n4762 878.823
R1063 vdd.n4766 vdd.n4758 878.823
R1064 vdd.n4768 vdd.n4764 878.823
R1065 vdd.n4778 vdd.n4768 878.823
R1066 vdd.n4832 vdd.n4804 878.823
R1067 vdd.n4839 vdd.n4804 878.823
R1068 vdd.n4811 vdd.n4807 878.823
R1069 vdd.n4811 vdd.n4803 878.823
R1070 vdd.n4813 vdd.n4809 878.823
R1071 vdd.n4823 vdd.n4813 878.823
R1072 vdd.n4878 vdd.n4850 878.823
R1073 vdd.n4885 vdd.n4850 878.823
R1074 vdd.n4857 vdd.n4853 878.823
R1075 vdd.n4857 vdd.n4849 878.823
R1076 vdd.n4859 vdd.n4855 878.823
R1077 vdd.n4869 vdd.n4859 878.823
R1078 vdd.n4929 vdd.n4901 878.823
R1079 vdd.n4936 vdd.n4901 878.823
R1080 vdd.n4908 vdd.n4904 878.823
R1081 vdd.n4908 vdd.n4900 878.823
R1082 vdd.n4910 vdd.n4906 878.823
R1083 vdd.n4920 vdd.n4910 878.823
R1084 vdd.n4975 vdd.n4947 878.823
R1085 vdd.n4982 vdd.n4947 878.823
R1086 vdd.n4954 vdd.n4950 878.823
R1087 vdd.n4954 vdd.n4946 878.823
R1088 vdd.n4956 vdd.n4952 878.823
R1089 vdd.n4966 vdd.n4956 878.823
R1090 vdd.n5023 vdd.n4995 878.823
R1091 vdd.n5030 vdd.n4995 878.823
R1092 vdd.n5002 vdd.n4998 878.823
R1093 vdd.n5002 vdd.n4994 878.823
R1094 vdd.n5004 vdd.n5000 878.823
R1095 vdd.n5014 vdd.n5004 878.823
R1096 vdd.n5069 vdd.n5041 878.823
R1097 vdd.n5076 vdd.n5041 878.823
R1098 vdd.n5048 vdd.n5044 878.823
R1099 vdd.n5048 vdd.n5040 878.823
R1100 vdd.n5050 vdd.n5046 878.823
R1101 vdd.n5060 vdd.n5050 878.823
R1102 vdd.n5114 vdd.n5086 878.823
R1103 vdd.n5121 vdd.n5086 878.823
R1104 vdd.n5093 vdd.n5089 878.823
R1105 vdd.n5093 vdd.n5085 878.823
R1106 vdd.n5095 vdd.n5091 878.823
R1107 vdd.n5105 vdd.n5095 878.823
R1108 vdd.n5164 vdd.n5136 878.823
R1109 vdd.n5171 vdd.n5136 878.823
R1110 vdd.n5143 vdd.n5139 878.823
R1111 vdd.n5143 vdd.n5135 878.823
R1112 vdd.n5145 vdd.n5141 878.823
R1113 vdd.n5155 vdd.n5145 878.823
R1114 vdd.n5210 vdd.n5182 878.823
R1115 vdd.n5217 vdd.n5182 878.823
R1116 vdd.n5189 vdd.n5185 878.823
R1117 vdd.n5189 vdd.n5181 878.823
R1118 vdd.n5191 vdd.n5187 878.823
R1119 vdd.n5201 vdd.n5191 878.823
R1120 vdd.n5258 vdd.n5230 878.823
R1121 vdd.n5265 vdd.n5230 878.823
R1122 vdd.n5237 vdd.n5233 878.823
R1123 vdd.n5237 vdd.n5229 878.823
R1124 vdd.n5239 vdd.n5235 878.823
R1125 vdd.n5249 vdd.n5239 878.823
R1126 vdd.n4217 vdd.n4198 878.823
R1127 vdd.n4224 vdd.n4198 878.823
R1128 vdd.n4203 vdd.n4202 878.823
R1129 vdd.n4202 vdd.n4194 878.823
R1130 vdd.n4209 vdd.n4192 878.823
R1131 vdd.n4231 vdd.n4192 878.823
R1132 vdd.n5305 vdd.n5277 878.823
R1133 vdd.n5312 vdd.n5277 878.823
R1134 vdd.n5284 vdd.n5280 878.823
R1135 vdd.n5284 vdd.n5276 878.823
R1136 vdd.n5286 vdd.n5282 878.823
R1137 vdd.n5296 vdd.n5286 878.823
R1138 vdd.n5350 vdd.n5322 878.823
R1139 vdd.n5357 vdd.n5322 878.823
R1140 vdd.n5329 vdd.n5325 878.823
R1141 vdd.n5329 vdd.n5321 878.823
R1142 vdd.n5331 vdd.n5327 878.823
R1143 vdd.n5341 vdd.n5331 878.823
R1144 vdd.n5400 vdd.n5372 878.823
R1145 vdd.n5407 vdd.n5372 878.823
R1146 vdd.n5379 vdd.n5375 878.823
R1147 vdd.n5379 vdd.n5371 878.823
R1148 vdd.n5381 vdd.n5377 878.823
R1149 vdd.n5391 vdd.n5381 878.823
R1150 vdd.n5446 vdd.n5418 878.823
R1151 vdd.n5453 vdd.n5418 878.823
R1152 vdd.n5425 vdd.n5421 878.823
R1153 vdd.n5425 vdd.n5417 878.823
R1154 vdd.n5427 vdd.n5423 878.823
R1155 vdd.n5437 vdd.n5427 878.823
R1156 vdd.n5494 vdd.n5466 878.823
R1157 vdd.n5501 vdd.n5466 878.823
R1158 vdd.n5473 vdd.n5469 878.823
R1159 vdd.n5473 vdd.n5465 878.823
R1160 vdd.n5475 vdd.n5471 878.823
R1161 vdd.n5485 vdd.n5475 878.823
R1162 vdd.n5611 vdd.n5603 878.823
R1163 vdd.n5612 vdd.n5611 878.823
R1164 vdd.n5624 vdd.n5614 878.823
R1165 vdd.n5614 vdd.n5610 878.823
R1166 vdd.n5638 vdd.n5604 878.823
R1167 vdd.n5638 vdd.n5637 878.823
R1168 vdd.n5565 vdd.n5557 878.823
R1169 vdd.n5566 vdd.n5565 878.823
R1170 vdd.n5578 vdd.n5568 878.823
R1171 vdd.n5568 vdd.n5564 878.823
R1172 vdd.n5592 vdd.n5558 878.823
R1173 vdd.n5592 vdd.n5591 878.823
R1174 vdd.n5658 vdd.n5650 878.823
R1175 vdd.n5659 vdd.n5658 878.823
R1176 vdd.n5671 vdd.n5661 878.823
R1177 vdd.n5661 vdd.n5657 878.823
R1178 vdd.n5685 vdd.n5651 878.823
R1179 vdd.n5685 vdd.n5684 878.823
R1180 vdd.n5706 vdd.n5698 878.823
R1181 vdd.n5707 vdd.n5706 878.823
R1182 vdd.n5719 vdd.n5709 878.823
R1183 vdd.n5709 vdd.n5705 878.823
R1184 vdd.n5733 vdd.n5699 878.823
R1185 vdd.n5733 vdd.n5732 878.823
R1186 vdd.n5752 vdd.n5744 878.823
R1187 vdd.n5753 vdd.n5752 878.823
R1188 vdd.n5765 vdd.n5755 878.823
R1189 vdd.n5755 vdd.n5751 878.823
R1190 vdd.n5779 vdd.n5745 878.823
R1191 vdd.n5779 vdd.n5778 878.823
R1192 vdd.n4011 vdd.n4008 878.823
R1193 vdd.n4012 vdd.n4011 878.823
R1194 vdd.n4016 vdd.n4007 878.823
R1195 vdd.n4017 vdd.n4016 878.823
R1196 vdd.n4038 vdd.n4037 878.823
R1197 vdd.n4037 vdd.n4002 878.823
R1198 vdd.n5894 vdd.n5886 878.823
R1199 vdd.n5895 vdd.n5894 878.823
R1200 vdd.n5907 vdd.n5897 878.823
R1201 vdd.n5897 vdd.n5893 878.823
R1202 vdd.n5921 vdd.n5887 878.823
R1203 vdd.n5921 vdd.n5920 878.823
R1204 vdd.n5847 vdd.n5839 878.823
R1205 vdd.n5848 vdd.n5847 878.823
R1206 vdd.n5860 vdd.n5850 878.823
R1207 vdd.n5850 vdd.n5846 878.823
R1208 vdd.n5874 vdd.n5840 878.823
R1209 vdd.n5874 vdd.n5873 878.823
R1210 vdd.n5801 vdd.n5793 878.823
R1211 vdd.n5802 vdd.n5801 878.823
R1212 vdd.n5814 vdd.n5804 878.823
R1213 vdd.n5804 vdd.n5800 878.823
R1214 vdd.n5828 vdd.n5794 878.823
R1215 vdd.n5828 vdd.n5827 878.823
R1216 vdd.n5941 vdd.n5933 878.823
R1217 vdd.n5942 vdd.n5941 878.823
R1218 vdd.n5954 vdd.n5944 878.823
R1219 vdd.n5944 vdd.n5940 878.823
R1220 vdd.n5968 vdd.n5934 878.823
R1221 vdd.n5968 vdd.n5967 878.823
R1222 vdd.n5989 vdd.n5981 878.823
R1223 vdd.n5990 vdd.n5989 878.823
R1224 vdd.n6002 vdd.n5992 878.823
R1225 vdd.n5992 vdd.n5988 878.823
R1226 vdd.n6016 vdd.n5982 878.823
R1227 vdd.n6016 vdd.n6015 878.823
R1228 vdd.n6035 vdd.n6027 878.823
R1229 vdd.n6036 vdd.n6035 878.823
R1230 vdd.n6048 vdd.n6038 878.823
R1231 vdd.n6038 vdd.n6034 878.823
R1232 vdd.n6062 vdd.n6028 878.823
R1233 vdd.n6062 vdd.n6061 878.823
R1234 vdd.n6129 vdd.n6121 878.823
R1235 vdd.n6130 vdd.n6129 878.823
R1236 vdd.n6142 vdd.n6132 878.823
R1237 vdd.n6132 vdd.n6128 878.823
R1238 vdd.n6156 vdd.n6122 878.823
R1239 vdd.n6156 vdd.n6155 878.823
R1240 vdd.n6083 vdd.n6075 878.823
R1241 vdd.n6084 vdd.n6083 878.823
R1242 vdd.n6096 vdd.n6086 878.823
R1243 vdd.n6086 vdd.n6082 878.823
R1244 vdd.n6110 vdd.n6076 878.823
R1245 vdd.n6110 vdd.n6109 878.823
R1246 vdd.n6176 vdd.n6168 878.823
R1247 vdd.n6177 vdd.n6176 878.823
R1248 vdd.n6189 vdd.n6179 878.823
R1249 vdd.n6179 vdd.n6175 878.823
R1250 vdd.n6203 vdd.n6169 878.823
R1251 vdd.n6203 vdd.n6202 878.823
R1252 vdd.n6224 vdd.n6216 878.823
R1253 vdd.n6225 vdd.n6224 878.823
R1254 vdd.n6237 vdd.n6227 878.823
R1255 vdd.n6227 vdd.n6223 878.823
R1256 vdd.n6251 vdd.n6217 878.823
R1257 vdd.n6251 vdd.n6250 878.823
R1258 vdd.n6270 vdd.n6262 878.823
R1259 vdd.n6271 vdd.n6270 878.823
R1260 vdd.n6283 vdd.n6273 878.823
R1261 vdd.n6273 vdd.n6269 878.823
R1262 vdd.n6297 vdd.n6263 878.823
R1263 vdd.n6297 vdd.n6296 878.823
R1264 vdd.n3775 vdd.n3772 878.823
R1265 vdd.n3776 vdd.n3775 878.823
R1266 vdd.n3780 vdd.n3771 878.823
R1267 vdd.n3781 vdd.n3780 878.823
R1268 vdd.n3802 vdd.n3801 878.823
R1269 vdd.n3801 vdd.n3766 878.823
R1270 vdd.n6365 vdd.n6357 878.823
R1271 vdd.n6366 vdd.n6365 878.823
R1272 vdd.n6378 vdd.n6368 878.823
R1273 vdd.n6368 vdd.n6364 878.823
R1274 vdd.n6392 vdd.n6358 878.823
R1275 vdd.n6392 vdd.n6391 878.823
R1276 vdd.n6319 vdd.n6311 878.823
R1277 vdd.n6320 vdd.n6319 878.823
R1278 vdd.n6332 vdd.n6322 878.823
R1279 vdd.n6322 vdd.n6318 878.823
R1280 vdd.n6346 vdd.n6312 878.823
R1281 vdd.n6346 vdd.n6345 878.823
R1282 vdd.n6412 vdd.n6404 878.823
R1283 vdd.n6413 vdd.n6412 878.823
R1284 vdd.n6425 vdd.n6415 878.823
R1285 vdd.n6415 vdd.n6411 878.823
R1286 vdd.n6439 vdd.n6405 878.823
R1287 vdd.n6439 vdd.n6438 878.823
R1288 vdd.n6460 vdd.n6452 878.823
R1289 vdd.n6461 vdd.n6460 878.823
R1290 vdd.n6473 vdd.n6463 878.823
R1291 vdd.n6463 vdd.n6459 878.823
R1292 vdd.n6487 vdd.n6453 878.823
R1293 vdd.n6487 vdd.n6486 878.823
R1294 vdd.n6506 vdd.n6498 878.823
R1295 vdd.n6507 vdd.n6506 878.823
R1296 vdd.n6519 vdd.n6509 878.823
R1297 vdd.n6509 vdd.n6505 878.823
R1298 vdd.n6533 vdd.n6499 878.823
R1299 vdd.n6533 vdd.n6532 878.823
R1300 vdd.n666 vdd.n658 878.823
R1301 vdd.n667 vdd.n666 878.823
R1302 vdd.n679 vdd.n669 878.823
R1303 vdd.n669 vdd.n665 878.823
R1304 vdd.n693 vdd.n659 878.823
R1305 vdd.n693 vdd.n692 878.823
R1306 vdd.n712 vdd.n704 878.823
R1307 vdd.n713 vdd.n712 878.823
R1308 vdd.n725 vdd.n715 878.823
R1309 vdd.n715 vdd.n711 878.823
R1310 vdd.n739 vdd.n705 878.823
R1311 vdd.n739 vdd.n738 878.823
R1312 vdd.n810 vdd.n802 878.823
R1313 vdd.n811 vdd.n810 878.823
R1314 vdd.n823 vdd.n813 878.823
R1315 vdd.n813 vdd.n809 878.823
R1316 vdd.n837 vdd.n803 878.823
R1317 vdd.n837 vdd.n836 878.823
R1318 vdd.n856 vdd.n848 878.823
R1319 vdd.n857 vdd.n856 878.823
R1320 vdd.n869 vdd.n859 878.823
R1321 vdd.n859 vdd.n855 878.823
R1322 vdd.n883 vdd.n849 878.823
R1323 vdd.n883 vdd.n882 878.823
R1324 vdd.n902 vdd.n894 878.823
R1325 vdd.n903 vdd.n902 878.823
R1326 vdd.n915 vdd.n905 878.823
R1327 vdd.n905 vdd.n901 878.823
R1328 vdd.n929 vdd.n895 878.823
R1329 vdd.n929 vdd.n928 878.823
R1330 vdd.n948 vdd.n940 878.823
R1331 vdd.n949 vdd.n948 878.823
R1332 vdd.n961 vdd.n951 878.823
R1333 vdd.n951 vdd.n947 878.823
R1334 vdd.n975 vdd.n941 878.823
R1335 vdd.n975 vdd.n974 878.823
R1336 vdd.n1046 vdd.n1038 878.823
R1337 vdd.n1047 vdd.n1046 878.823
R1338 vdd.n1059 vdd.n1049 878.823
R1339 vdd.n1049 vdd.n1045 878.823
R1340 vdd.n1073 vdd.n1039 878.823
R1341 vdd.n1073 vdd.n1072 878.823
R1342 vdd.n2504 vdd.n2496 878.823
R1343 vdd.n2505 vdd.n2504 878.823
R1344 vdd.n2517 vdd.n2507 878.823
R1345 vdd.n2507 vdd.n2503 878.823
R1346 vdd.n2531 vdd.n2497 878.823
R1347 vdd.n2531 vdd.n2530 878.823
R1348 vdd.n1115 vdd.n1087 878.823
R1349 vdd.n1122 vdd.n1087 878.823
R1350 vdd.n1094 vdd.n1090 878.823
R1351 vdd.n1094 vdd.n1086 878.823
R1352 vdd.n1096 vdd.n1092 878.823
R1353 vdd.n1106 vdd.n1096 878.823
R1354 vdd.n1161 vdd.n1133 878.823
R1355 vdd.n1168 vdd.n1133 878.823
R1356 vdd.n1140 vdd.n1136 878.823
R1357 vdd.n1140 vdd.n1132 878.823
R1358 vdd.n1142 vdd.n1138 878.823
R1359 vdd.n1152 vdd.n1142 878.823
R1360 vdd.n1258 vdd.n1230 878.823
R1361 vdd.n1265 vdd.n1230 878.823
R1362 vdd.n1237 vdd.n1233 878.823
R1363 vdd.n1237 vdd.n1229 878.823
R1364 vdd.n1239 vdd.n1235 878.823
R1365 vdd.n1249 vdd.n1239 878.823
R1366 vdd.n1304 vdd.n1276 878.823
R1367 vdd.n1311 vdd.n1276 878.823
R1368 vdd.n1283 vdd.n1279 878.823
R1369 vdd.n1283 vdd.n1275 878.823
R1370 vdd.n1285 vdd.n1281 878.823
R1371 vdd.n1295 vdd.n1285 878.823
R1372 vdd.n1350 vdd.n1322 878.823
R1373 vdd.n1357 vdd.n1322 878.823
R1374 vdd.n1329 vdd.n1325 878.823
R1375 vdd.n1329 vdd.n1321 878.823
R1376 vdd.n1331 vdd.n1327 878.823
R1377 vdd.n1341 vdd.n1331 878.823
R1378 vdd.n1396 vdd.n1368 878.823
R1379 vdd.n1403 vdd.n1368 878.823
R1380 vdd.n1375 vdd.n1371 878.823
R1381 vdd.n1375 vdd.n1367 878.823
R1382 vdd.n1377 vdd.n1373 878.823
R1383 vdd.n1387 vdd.n1377 878.823
R1384 vdd.n1493 vdd.n1465 878.823
R1385 vdd.n1500 vdd.n1465 878.823
R1386 vdd.n1472 vdd.n1468 878.823
R1387 vdd.n1472 vdd.n1464 878.823
R1388 vdd.n1474 vdd.n1470 878.823
R1389 vdd.n1484 vdd.n1474 878.823
R1390 vdd.n642 vdd.n614 878.823
R1391 vdd.n649 vdd.n614 878.823
R1392 vdd.n621 vdd.n617 878.823
R1393 vdd.n621 vdd.n613 878.823
R1394 vdd.n623 vdd.n619 878.823
R1395 vdd.n633 vdd.n623 878.823
R1396 vdd.n1537 vdd.n1509 878.823
R1397 vdd.n1544 vdd.n1509 878.823
R1398 vdd.n1516 vdd.n1512 878.823
R1399 vdd.n1516 vdd.n1508 878.823
R1400 vdd.n1518 vdd.n1514 878.823
R1401 vdd.n1528 vdd.n1518 878.823
R1402 vdd.n1582 vdd.n1554 878.823
R1403 vdd.n1589 vdd.n1554 878.823
R1404 vdd.n1561 vdd.n1557 878.823
R1405 vdd.n1561 vdd.n1553 878.823
R1406 vdd.n1563 vdd.n1559 878.823
R1407 vdd.n1573 vdd.n1563 878.823
R1408 vdd.n1632 vdd.n1604 878.823
R1409 vdd.n1639 vdd.n1604 878.823
R1410 vdd.n1611 vdd.n1607 878.823
R1411 vdd.n1611 vdd.n1603 878.823
R1412 vdd.n1613 vdd.n1609 878.823
R1413 vdd.n1623 vdd.n1613 878.823
R1414 vdd.n1678 vdd.n1650 878.823
R1415 vdd.n1685 vdd.n1650 878.823
R1416 vdd.n1657 vdd.n1653 878.823
R1417 vdd.n1657 vdd.n1649 878.823
R1418 vdd.n1659 vdd.n1655 878.823
R1419 vdd.n1669 vdd.n1659 878.823
R1420 vdd.n1726 vdd.n1698 878.823
R1421 vdd.n1733 vdd.n1698 878.823
R1422 vdd.n1705 vdd.n1701 878.823
R1423 vdd.n1705 vdd.n1697 878.823
R1424 vdd.n1707 vdd.n1703 878.823
R1425 vdd.n1717 vdd.n1707 878.823
R1426 vdd.n1438 vdd.n1419 878.823
R1427 vdd.n1445 vdd.n1419 878.823
R1428 vdd.n1424 vdd.n1423 878.823
R1429 vdd.n1423 vdd.n1415 878.823
R1430 vdd.n1430 vdd.n1413 878.823
R1431 vdd.n1452 vdd.n1413 878.823
R1432 vdd.n1773 vdd.n1745 878.823
R1433 vdd.n1780 vdd.n1745 878.823
R1434 vdd.n1752 vdd.n1748 878.823
R1435 vdd.n1752 vdd.n1744 878.823
R1436 vdd.n1754 vdd.n1750 878.823
R1437 vdd.n1764 vdd.n1754 878.823
R1438 vdd.n1818 vdd.n1790 878.823
R1439 vdd.n1825 vdd.n1790 878.823
R1440 vdd.n1797 vdd.n1793 878.823
R1441 vdd.n1797 vdd.n1789 878.823
R1442 vdd.n1799 vdd.n1795 878.823
R1443 vdd.n1809 vdd.n1799 878.823
R1444 vdd.n1864 vdd.n1836 878.823
R1445 vdd.n1871 vdd.n1836 878.823
R1446 vdd.n1843 vdd.n1839 878.823
R1447 vdd.n1843 vdd.n1835 878.823
R1448 vdd.n1845 vdd.n1841 878.823
R1449 vdd.n1855 vdd.n1845 878.823
R1450 vdd.n1915 vdd.n1887 878.823
R1451 vdd.n1922 vdd.n1887 878.823
R1452 vdd.n1894 vdd.n1890 878.823
R1453 vdd.n1894 vdd.n1886 878.823
R1454 vdd.n1896 vdd.n1892 878.823
R1455 vdd.n1906 vdd.n1896 878.823
R1456 vdd.n1961 vdd.n1933 878.823
R1457 vdd.n1968 vdd.n1933 878.823
R1458 vdd.n1940 vdd.n1936 878.823
R1459 vdd.n1940 vdd.n1932 878.823
R1460 vdd.n1942 vdd.n1938 878.823
R1461 vdd.n1952 vdd.n1942 878.823
R1462 vdd.n2009 vdd.n1981 878.823
R1463 vdd.n2016 vdd.n1981 878.823
R1464 vdd.n1988 vdd.n1984 878.823
R1465 vdd.n1988 vdd.n1980 878.823
R1466 vdd.n1990 vdd.n1986 878.823
R1467 vdd.n2000 vdd.n1990 878.823
R1468 vdd.n2055 vdd.n2027 878.823
R1469 vdd.n2062 vdd.n2027 878.823
R1470 vdd.n2034 vdd.n2030 878.823
R1471 vdd.n2034 vdd.n2026 878.823
R1472 vdd.n2036 vdd.n2032 878.823
R1473 vdd.n2046 vdd.n2036 878.823
R1474 vdd.n2100 vdd.n2072 878.823
R1475 vdd.n2107 vdd.n2072 878.823
R1476 vdd.n2079 vdd.n2075 878.823
R1477 vdd.n2079 vdd.n2071 878.823
R1478 vdd.n2081 vdd.n2077 878.823
R1479 vdd.n2091 vdd.n2081 878.823
R1480 vdd.n2150 vdd.n2122 878.823
R1481 vdd.n2157 vdd.n2122 878.823
R1482 vdd.n2129 vdd.n2125 878.823
R1483 vdd.n2129 vdd.n2121 878.823
R1484 vdd.n2131 vdd.n2127 878.823
R1485 vdd.n2141 vdd.n2131 878.823
R1486 vdd.n2196 vdd.n2168 878.823
R1487 vdd.n2203 vdd.n2168 878.823
R1488 vdd.n2175 vdd.n2171 878.823
R1489 vdd.n2175 vdd.n2167 878.823
R1490 vdd.n2177 vdd.n2173 878.823
R1491 vdd.n2187 vdd.n2177 878.823
R1492 vdd.n2244 vdd.n2216 878.823
R1493 vdd.n2251 vdd.n2216 878.823
R1494 vdd.n2223 vdd.n2219 878.823
R1495 vdd.n2223 vdd.n2215 878.823
R1496 vdd.n2225 vdd.n2221 878.823
R1497 vdd.n2235 vdd.n2225 878.823
R1498 vdd.n1203 vdd.n1184 878.823
R1499 vdd.n1210 vdd.n1184 878.823
R1500 vdd.n1189 vdd.n1188 878.823
R1501 vdd.n1188 vdd.n1180 878.823
R1502 vdd.n1195 vdd.n1178 878.823
R1503 vdd.n1217 vdd.n1178 878.823
R1504 vdd.n2291 vdd.n2263 878.823
R1505 vdd.n2298 vdd.n2263 878.823
R1506 vdd.n2270 vdd.n2266 878.823
R1507 vdd.n2270 vdd.n2262 878.823
R1508 vdd.n2272 vdd.n2268 878.823
R1509 vdd.n2282 vdd.n2272 878.823
R1510 vdd.n2336 vdd.n2308 878.823
R1511 vdd.n2343 vdd.n2308 878.823
R1512 vdd.n2315 vdd.n2311 878.823
R1513 vdd.n2315 vdd.n2307 878.823
R1514 vdd.n2317 vdd.n2313 878.823
R1515 vdd.n2327 vdd.n2317 878.823
R1516 vdd.n2386 vdd.n2358 878.823
R1517 vdd.n2393 vdd.n2358 878.823
R1518 vdd.n2365 vdd.n2361 878.823
R1519 vdd.n2365 vdd.n2357 878.823
R1520 vdd.n2367 vdd.n2363 878.823
R1521 vdd.n2377 vdd.n2367 878.823
R1522 vdd.n2432 vdd.n2404 878.823
R1523 vdd.n2439 vdd.n2404 878.823
R1524 vdd.n2411 vdd.n2407 878.823
R1525 vdd.n2411 vdd.n2403 878.823
R1526 vdd.n2413 vdd.n2409 878.823
R1527 vdd.n2423 vdd.n2413 878.823
R1528 vdd.n2480 vdd.n2452 878.823
R1529 vdd.n2487 vdd.n2452 878.823
R1530 vdd.n2459 vdd.n2455 878.823
R1531 vdd.n2459 vdd.n2451 878.823
R1532 vdd.n2461 vdd.n2457 878.823
R1533 vdd.n2471 vdd.n2461 878.823
R1534 vdd.n2597 vdd.n2589 878.823
R1535 vdd.n2598 vdd.n2597 878.823
R1536 vdd.n2610 vdd.n2600 878.823
R1537 vdd.n2600 vdd.n2596 878.823
R1538 vdd.n2624 vdd.n2590 878.823
R1539 vdd.n2624 vdd.n2623 878.823
R1540 vdd.n2551 vdd.n2543 878.823
R1541 vdd.n2552 vdd.n2551 878.823
R1542 vdd.n2564 vdd.n2554 878.823
R1543 vdd.n2554 vdd.n2550 878.823
R1544 vdd.n2578 vdd.n2544 878.823
R1545 vdd.n2578 vdd.n2577 878.823
R1546 vdd.n2644 vdd.n2636 878.823
R1547 vdd.n2645 vdd.n2644 878.823
R1548 vdd.n2657 vdd.n2647 878.823
R1549 vdd.n2647 vdd.n2643 878.823
R1550 vdd.n2671 vdd.n2637 878.823
R1551 vdd.n2671 vdd.n2670 878.823
R1552 vdd.n2692 vdd.n2684 878.823
R1553 vdd.n2693 vdd.n2692 878.823
R1554 vdd.n2705 vdd.n2695 878.823
R1555 vdd.n2695 vdd.n2691 878.823
R1556 vdd.n2719 vdd.n2685 878.823
R1557 vdd.n2719 vdd.n2718 878.823
R1558 vdd.n2738 vdd.n2730 878.823
R1559 vdd.n2739 vdd.n2738 878.823
R1560 vdd.n2751 vdd.n2741 878.823
R1561 vdd.n2741 vdd.n2737 878.823
R1562 vdd.n2765 vdd.n2731 878.823
R1563 vdd.n2765 vdd.n2764 878.823
R1564 vdd.n997 vdd.n994 878.823
R1565 vdd.n998 vdd.n997 878.823
R1566 vdd.n1002 vdd.n993 878.823
R1567 vdd.n1003 vdd.n1002 878.823
R1568 vdd.n1024 vdd.n1023 878.823
R1569 vdd.n1023 vdd.n988 878.823
R1570 vdd.n2880 vdd.n2872 878.823
R1571 vdd.n2881 vdd.n2880 878.823
R1572 vdd.n2893 vdd.n2883 878.823
R1573 vdd.n2883 vdd.n2879 878.823
R1574 vdd.n2907 vdd.n2873 878.823
R1575 vdd.n2907 vdd.n2906 878.823
R1576 vdd.n2833 vdd.n2825 878.823
R1577 vdd.n2834 vdd.n2833 878.823
R1578 vdd.n2846 vdd.n2836 878.823
R1579 vdd.n2836 vdd.n2832 878.823
R1580 vdd.n2860 vdd.n2826 878.823
R1581 vdd.n2860 vdd.n2859 878.823
R1582 vdd.n2787 vdd.n2779 878.823
R1583 vdd.n2788 vdd.n2787 878.823
R1584 vdd.n2800 vdd.n2790 878.823
R1585 vdd.n2790 vdd.n2786 878.823
R1586 vdd.n2814 vdd.n2780 878.823
R1587 vdd.n2814 vdd.n2813 878.823
R1588 vdd.n2927 vdd.n2919 878.823
R1589 vdd.n2928 vdd.n2927 878.823
R1590 vdd.n2940 vdd.n2930 878.823
R1591 vdd.n2930 vdd.n2926 878.823
R1592 vdd.n2954 vdd.n2920 878.823
R1593 vdd.n2954 vdd.n2953 878.823
R1594 vdd.n2975 vdd.n2967 878.823
R1595 vdd.n2976 vdd.n2975 878.823
R1596 vdd.n2988 vdd.n2978 878.823
R1597 vdd.n2978 vdd.n2974 878.823
R1598 vdd.n3002 vdd.n2968 878.823
R1599 vdd.n3002 vdd.n3001 878.823
R1600 vdd.n3021 vdd.n3013 878.823
R1601 vdd.n3022 vdd.n3021 878.823
R1602 vdd.n3034 vdd.n3024 878.823
R1603 vdd.n3024 vdd.n3020 878.823
R1604 vdd.n3048 vdd.n3014 878.823
R1605 vdd.n3048 vdd.n3047 878.823
R1606 vdd.n3115 vdd.n3107 878.823
R1607 vdd.n3116 vdd.n3115 878.823
R1608 vdd.n3128 vdd.n3118 878.823
R1609 vdd.n3118 vdd.n3114 878.823
R1610 vdd.n3142 vdd.n3108 878.823
R1611 vdd.n3142 vdd.n3141 878.823
R1612 vdd.n3069 vdd.n3061 878.823
R1613 vdd.n3070 vdd.n3069 878.823
R1614 vdd.n3082 vdd.n3072 878.823
R1615 vdd.n3072 vdd.n3068 878.823
R1616 vdd.n3096 vdd.n3062 878.823
R1617 vdd.n3096 vdd.n3095 878.823
R1618 vdd.n3162 vdd.n3154 878.823
R1619 vdd.n3163 vdd.n3162 878.823
R1620 vdd.n3175 vdd.n3165 878.823
R1621 vdd.n3165 vdd.n3161 878.823
R1622 vdd.n3189 vdd.n3155 878.823
R1623 vdd.n3189 vdd.n3188 878.823
R1624 vdd.n3210 vdd.n3202 878.823
R1625 vdd.n3211 vdd.n3210 878.823
R1626 vdd.n3223 vdd.n3213 878.823
R1627 vdd.n3213 vdd.n3209 878.823
R1628 vdd.n3237 vdd.n3203 878.823
R1629 vdd.n3237 vdd.n3236 878.823
R1630 vdd.n3256 vdd.n3248 878.823
R1631 vdd.n3257 vdd.n3256 878.823
R1632 vdd.n3269 vdd.n3259 878.823
R1633 vdd.n3259 vdd.n3255 878.823
R1634 vdd.n3283 vdd.n3249 878.823
R1635 vdd.n3283 vdd.n3282 878.823
R1636 vdd.n761 vdd.n758 878.823
R1637 vdd.n762 vdd.n761 878.823
R1638 vdd.n766 vdd.n757 878.823
R1639 vdd.n767 vdd.n766 878.823
R1640 vdd.n788 vdd.n787 878.823
R1641 vdd.n787 vdd.n752 878.823
R1642 vdd.n3351 vdd.n3343 878.823
R1643 vdd.n3352 vdd.n3351 878.823
R1644 vdd.n3364 vdd.n3354 878.823
R1645 vdd.n3354 vdd.n3350 878.823
R1646 vdd.n3378 vdd.n3344 878.823
R1647 vdd.n3378 vdd.n3377 878.823
R1648 vdd.n3305 vdd.n3297 878.823
R1649 vdd.n3306 vdd.n3305 878.823
R1650 vdd.n3318 vdd.n3308 878.823
R1651 vdd.n3308 vdd.n3304 878.823
R1652 vdd.n3332 vdd.n3298 878.823
R1653 vdd.n3332 vdd.n3331 878.823
R1654 vdd.n3398 vdd.n3390 878.823
R1655 vdd.n3399 vdd.n3398 878.823
R1656 vdd.n3411 vdd.n3401 878.823
R1657 vdd.n3401 vdd.n3397 878.823
R1658 vdd.n3425 vdd.n3391 878.823
R1659 vdd.n3425 vdd.n3424 878.823
R1660 vdd.n3446 vdd.n3438 878.823
R1661 vdd.n3447 vdd.n3446 878.823
R1662 vdd.n3459 vdd.n3449 878.823
R1663 vdd.n3449 vdd.n3445 878.823
R1664 vdd.n3473 vdd.n3439 878.823
R1665 vdd.n3473 vdd.n3472 878.823
R1666 vdd.n3492 vdd.n3484 878.823
R1667 vdd.n3493 vdd.n3492 878.823
R1668 vdd.n3505 vdd.n3495 878.823
R1669 vdd.n3495 vdd.n3491 878.823
R1670 vdd.n3519 vdd.n3485 878.823
R1671 vdd.n3519 vdd.n3518 878.823
R1672 vdd.n574 vdd.n566 878.823
R1673 vdd.n575 vdd.n574 878.823
R1674 vdd.n587 vdd.n577 878.823
R1675 vdd.n577 vdd.n573 878.823
R1676 vdd.n601 vdd.n567 878.823
R1677 vdd.n601 vdd.n600 878.823
R1678 vdd.n3587 vdd.n3579 878.823
R1679 vdd.n3588 vdd.n3587 878.823
R1680 vdd.n3600 vdd.n3590 878.823
R1681 vdd.n3590 vdd.n3586 878.823
R1682 vdd.n3614 vdd.n3580 878.823
R1683 vdd.n3614 vdd.n3613 878.823
R1684 vdd.n3541 vdd.n3533 878.823
R1685 vdd.n3542 vdd.n3541 878.823
R1686 vdd.n3554 vdd.n3544 878.823
R1687 vdd.n3544 vdd.n3540 878.823
R1688 vdd.n3568 vdd.n3534 878.823
R1689 vdd.n3568 vdd.n3567 878.823
R1690 vdd.n6601 vdd.n6593 878.823
R1691 vdd.n6602 vdd.n6601 878.823
R1692 vdd.n6614 vdd.n6604 878.823
R1693 vdd.n6604 vdd.n6600 878.823
R1694 vdd.n6628 vdd.n6594 878.823
R1695 vdd.n6628 vdd.n6627 878.823
R1696 vdd.n6555 vdd.n6547 878.823
R1697 vdd.n6556 vdd.n6555 878.823
R1698 vdd.n6568 vdd.n6558 878.823
R1699 vdd.n6558 vdd.n6554 878.823
R1700 vdd.n6582 vdd.n6548 878.823
R1701 vdd.n6582 vdd.n6581 878.823
R1702 vdd.n9615 vdd.n9607 878.823
R1703 vdd.n9616 vdd.n9615 878.823
R1704 vdd.n9628 vdd.n9618 878.823
R1705 vdd.n9618 vdd.n9614 878.823
R1706 vdd.n9642 vdd.n9608 878.823
R1707 vdd.n9642 vdd.n9641 878.823
R1708 vdd.n9569 vdd.n9561 878.823
R1709 vdd.n9570 vdd.n9569 878.823
R1710 vdd.n9582 vdd.n9572 878.823
R1711 vdd.n9572 vdd.n9568 878.823
R1712 vdd.n9596 vdd.n9562 878.823
R1713 vdd.n9596 vdd.n9595 878.823
R1714 vdd.n9661 vdd.n9653 878.823
R1715 vdd.n9662 vdd.n9661 878.823
R1716 vdd.n9674 vdd.n9664 878.823
R1717 vdd.n9664 vdd.n9660 878.823
R1718 vdd.n9688 vdd.n9654 878.823
R1719 vdd.n9688 vdd.n9687 878.823
R1720 vdd.n9707 vdd.n9699 878.823
R1721 vdd.n9708 vdd.n9707 878.823
R1722 vdd.n9720 vdd.n9710 878.823
R1723 vdd.n9710 vdd.n9706 878.823
R1724 vdd.n9734 vdd.n9700 878.823
R1725 vdd.n9734 vdd.n9733 878.823
R1726 vdd.n9805 vdd.n9797 878.823
R1727 vdd.n9806 vdd.n9805 878.823
R1728 vdd.n9818 vdd.n9808 878.823
R1729 vdd.n9808 vdd.n9804 878.823
R1730 vdd.n9832 vdd.n9798 878.823
R1731 vdd.n9832 vdd.n9831 878.823
R1732 vdd.n9851 vdd.n9843 878.823
R1733 vdd.n9852 vdd.n9851 878.823
R1734 vdd.n9864 vdd.n9854 878.823
R1735 vdd.n9854 vdd.n9850 878.823
R1736 vdd.n9878 vdd.n9844 878.823
R1737 vdd.n9878 vdd.n9877 878.823
R1738 vdd.n9897 vdd.n9889 878.823
R1739 vdd.n9898 vdd.n9897 878.823
R1740 vdd.n9910 vdd.n9900 878.823
R1741 vdd.n9900 vdd.n9896 878.823
R1742 vdd.n9924 vdd.n9890 878.823
R1743 vdd.n9924 vdd.n9923 878.823
R1744 vdd.n9943 vdd.n9935 878.823
R1745 vdd.n9944 vdd.n9943 878.823
R1746 vdd.n9956 vdd.n9946 878.823
R1747 vdd.n9946 vdd.n9942 878.823
R1748 vdd.n9970 vdd.n9936 878.823
R1749 vdd.n9970 vdd.n9969 878.823
R1750 vdd.n10041 vdd.n10033 878.823
R1751 vdd.n10042 vdd.n10041 878.823
R1752 vdd.n10054 vdd.n10044 878.823
R1753 vdd.n10044 vdd.n10040 878.823
R1754 vdd.n10068 vdd.n10034 878.823
R1755 vdd.n10068 vdd.n10067 878.823
R1756 vdd.n57 vdd.n49 878.823
R1757 vdd.n58 vdd.n57 878.823
R1758 vdd.n70 vdd.n60 878.823
R1759 vdd.n60 vdd.n56 878.823
R1760 vdd.n84 vdd.n50 878.823
R1761 vdd.n84 vdd.n83 878.823
R1762 vdd.n11 vdd.n3 878.823
R1763 vdd.n12 vdd.n11 878.823
R1764 vdd.n24 vdd.n14 878.823
R1765 vdd.n14 vdd.n10 878.823
R1766 vdd.n38 vdd.n4 878.823
R1767 vdd.n38 vdd.n37 878.823
R1768 vdd.n10087 vdd.n10079 878.823
R1769 vdd.n10088 vdd.n10087 878.823
R1770 vdd.n10100 vdd.n10090 878.823
R1771 vdd.n10090 vdd.n10086 878.823
R1772 vdd.n10114 vdd.n10080 878.823
R1773 vdd.n10114 vdd.n10113 878.823
R1774 vdd.n10135 vdd.n10127 878.823
R1775 vdd.n10136 vdd.n10135 878.823
R1776 vdd.n10148 vdd.n10138 878.823
R1777 vdd.n10138 vdd.n10134 878.823
R1778 vdd.n10162 vdd.n10128 878.823
R1779 vdd.n10162 vdd.n10161 878.823
R1780 vdd.n10181 vdd.n10173 878.823
R1781 vdd.n10182 vdd.n10181 878.823
R1782 vdd.n10194 vdd.n10184 878.823
R1783 vdd.n10184 vdd.n10180 878.823
R1784 vdd.n10208 vdd.n10174 878.823
R1785 vdd.n10208 vdd.n10207 878.823
R1786 vdd.n9992 vdd.n9989 878.823
R1787 vdd.n9993 vdd.n9992 878.823
R1788 vdd.n9997 vdd.n9988 878.823
R1789 vdd.n9998 vdd.n9997 878.823
R1790 vdd.n10019 vdd.n10018 878.823
R1791 vdd.n10018 vdd.n9983 878.823
R1792 vdd.n10323 vdd.n10315 878.823
R1793 vdd.n10324 vdd.n10323 878.823
R1794 vdd.n10336 vdd.n10326 878.823
R1795 vdd.n10326 vdd.n10322 878.823
R1796 vdd.n10350 vdd.n10316 878.823
R1797 vdd.n10350 vdd.n10349 878.823
R1798 vdd.n10276 vdd.n10268 878.823
R1799 vdd.n10277 vdd.n10276 878.823
R1800 vdd.n10289 vdd.n10279 878.823
R1801 vdd.n10279 vdd.n10275 878.823
R1802 vdd.n10303 vdd.n10269 878.823
R1803 vdd.n10303 vdd.n10302 878.823
R1804 vdd.n10230 vdd.n10222 878.823
R1805 vdd.n10231 vdd.n10230 878.823
R1806 vdd.n10243 vdd.n10233 878.823
R1807 vdd.n10233 vdd.n10229 878.823
R1808 vdd.n10257 vdd.n10223 878.823
R1809 vdd.n10257 vdd.n10256 878.823
R1810 vdd.n10370 vdd.n10362 878.823
R1811 vdd.n10371 vdd.n10370 878.823
R1812 vdd.n10383 vdd.n10373 878.823
R1813 vdd.n10373 vdd.n10369 878.823
R1814 vdd.n10397 vdd.n10363 878.823
R1815 vdd.n10397 vdd.n10396 878.823
R1816 vdd.n10418 vdd.n10410 878.823
R1817 vdd.n10419 vdd.n10418 878.823
R1818 vdd.n10431 vdd.n10421 878.823
R1819 vdd.n10421 vdd.n10417 878.823
R1820 vdd.n10445 vdd.n10411 878.823
R1821 vdd.n10445 vdd.n10444 878.823
R1822 vdd.n10464 vdd.n10456 878.823
R1823 vdd.n10465 vdd.n10464 878.823
R1824 vdd.n10477 vdd.n10467 878.823
R1825 vdd.n10467 vdd.n10463 878.823
R1826 vdd.n10491 vdd.n10457 878.823
R1827 vdd.n10491 vdd.n10490 878.823
R1828 vdd.n10558 vdd.n10550 878.823
R1829 vdd.n10559 vdd.n10558 878.823
R1830 vdd.n10571 vdd.n10561 878.823
R1831 vdd.n10561 vdd.n10557 878.823
R1832 vdd.n10585 vdd.n10551 878.823
R1833 vdd.n10585 vdd.n10584 878.823
R1834 vdd.n10512 vdd.n10504 878.823
R1835 vdd.n10513 vdd.n10512 878.823
R1836 vdd.n10525 vdd.n10515 878.823
R1837 vdd.n10515 vdd.n10511 878.823
R1838 vdd.n10539 vdd.n10505 878.823
R1839 vdd.n10539 vdd.n10538 878.823
R1840 vdd.n10605 vdd.n10597 878.823
R1841 vdd.n10606 vdd.n10605 878.823
R1842 vdd.n10618 vdd.n10608 878.823
R1843 vdd.n10608 vdd.n10604 878.823
R1844 vdd.n10632 vdd.n10598 878.823
R1845 vdd.n10632 vdd.n10631 878.823
R1846 vdd.n10653 vdd.n10645 878.823
R1847 vdd.n10654 vdd.n10653 878.823
R1848 vdd.n10666 vdd.n10656 878.823
R1849 vdd.n10656 vdd.n10652 878.823
R1850 vdd.n10680 vdd.n10646 878.823
R1851 vdd.n10680 vdd.n10679 878.823
R1852 vdd.n10699 vdd.n10691 878.823
R1853 vdd.n10700 vdd.n10699 878.823
R1854 vdd.n10712 vdd.n10702 878.823
R1855 vdd.n10702 vdd.n10698 878.823
R1856 vdd.n10726 vdd.n10692 878.823
R1857 vdd.n10726 vdd.n10725 878.823
R1858 vdd.n9756 vdd.n9753 878.823
R1859 vdd.n9757 vdd.n9756 878.823
R1860 vdd.n9761 vdd.n9752 878.823
R1861 vdd.n9762 vdd.n9761 878.823
R1862 vdd.n9783 vdd.n9782 878.823
R1863 vdd.n9782 vdd.n9747 878.823
R1864 vdd.n10794 vdd.n10786 878.823
R1865 vdd.n10795 vdd.n10794 878.823
R1866 vdd.n10807 vdd.n10797 878.823
R1867 vdd.n10797 vdd.n10793 878.823
R1868 vdd.n10821 vdd.n10787 878.823
R1869 vdd.n10821 vdd.n10820 878.823
R1870 vdd.n10748 vdd.n10740 878.823
R1871 vdd.n10749 vdd.n10748 878.823
R1872 vdd.n10761 vdd.n10751 878.823
R1873 vdd.n10751 vdd.n10747 878.823
R1874 vdd.n10775 vdd.n10741 878.823
R1875 vdd.n10775 vdd.n10774 878.823
R1876 vdd.n10841 vdd.n10833 878.823
R1877 vdd.n10842 vdd.n10841 878.823
R1878 vdd.n10854 vdd.n10844 878.823
R1879 vdd.n10844 vdd.n10840 878.823
R1880 vdd.n10868 vdd.n10834 878.823
R1881 vdd.n10868 vdd.n10867 878.823
R1882 vdd.n10889 vdd.n10881 878.823
R1883 vdd.n10890 vdd.n10889 878.823
R1884 vdd.n10902 vdd.n10892 878.823
R1885 vdd.n10892 vdd.n10888 878.823
R1886 vdd.n10916 vdd.n10882 878.823
R1887 vdd.n10916 vdd.n10915 878.823
R1888 vdd.n10935 vdd.n10927 878.823
R1889 vdd.n10936 vdd.n10935 878.823
R1890 vdd.n10948 vdd.n10938 878.823
R1891 vdd.n10938 vdd.n10934 878.823
R1892 vdd.n10962 vdd.n10928 878.823
R1893 vdd.n10962 vdd.n10961 878.823
R1894 vdd.n11005 vdd.n10977 878.823
R1895 vdd.n11012 vdd.n10977 878.823
R1896 vdd.n10984 vdd.n10980 878.823
R1897 vdd.n10984 vdd.n10976 878.823
R1898 vdd.n10986 vdd.n10982 878.823
R1899 vdd.n10996 vdd.n10986 878.823
R1900 vdd.n11050 vdd.n11022 878.823
R1901 vdd.n11057 vdd.n11022 878.823
R1902 vdd.n11029 vdd.n11025 878.823
R1903 vdd.n11029 vdd.n11021 878.823
R1904 vdd.n11031 vdd.n11027 878.823
R1905 vdd.n11041 vdd.n11031 878.823
R1906 vdd.n11100 vdd.n11072 878.823
R1907 vdd.n11107 vdd.n11072 878.823
R1908 vdd.n11079 vdd.n11075 878.823
R1909 vdd.n11079 vdd.n11071 878.823
R1910 vdd.n11081 vdd.n11077 878.823
R1911 vdd.n11091 vdd.n11081 878.823
R1912 vdd.n11146 vdd.n11118 878.823
R1913 vdd.n11153 vdd.n11118 878.823
R1914 vdd.n11125 vdd.n11121 878.823
R1915 vdd.n11125 vdd.n11117 878.823
R1916 vdd.n11127 vdd.n11123 878.823
R1917 vdd.n11137 vdd.n11127 878.823
R1918 vdd.n11194 vdd.n11166 878.823
R1919 vdd.n11201 vdd.n11166 878.823
R1920 vdd.n11173 vdd.n11169 878.823
R1921 vdd.n11173 vdd.n11165 878.823
R1922 vdd.n11175 vdd.n11171 878.823
R1923 vdd.n11185 vdd.n11175 878.823
R1924 vdd.n450 vdd.n431 878.823
R1925 vdd.n457 vdd.n431 878.823
R1926 vdd.n436 vdd.n435 878.823
R1927 vdd.n435 vdd.n427 878.823
R1928 vdd.n442 vdd.n425 878.823
R1929 vdd.n464 vdd.n425 878.823
R1930 vdd.n11241 vdd.n11213 878.823
R1931 vdd.n11248 vdd.n11213 878.823
R1932 vdd.n11220 vdd.n11216 878.823
R1933 vdd.n11220 vdd.n11212 878.823
R1934 vdd.n11222 vdd.n11218 878.823
R1935 vdd.n11232 vdd.n11222 878.823
R1936 vdd.n11286 vdd.n11258 878.823
R1937 vdd.n11293 vdd.n11258 878.823
R1938 vdd.n11265 vdd.n11261 878.823
R1939 vdd.n11265 vdd.n11257 878.823
R1940 vdd.n11267 vdd.n11263 878.823
R1941 vdd.n11277 vdd.n11267 878.823
R1942 vdd.n11332 vdd.n11304 878.823
R1943 vdd.n11339 vdd.n11304 878.823
R1944 vdd.n11311 vdd.n11307 878.823
R1945 vdd.n11311 vdd.n11303 878.823
R1946 vdd.n11313 vdd.n11309 878.823
R1947 vdd.n11323 vdd.n11313 878.823
R1948 vdd.n11383 vdd.n11355 878.823
R1949 vdd.n11390 vdd.n11355 878.823
R1950 vdd.n11362 vdd.n11358 878.823
R1951 vdd.n11362 vdd.n11354 878.823
R1952 vdd.n11364 vdd.n11360 878.823
R1953 vdd.n11374 vdd.n11364 878.823
R1954 vdd.n11429 vdd.n11401 878.823
R1955 vdd.n11436 vdd.n11401 878.823
R1956 vdd.n11408 vdd.n11404 878.823
R1957 vdd.n11408 vdd.n11400 878.823
R1958 vdd.n11410 vdd.n11406 878.823
R1959 vdd.n11420 vdd.n11410 878.823
R1960 vdd.n11477 vdd.n11449 878.823
R1961 vdd.n11484 vdd.n11449 878.823
R1962 vdd.n11456 vdd.n11452 878.823
R1963 vdd.n11456 vdd.n11448 878.823
R1964 vdd.n11458 vdd.n11454 878.823
R1965 vdd.n11468 vdd.n11458 878.823
R1966 vdd.n11523 vdd.n11495 878.823
R1967 vdd.n11530 vdd.n11495 878.823
R1968 vdd.n11502 vdd.n11498 878.823
R1969 vdd.n11502 vdd.n11494 878.823
R1970 vdd.n11504 vdd.n11500 878.823
R1971 vdd.n11514 vdd.n11504 878.823
R1972 vdd.n11568 vdd.n11540 878.823
R1973 vdd.n11575 vdd.n11540 878.823
R1974 vdd.n11547 vdd.n11543 878.823
R1975 vdd.n11547 vdd.n11539 878.823
R1976 vdd.n11549 vdd.n11545 878.823
R1977 vdd.n11559 vdd.n11549 878.823
R1978 vdd.n11618 vdd.n11590 878.823
R1979 vdd.n11625 vdd.n11590 878.823
R1980 vdd.n11597 vdd.n11593 878.823
R1981 vdd.n11597 vdd.n11589 878.823
R1982 vdd.n11599 vdd.n11595 878.823
R1983 vdd.n11609 vdd.n11599 878.823
R1984 vdd.n11664 vdd.n11636 878.823
R1985 vdd.n11671 vdd.n11636 878.823
R1986 vdd.n11643 vdd.n11639 878.823
R1987 vdd.n11643 vdd.n11635 878.823
R1988 vdd.n11645 vdd.n11641 878.823
R1989 vdd.n11655 vdd.n11645 878.823
R1990 vdd.n11712 vdd.n11684 878.823
R1991 vdd.n11719 vdd.n11684 878.823
R1992 vdd.n11691 vdd.n11687 878.823
R1993 vdd.n11691 vdd.n11683 878.823
R1994 vdd.n11693 vdd.n11689 878.823
R1995 vdd.n11703 vdd.n11693 878.823
R1996 vdd.n215 vdd.n196 878.823
R1997 vdd.n222 vdd.n196 878.823
R1998 vdd.n201 vdd.n200 878.823
R1999 vdd.n200 vdd.n192 878.823
R2000 vdd.n207 vdd.n190 878.823
R2001 vdd.n229 vdd.n190 878.823
R2002 vdd.n11759 vdd.n11731 878.823
R2003 vdd.n11766 vdd.n11731 878.823
R2004 vdd.n11738 vdd.n11734 878.823
R2005 vdd.n11738 vdd.n11730 878.823
R2006 vdd.n11740 vdd.n11736 878.823
R2007 vdd.n11750 vdd.n11740 878.823
R2008 vdd.n11804 vdd.n11776 878.823
R2009 vdd.n11811 vdd.n11776 878.823
R2010 vdd.n11783 vdd.n11779 878.823
R2011 vdd.n11783 vdd.n11775 878.823
R2012 vdd.n11785 vdd.n11781 878.823
R2013 vdd.n11795 vdd.n11785 878.823
R2014 vdd.n11854 vdd.n11826 878.823
R2015 vdd.n11861 vdd.n11826 878.823
R2016 vdd.n11833 vdd.n11829 878.823
R2017 vdd.n11833 vdd.n11825 878.823
R2018 vdd.n11835 vdd.n11831 878.823
R2019 vdd.n11845 vdd.n11835 878.823
R2020 vdd.n11900 vdd.n11872 878.823
R2021 vdd.n11907 vdd.n11872 878.823
R2022 vdd.n11879 vdd.n11875 878.823
R2023 vdd.n11879 vdd.n11871 878.823
R2024 vdd.n11881 vdd.n11877 878.823
R2025 vdd.n11891 vdd.n11881 878.823
R2026 vdd.n11948 vdd.n11920 878.823
R2027 vdd.n11955 vdd.n11920 878.823
R2028 vdd.n11927 vdd.n11923 878.823
R2029 vdd.n11927 vdd.n11919 878.823
R2030 vdd.n11929 vdd.n11925 878.823
R2031 vdd.n11939 vdd.n11929 878.823
R2032 vdd.n11982 vdd.n11976 681.178
R2033 vdd.n12002 vdd.n11995 681.178
R2034 vdd.n12002 vdd.n11996 681.178
R2035 vdd.n11981 vdd.n11977 681.178
R2036 vdd.n11981 vdd.n11978 681.178
R2037 vdd.n12001 vdd.n11997 681.178
R2038 vdd.n111 vdd.n104 681.178
R2039 vdd.n120 vdd.n104 681.178
R2040 vdd.n120 vdd.n102 681.178
R2041 vdd.n126 vdd.n102 681.178
R2042 vdd.n127 vdd.n126 681.178
R2043 vdd.n129 vdd.n127 681.178
R2044 vdd.n118 vdd.n117 681.178
R2045 vdd.n119 vdd.n118 681.178
R2046 vdd.n119 vdd.n98 681.178
R2047 vdd.n135 vdd.n98 681.178
R2048 vdd.n135 vdd.n134 681.178
R2049 vdd.n134 vdd.n133 681.178
R2050 vdd.n157 vdd.n150 681.178
R2051 vdd.n166 vdd.n150 681.178
R2052 vdd.n166 vdd.n148 681.178
R2053 vdd.n172 vdd.n148 681.178
R2054 vdd.n173 vdd.n172 681.178
R2055 vdd.n175 vdd.n173 681.178
R2056 vdd.n164 vdd.n163 681.178
R2057 vdd.n165 vdd.n164 681.178
R2058 vdd.n165 vdd.n144 681.178
R2059 vdd.n181 vdd.n144 681.178
R2060 vdd.n181 vdd.n180 681.178
R2061 vdd.n180 vdd.n179 681.178
R2062 vdd.n254 vdd.n247 681.178
R2063 vdd.n263 vdd.n247 681.178
R2064 vdd.n263 vdd.n245 681.178
R2065 vdd.n269 vdd.n245 681.178
R2066 vdd.n270 vdd.n269 681.178
R2067 vdd.n272 vdd.n270 681.178
R2068 vdd.n261 vdd.n260 681.178
R2069 vdd.n262 vdd.n261 681.178
R2070 vdd.n262 vdd.n241 681.178
R2071 vdd.n278 vdd.n241 681.178
R2072 vdd.n278 vdd.n277 681.178
R2073 vdd.n277 vdd.n276 681.178
R2074 vdd.n300 vdd.n293 681.178
R2075 vdd.n309 vdd.n293 681.178
R2076 vdd.n309 vdd.n291 681.178
R2077 vdd.n315 vdd.n291 681.178
R2078 vdd.n316 vdd.n315 681.178
R2079 vdd.n318 vdd.n316 681.178
R2080 vdd.n307 vdd.n306 681.178
R2081 vdd.n308 vdd.n307 681.178
R2082 vdd.n308 vdd.n287 681.178
R2083 vdd.n324 vdd.n287 681.178
R2084 vdd.n324 vdd.n323 681.178
R2085 vdd.n323 vdd.n322 681.178
R2086 vdd.n346 vdd.n339 681.178
R2087 vdd.n355 vdd.n339 681.178
R2088 vdd.n355 vdd.n337 681.178
R2089 vdd.n361 vdd.n337 681.178
R2090 vdd.n362 vdd.n361 681.178
R2091 vdd.n364 vdd.n362 681.178
R2092 vdd.n353 vdd.n352 681.178
R2093 vdd.n354 vdd.n353 681.178
R2094 vdd.n354 vdd.n333 681.178
R2095 vdd.n370 vdd.n333 681.178
R2096 vdd.n370 vdd.n369 681.178
R2097 vdd.n369 vdd.n368 681.178
R2098 vdd.n392 vdd.n385 681.178
R2099 vdd.n401 vdd.n385 681.178
R2100 vdd.n401 vdd.n383 681.178
R2101 vdd.n407 vdd.n383 681.178
R2102 vdd.n408 vdd.n407 681.178
R2103 vdd.n410 vdd.n408 681.178
R2104 vdd.n399 vdd.n398 681.178
R2105 vdd.n400 vdd.n399 681.178
R2106 vdd.n400 vdd.n379 681.178
R2107 vdd.n416 vdd.n379 681.178
R2108 vdd.n416 vdd.n415 681.178
R2109 vdd.n415 vdd.n414 681.178
R2110 vdd.n489 vdd.n482 681.178
R2111 vdd.n498 vdd.n482 681.178
R2112 vdd.n498 vdd.n480 681.178
R2113 vdd.n504 vdd.n480 681.178
R2114 vdd.n505 vdd.n504 681.178
R2115 vdd.n507 vdd.n505 681.178
R2116 vdd.n496 vdd.n495 681.178
R2117 vdd.n497 vdd.n496 681.178
R2118 vdd.n497 vdd.n476 681.178
R2119 vdd.n513 vdd.n476 681.178
R2120 vdd.n513 vdd.n512 681.178
R2121 vdd.n512 vdd.n511 681.178
R2122 vdd.n535 vdd.n528 681.178
R2123 vdd.n544 vdd.n528 681.178
R2124 vdd.n544 vdd.n526 681.178
R2125 vdd.n550 vdd.n526 681.178
R2126 vdd.n551 vdd.n550 681.178
R2127 vdd.n553 vdd.n551 681.178
R2128 vdd.n542 vdd.n541 681.178
R2129 vdd.n543 vdd.n542 681.178
R2130 vdd.n543 vdd.n522 681.178
R2131 vdd.n559 vdd.n522 681.178
R2132 vdd.n559 vdd.n558 681.178
R2133 vdd.n558 vdd.n557 681.178
R2134 vdd.n6707 vdd.n6706 681.178
R2135 vdd.n6708 vdd.n6707 681.178
R2136 vdd.n6708 vdd.n6686 681.178
R2137 vdd.n6723 vdd.n6686 681.178
R2138 vdd.n6723 vdd.n6687 681.178
R2139 vdd.n6715 vdd.n6687 681.178
R2140 vdd.n6700 vdd.n6693 681.178
R2141 vdd.n6709 vdd.n6693 681.178
R2142 vdd.n6709 vdd.n6695 681.178
R2143 vdd.n6695 vdd.n6689 681.178
R2144 vdd.n6720 vdd.n6689 681.178
R2145 vdd.n6720 vdd.n6719 681.178
R2146 vdd.n6753 vdd.n6752 681.178
R2147 vdd.n6754 vdd.n6753 681.178
R2148 vdd.n6754 vdd.n6732 681.178
R2149 vdd.n6769 vdd.n6732 681.178
R2150 vdd.n6769 vdd.n6733 681.178
R2151 vdd.n6761 vdd.n6733 681.178
R2152 vdd.n6746 vdd.n6739 681.178
R2153 vdd.n6755 vdd.n6739 681.178
R2154 vdd.n6755 vdd.n6741 681.178
R2155 vdd.n6741 vdd.n6735 681.178
R2156 vdd.n6766 vdd.n6735 681.178
R2157 vdd.n6766 vdd.n6765 681.178
R2158 vdd.n6851 vdd.n6850 681.178
R2159 vdd.n6852 vdd.n6851 681.178
R2160 vdd.n6852 vdd.n6830 681.178
R2161 vdd.n6867 vdd.n6830 681.178
R2162 vdd.n6867 vdd.n6831 681.178
R2163 vdd.n6859 vdd.n6831 681.178
R2164 vdd.n6844 vdd.n6837 681.178
R2165 vdd.n6853 vdd.n6837 681.178
R2166 vdd.n6853 vdd.n6839 681.178
R2167 vdd.n6839 vdd.n6833 681.178
R2168 vdd.n6864 vdd.n6833 681.178
R2169 vdd.n6864 vdd.n6863 681.178
R2170 vdd.n6897 vdd.n6896 681.178
R2171 vdd.n6898 vdd.n6897 681.178
R2172 vdd.n6898 vdd.n6876 681.178
R2173 vdd.n6913 vdd.n6876 681.178
R2174 vdd.n6913 vdd.n6877 681.178
R2175 vdd.n6905 vdd.n6877 681.178
R2176 vdd.n6890 vdd.n6883 681.178
R2177 vdd.n6899 vdd.n6883 681.178
R2178 vdd.n6899 vdd.n6885 681.178
R2179 vdd.n6885 vdd.n6879 681.178
R2180 vdd.n6910 vdd.n6879 681.178
R2181 vdd.n6910 vdd.n6909 681.178
R2182 vdd.n6943 vdd.n6942 681.178
R2183 vdd.n6944 vdd.n6943 681.178
R2184 vdd.n6944 vdd.n6922 681.178
R2185 vdd.n6959 vdd.n6922 681.178
R2186 vdd.n6959 vdd.n6923 681.178
R2187 vdd.n6951 vdd.n6923 681.178
R2188 vdd.n6936 vdd.n6929 681.178
R2189 vdd.n6945 vdd.n6929 681.178
R2190 vdd.n6945 vdd.n6931 681.178
R2191 vdd.n6931 vdd.n6925 681.178
R2192 vdd.n6956 vdd.n6925 681.178
R2193 vdd.n6956 vdd.n6955 681.178
R2194 vdd.n6989 vdd.n6988 681.178
R2195 vdd.n6990 vdd.n6989 681.178
R2196 vdd.n6990 vdd.n6968 681.178
R2197 vdd.n7005 vdd.n6968 681.178
R2198 vdd.n7005 vdd.n6969 681.178
R2199 vdd.n6997 vdd.n6969 681.178
R2200 vdd.n6982 vdd.n6975 681.178
R2201 vdd.n6991 vdd.n6975 681.178
R2202 vdd.n6991 vdd.n6977 681.178
R2203 vdd.n6977 vdd.n6971 681.178
R2204 vdd.n7002 vdd.n6971 681.178
R2205 vdd.n7002 vdd.n7001 681.178
R2206 vdd.n7087 vdd.n7086 681.178
R2207 vdd.n7088 vdd.n7087 681.178
R2208 vdd.n7088 vdd.n7066 681.178
R2209 vdd.n7103 vdd.n7066 681.178
R2210 vdd.n7103 vdd.n7067 681.178
R2211 vdd.n7095 vdd.n7067 681.178
R2212 vdd.n7080 vdd.n7073 681.178
R2213 vdd.n7089 vdd.n7073 681.178
R2214 vdd.n7089 vdd.n7075 681.178
R2215 vdd.n7075 vdd.n7069 681.178
R2216 vdd.n7100 vdd.n7069 681.178
R2217 vdd.n7100 vdd.n7099 681.178
R2218 vdd.n8545 vdd.n8544 681.178
R2219 vdd.n8546 vdd.n8545 681.178
R2220 vdd.n8546 vdd.n8524 681.178
R2221 vdd.n8561 vdd.n8524 681.178
R2222 vdd.n8561 vdd.n8525 681.178
R2223 vdd.n8553 vdd.n8525 681.178
R2224 vdd.n8538 vdd.n8531 681.178
R2225 vdd.n8547 vdd.n8531 681.178
R2226 vdd.n8547 vdd.n8533 681.178
R2227 vdd.n8533 vdd.n8527 681.178
R2228 vdd.n8558 vdd.n8527 681.178
R2229 vdd.n8558 vdd.n8557 681.178
R2230 vdd.n7127 vdd.n7120 681.178
R2231 vdd.n7136 vdd.n7120 681.178
R2232 vdd.n7136 vdd.n7118 681.178
R2233 vdd.n7142 vdd.n7118 681.178
R2234 vdd.n7143 vdd.n7142 681.178
R2235 vdd.n7145 vdd.n7143 681.178
R2236 vdd.n7134 vdd.n7133 681.178
R2237 vdd.n7135 vdd.n7134 681.178
R2238 vdd.n7135 vdd.n7114 681.178
R2239 vdd.n7151 vdd.n7114 681.178
R2240 vdd.n7151 vdd.n7150 681.178
R2241 vdd.n7150 vdd.n7149 681.178
R2242 vdd.n7173 vdd.n7166 681.178
R2243 vdd.n7182 vdd.n7166 681.178
R2244 vdd.n7182 vdd.n7164 681.178
R2245 vdd.n7188 vdd.n7164 681.178
R2246 vdd.n7189 vdd.n7188 681.178
R2247 vdd.n7191 vdd.n7189 681.178
R2248 vdd.n7180 vdd.n7179 681.178
R2249 vdd.n7181 vdd.n7180 681.178
R2250 vdd.n7181 vdd.n7160 681.178
R2251 vdd.n7197 vdd.n7160 681.178
R2252 vdd.n7197 vdd.n7196 681.178
R2253 vdd.n7196 vdd.n7195 681.178
R2254 vdd.n7270 vdd.n7263 681.178
R2255 vdd.n7279 vdd.n7263 681.178
R2256 vdd.n7279 vdd.n7261 681.178
R2257 vdd.n7285 vdd.n7261 681.178
R2258 vdd.n7286 vdd.n7285 681.178
R2259 vdd.n7288 vdd.n7286 681.178
R2260 vdd.n7277 vdd.n7276 681.178
R2261 vdd.n7278 vdd.n7277 681.178
R2262 vdd.n7278 vdd.n7257 681.178
R2263 vdd.n7294 vdd.n7257 681.178
R2264 vdd.n7294 vdd.n7293 681.178
R2265 vdd.n7293 vdd.n7292 681.178
R2266 vdd.n7316 vdd.n7309 681.178
R2267 vdd.n7325 vdd.n7309 681.178
R2268 vdd.n7325 vdd.n7307 681.178
R2269 vdd.n7331 vdd.n7307 681.178
R2270 vdd.n7332 vdd.n7331 681.178
R2271 vdd.n7334 vdd.n7332 681.178
R2272 vdd.n7323 vdd.n7322 681.178
R2273 vdd.n7324 vdd.n7323 681.178
R2274 vdd.n7324 vdd.n7303 681.178
R2275 vdd.n7340 vdd.n7303 681.178
R2276 vdd.n7340 vdd.n7339 681.178
R2277 vdd.n7339 vdd.n7338 681.178
R2278 vdd.n7362 vdd.n7355 681.178
R2279 vdd.n7371 vdd.n7355 681.178
R2280 vdd.n7371 vdd.n7353 681.178
R2281 vdd.n7377 vdd.n7353 681.178
R2282 vdd.n7378 vdd.n7377 681.178
R2283 vdd.n7380 vdd.n7378 681.178
R2284 vdd.n7369 vdd.n7368 681.178
R2285 vdd.n7370 vdd.n7369 681.178
R2286 vdd.n7370 vdd.n7349 681.178
R2287 vdd.n7386 vdd.n7349 681.178
R2288 vdd.n7386 vdd.n7385 681.178
R2289 vdd.n7385 vdd.n7384 681.178
R2290 vdd.n7408 vdd.n7401 681.178
R2291 vdd.n7417 vdd.n7401 681.178
R2292 vdd.n7417 vdd.n7399 681.178
R2293 vdd.n7423 vdd.n7399 681.178
R2294 vdd.n7424 vdd.n7423 681.178
R2295 vdd.n7426 vdd.n7424 681.178
R2296 vdd.n7415 vdd.n7414 681.178
R2297 vdd.n7416 vdd.n7415 681.178
R2298 vdd.n7416 vdd.n7395 681.178
R2299 vdd.n7432 vdd.n7395 681.178
R2300 vdd.n7432 vdd.n7431 681.178
R2301 vdd.n7431 vdd.n7430 681.178
R2302 vdd.n7505 vdd.n7498 681.178
R2303 vdd.n7514 vdd.n7498 681.178
R2304 vdd.n7514 vdd.n7496 681.178
R2305 vdd.n7520 vdd.n7496 681.178
R2306 vdd.n7521 vdd.n7520 681.178
R2307 vdd.n7523 vdd.n7521 681.178
R2308 vdd.n7512 vdd.n7511 681.178
R2309 vdd.n7513 vdd.n7512 681.178
R2310 vdd.n7513 vdd.n7492 681.178
R2311 vdd.n7529 vdd.n7492 681.178
R2312 vdd.n7529 vdd.n7528 681.178
R2313 vdd.n7528 vdd.n7527 681.178
R2314 vdd.n6654 vdd.n6647 681.178
R2315 vdd.n6663 vdd.n6647 681.178
R2316 vdd.n6663 vdd.n6645 681.178
R2317 vdd.n6669 vdd.n6645 681.178
R2318 vdd.n6670 vdd.n6669 681.178
R2319 vdd.n6672 vdd.n6670 681.178
R2320 vdd.n6661 vdd.n6660 681.178
R2321 vdd.n6662 vdd.n6661 681.178
R2322 vdd.n6662 vdd.n6641 681.178
R2323 vdd.n6678 vdd.n6641 681.178
R2324 vdd.n6678 vdd.n6677 681.178
R2325 vdd.n6677 vdd.n6676 681.178
R2326 vdd.n7549 vdd.n7542 681.178
R2327 vdd.n7558 vdd.n7542 681.178
R2328 vdd.n7558 vdd.n7540 681.178
R2329 vdd.n7564 vdd.n7540 681.178
R2330 vdd.n7565 vdd.n7564 681.178
R2331 vdd.n7567 vdd.n7565 681.178
R2332 vdd.n7556 vdd.n7555 681.178
R2333 vdd.n7557 vdd.n7556 681.178
R2334 vdd.n7557 vdd.n7536 681.178
R2335 vdd.n7573 vdd.n7536 681.178
R2336 vdd.n7573 vdd.n7572 681.178
R2337 vdd.n7572 vdd.n7571 681.178
R2338 vdd.n7594 vdd.n7587 681.178
R2339 vdd.n7603 vdd.n7587 681.178
R2340 vdd.n7603 vdd.n7585 681.178
R2341 vdd.n7609 vdd.n7585 681.178
R2342 vdd.n7610 vdd.n7609 681.178
R2343 vdd.n7612 vdd.n7610 681.178
R2344 vdd.n7601 vdd.n7600 681.178
R2345 vdd.n7602 vdd.n7601 681.178
R2346 vdd.n7602 vdd.n7581 681.178
R2347 vdd.n7618 vdd.n7581 681.178
R2348 vdd.n7618 vdd.n7617 681.178
R2349 vdd.n7617 vdd.n7616 681.178
R2350 vdd.n7644 vdd.n7637 681.178
R2351 vdd.n7653 vdd.n7637 681.178
R2352 vdd.n7653 vdd.n7635 681.178
R2353 vdd.n7659 vdd.n7635 681.178
R2354 vdd.n7660 vdd.n7659 681.178
R2355 vdd.n7662 vdd.n7660 681.178
R2356 vdd.n7651 vdd.n7650 681.178
R2357 vdd.n7652 vdd.n7651 681.178
R2358 vdd.n7652 vdd.n7631 681.178
R2359 vdd.n7668 vdd.n7631 681.178
R2360 vdd.n7668 vdd.n7667 681.178
R2361 vdd.n7667 vdd.n7666 681.178
R2362 vdd.n7690 vdd.n7683 681.178
R2363 vdd.n7699 vdd.n7683 681.178
R2364 vdd.n7699 vdd.n7681 681.178
R2365 vdd.n7705 vdd.n7681 681.178
R2366 vdd.n7706 vdd.n7705 681.178
R2367 vdd.n7708 vdd.n7706 681.178
R2368 vdd.n7697 vdd.n7696 681.178
R2369 vdd.n7698 vdd.n7697 681.178
R2370 vdd.n7698 vdd.n7677 681.178
R2371 vdd.n7714 vdd.n7677 681.178
R2372 vdd.n7714 vdd.n7713 681.178
R2373 vdd.n7713 vdd.n7712 681.178
R2374 vdd.n7738 vdd.n7731 681.178
R2375 vdd.n7747 vdd.n7731 681.178
R2376 vdd.n7747 vdd.n7729 681.178
R2377 vdd.n7753 vdd.n7729 681.178
R2378 vdd.n7754 vdd.n7753 681.178
R2379 vdd.n7756 vdd.n7754 681.178
R2380 vdd.n7745 vdd.n7744 681.178
R2381 vdd.n7746 vdd.n7745 681.178
R2382 vdd.n7746 vdd.n7725 681.178
R2383 vdd.n7762 vdd.n7725 681.178
R2384 vdd.n7762 vdd.n7761 681.178
R2385 vdd.n7761 vdd.n7760 681.178
R2386 vdd.n7458 vdd.n7457 681.178
R2387 vdd.n7459 vdd.n7458 681.178
R2388 vdd.n7459 vdd.n7452 681.178
R2389 vdd.n7465 vdd.n7452 681.178
R2390 vdd.n7466 vdd.n7465 681.178
R2391 vdd.n7468 vdd.n7466 681.178
R2392 vdd.n7481 vdd.n7480 681.178
R2393 vdd.n7480 vdd.n7479 681.178
R2394 vdd.n7479 vdd.n7443 681.178
R2395 vdd.n7474 vdd.n7443 681.178
R2396 vdd.n7474 vdd.n7473 681.178
R2397 vdd.n7473 vdd.n7472 681.178
R2398 vdd.n7785 vdd.n7778 681.178
R2399 vdd.n7794 vdd.n7778 681.178
R2400 vdd.n7794 vdd.n7776 681.178
R2401 vdd.n7800 vdd.n7776 681.178
R2402 vdd.n7801 vdd.n7800 681.178
R2403 vdd.n7803 vdd.n7801 681.178
R2404 vdd.n7792 vdd.n7791 681.178
R2405 vdd.n7793 vdd.n7792 681.178
R2406 vdd.n7793 vdd.n7772 681.178
R2407 vdd.n7809 vdd.n7772 681.178
R2408 vdd.n7809 vdd.n7808 681.178
R2409 vdd.n7808 vdd.n7807 681.178
R2410 vdd.n7830 vdd.n7823 681.178
R2411 vdd.n7839 vdd.n7823 681.178
R2412 vdd.n7839 vdd.n7821 681.178
R2413 vdd.n7845 vdd.n7821 681.178
R2414 vdd.n7846 vdd.n7845 681.178
R2415 vdd.n7848 vdd.n7846 681.178
R2416 vdd.n7837 vdd.n7836 681.178
R2417 vdd.n7838 vdd.n7837 681.178
R2418 vdd.n7838 vdd.n7817 681.178
R2419 vdd.n7854 vdd.n7817 681.178
R2420 vdd.n7854 vdd.n7853 681.178
R2421 vdd.n7853 vdd.n7852 681.178
R2422 vdd.n7876 vdd.n7869 681.178
R2423 vdd.n7885 vdd.n7869 681.178
R2424 vdd.n7885 vdd.n7867 681.178
R2425 vdd.n7891 vdd.n7867 681.178
R2426 vdd.n7892 vdd.n7891 681.178
R2427 vdd.n7894 vdd.n7892 681.178
R2428 vdd.n7883 vdd.n7882 681.178
R2429 vdd.n7884 vdd.n7883 681.178
R2430 vdd.n7884 vdd.n7863 681.178
R2431 vdd.n7900 vdd.n7863 681.178
R2432 vdd.n7900 vdd.n7899 681.178
R2433 vdd.n7899 vdd.n7898 681.178
R2434 vdd.n7927 vdd.n7920 681.178
R2435 vdd.n7936 vdd.n7920 681.178
R2436 vdd.n7936 vdd.n7918 681.178
R2437 vdd.n7942 vdd.n7918 681.178
R2438 vdd.n7943 vdd.n7942 681.178
R2439 vdd.n7945 vdd.n7943 681.178
R2440 vdd.n7934 vdd.n7933 681.178
R2441 vdd.n7935 vdd.n7934 681.178
R2442 vdd.n7935 vdd.n7914 681.178
R2443 vdd.n7951 vdd.n7914 681.178
R2444 vdd.n7951 vdd.n7950 681.178
R2445 vdd.n7950 vdd.n7949 681.178
R2446 vdd.n7973 vdd.n7966 681.178
R2447 vdd.n7982 vdd.n7966 681.178
R2448 vdd.n7982 vdd.n7964 681.178
R2449 vdd.n7988 vdd.n7964 681.178
R2450 vdd.n7989 vdd.n7988 681.178
R2451 vdd.n7991 vdd.n7989 681.178
R2452 vdd.n7980 vdd.n7979 681.178
R2453 vdd.n7981 vdd.n7980 681.178
R2454 vdd.n7981 vdd.n7960 681.178
R2455 vdd.n7997 vdd.n7960 681.178
R2456 vdd.n7997 vdd.n7996 681.178
R2457 vdd.n7996 vdd.n7995 681.178
R2458 vdd.n8021 vdd.n8014 681.178
R2459 vdd.n8030 vdd.n8014 681.178
R2460 vdd.n8030 vdd.n8012 681.178
R2461 vdd.n8036 vdd.n8012 681.178
R2462 vdd.n8037 vdd.n8036 681.178
R2463 vdd.n8039 vdd.n8037 681.178
R2464 vdd.n8028 vdd.n8027 681.178
R2465 vdd.n8029 vdd.n8028 681.178
R2466 vdd.n8029 vdd.n8008 681.178
R2467 vdd.n8045 vdd.n8008 681.178
R2468 vdd.n8045 vdd.n8044 681.178
R2469 vdd.n8044 vdd.n8043 681.178
R2470 vdd.n8067 vdd.n8060 681.178
R2471 vdd.n8076 vdd.n8060 681.178
R2472 vdd.n8076 vdd.n8058 681.178
R2473 vdd.n8082 vdd.n8058 681.178
R2474 vdd.n8083 vdd.n8082 681.178
R2475 vdd.n8085 vdd.n8083 681.178
R2476 vdd.n8074 vdd.n8073 681.178
R2477 vdd.n8075 vdd.n8074 681.178
R2478 vdd.n8075 vdd.n8054 681.178
R2479 vdd.n8091 vdd.n8054 681.178
R2480 vdd.n8091 vdd.n8090 681.178
R2481 vdd.n8090 vdd.n8089 681.178
R2482 vdd.n8112 vdd.n8105 681.178
R2483 vdd.n8121 vdd.n8105 681.178
R2484 vdd.n8121 vdd.n8103 681.178
R2485 vdd.n8127 vdd.n8103 681.178
R2486 vdd.n8128 vdd.n8127 681.178
R2487 vdd.n8130 vdd.n8128 681.178
R2488 vdd.n8119 vdd.n8118 681.178
R2489 vdd.n8120 vdd.n8119 681.178
R2490 vdd.n8120 vdd.n8099 681.178
R2491 vdd.n8136 vdd.n8099 681.178
R2492 vdd.n8136 vdd.n8135 681.178
R2493 vdd.n8135 vdd.n8134 681.178
R2494 vdd.n8162 vdd.n8155 681.178
R2495 vdd.n8171 vdd.n8155 681.178
R2496 vdd.n8171 vdd.n8153 681.178
R2497 vdd.n8177 vdd.n8153 681.178
R2498 vdd.n8178 vdd.n8177 681.178
R2499 vdd.n8180 vdd.n8178 681.178
R2500 vdd.n8169 vdd.n8168 681.178
R2501 vdd.n8170 vdd.n8169 681.178
R2502 vdd.n8170 vdd.n8149 681.178
R2503 vdd.n8186 vdd.n8149 681.178
R2504 vdd.n8186 vdd.n8185 681.178
R2505 vdd.n8185 vdd.n8184 681.178
R2506 vdd.n8208 vdd.n8201 681.178
R2507 vdd.n8217 vdd.n8201 681.178
R2508 vdd.n8217 vdd.n8199 681.178
R2509 vdd.n8223 vdd.n8199 681.178
R2510 vdd.n8224 vdd.n8223 681.178
R2511 vdd.n8226 vdd.n8224 681.178
R2512 vdd.n8215 vdd.n8214 681.178
R2513 vdd.n8216 vdd.n8215 681.178
R2514 vdd.n8216 vdd.n8195 681.178
R2515 vdd.n8232 vdd.n8195 681.178
R2516 vdd.n8232 vdd.n8231 681.178
R2517 vdd.n8231 vdd.n8230 681.178
R2518 vdd.n8256 vdd.n8249 681.178
R2519 vdd.n8265 vdd.n8249 681.178
R2520 vdd.n8265 vdd.n8247 681.178
R2521 vdd.n8271 vdd.n8247 681.178
R2522 vdd.n8272 vdd.n8271 681.178
R2523 vdd.n8274 vdd.n8272 681.178
R2524 vdd.n8263 vdd.n8262 681.178
R2525 vdd.n8264 vdd.n8263 681.178
R2526 vdd.n8264 vdd.n8243 681.178
R2527 vdd.n8280 vdd.n8243 681.178
R2528 vdd.n8280 vdd.n8279 681.178
R2529 vdd.n8279 vdd.n8278 681.178
R2530 vdd.n7223 vdd.n7222 681.178
R2531 vdd.n7224 vdd.n7223 681.178
R2532 vdd.n7224 vdd.n7217 681.178
R2533 vdd.n7230 vdd.n7217 681.178
R2534 vdd.n7231 vdd.n7230 681.178
R2535 vdd.n7233 vdd.n7231 681.178
R2536 vdd.n7246 vdd.n7245 681.178
R2537 vdd.n7245 vdd.n7244 681.178
R2538 vdd.n7244 vdd.n7208 681.178
R2539 vdd.n7239 vdd.n7208 681.178
R2540 vdd.n7239 vdd.n7238 681.178
R2541 vdd.n7238 vdd.n7237 681.178
R2542 vdd.n8303 vdd.n8296 681.178
R2543 vdd.n8312 vdd.n8296 681.178
R2544 vdd.n8312 vdd.n8294 681.178
R2545 vdd.n8318 vdd.n8294 681.178
R2546 vdd.n8319 vdd.n8318 681.178
R2547 vdd.n8321 vdd.n8319 681.178
R2548 vdd.n8310 vdd.n8309 681.178
R2549 vdd.n8311 vdd.n8310 681.178
R2550 vdd.n8311 vdd.n8290 681.178
R2551 vdd.n8327 vdd.n8290 681.178
R2552 vdd.n8327 vdd.n8326 681.178
R2553 vdd.n8326 vdd.n8325 681.178
R2554 vdd.n8348 vdd.n8341 681.178
R2555 vdd.n8357 vdd.n8341 681.178
R2556 vdd.n8357 vdd.n8339 681.178
R2557 vdd.n8363 vdd.n8339 681.178
R2558 vdd.n8364 vdd.n8363 681.178
R2559 vdd.n8366 vdd.n8364 681.178
R2560 vdd.n8355 vdd.n8354 681.178
R2561 vdd.n8356 vdd.n8355 681.178
R2562 vdd.n8356 vdd.n8335 681.178
R2563 vdd.n8372 vdd.n8335 681.178
R2564 vdd.n8372 vdd.n8371 681.178
R2565 vdd.n8371 vdd.n8370 681.178
R2566 vdd.n8398 vdd.n8391 681.178
R2567 vdd.n8407 vdd.n8391 681.178
R2568 vdd.n8407 vdd.n8389 681.178
R2569 vdd.n8413 vdd.n8389 681.178
R2570 vdd.n8414 vdd.n8413 681.178
R2571 vdd.n8416 vdd.n8414 681.178
R2572 vdd.n8405 vdd.n8404 681.178
R2573 vdd.n8406 vdd.n8405 681.178
R2574 vdd.n8406 vdd.n8385 681.178
R2575 vdd.n8422 vdd.n8385 681.178
R2576 vdd.n8422 vdd.n8421 681.178
R2577 vdd.n8421 vdd.n8420 681.178
R2578 vdd.n8444 vdd.n8437 681.178
R2579 vdd.n8453 vdd.n8437 681.178
R2580 vdd.n8453 vdd.n8435 681.178
R2581 vdd.n8459 vdd.n8435 681.178
R2582 vdd.n8460 vdd.n8459 681.178
R2583 vdd.n8462 vdd.n8460 681.178
R2584 vdd.n8451 vdd.n8450 681.178
R2585 vdd.n8452 vdd.n8451 681.178
R2586 vdd.n8452 vdd.n8431 681.178
R2587 vdd.n8468 vdd.n8431 681.178
R2588 vdd.n8468 vdd.n8467 681.178
R2589 vdd.n8467 vdd.n8466 681.178
R2590 vdd.n8492 vdd.n8485 681.178
R2591 vdd.n8501 vdd.n8485 681.178
R2592 vdd.n8501 vdd.n8483 681.178
R2593 vdd.n8507 vdd.n8483 681.178
R2594 vdd.n8508 vdd.n8507 681.178
R2595 vdd.n8510 vdd.n8508 681.178
R2596 vdd.n8499 vdd.n8498 681.178
R2597 vdd.n8500 vdd.n8499 681.178
R2598 vdd.n8500 vdd.n8479 681.178
R2599 vdd.n8516 vdd.n8479 681.178
R2600 vdd.n8516 vdd.n8515 681.178
R2601 vdd.n8515 vdd.n8514 681.178
R2602 vdd.n8638 vdd.n8637 681.178
R2603 vdd.n8639 vdd.n8638 681.178
R2604 vdd.n8639 vdd.n8617 681.178
R2605 vdd.n8654 vdd.n8617 681.178
R2606 vdd.n8654 vdd.n8618 681.178
R2607 vdd.n8646 vdd.n8618 681.178
R2608 vdd.n8631 vdd.n8624 681.178
R2609 vdd.n8640 vdd.n8624 681.178
R2610 vdd.n8640 vdd.n8626 681.178
R2611 vdd.n8626 vdd.n8620 681.178
R2612 vdd.n8651 vdd.n8620 681.178
R2613 vdd.n8651 vdd.n8650 681.178
R2614 vdd.n8592 vdd.n8591 681.178
R2615 vdd.n8593 vdd.n8592 681.178
R2616 vdd.n8593 vdd.n8571 681.178
R2617 vdd.n8608 vdd.n8571 681.178
R2618 vdd.n8608 vdd.n8572 681.178
R2619 vdd.n8600 vdd.n8572 681.178
R2620 vdd.n8585 vdd.n8578 681.178
R2621 vdd.n8594 vdd.n8578 681.178
R2622 vdd.n8594 vdd.n8580 681.178
R2623 vdd.n8580 vdd.n8574 681.178
R2624 vdd.n8605 vdd.n8574 681.178
R2625 vdd.n8605 vdd.n8604 681.178
R2626 vdd.n8685 vdd.n8684 681.178
R2627 vdd.n8686 vdd.n8685 681.178
R2628 vdd.n8686 vdd.n8664 681.178
R2629 vdd.n8701 vdd.n8664 681.178
R2630 vdd.n8701 vdd.n8665 681.178
R2631 vdd.n8693 vdd.n8665 681.178
R2632 vdd.n8678 vdd.n8671 681.178
R2633 vdd.n8687 vdd.n8671 681.178
R2634 vdd.n8687 vdd.n8673 681.178
R2635 vdd.n8673 vdd.n8667 681.178
R2636 vdd.n8698 vdd.n8667 681.178
R2637 vdd.n8698 vdd.n8697 681.178
R2638 vdd.n8733 vdd.n8732 681.178
R2639 vdd.n8734 vdd.n8733 681.178
R2640 vdd.n8734 vdd.n8712 681.178
R2641 vdd.n8749 vdd.n8712 681.178
R2642 vdd.n8749 vdd.n8713 681.178
R2643 vdd.n8741 vdd.n8713 681.178
R2644 vdd.n8726 vdd.n8719 681.178
R2645 vdd.n8735 vdd.n8719 681.178
R2646 vdd.n8735 vdd.n8721 681.178
R2647 vdd.n8721 vdd.n8715 681.178
R2648 vdd.n8746 vdd.n8715 681.178
R2649 vdd.n8746 vdd.n8745 681.178
R2650 vdd.n8779 vdd.n8778 681.178
R2651 vdd.n8780 vdd.n8779 681.178
R2652 vdd.n8780 vdd.n8758 681.178
R2653 vdd.n8795 vdd.n8758 681.178
R2654 vdd.n8795 vdd.n8759 681.178
R2655 vdd.n8787 vdd.n8759 681.178
R2656 vdd.n8772 vdd.n8765 681.178
R2657 vdd.n8781 vdd.n8765 681.178
R2658 vdd.n8781 vdd.n8767 681.178
R2659 vdd.n8767 vdd.n8761 681.178
R2660 vdd.n8792 vdd.n8761 681.178
R2661 vdd.n8792 vdd.n8791 681.178
R2662 vdd.n7033 vdd.n7021 681.178
R2663 vdd.n7043 vdd.n7021 681.178
R2664 vdd.n7043 vdd.n7022 681.178
R2665 vdd.n7022 vdd.n7018 681.178
R2666 vdd.n7052 vdd.n7018 681.178
R2667 vdd.n7053 vdd.n7052 681.178
R2668 vdd.n7035 vdd.n7031 681.178
R2669 vdd.n7031 vdd.n7024 681.178
R2670 vdd.n7026 vdd.n7024 681.178
R2671 vdd.n7041 vdd.n7026 681.178
R2672 vdd.n7041 vdd.n7016 681.178
R2673 vdd.n7055 vdd.n7016 681.178
R2674 vdd.n8921 vdd.n8920 681.178
R2675 vdd.n8922 vdd.n8921 681.178
R2676 vdd.n8922 vdd.n8900 681.178
R2677 vdd.n8937 vdd.n8900 681.178
R2678 vdd.n8937 vdd.n8901 681.178
R2679 vdd.n8929 vdd.n8901 681.178
R2680 vdd.n8914 vdd.n8907 681.178
R2681 vdd.n8923 vdd.n8907 681.178
R2682 vdd.n8923 vdd.n8909 681.178
R2683 vdd.n8909 vdd.n8903 681.178
R2684 vdd.n8934 vdd.n8903 681.178
R2685 vdd.n8934 vdd.n8933 681.178
R2686 vdd.n8874 vdd.n8873 681.178
R2687 vdd.n8875 vdd.n8874 681.178
R2688 vdd.n8875 vdd.n8853 681.178
R2689 vdd.n8890 vdd.n8853 681.178
R2690 vdd.n8890 vdd.n8854 681.178
R2691 vdd.n8882 vdd.n8854 681.178
R2692 vdd.n8867 vdd.n8860 681.178
R2693 vdd.n8876 vdd.n8860 681.178
R2694 vdd.n8876 vdd.n8862 681.178
R2695 vdd.n8862 vdd.n8856 681.178
R2696 vdd.n8887 vdd.n8856 681.178
R2697 vdd.n8887 vdd.n8886 681.178
R2698 vdd.n8828 vdd.n8827 681.178
R2699 vdd.n8829 vdd.n8828 681.178
R2700 vdd.n8829 vdd.n8807 681.178
R2701 vdd.n8844 vdd.n8807 681.178
R2702 vdd.n8844 vdd.n8808 681.178
R2703 vdd.n8836 vdd.n8808 681.178
R2704 vdd.n8821 vdd.n8814 681.178
R2705 vdd.n8830 vdd.n8814 681.178
R2706 vdd.n8830 vdd.n8816 681.178
R2707 vdd.n8816 vdd.n8810 681.178
R2708 vdd.n8841 vdd.n8810 681.178
R2709 vdd.n8841 vdd.n8840 681.178
R2710 vdd.n8968 vdd.n8967 681.178
R2711 vdd.n8969 vdd.n8968 681.178
R2712 vdd.n8969 vdd.n8947 681.178
R2713 vdd.n8984 vdd.n8947 681.178
R2714 vdd.n8984 vdd.n8948 681.178
R2715 vdd.n8976 vdd.n8948 681.178
R2716 vdd.n8961 vdd.n8954 681.178
R2717 vdd.n8970 vdd.n8954 681.178
R2718 vdd.n8970 vdd.n8956 681.178
R2719 vdd.n8956 vdd.n8950 681.178
R2720 vdd.n8981 vdd.n8950 681.178
R2721 vdd.n8981 vdd.n8980 681.178
R2722 vdd.n9016 vdd.n9015 681.178
R2723 vdd.n9017 vdd.n9016 681.178
R2724 vdd.n9017 vdd.n8995 681.178
R2725 vdd.n9032 vdd.n8995 681.178
R2726 vdd.n9032 vdd.n8996 681.178
R2727 vdd.n9024 vdd.n8996 681.178
R2728 vdd.n9009 vdd.n9002 681.178
R2729 vdd.n9018 vdd.n9002 681.178
R2730 vdd.n9018 vdd.n9004 681.178
R2731 vdd.n9004 vdd.n8998 681.178
R2732 vdd.n9029 vdd.n8998 681.178
R2733 vdd.n9029 vdd.n9028 681.178
R2734 vdd.n9062 vdd.n9061 681.178
R2735 vdd.n9063 vdd.n9062 681.178
R2736 vdd.n9063 vdd.n9041 681.178
R2737 vdd.n9078 vdd.n9041 681.178
R2738 vdd.n9078 vdd.n9042 681.178
R2739 vdd.n9070 vdd.n9042 681.178
R2740 vdd.n9055 vdd.n9048 681.178
R2741 vdd.n9064 vdd.n9048 681.178
R2742 vdd.n9064 vdd.n9050 681.178
R2743 vdd.n9050 vdd.n9044 681.178
R2744 vdd.n9075 vdd.n9044 681.178
R2745 vdd.n9075 vdd.n9074 681.178
R2746 vdd.n9156 vdd.n9155 681.178
R2747 vdd.n9157 vdd.n9156 681.178
R2748 vdd.n9157 vdd.n9135 681.178
R2749 vdd.n9172 vdd.n9135 681.178
R2750 vdd.n9172 vdd.n9136 681.178
R2751 vdd.n9164 vdd.n9136 681.178
R2752 vdd.n9149 vdd.n9142 681.178
R2753 vdd.n9158 vdd.n9142 681.178
R2754 vdd.n9158 vdd.n9144 681.178
R2755 vdd.n9144 vdd.n9138 681.178
R2756 vdd.n9169 vdd.n9138 681.178
R2757 vdd.n9169 vdd.n9168 681.178
R2758 vdd.n9110 vdd.n9109 681.178
R2759 vdd.n9111 vdd.n9110 681.178
R2760 vdd.n9111 vdd.n9089 681.178
R2761 vdd.n9126 vdd.n9089 681.178
R2762 vdd.n9126 vdd.n9090 681.178
R2763 vdd.n9118 vdd.n9090 681.178
R2764 vdd.n9103 vdd.n9096 681.178
R2765 vdd.n9112 vdd.n9096 681.178
R2766 vdd.n9112 vdd.n9098 681.178
R2767 vdd.n9098 vdd.n9092 681.178
R2768 vdd.n9123 vdd.n9092 681.178
R2769 vdd.n9123 vdd.n9122 681.178
R2770 vdd.n9203 vdd.n9202 681.178
R2771 vdd.n9204 vdd.n9203 681.178
R2772 vdd.n9204 vdd.n9182 681.178
R2773 vdd.n9219 vdd.n9182 681.178
R2774 vdd.n9219 vdd.n9183 681.178
R2775 vdd.n9211 vdd.n9183 681.178
R2776 vdd.n9196 vdd.n9189 681.178
R2777 vdd.n9205 vdd.n9189 681.178
R2778 vdd.n9205 vdd.n9191 681.178
R2779 vdd.n9191 vdd.n9185 681.178
R2780 vdd.n9216 vdd.n9185 681.178
R2781 vdd.n9216 vdd.n9215 681.178
R2782 vdd.n9251 vdd.n9250 681.178
R2783 vdd.n9252 vdd.n9251 681.178
R2784 vdd.n9252 vdd.n9230 681.178
R2785 vdd.n9267 vdd.n9230 681.178
R2786 vdd.n9267 vdd.n9231 681.178
R2787 vdd.n9259 vdd.n9231 681.178
R2788 vdd.n9244 vdd.n9237 681.178
R2789 vdd.n9253 vdd.n9237 681.178
R2790 vdd.n9253 vdd.n9239 681.178
R2791 vdd.n9239 vdd.n9233 681.178
R2792 vdd.n9264 vdd.n9233 681.178
R2793 vdd.n9264 vdd.n9263 681.178
R2794 vdd.n9297 vdd.n9296 681.178
R2795 vdd.n9298 vdd.n9297 681.178
R2796 vdd.n9298 vdd.n9276 681.178
R2797 vdd.n9313 vdd.n9276 681.178
R2798 vdd.n9313 vdd.n9277 681.178
R2799 vdd.n9305 vdd.n9277 681.178
R2800 vdd.n9290 vdd.n9283 681.178
R2801 vdd.n9299 vdd.n9283 681.178
R2802 vdd.n9299 vdd.n9285 681.178
R2803 vdd.n9285 vdd.n9279 681.178
R2804 vdd.n9310 vdd.n9279 681.178
R2805 vdd.n9310 vdd.n9309 681.178
R2806 vdd.n6797 vdd.n6785 681.178
R2807 vdd.n6807 vdd.n6785 681.178
R2808 vdd.n6807 vdd.n6786 681.178
R2809 vdd.n6786 vdd.n6782 681.178
R2810 vdd.n6816 vdd.n6782 681.178
R2811 vdd.n6817 vdd.n6816 681.178
R2812 vdd.n6799 vdd.n6795 681.178
R2813 vdd.n6795 vdd.n6788 681.178
R2814 vdd.n6790 vdd.n6788 681.178
R2815 vdd.n6805 vdd.n6790 681.178
R2816 vdd.n6805 vdd.n6780 681.178
R2817 vdd.n6819 vdd.n6780 681.178
R2818 vdd.n9392 vdd.n9391 681.178
R2819 vdd.n9393 vdd.n9392 681.178
R2820 vdd.n9393 vdd.n9371 681.178
R2821 vdd.n9408 vdd.n9371 681.178
R2822 vdd.n9408 vdd.n9372 681.178
R2823 vdd.n9400 vdd.n9372 681.178
R2824 vdd.n9385 vdd.n9378 681.178
R2825 vdd.n9394 vdd.n9378 681.178
R2826 vdd.n9394 vdd.n9380 681.178
R2827 vdd.n9380 vdd.n9374 681.178
R2828 vdd.n9405 vdd.n9374 681.178
R2829 vdd.n9405 vdd.n9404 681.178
R2830 vdd.n9346 vdd.n9345 681.178
R2831 vdd.n9347 vdd.n9346 681.178
R2832 vdd.n9347 vdd.n9325 681.178
R2833 vdd.n9362 vdd.n9325 681.178
R2834 vdd.n9362 vdd.n9326 681.178
R2835 vdd.n9354 vdd.n9326 681.178
R2836 vdd.n9339 vdd.n9332 681.178
R2837 vdd.n9348 vdd.n9332 681.178
R2838 vdd.n9348 vdd.n9334 681.178
R2839 vdd.n9334 vdd.n9328 681.178
R2840 vdd.n9359 vdd.n9328 681.178
R2841 vdd.n9359 vdd.n9358 681.178
R2842 vdd.n9439 vdd.n9438 681.178
R2843 vdd.n9440 vdd.n9439 681.178
R2844 vdd.n9440 vdd.n9418 681.178
R2845 vdd.n9455 vdd.n9418 681.178
R2846 vdd.n9455 vdd.n9419 681.178
R2847 vdd.n9447 vdd.n9419 681.178
R2848 vdd.n9432 vdd.n9425 681.178
R2849 vdd.n9441 vdd.n9425 681.178
R2850 vdd.n9441 vdd.n9427 681.178
R2851 vdd.n9427 vdd.n9421 681.178
R2852 vdd.n9452 vdd.n9421 681.178
R2853 vdd.n9452 vdd.n9451 681.178
R2854 vdd.n9487 vdd.n9486 681.178
R2855 vdd.n9488 vdd.n9487 681.178
R2856 vdd.n9488 vdd.n9466 681.178
R2857 vdd.n9503 vdd.n9466 681.178
R2858 vdd.n9503 vdd.n9467 681.178
R2859 vdd.n9495 vdd.n9467 681.178
R2860 vdd.n9480 vdd.n9473 681.178
R2861 vdd.n9489 vdd.n9473 681.178
R2862 vdd.n9489 vdd.n9475 681.178
R2863 vdd.n9475 vdd.n9469 681.178
R2864 vdd.n9500 vdd.n9469 681.178
R2865 vdd.n9500 vdd.n9499 681.178
R2866 vdd.n9533 vdd.n9532 681.178
R2867 vdd.n9534 vdd.n9533 681.178
R2868 vdd.n9534 vdd.n9512 681.178
R2869 vdd.n9549 vdd.n9512 681.178
R2870 vdd.n9549 vdd.n9513 681.178
R2871 vdd.n9541 vdd.n9513 681.178
R2872 vdd.n9526 vdd.n9519 681.178
R2873 vdd.n9535 vdd.n9519 681.178
R2874 vdd.n9535 vdd.n9521 681.178
R2875 vdd.n9521 vdd.n9515 681.178
R2876 vdd.n9546 vdd.n9515 681.178
R2877 vdd.n9546 vdd.n9545 681.178
R2878 vdd.n3693 vdd.n3692 681.178
R2879 vdd.n3694 vdd.n3693 681.178
R2880 vdd.n3694 vdd.n3672 681.178
R2881 vdd.n3709 vdd.n3672 681.178
R2882 vdd.n3709 vdd.n3673 681.178
R2883 vdd.n3701 vdd.n3673 681.178
R2884 vdd.n3686 vdd.n3679 681.178
R2885 vdd.n3695 vdd.n3679 681.178
R2886 vdd.n3695 vdd.n3681 681.178
R2887 vdd.n3681 vdd.n3675 681.178
R2888 vdd.n3706 vdd.n3675 681.178
R2889 vdd.n3706 vdd.n3705 681.178
R2890 vdd.n3739 vdd.n3738 681.178
R2891 vdd.n3740 vdd.n3739 681.178
R2892 vdd.n3740 vdd.n3718 681.178
R2893 vdd.n3755 vdd.n3718 681.178
R2894 vdd.n3755 vdd.n3719 681.178
R2895 vdd.n3747 vdd.n3719 681.178
R2896 vdd.n3732 vdd.n3725 681.178
R2897 vdd.n3741 vdd.n3725 681.178
R2898 vdd.n3741 vdd.n3727 681.178
R2899 vdd.n3727 vdd.n3721 681.178
R2900 vdd.n3752 vdd.n3721 681.178
R2901 vdd.n3752 vdd.n3751 681.178
R2902 vdd.n3837 vdd.n3836 681.178
R2903 vdd.n3838 vdd.n3837 681.178
R2904 vdd.n3838 vdd.n3816 681.178
R2905 vdd.n3853 vdd.n3816 681.178
R2906 vdd.n3853 vdd.n3817 681.178
R2907 vdd.n3845 vdd.n3817 681.178
R2908 vdd.n3830 vdd.n3823 681.178
R2909 vdd.n3839 vdd.n3823 681.178
R2910 vdd.n3839 vdd.n3825 681.178
R2911 vdd.n3825 vdd.n3819 681.178
R2912 vdd.n3850 vdd.n3819 681.178
R2913 vdd.n3850 vdd.n3849 681.178
R2914 vdd.n3883 vdd.n3882 681.178
R2915 vdd.n3884 vdd.n3883 681.178
R2916 vdd.n3884 vdd.n3862 681.178
R2917 vdd.n3899 vdd.n3862 681.178
R2918 vdd.n3899 vdd.n3863 681.178
R2919 vdd.n3891 vdd.n3863 681.178
R2920 vdd.n3876 vdd.n3869 681.178
R2921 vdd.n3885 vdd.n3869 681.178
R2922 vdd.n3885 vdd.n3871 681.178
R2923 vdd.n3871 vdd.n3865 681.178
R2924 vdd.n3896 vdd.n3865 681.178
R2925 vdd.n3896 vdd.n3895 681.178
R2926 vdd.n3929 vdd.n3928 681.178
R2927 vdd.n3930 vdd.n3929 681.178
R2928 vdd.n3930 vdd.n3908 681.178
R2929 vdd.n3945 vdd.n3908 681.178
R2930 vdd.n3945 vdd.n3909 681.178
R2931 vdd.n3937 vdd.n3909 681.178
R2932 vdd.n3922 vdd.n3915 681.178
R2933 vdd.n3931 vdd.n3915 681.178
R2934 vdd.n3931 vdd.n3917 681.178
R2935 vdd.n3917 vdd.n3911 681.178
R2936 vdd.n3942 vdd.n3911 681.178
R2937 vdd.n3942 vdd.n3941 681.178
R2938 vdd.n3975 vdd.n3974 681.178
R2939 vdd.n3976 vdd.n3975 681.178
R2940 vdd.n3976 vdd.n3954 681.178
R2941 vdd.n3991 vdd.n3954 681.178
R2942 vdd.n3991 vdd.n3955 681.178
R2943 vdd.n3983 vdd.n3955 681.178
R2944 vdd.n3968 vdd.n3961 681.178
R2945 vdd.n3977 vdd.n3961 681.178
R2946 vdd.n3977 vdd.n3963 681.178
R2947 vdd.n3963 vdd.n3957 681.178
R2948 vdd.n3988 vdd.n3957 681.178
R2949 vdd.n3988 vdd.n3987 681.178
R2950 vdd.n4073 vdd.n4072 681.178
R2951 vdd.n4074 vdd.n4073 681.178
R2952 vdd.n4074 vdd.n4052 681.178
R2953 vdd.n4089 vdd.n4052 681.178
R2954 vdd.n4089 vdd.n4053 681.178
R2955 vdd.n4081 vdd.n4053 681.178
R2956 vdd.n4066 vdd.n4059 681.178
R2957 vdd.n4075 vdd.n4059 681.178
R2958 vdd.n4075 vdd.n4061 681.178
R2959 vdd.n4061 vdd.n4055 681.178
R2960 vdd.n4086 vdd.n4055 681.178
R2961 vdd.n4086 vdd.n4085 681.178
R2962 vdd.n5531 vdd.n5530 681.178
R2963 vdd.n5532 vdd.n5531 681.178
R2964 vdd.n5532 vdd.n5510 681.178
R2965 vdd.n5547 vdd.n5510 681.178
R2966 vdd.n5547 vdd.n5511 681.178
R2967 vdd.n5539 vdd.n5511 681.178
R2968 vdd.n5524 vdd.n5517 681.178
R2969 vdd.n5533 vdd.n5517 681.178
R2970 vdd.n5533 vdd.n5519 681.178
R2971 vdd.n5519 vdd.n5513 681.178
R2972 vdd.n5544 vdd.n5513 681.178
R2973 vdd.n5544 vdd.n5543 681.178
R2974 vdd.n4113 vdd.n4106 681.178
R2975 vdd.n4122 vdd.n4106 681.178
R2976 vdd.n4122 vdd.n4104 681.178
R2977 vdd.n4128 vdd.n4104 681.178
R2978 vdd.n4129 vdd.n4128 681.178
R2979 vdd.n4131 vdd.n4129 681.178
R2980 vdd.n4120 vdd.n4119 681.178
R2981 vdd.n4121 vdd.n4120 681.178
R2982 vdd.n4121 vdd.n4100 681.178
R2983 vdd.n4137 vdd.n4100 681.178
R2984 vdd.n4137 vdd.n4136 681.178
R2985 vdd.n4136 vdd.n4135 681.178
R2986 vdd.n4159 vdd.n4152 681.178
R2987 vdd.n4168 vdd.n4152 681.178
R2988 vdd.n4168 vdd.n4150 681.178
R2989 vdd.n4174 vdd.n4150 681.178
R2990 vdd.n4175 vdd.n4174 681.178
R2991 vdd.n4177 vdd.n4175 681.178
R2992 vdd.n4166 vdd.n4165 681.178
R2993 vdd.n4167 vdd.n4166 681.178
R2994 vdd.n4167 vdd.n4146 681.178
R2995 vdd.n4183 vdd.n4146 681.178
R2996 vdd.n4183 vdd.n4182 681.178
R2997 vdd.n4182 vdd.n4181 681.178
R2998 vdd.n4256 vdd.n4249 681.178
R2999 vdd.n4265 vdd.n4249 681.178
R3000 vdd.n4265 vdd.n4247 681.178
R3001 vdd.n4271 vdd.n4247 681.178
R3002 vdd.n4272 vdd.n4271 681.178
R3003 vdd.n4274 vdd.n4272 681.178
R3004 vdd.n4263 vdd.n4262 681.178
R3005 vdd.n4264 vdd.n4263 681.178
R3006 vdd.n4264 vdd.n4243 681.178
R3007 vdd.n4280 vdd.n4243 681.178
R3008 vdd.n4280 vdd.n4279 681.178
R3009 vdd.n4279 vdd.n4278 681.178
R3010 vdd.n4302 vdd.n4295 681.178
R3011 vdd.n4311 vdd.n4295 681.178
R3012 vdd.n4311 vdd.n4293 681.178
R3013 vdd.n4317 vdd.n4293 681.178
R3014 vdd.n4318 vdd.n4317 681.178
R3015 vdd.n4320 vdd.n4318 681.178
R3016 vdd.n4309 vdd.n4308 681.178
R3017 vdd.n4310 vdd.n4309 681.178
R3018 vdd.n4310 vdd.n4289 681.178
R3019 vdd.n4326 vdd.n4289 681.178
R3020 vdd.n4326 vdd.n4325 681.178
R3021 vdd.n4325 vdd.n4324 681.178
R3022 vdd.n4348 vdd.n4341 681.178
R3023 vdd.n4357 vdd.n4341 681.178
R3024 vdd.n4357 vdd.n4339 681.178
R3025 vdd.n4363 vdd.n4339 681.178
R3026 vdd.n4364 vdd.n4363 681.178
R3027 vdd.n4366 vdd.n4364 681.178
R3028 vdd.n4355 vdd.n4354 681.178
R3029 vdd.n4356 vdd.n4355 681.178
R3030 vdd.n4356 vdd.n4335 681.178
R3031 vdd.n4372 vdd.n4335 681.178
R3032 vdd.n4372 vdd.n4371 681.178
R3033 vdd.n4371 vdd.n4370 681.178
R3034 vdd.n4394 vdd.n4387 681.178
R3035 vdd.n4403 vdd.n4387 681.178
R3036 vdd.n4403 vdd.n4385 681.178
R3037 vdd.n4409 vdd.n4385 681.178
R3038 vdd.n4410 vdd.n4409 681.178
R3039 vdd.n4412 vdd.n4410 681.178
R3040 vdd.n4401 vdd.n4400 681.178
R3041 vdd.n4402 vdd.n4401 681.178
R3042 vdd.n4402 vdd.n4381 681.178
R3043 vdd.n4418 vdd.n4381 681.178
R3044 vdd.n4418 vdd.n4417 681.178
R3045 vdd.n4417 vdd.n4416 681.178
R3046 vdd.n4491 vdd.n4484 681.178
R3047 vdd.n4500 vdd.n4484 681.178
R3048 vdd.n4500 vdd.n4482 681.178
R3049 vdd.n4506 vdd.n4482 681.178
R3050 vdd.n4507 vdd.n4506 681.178
R3051 vdd.n4509 vdd.n4507 681.178
R3052 vdd.n4498 vdd.n4497 681.178
R3053 vdd.n4499 vdd.n4498 681.178
R3054 vdd.n4499 vdd.n4478 681.178
R3055 vdd.n4515 vdd.n4478 681.178
R3056 vdd.n4515 vdd.n4514 681.178
R3057 vdd.n4514 vdd.n4513 681.178
R3058 vdd.n3640 vdd.n3633 681.178
R3059 vdd.n3649 vdd.n3633 681.178
R3060 vdd.n3649 vdd.n3631 681.178
R3061 vdd.n3655 vdd.n3631 681.178
R3062 vdd.n3656 vdd.n3655 681.178
R3063 vdd.n3658 vdd.n3656 681.178
R3064 vdd.n3647 vdd.n3646 681.178
R3065 vdd.n3648 vdd.n3647 681.178
R3066 vdd.n3648 vdd.n3627 681.178
R3067 vdd.n3664 vdd.n3627 681.178
R3068 vdd.n3664 vdd.n3663 681.178
R3069 vdd.n3663 vdd.n3662 681.178
R3070 vdd.n4535 vdd.n4528 681.178
R3071 vdd.n4544 vdd.n4528 681.178
R3072 vdd.n4544 vdd.n4526 681.178
R3073 vdd.n4550 vdd.n4526 681.178
R3074 vdd.n4551 vdd.n4550 681.178
R3075 vdd.n4553 vdd.n4551 681.178
R3076 vdd.n4542 vdd.n4541 681.178
R3077 vdd.n4543 vdd.n4542 681.178
R3078 vdd.n4543 vdd.n4522 681.178
R3079 vdd.n4559 vdd.n4522 681.178
R3080 vdd.n4559 vdd.n4558 681.178
R3081 vdd.n4558 vdd.n4557 681.178
R3082 vdd.n4580 vdd.n4573 681.178
R3083 vdd.n4589 vdd.n4573 681.178
R3084 vdd.n4589 vdd.n4571 681.178
R3085 vdd.n4595 vdd.n4571 681.178
R3086 vdd.n4596 vdd.n4595 681.178
R3087 vdd.n4598 vdd.n4596 681.178
R3088 vdd.n4587 vdd.n4586 681.178
R3089 vdd.n4588 vdd.n4587 681.178
R3090 vdd.n4588 vdd.n4567 681.178
R3091 vdd.n4604 vdd.n4567 681.178
R3092 vdd.n4604 vdd.n4603 681.178
R3093 vdd.n4603 vdd.n4602 681.178
R3094 vdd.n4630 vdd.n4623 681.178
R3095 vdd.n4639 vdd.n4623 681.178
R3096 vdd.n4639 vdd.n4621 681.178
R3097 vdd.n4645 vdd.n4621 681.178
R3098 vdd.n4646 vdd.n4645 681.178
R3099 vdd.n4648 vdd.n4646 681.178
R3100 vdd.n4637 vdd.n4636 681.178
R3101 vdd.n4638 vdd.n4637 681.178
R3102 vdd.n4638 vdd.n4617 681.178
R3103 vdd.n4654 vdd.n4617 681.178
R3104 vdd.n4654 vdd.n4653 681.178
R3105 vdd.n4653 vdd.n4652 681.178
R3106 vdd.n4676 vdd.n4669 681.178
R3107 vdd.n4685 vdd.n4669 681.178
R3108 vdd.n4685 vdd.n4667 681.178
R3109 vdd.n4691 vdd.n4667 681.178
R3110 vdd.n4692 vdd.n4691 681.178
R3111 vdd.n4694 vdd.n4692 681.178
R3112 vdd.n4683 vdd.n4682 681.178
R3113 vdd.n4684 vdd.n4683 681.178
R3114 vdd.n4684 vdd.n4663 681.178
R3115 vdd.n4700 vdd.n4663 681.178
R3116 vdd.n4700 vdd.n4699 681.178
R3117 vdd.n4699 vdd.n4698 681.178
R3118 vdd.n4724 vdd.n4717 681.178
R3119 vdd.n4733 vdd.n4717 681.178
R3120 vdd.n4733 vdd.n4715 681.178
R3121 vdd.n4739 vdd.n4715 681.178
R3122 vdd.n4740 vdd.n4739 681.178
R3123 vdd.n4742 vdd.n4740 681.178
R3124 vdd.n4731 vdd.n4730 681.178
R3125 vdd.n4732 vdd.n4731 681.178
R3126 vdd.n4732 vdd.n4711 681.178
R3127 vdd.n4748 vdd.n4711 681.178
R3128 vdd.n4748 vdd.n4747 681.178
R3129 vdd.n4747 vdd.n4746 681.178
R3130 vdd.n4444 vdd.n4443 681.178
R3131 vdd.n4445 vdd.n4444 681.178
R3132 vdd.n4445 vdd.n4438 681.178
R3133 vdd.n4451 vdd.n4438 681.178
R3134 vdd.n4452 vdd.n4451 681.178
R3135 vdd.n4454 vdd.n4452 681.178
R3136 vdd.n4467 vdd.n4466 681.178
R3137 vdd.n4466 vdd.n4465 681.178
R3138 vdd.n4465 vdd.n4429 681.178
R3139 vdd.n4460 vdd.n4429 681.178
R3140 vdd.n4460 vdd.n4459 681.178
R3141 vdd.n4459 vdd.n4458 681.178
R3142 vdd.n4771 vdd.n4764 681.178
R3143 vdd.n4780 vdd.n4764 681.178
R3144 vdd.n4780 vdd.n4762 681.178
R3145 vdd.n4786 vdd.n4762 681.178
R3146 vdd.n4787 vdd.n4786 681.178
R3147 vdd.n4789 vdd.n4787 681.178
R3148 vdd.n4778 vdd.n4777 681.178
R3149 vdd.n4779 vdd.n4778 681.178
R3150 vdd.n4779 vdd.n4758 681.178
R3151 vdd.n4795 vdd.n4758 681.178
R3152 vdd.n4795 vdd.n4794 681.178
R3153 vdd.n4794 vdd.n4793 681.178
R3154 vdd.n4816 vdd.n4809 681.178
R3155 vdd.n4825 vdd.n4809 681.178
R3156 vdd.n4825 vdd.n4807 681.178
R3157 vdd.n4831 vdd.n4807 681.178
R3158 vdd.n4832 vdd.n4831 681.178
R3159 vdd.n4834 vdd.n4832 681.178
R3160 vdd.n4823 vdd.n4822 681.178
R3161 vdd.n4824 vdd.n4823 681.178
R3162 vdd.n4824 vdd.n4803 681.178
R3163 vdd.n4840 vdd.n4803 681.178
R3164 vdd.n4840 vdd.n4839 681.178
R3165 vdd.n4839 vdd.n4838 681.178
R3166 vdd.n4862 vdd.n4855 681.178
R3167 vdd.n4871 vdd.n4855 681.178
R3168 vdd.n4871 vdd.n4853 681.178
R3169 vdd.n4877 vdd.n4853 681.178
R3170 vdd.n4878 vdd.n4877 681.178
R3171 vdd.n4880 vdd.n4878 681.178
R3172 vdd.n4869 vdd.n4868 681.178
R3173 vdd.n4870 vdd.n4869 681.178
R3174 vdd.n4870 vdd.n4849 681.178
R3175 vdd.n4886 vdd.n4849 681.178
R3176 vdd.n4886 vdd.n4885 681.178
R3177 vdd.n4885 vdd.n4884 681.178
R3178 vdd.n4913 vdd.n4906 681.178
R3179 vdd.n4922 vdd.n4906 681.178
R3180 vdd.n4922 vdd.n4904 681.178
R3181 vdd.n4928 vdd.n4904 681.178
R3182 vdd.n4929 vdd.n4928 681.178
R3183 vdd.n4931 vdd.n4929 681.178
R3184 vdd.n4920 vdd.n4919 681.178
R3185 vdd.n4921 vdd.n4920 681.178
R3186 vdd.n4921 vdd.n4900 681.178
R3187 vdd.n4937 vdd.n4900 681.178
R3188 vdd.n4937 vdd.n4936 681.178
R3189 vdd.n4936 vdd.n4935 681.178
R3190 vdd.n4959 vdd.n4952 681.178
R3191 vdd.n4968 vdd.n4952 681.178
R3192 vdd.n4968 vdd.n4950 681.178
R3193 vdd.n4974 vdd.n4950 681.178
R3194 vdd.n4975 vdd.n4974 681.178
R3195 vdd.n4977 vdd.n4975 681.178
R3196 vdd.n4966 vdd.n4965 681.178
R3197 vdd.n4967 vdd.n4966 681.178
R3198 vdd.n4967 vdd.n4946 681.178
R3199 vdd.n4983 vdd.n4946 681.178
R3200 vdd.n4983 vdd.n4982 681.178
R3201 vdd.n4982 vdd.n4981 681.178
R3202 vdd.n5007 vdd.n5000 681.178
R3203 vdd.n5016 vdd.n5000 681.178
R3204 vdd.n5016 vdd.n4998 681.178
R3205 vdd.n5022 vdd.n4998 681.178
R3206 vdd.n5023 vdd.n5022 681.178
R3207 vdd.n5025 vdd.n5023 681.178
R3208 vdd.n5014 vdd.n5013 681.178
R3209 vdd.n5015 vdd.n5014 681.178
R3210 vdd.n5015 vdd.n4994 681.178
R3211 vdd.n5031 vdd.n4994 681.178
R3212 vdd.n5031 vdd.n5030 681.178
R3213 vdd.n5030 vdd.n5029 681.178
R3214 vdd.n5053 vdd.n5046 681.178
R3215 vdd.n5062 vdd.n5046 681.178
R3216 vdd.n5062 vdd.n5044 681.178
R3217 vdd.n5068 vdd.n5044 681.178
R3218 vdd.n5069 vdd.n5068 681.178
R3219 vdd.n5071 vdd.n5069 681.178
R3220 vdd.n5060 vdd.n5059 681.178
R3221 vdd.n5061 vdd.n5060 681.178
R3222 vdd.n5061 vdd.n5040 681.178
R3223 vdd.n5077 vdd.n5040 681.178
R3224 vdd.n5077 vdd.n5076 681.178
R3225 vdd.n5076 vdd.n5075 681.178
R3226 vdd.n5098 vdd.n5091 681.178
R3227 vdd.n5107 vdd.n5091 681.178
R3228 vdd.n5107 vdd.n5089 681.178
R3229 vdd.n5113 vdd.n5089 681.178
R3230 vdd.n5114 vdd.n5113 681.178
R3231 vdd.n5116 vdd.n5114 681.178
R3232 vdd.n5105 vdd.n5104 681.178
R3233 vdd.n5106 vdd.n5105 681.178
R3234 vdd.n5106 vdd.n5085 681.178
R3235 vdd.n5122 vdd.n5085 681.178
R3236 vdd.n5122 vdd.n5121 681.178
R3237 vdd.n5121 vdd.n5120 681.178
R3238 vdd.n5148 vdd.n5141 681.178
R3239 vdd.n5157 vdd.n5141 681.178
R3240 vdd.n5157 vdd.n5139 681.178
R3241 vdd.n5163 vdd.n5139 681.178
R3242 vdd.n5164 vdd.n5163 681.178
R3243 vdd.n5166 vdd.n5164 681.178
R3244 vdd.n5155 vdd.n5154 681.178
R3245 vdd.n5156 vdd.n5155 681.178
R3246 vdd.n5156 vdd.n5135 681.178
R3247 vdd.n5172 vdd.n5135 681.178
R3248 vdd.n5172 vdd.n5171 681.178
R3249 vdd.n5171 vdd.n5170 681.178
R3250 vdd.n5194 vdd.n5187 681.178
R3251 vdd.n5203 vdd.n5187 681.178
R3252 vdd.n5203 vdd.n5185 681.178
R3253 vdd.n5209 vdd.n5185 681.178
R3254 vdd.n5210 vdd.n5209 681.178
R3255 vdd.n5212 vdd.n5210 681.178
R3256 vdd.n5201 vdd.n5200 681.178
R3257 vdd.n5202 vdd.n5201 681.178
R3258 vdd.n5202 vdd.n5181 681.178
R3259 vdd.n5218 vdd.n5181 681.178
R3260 vdd.n5218 vdd.n5217 681.178
R3261 vdd.n5217 vdd.n5216 681.178
R3262 vdd.n5242 vdd.n5235 681.178
R3263 vdd.n5251 vdd.n5235 681.178
R3264 vdd.n5251 vdd.n5233 681.178
R3265 vdd.n5257 vdd.n5233 681.178
R3266 vdd.n5258 vdd.n5257 681.178
R3267 vdd.n5260 vdd.n5258 681.178
R3268 vdd.n5249 vdd.n5248 681.178
R3269 vdd.n5250 vdd.n5249 681.178
R3270 vdd.n5250 vdd.n5229 681.178
R3271 vdd.n5266 vdd.n5229 681.178
R3272 vdd.n5266 vdd.n5265 681.178
R3273 vdd.n5265 vdd.n5264 681.178
R3274 vdd.n4209 vdd.n4208 681.178
R3275 vdd.n4210 vdd.n4209 681.178
R3276 vdd.n4210 vdd.n4203 681.178
R3277 vdd.n4216 vdd.n4203 681.178
R3278 vdd.n4217 vdd.n4216 681.178
R3279 vdd.n4219 vdd.n4217 681.178
R3280 vdd.n4232 vdd.n4231 681.178
R3281 vdd.n4231 vdd.n4230 681.178
R3282 vdd.n4230 vdd.n4194 681.178
R3283 vdd.n4225 vdd.n4194 681.178
R3284 vdd.n4225 vdd.n4224 681.178
R3285 vdd.n4224 vdd.n4223 681.178
R3286 vdd.n5289 vdd.n5282 681.178
R3287 vdd.n5298 vdd.n5282 681.178
R3288 vdd.n5298 vdd.n5280 681.178
R3289 vdd.n5304 vdd.n5280 681.178
R3290 vdd.n5305 vdd.n5304 681.178
R3291 vdd.n5307 vdd.n5305 681.178
R3292 vdd.n5296 vdd.n5295 681.178
R3293 vdd.n5297 vdd.n5296 681.178
R3294 vdd.n5297 vdd.n5276 681.178
R3295 vdd.n5313 vdd.n5276 681.178
R3296 vdd.n5313 vdd.n5312 681.178
R3297 vdd.n5312 vdd.n5311 681.178
R3298 vdd.n5334 vdd.n5327 681.178
R3299 vdd.n5343 vdd.n5327 681.178
R3300 vdd.n5343 vdd.n5325 681.178
R3301 vdd.n5349 vdd.n5325 681.178
R3302 vdd.n5350 vdd.n5349 681.178
R3303 vdd.n5352 vdd.n5350 681.178
R3304 vdd.n5341 vdd.n5340 681.178
R3305 vdd.n5342 vdd.n5341 681.178
R3306 vdd.n5342 vdd.n5321 681.178
R3307 vdd.n5358 vdd.n5321 681.178
R3308 vdd.n5358 vdd.n5357 681.178
R3309 vdd.n5357 vdd.n5356 681.178
R3310 vdd.n5384 vdd.n5377 681.178
R3311 vdd.n5393 vdd.n5377 681.178
R3312 vdd.n5393 vdd.n5375 681.178
R3313 vdd.n5399 vdd.n5375 681.178
R3314 vdd.n5400 vdd.n5399 681.178
R3315 vdd.n5402 vdd.n5400 681.178
R3316 vdd.n5391 vdd.n5390 681.178
R3317 vdd.n5392 vdd.n5391 681.178
R3318 vdd.n5392 vdd.n5371 681.178
R3319 vdd.n5408 vdd.n5371 681.178
R3320 vdd.n5408 vdd.n5407 681.178
R3321 vdd.n5407 vdd.n5406 681.178
R3322 vdd.n5430 vdd.n5423 681.178
R3323 vdd.n5439 vdd.n5423 681.178
R3324 vdd.n5439 vdd.n5421 681.178
R3325 vdd.n5445 vdd.n5421 681.178
R3326 vdd.n5446 vdd.n5445 681.178
R3327 vdd.n5448 vdd.n5446 681.178
R3328 vdd.n5437 vdd.n5436 681.178
R3329 vdd.n5438 vdd.n5437 681.178
R3330 vdd.n5438 vdd.n5417 681.178
R3331 vdd.n5454 vdd.n5417 681.178
R3332 vdd.n5454 vdd.n5453 681.178
R3333 vdd.n5453 vdd.n5452 681.178
R3334 vdd.n5478 vdd.n5471 681.178
R3335 vdd.n5487 vdd.n5471 681.178
R3336 vdd.n5487 vdd.n5469 681.178
R3337 vdd.n5493 vdd.n5469 681.178
R3338 vdd.n5494 vdd.n5493 681.178
R3339 vdd.n5496 vdd.n5494 681.178
R3340 vdd.n5485 vdd.n5484 681.178
R3341 vdd.n5486 vdd.n5485 681.178
R3342 vdd.n5486 vdd.n5465 681.178
R3343 vdd.n5502 vdd.n5465 681.178
R3344 vdd.n5502 vdd.n5501 681.178
R3345 vdd.n5501 vdd.n5500 681.178
R3346 vdd.n5624 vdd.n5623 681.178
R3347 vdd.n5625 vdd.n5624 681.178
R3348 vdd.n5625 vdd.n5603 681.178
R3349 vdd.n5640 vdd.n5603 681.178
R3350 vdd.n5640 vdd.n5604 681.178
R3351 vdd.n5632 vdd.n5604 681.178
R3352 vdd.n5617 vdd.n5610 681.178
R3353 vdd.n5626 vdd.n5610 681.178
R3354 vdd.n5626 vdd.n5612 681.178
R3355 vdd.n5612 vdd.n5606 681.178
R3356 vdd.n5637 vdd.n5606 681.178
R3357 vdd.n5637 vdd.n5636 681.178
R3358 vdd.n5578 vdd.n5577 681.178
R3359 vdd.n5579 vdd.n5578 681.178
R3360 vdd.n5579 vdd.n5557 681.178
R3361 vdd.n5594 vdd.n5557 681.178
R3362 vdd.n5594 vdd.n5558 681.178
R3363 vdd.n5586 vdd.n5558 681.178
R3364 vdd.n5571 vdd.n5564 681.178
R3365 vdd.n5580 vdd.n5564 681.178
R3366 vdd.n5580 vdd.n5566 681.178
R3367 vdd.n5566 vdd.n5560 681.178
R3368 vdd.n5591 vdd.n5560 681.178
R3369 vdd.n5591 vdd.n5590 681.178
R3370 vdd.n5671 vdd.n5670 681.178
R3371 vdd.n5672 vdd.n5671 681.178
R3372 vdd.n5672 vdd.n5650 681.178
R3373 vdd.n5687 vdd.n5650 681.178
R3374 vdd.n5687 vdd.n5651 681.178
R3375 vdd.n5679 vdd.n5651 681.178
R3376 vdd.n5664 vdd.n5657 681.178
R3377 vdd.n5673 vdd.n5657 681.178
R3378 vdd.n5673 vdd.n5659 681.178
R3379 vdd.n5659 vdd.n5653 681.178
R3380 vdd.n5684 vdd.n5653 681.178
R3381 vdd.n5684 vdd.n5683 681.178
R3382 vdd.n5719 vdd.n5718 681.178
R3383 vdd.n5720 vdd.n5719 681.178
R3384 vdd.n5720 vdd.n5698 681.178
R3385 vdd.n5735 vdd.n5698 681.178
R3386 vdd.n5735 vdd.n5699 681.178
R3387 vdd.n5727 vdd.n5699 681.178
R3388 vdd.n5712 vdd.n5705 681.178
R3389 vdd.n5721 vdd.n5705 681.178
R3390 vdd.n5721 vdd.n5707 681.178
R3391 vdd.n5707 vdd.n5701 681.178
R3392 vdd.n5732 vdd.n5701 681.178
R3393 vdd.n5732 vdd.n5731 681.178
R3394 vdd.n5765 vdd.n5764 681.178
R3395 vdd.n5766 vdd.n5765 681.178
R3396 vdd.n5766 vdd.n5744 681.178
R3397 vdd.n5781 vdd.n5744 681.178
R3398 vdd.n5781 vdd.n5745 681.178
R3399 vdd.n5773 vdd.n5745 681.178
R3400 vdd.n5758 vdd.n5751 681.178
R3401 vdd.n5767 vdd.n5751 681.178
R3402 vdd.n5767 vdd.n5753 681.178
R3403 vdd.n5753 vdd.n5747 681.178
R3404 vdd.n5778 vdd.n5747 681.178
R3405 vdd.n5778 vdd.n5777 681.178
R3406 vdd.n4019 vdd.n4007 681.178
R3407 vdd.n4029 vdd.n4007 681.178
R3408 vdd.n4029 vdd.n4008 681.178
R3409 vdd.n4008 vdd.n4004 681.178
R3410 vdd.n4038 vdd.n4004 681.178
R3411 vdd.n4039 vdd.n4038 681.178
R3412 vdd.n4021 vdd.n4017 681.178
R3413 vdd.n4017 vdd.n4010 681.178
R3414 vdd.n4012 vdd.n4010 681.178
R3415 vdd.n4027 vdd.n4012 681.178
R3416 vdd.n4027 vdd.n4002 681.178
R3417 vdd.n4041 vdd.n4002 681.178
R3418 vdd.n5907 vdd.n5906 681.178
R3419 vdd.n5908 vdd.n5907 681.178
R3420 vdd.n5908 vdd.n5886 681.178
R3421 vdd.n5923 vdd.n5886 681.178
R3422 vdd.n5923 vdd.n5887 681.178
R3423 vdd.n5915 vdd.n5887 681.178
R3424 vdd.n5900 vdd.n5893 681.178
R3425 vdd.n5909 vdd.n5893 681.178
R3426 vdd.n5909 vdd.n5895 681.178
R3427 vdd.n5895 vdd.n5889 681.178
R3428 vdd.n5920 vdd.n5889 681.178
R3429 vdd.n5920 vdd.n5919 681.178
R3430 vdd.n5860 vdd.n5859 681.178
R3431 vdd.n5861 vdd.n5860 681.178
R3432 vdd.n5861 vdd.n5839 681.178
R3433 vdd.n5876 vdd.n5839 681.178
R3434 vdd.n5876 vdd.n5840 681.178
R3435 vdd.n5868 vdd.n5840 681.178
R3436 vdd.n5853 vdd.n5846 681.178
R3437 vdd.n5862 vdd.n5846 681.178
R3438 vdd.n5862 vdd.n5848 681.178
R3439 vdd.n5848 vdd.n5842 681.178
R3440 vdd.n5873 vdd.n5842 681.178
R3441 vdd.n5873 vdd.n5872 681.178
R3442 vdd.n5814 vdd.n5813 681.178
R3443 vdd.n5815 vdd.n5814 681.178
R3444 vdd.n5815 vdd.n5793 681.178
R3445 vdd.n5830 vdd.n5793 681.178
R3446 vdd.n5830 vdd.n5794 681.178
R3447 vdd.n5822 vdd.n5794 681.178
R3448 vdd.n5807 vdd.n5800 681.178
R3449 vdd.n5816 vdd.n5800 681.178
R3450 vdd.n5816 vdd.n5802 681.178
R3451 vdd.n5802 vdd.n5796 681.178
R3452 vdd.n5827 vdd.n5796 681.178
R3453 vdd.n5827 vdd.n5826 681.178
R3454 vdd.n5954 vdd.n5953 681.178
R3455 vdd.n5955 vdd.n5954 681.178
R3456 vdd.n5955 vdd.n5933 681.178
R3457 vdd.n5970 vdd.n5933 681.178
R3458 vdd.n5970 vdd.n5934 681.178
R3459 vdd.n5962 vdd.n5934 681.178
R3460 vdd.n5947 vdd.n5940 681.178
R3461 vdd.n5956 vdd.n5940 681.178
R3462 vdd.n5956 vdd.n5942 681.178
R3463 vdd.n5942 vdd.n5936 681.178
R3464 vdd.n5967 vdd.n5936 681.178
R3465 vdd.n5967 vdd.n5966 681.178
R3466 vdd.n6002 vdd.n6001 681.178
R3467 vdd.n6003 vdd.n6002 681.178
R3468 vdd.n6003 vdd.n5981 681.178
R3469 vdd.n6018 vdd.n5981 681.178
R3470 vdd.n6018 vdd.n5982 681.178
R3471 vdd.n6010 vdd.n5982 681.178
R3472 vdd.n5995 vdd.n5988 681.178
R3473 vdd.n6004 vdd.n5988 681.178
R3474 vdd.n6004 vdd.n5990 681.178
R3475 vdd.n5990 vdd.n5984 681.178
R3476 vdd.n6015 vdd.n5984 681.178
R3477 vdd.n6015 vdd.n6014 681.178
R3478 vdd.n6048 vdd.n6047 681.178
R3479 vdd.n6049 vdd.n6048 681.178
R3480 vdd.n6049 vdd.n6027 681.178
R3481 vdd.n6064 vdd.n6027 681.178
R3482 vdd.n6064 vdd.n6028 681.178
R3483 vdd.n6056 vdd.n6028 681.178
R3484 vdd.n6041 vdd.n6034 681.178
R3485 vdd.n6050 vdd.n6034 681.178
R3486 vdd.n6050 vdd.n6036 681.178
R3487 vdd.n6036 vdd.n6030 681.178
R3488 vdd.n6061 vdd.n6030 681.178
R3489 vdd.n6061 vdd.n6060 681.178
R3490 vdd.n6142 vdd.n6141 681.178
R3491 vdd.n6143 vdd.n6142 681.178
R3492 vdd.n6143 vdd.n6121 681.178
R3493 vdd.n6158 vdd.n6121 681.178
R3494 vdd.n6158 vdd.n6122 681.178
R3495 vdd.n6150 vdd.n6122 681.178
R3496 vdd.n6135 vdd.n6128 681.178
R3497 vdd.n6144 vdd.n6128 681.178
R3498 vdd.n6144 vdd.n6130 681.178
R3499 vdd.n6130 vdd.n6124 681.178
R3500 vdd.n6155 vdd.n6124 681.178
R3501 vdd.n6155 vdd.n6154 681.178
R3502 vdd.n6096 vdd.n6095 681.178
R3503 vdd.n6097 vdd.n6096 681.178
R3504 vdd.n6097 vdd.n6075 681.178
R3505 vdd.n6112 vdd.n6075 681.178
R3506 vdd.n6112 vdd.n6076 681.178
R3507 vdd.n6104 vdd.n6076 681.178
R3508 vdd.n6089 vdd.n6082 681.178
R3509 vdd.n6098 vdd.n6082 681.178
R3510 vdd.n6098 vdd.n6084 681.178
R3511 vdd.n6084 vdd.n6078 681.178
R3512 vdd.n6109 vdd.n6078 681.178
R3513 vdd.n6109 vdd.n6108 681.178
R3514 vdd.n6189 vdd.n6188 681.178
R3515 vdd.n6190 vdd.n6189 681.178
R3516 vdd.n6190 vdd.n6168 681.178
R3517 vdd.n6205 vdd.n6168 681.178
R3518 vdd.n6205 vdd.n6169 681.178
R3519 vdd.n6197 vdd.n6169 681.178
R3520 vdd.n6182 vdd.n6175 681.178
R3521 vdd.n6191 vdd.n6175 681.178
R3522 vdd.n6191 vdd.n6177 681.178
R3523 vdd.n6177 vdd.n6171 681.178
R3524 vdd.n6202 vdd.n6171 681.178
R3525 vdd.n6202 vdd.n6201 681.178
R3526 vdd.n6237 vdd.n6236 681.178
R3527 vdd.n6238 vdd.n6237 681.178
R3528 vdd.n6238 vdd.n6216 681.178
R3529 vdd.n6253 vdd.n6216 681.178
R3530 vdd.n6253 vdd.n6217 681.178
R3531 vdd.n6245 vdd.n6217 681.178
R3532 vdd.n6230 vdd.n6223 681.178
R3533 vdd.n6239 vdd.n6223 681.178
R3534 vdd.n6239 vdd.n6225 681.178
R3535 vdd.n6225 vdd.n6219 681.178
R3536 vdd.n6250 vdd.n6219 681.178
R3537 vdd.n6250 vdd.n6249 681.178
R3538 vdd.n6283 vdd.n6282 681.178
R3539 vdd.n6284 vdd.n6283 681.178
R3540 vdd.n6284 vdd.n6262 681.178
R3541 vdd.n6299 vdd.n6262 681.178
R3542 vdd.n6299 vdd.n6263 681.178
R3543 vdd.n6291 vdd.n6263 681.178
R3544 vdd.n6276 vdd.n6269 681.178
R3545 vdd.n6285 vdd.n6269 681.178
R3546 vdd.n6285 vdd.n6271 681.178
R3547 vdd.n6271 vdd.n6265 681.178
R3548 vdd.n6296 vdd.n6265 681.178
R3549 vdd.n6296 vdd.n6295 681.178
R3550 vdd.n3783 vdd.n3771 681.178
R3551 vdd.n3793 vdd.n3771 681.178
R3552 vdd.n3793 vdd.n3772 681.178
R3553 vdd.n3772 vdd.n3768 681.178
R3554 vdd.n3802 vdd.n3768 681.178
R3555 vdd.n3803 vdd.n3802 681.178
R3556 vdd.n3785 vdd.n3781 681.178
R3557 vdd.n3781 vdd.n3774 681.178
R3558 vdd.n3776 vdd.n3774 681.178
R3559 vdd.n3791 vdd.n3776 681.178
R3560 vdd.n3791 vdd.n3766 681.178
R3561 vdd.n3805 vdd.n3766 681.178
R3562 vdd.n6378 vdd.n6377 681.178
R3563 vdd.n6379 vdd.n6378 681.178
R3564 vdd.n6379 vdd.n6357 681.178
R3565 vdd.n6394 vdd.n6357 681.178
R3566 vdd.n6394 vdd.n6358 681.178
R3567 vdd.n6386 vdd.n6358 681.178
R3568 vdd.n6371 vdd.n6364 681.178
R3569 vdd.n6380 vdd.n6364 681.178
R3570 vdd.n6380 vdd.n6366 681.178
R3571 vdd.n6366 vdd.n6360 681.178
R3572 vdd.n6391 vdd.n6360 681.178
R3573 vdd.n6391 vdd.n6390 681.178
R3574 vdd.n6332 vdd.n6331 681.178
R3575 vdd.n6333 vdd.n6332 681.178
R3576 vdd.n6333 vdd.n6311 681.178
R3577 vdd.n6348 vdd.n6311 681.178
R3578 vdd.n6348 vdd.n6312 681.178
R3579 vdd.n6340 vdd.n6312 681.178
R3580 vdd.n6325 vdd.n6318 681.178
R3581 vdd.n6334 vdd.n6318 681.178
R3582 vdd.n6334 vdd.n6320 681.178
R3583 vdd.n6320 vdd.n6314 681.178
R3584 vdd.n6345 vdd.n6314 681.178
R3585 vdd.n6345 vdd.n6344 681.178
R3586 vdd.n6425 vdd.n6424 681.178
R3587 vdd.n6426 vdd.n6425 681.178
R3588 vdd.n6426 vdd.n6404 681.178
R3589 vdd.n6441 vdd.n6404 681.178
R3590 vdd.n6441 vdd.n6405 681.178
R3591 vdd.n6433 vdd.n6405 681.178
R3592 vdd.n6418 vdd.n6411 681.178
R3593 vdd.n6427 vdd.n6411 681.178
R3594 vdd.n6427 vdd.n6413 681.178
R3595 vdd.n6413 vdd.n6407 681.178
R3596 vdd.n6438 vdd.n6407 681.178
R3597 vdd.n6438 vdd.n6437 681.178
R3598 vdd.n6473 vdd.n6472 681.178
R3599 vdd.n6474 vdd.n6473 681.178
R3600 vdd.n6474 vdd.n6452 681.178
R3601 vdd.n6489 vdd.n6452 681.178
R3602 vdd.n6489 vdd.n6453 681.178
R3603 vdd.n6481 vdd.n6453 681.178
R3604 vdd.n6466 vdd.n6459 681.178
R3605 vdd.n6475 vdd.n6459 681.178
R3606 vdd.n6475 vdd.n6461 681.178
R3607 vdd.n6461 vdd.n6455 681.178
R3608 vdd.n6486 vdd.n6455 681.178
R3609 vdd.n6486 vdd.n6485 681.178
R3610 vdd.n6519 vdd.n6518 681.178
R3611 vdd.n6520 vdd.n6519 681.178
R3612 vdd.n6520 vdd.n6498 681.178
R3613 vdd.n6535 vdd.n6498 681.178
R3614 vdd.n6535 vdd.n6499 681.178
R3615 vdd.n6527 vdd.n6499 681.178
R3616 vdd.n6512 vdd.n6505 681.178
R3617 vdd.n6521 vdd.n6505 681.178
R3618 vdd.n6521 vdd.n6507 681.178
R3619 vdd.n6507 vdd.n6501 681.178
R3620 vdd.n6532 vdd.n6501 681.178
R3621 vdd.n6532 vdd.n6531 681.178
R3622 vdd.n679 vdd.n678 681.178
R3623 vdd.n680 vdd.n679 681.178
R3624 vdd.n680 vdd.n658 681.178
R3625 vdd.n695 vdd.n658 681.178
R3626 vdd.n695 vdd.n659 681.178
R3627 vdd.n687 vdd.n659 681.178
R3628 vdd.n672 vdd.n665 681.178
R3629 vdd.n681 vdd.n665 681.178
R3630 vdd.n681 vdd.n667 681.178
R3631 vdd.n667 vdd.n661 681.178
R3632 vdd.n692 vdd.n661 681.178
R3633 vdd.n692 vdd.n691 681.178
R3634 vdd.n725 vdd.n724 681.178
R3635 vdd.n726 vdd.n725 681.178
R3636 vdd.n726 vdd.n704 681.178
R3637 vdd.n741 vdd.n704 681.178
R3638 vdd.n741 vdd.n705 681.178
R3639 vdd.n733 vdd.n705 681.178
R3640 vdd.n718 vdd.n711 681.178
R3641 vdd.n727 vdd.n711 681.178
R3642 vdd.n727 vdd.n713 681.178
R3643 vdd.n713 vdd.n707 681.178
R3644 vdd.n738 vdd.n707 681.178
R3645 vdd.n738 vdd.n737 681.178
R3646 vdd.n823 vdd.n822 681.178
R3647 vdd.n824 vdd.n823 681.178
R3648 vdd.n824 vdd.n802 681.178
R3649 vdd.n839 vdd.n802 681.178
R3650 vdd.n839 vdd.n803 681.178
R3651 vdd.n831 vdd.n803 681.178
R3652 vdd.n816 vdd.n809 681.178
R3653 vdd.n825 vdd.n809 681.178
R3654 vdd.n825 vdd.n811 681.178
R3655 vdd.n811 vdd.n805 681.178
R3656 vdd.n836 vdd.n805 681.178
R3657 vdd.n836 vdd.n835 681.178
R3658 vdd.n869 vdd.n868 681.178
R3659 vdd.n870 vdd.n869 681.178
R3660 vdd.n870 vdd.n848 681.178
R3661 vdd.n885 vdd.n848 681.178
R3662 vdd.n885 vdd.n849 681.178
R3663 vdd.n877 vdd.n849 681.178
R3664 vdd.n862 vdd.n855 681.178
R3665 vdd.n871 vdd.n855 681.178
R3666 vdd.n871 vdd.n857 681.178
R3667 vdd.n857 vdd.n851 681.178
R3668 vdd.n882 vdd.n851 681.178
R3669 vdd.n882 vdd.n881 681.178
R3670 vdd.n915 vdd.n914 681.178
R3671 vdd.n916 vdd.n915 681.178
R3672 vdd.n916 vdd.n894 681.178
R3673 vdd.n931 vdd.n894 681.178
R3674 vdd.n931 vdd.n895 681.178
R3675 vdd.n923 vdd.n895 681.178
R3676 vdd.n908 vdd.n901 681.178
R3677 vdd.n917 vdd.n901 681.178
R3678 vdd.n917 vdd.n903 681.178
R3679 vdd.n903 vdd.n897 681.178
R3680 vdd.n928 vdd.n897 681.178
R3681 vdd.n928 vdd.n927 681.178
R3682 vdd.n961 vdd.n960 681.178
R3683 vdd.n962 vdd.n961 681.178
R3684 vdd.n962 vdd.n940 681.178
R3685 vdd.n977 vdd.n940 681.178
R3686 vdd.n977 vdd.n941 681.178
R3687 vdd.n969 vdd.n941 681.178
R3688 vdd.n954 vdd.n947 681.178
R3689 vdd.n963 vdd.n947 681.178
R3690 vdd.n963 vdd.n949 681.178
R3691 vdd.n949 vdd.n943 681.178
R3692 vdd.n974 vdd.n943 681.178
R3693 vdd.n974 vdd.n973 681.178
R3694 vdd.n1059 vdd.n1058 681.178
R3695 vdd.n1060 vdd.n1059 681.178
R3696 vdd.n1060 vdd.n1038 681.178
R3697 vdd.n1075 vdd.n1038 681.178
R3698 vdd.n1075 vdd.n1039 681.178
R3699 vdd.n1067 vdd.n1039 681.178
R3700 vdd.n1052 vdd.n1045 681.178
R3701 vdd.n1061 vdd.n1045 681.178
R3702 vdd.n1061 vdd.n1047 681.178
R3703 vdd.n1047 vdd.n1041 681.178
R3704 vdd.n1072 vdd.n1041 681.178
R3705 vdd.n1072 vdd.n1071 681.178
R3706 vdd.n2517 vdd.n2516 681.178
R3707 vdd.n2518 vdd.n2517 681.178
R3708 vdd.n2518 vdd.n2496 681.178
R3709 vdd.n2533 vdd.n2496 681.178
R3710 vdd.n2533 vdd.n2497 681.178
R3711 vdd.n2525 vdd.n2497 681.178
R3712 vdd.n2510 vdd.n2503 681.178
R3713 vdd.n2519 vdd.n2503 681.178
R3714 vdd.n2519 vdd.n2505 681.178
R3715 vdd.n2505 vdd.n2499 681.178
R3716 vdd.n2530 vdd.n2499 681.178
R3717 vdd.n2530 vdd.n2529 681.178
R3718 vdd.n1099 vdd.n1092 681.178
R3719 vdd.n1108 vdd.n1092 681.178
R3720 vdd.n1108 vdd.n1090 681.178
R3721 vdd.n1114 vdd.n1090 681.178
R3722 vdd.n1115 vdd.n1114 681.178
R3723 vdd.n1117 vdd.n1115 681.178
R3724 vdd.n1106 vdd.n1105 681.178
R3725 vdd.n1107 vdd.n1106 681.178
R3726 vdd.n1107 vdd.n1086 681.178
R3727 vdd.n1123 vdd.n1086 681.178
R3728 vdd.n1123 vdd.n1122 681.178
R3729 vdd.n1122 vdd.n1121 681.178
R3730 vdd.n1145 vdd.n1138 681.178
R3731 vdd.n1154 vdd.n1138 681.178
R3732 vdd.n1154 vdd.n1136 681.178
R3733 vdd.n1160 vdd.n1136 681.178
R3734 vdd.n1161 vdd.n1160 681.178
R3735 vdd.n1163 vdd.n1161 681.178
R3736 vdd.n1152 vdd.n1151 681.178
R3737 vdd.n1153 vdd.n1152 681.178
R3738 vdd.n1153 vdd.n1132 681.178
R3739 vdd.n1169 vdd.n1132 681.178
R3740 vdd.n1169 vdd.n1168 681.178
R3741 vdd.n1168 vdd.n1167 681.178
R3742 vdd.n1242 vdd.n1235 681.178
R3743 vdd.n1251 vdd.n1235 681.178
R3744 vdd.n1251 vdd.n1233 681.178
R3745 vdd.n1257 vdd.n1233 681.178
R3746 vdd.n1258 vdd.n1257 681.178
R3747 vdd.n1260 vdd.n1258 681.178
R3748 vdd.n1249 vdd.n1248 681.178
R3749 vdd.n1250 vdd.n1249 681.178
R3750 vdd.n1250 vdd.n1229 681.178
R3751 vdd.n1266 vdd.n1229 681.178
R3752 vdd.n1266 vdd.n1265 681.178
R3753 vdd.n1265 vdd.n1264 681.178
R3754 vdd.n1288 vdd.n1281 681.178
R3755 vdd.n1297 vdd.n1281 681.178
R3756 vdd.n1297 vdd.n1279 681.178
R3757 vdd.n1303 vdd.n1279 681.178
R3758 vdd.n1304 vdd.n1303 681.178
R3759 vdd.n1306 vdd.n1304 681.178
R3760 vdd.n1295 vdd.n1294 681.178
R3761 vdd.n1296 vdd.n1295 681.178
R3762 vdd.n1296 vdd.n1275 681.178
R3763 vdd.n1312 vdd.n1275 681.178
R3764 vdd.n1312 vdd.n1311 681.178
R3765 vdd.n1311 vdd.n1310 681.178
R3766 vdd.n1334 vdd.n1327 681.178
R3767 vdd.n1343 vdd.n1327 681.178
R3768 vdd.n1343 vdd.n1325 681.178
R3769 vdd.n1349 vdd.n1325 681.178
R3770 vdd.n1350 vdd.n1349 681.178
R3771 vdd.n1352 vdd.n1350 681.178
R3772 vdd.n1341 vdd.n1340 681.178
R3773 vdd.n1342 vdd.n1341 681.178
R3774 vdd.n1342 vdd.n1321 681.178
R3775 vdd.n1358 vdd.n1321 681.178
R3776 vdd.n1358 vdd.n1357 681.178
R3777 vdd.n1357 vdd.n1356 681.178
R3778 vdd.n1380 vdd.n1373 681.178
R3779 vdd.n1389 vdd.n1373 681.178
R3780 vdd.n1389 vdd.n1371 681.178
R3781 vdd.n1395 vdd.n1371 681.178
R3782 vdd.n1396 vdd.n1395 681.178
R3783 vdd.n1398 vdd.n1396 681.178
R3784 vdd.n1387 vdd.n1386 681.178
R3785 vdd.n1388 vdd.n1387 681.178
R3786 vdd.n1388 vdd.n1367 681.178
R3787 vdd.n1404 vdd.n1367 681.178
R3788 vdd.n1404 vdd.n1403 681.178
R3789 vdd.n1403 vdd.n1402 681.178
R3790 vdd.n1477 vdd.n1470 681.178
R3791 vdd.n1486 vdd.n1470 681.178
R3792 vdd.n1486 vdd.n1468 681.178
R3793 vdd.n1492 vdd.n1468 681.178
R3794 vdd.n1493 vdd.n1492 681.178
R3795 vdd.n1495 vdd.n1493 681.178
R3796 vdd.n1484 vdd.n1483 681.178
R3797 vdd.n1485 vdd.n1484 681.178
R3798 vdd.n1485 vdd.n1464 681.178
R3799 vdd.n1501 vdd.n1464 681.178
R3800 vdd.n1501 vdd.n1500 681.178
R3801 vdd.n1500 vdd.n1499 681.178
R3802 vdd.n626 vdd.n619 681.178
R3803 vdd.n635 vdd.n619 681.178
R3804 vdd.n635 vdd.n617 681.178
R3805 vdd.n641 vdd.n617 681.178
R3806 vdd.n642 vdd.n641 681.178
R3807 vdd.n644 vdd.n642 681.178
R3808 vdd.n633 vdd.n632 681.178
R3809 vdd.n634 vdd.n633 681.178
R3810 vdd.n634 vdd.n613 681.178
R3811 vdd.n650 vdd.n613 681.178
R3812 vdd.n650 vdd.n649 681.178
R3813 vdd.n649 vdd.n648 681.178
R3814 vdd.n1521 vdd.n1514 681.178
R3815 vdd.n1530 vdd.n1514 681.178
R3816 vdd.n1530 vdd.n1512 681.178
R3817 vdd.n1536 vdd.n1512 681.178
R3818 vdd.n1537 vdd.n1536 681.178
R3819 vdd.n1539 vdd.n1537 681.178
R3820 vdd.n1528 vdd.n1527 681.178
R3821 vdd.n1529 vdd.n1528 681.178
R3822 vdd.n1529 vdd.n1508 681.178
R3823 vdd.n1545 vdd.n1508 681.178
R3824 vdd.n1545 vdd.n1544 681.178
R3825 vdd.n1544 vdd.n1543 681.178
R3826 vdd.n1566 vdd.n1559 681.178
R3827 vdd.n1575 vdd.n1559 681.178
R3828 vdd.n1575 vdd.n1557 681.178
R3829 vdd.n1581 vdd.n1557 681.178
R3830 vdd.n1582 vdd.n1581 681.178
R3831 vdd.n1584 vdd.n1582 681.178
R3832 vdd.n1573 vdd.n1572 681.178
R3833 vdd.n1574 vdd.n1573 681.178
R3834 vdd.n1574 vdd.n1553 681.178
R3835 vdd.n1590 vdd.n1553 681.178
R3836 vdd.n1590 vdd.n1589 681.178
R3837 vdd.n1589 vdd.n1588 681.178
R3838 vdd.n1616 vdd.n1609 681.178
R3839 vdd.n1625 vdd.n1609 681.178
R3840 vdd.n1625 vdd.n1607 681.178
R3841 vdd.n1631 vdd.n1607 681.178
R3842 vdd.n1632 vdd.n1631 681.178
R3843 vdd.n1634 vdd.n1632 681.178
R3844 vdd.n1623 vdd.n1622 681.178
R3845 vdd.n1624 vdd.n1623 681.178
R3846 vdd.n1624 vdd.n1603 681.178
R3847 vdd.n1640 vdd.n1603 681.178
R3848 vdd.n1640 vdd.n1639 681.178
R3849 vdd.n1639 vdd.n1638 681.178
R3850 vdd.n1662 vdd.n1655 681.178
R3851 vdd.n1671 vdd.n1655 681.178
R3852 vdd.n1671 vdd.n1653 681.178
R3853 vdd.n1677 vdd.n1653 681.178
R3854 vdd.n1678 vdd.n1677 681.178
R3855 vdd.n1680 vdd.n1678 681.178
R3856 vdd.n1669 vdd.n1668 681.178
R3857 vdd.n1670 vdd.n1669 681.178
R3858 vdd.n1670 vdd.n1649 681.178
R3859 vdd.n1686 vdd.n1649 681.178
R3860 vdd.n1686 vdd.n1685 681.178
R3861 vdd.n1685 vdd.n1684 681.178
R3862 vdd.n1710 vdd.n1703 681.178
R3863 vdd.n1719 vdd.n1703 681.178
R3864 vdd.n1719 vdd.n1701 681.178
R3865 vdd.n1725 vdd.n1701 681.178
R3866 vdd.n1726 vdd.n1725 681.178
R3867 vdd.n1728 vdd.n1726 681.178
R3868 vdd.n1717 vdd.n1716 681.178
R3869 vdd.n1718 vdd.n1717 681.178
R3870 vdd.n1718 vdd.n1697 681.178
R3871 vdd.n1734 vdd.n1697 681.178
R3872 vdd.n1734 vdd.n1733 681.178
R3873 vdd.n1733 vdd.n1732 681.178
R3874 vdd.n1430 vdd.n1429 681.178
R3875 vdd.n1431 vdd.n1430 681.178
R3876 vdd.n1431 vdd.n1424 681.178
R3877 vdd.n1437 vdd.n1424 681.178
R3878 vdd.n1438 vdd.n1437 681.178
R3879 vdd.n1440 vdd.n1438 681.178
R3880 vdd.n1453 vdd.n1452 681.178
R3881 vdd.n1452 vdd.n1451 681.178
R3882 vdd.n1451 vdd.n1415 681.178
R3883 vdd.n1446 vdd.n1415 681.178
R3884 vdd.n1446 vdd.n1445 681.178
R3885 vdd.n1445 vdd.n1444 681.178
R3886 vdd.n1757 vdd.n1750 681.178
R3887 vdd.n1766 vdd.n1750 681.178
R3888 vdd.n1766 vdd.n1748 681.178
R3889 vdd.n1772 vdd.n1748 681.178
R3890 vdd.n1773 vdd.n1772 681.178
R3891 vdd.n1775 vdd.n1773 681.178
R3892 vdd.n1764 vdd.n1763 681.178
R3893 vdd.n1765 vdd.n1764 681.178
R3894 vdd.n1765 vdd.n1744 681.178
R3895 vdd.n1781 vdd.n1744 681.178
R3896 vdd.n1781 vdd.n1780 681.178
R3897 vdd.n1780 vdd.n1779 681.178
R3898 vdd.n1802 vdd.n1795 681.178
R3899 vdd.n1811 vdd.n1795 681.178
R3900 vdd.n1811 vdd.n1793 681.178
R3901 vdd.n1817 vdd.n1793 681.178
R3902 vdd.n1818 vdd.n1817 681.178
R3903 vdd.n1820 vdd.n1818 681.178
R3904 vdd.n1809 vdd.n1808 681.178
R3905 vdd.n1810 vdd.n1809 681.178
R3906 vdd.n1810 vdd.n1789 681.178
R3907 vdd.n1826 vdd.n1789 681.178
R3908 vdd.n1826 vdd.n1825 681.178
R3909 vdd.n1825 vdd.n1824 681.178
R3910 vdd.n1848 vdd.n1841 681.178
R3911 vdd.n1857 vdd.n1841 681.178
R3912 vdd.n1857 vdd.n1839 681.178
R3913 vdd.n1863 vdd.n1839 681.178
R3914 vdd.n1864 vdd.n1863 681.178
R3915 vdd.n1866 vdd.n1864 681.178
R3916 vdd.n1855 vdd.n1854 681.178
R3917 vdd.n1856 vdd.n1855 681.178
R3918 vdd.n1856 vdd.n1835 681.178
R3919 vdd.n1872 vdd.n1835 681.178
R3920 vdd.n1872 vdd.n1871 681.178
R3921 vdd.n1871 vdd.n1870 681.178
R3922 vdd.n1899 vdd.n1892 681.178
R3923 vdd.n1908 vdd.n1892 681.178
R3924 vdd.n1908 vdd.n1890 681.178
R3925 vdd.n1914 vdd.n1890 681.178
R3926 vdd.n1915 vdd.n1914 681.178
R3927 vdd.n1917 vdd.n1915 681.178
R3928 vdd.n1906 vdd.n1905 681.178
R3929 vdd.n1907 vdd.n1906 681.178
R3930 vdd.n1907 vdd.n1886 681.178
R3931 vdd.n1923 vdd.n1886 681.178
R3932 vdd.n1923 vdd.n1922 681.178
R3933 vdd.n1922 vdd.n1921 681.178
R3934 vdd.n1945 vdd.n1938 681.178
R3935 vdd.n1954 vdd.n1938 681.178
R3936 vdd.n1954 vdd.n1936 681.178
R3937 vdd.n1960 vdd.n1936 681.178
R3938 vdd.n1961 vdd.n1960 681.178
R3939 vdd.n1963 vdd.n1961 681.178
R3940 vdd.n1952 vdd.n1951 681.178
R3941 vdd.n1953 vdd.n1952 681.178
R3942 vdd.n1953 vdd.n1932 681.178
R3943 vdd.n1969 vdd.n1932 681.178
R3944 vdd.n1969 vdd.n1968 681.178
R3945 vdd.n1968 vdd.n1967 681.178
R3946 vdd.n1993 vdd.n1986 681.178
R3947 vdd.n2002 vdd.n1986 681.178
R3948 vdd.n2002 vdd.n1984 681.178
R3949 vdd.n2008 vdd.n1984 681.178
R3950 vdd.n2009 vdd.n2008 681.178
R3951 vdd.n2011 vdd.n2009 681.178
R3952 vdd.n2000 vdd.n1999 681.178
R3953 vdd.n2001 vdd.n2000 681.178
R3954 vdd.n2001 vdd.n1980 681.178
R3955 vdd.n2017 vdd.n1980 681.178
R3956 vdd.n2017 vdd.n2016 681.178
R3957 vdd.n2016 vdd.n2015 681.178
R3958 vdd.n2039 vdd.n2032 681.178
R3959 vdd.n2048 vdd.n2032 681.178
R3960 vdd.n2048 vdd.n2030 681.178
R3961 vdd.n2054 vdd.n2030 681.178
R3962 vdd.n2055 vdd.n2054 681.178
R3963 vdd.n2057 vdd.n2055 681.178
R3964 vdd.n2046 vdd.n2045 681.178
R3965 vdd.n2047 vdd.n2046 681.178
R3966 vdd.n2047 vdd.n2026 681.178
R3967 vdd.n2063 vdd.n2026 681.178
R3968 vdd.n2063 vdd.n2062 681.178
R3969 vdd.n2062 vdd.n2061 681.178
R3970 vdd.n2084 vdd.n2077 681.178
R3971 vdd.n2093 vdd.n2077 681.178
R3972 vdd.n2093 vdd.n2075 681.178
R3973 vdd.n2099 vdd.n2075 681.178
R3974 vdd.n2100 vdd.n2099 681.178
R3975 vdd.n2102 vdd.n2100 681.178
R3976 vdd.n2091 vdd.n2090 681.178
R3977 vdd.n2092 vdd.n2091 681.178
R3978 vdd.n2092 vdd.n2071 681.178
R3979 vdd.n2108 vdd.n2071 681.178
R3980 vdd.n2108 vdd.n2107 681.178
R3981 vdd.n2107 vdd.n2106 681.178
R3982 vdd.n2134 vdd.n2127 681.178
R3983 vdd.n2143 vdd.n2127 681.178
R3984 vdd.n2143 vdd.n2125 681.178
R3985 vdd.n2149 vdd.n2125 681.178
R3986 vdd.n2150 vdd.n2149 681.178
R3987 vdd.n2152 vdd.n2150 681.178
R3988 vdd.n2141 vdd.n2140 681.178
R3989 vdd.n2142 vdd.n2141 681.178
R3990 vdd.n2142 vdd.n2121 681.178
R3991 vdd.n2158 vdd.n2121 681.178
R3992 vdd.n2158 vdd.n2157 681.178
R3993 vdd.n2157 vdd.n2156 681.178
R3994 vdd.n2180 vdd.n2173 681.178
R3995 vdd.n2189 vdd.n2173 681.178
R3996 vdd.n2189 vdd.n2171 681.178
R3997 vdd.n2195 vdd.n2171 681.178
R3998 vdd.n2196 vdd.n2195 681.178
R3999 vdd.n2198 vdd.n2196 681.178
R4000 vdd.n2187 vdd.n2186 681.178
R4001 vdd.n2188 vdd.n2187 681.178
R4002 vdd.n2188 vdd.n2167 681.178
R4003 vdd.n2204 vdd.n2167 681.178
R4004 vdd.n2204 vdd.n2203 681.178
R4005 vdd.n2203 vdd.n2202 681.178
R4006 vdd.n2228 vdd.n2221 681.178
R4007 vdd.n2237 vdd.n2221 681.178
R4008 vdd.n2237 vdd.n2219 681.178
R4009 vdd.n2243 vdd.n2219 681.178
R4010 vdd.n2244 vdd.n2243 681.178
R4011 vdd.n2246 vdd.n2244 681.178
R4012 vdd.n2235 vdd.n2234 681.178
R4013 vdd.n2236 vdd.n2235 681.178
R4014 vdd.n2236 vdd.n2215 681.178
R4015 vdd.n2252 vdd.n2215 681.178
R4016 vdd.n2252 vdd.n2251 681.178
R4017 vdd.n2251 vdd.n2250 681.178
R4018 vdd.n1195 vdd.n1194 681.178
R4019 vdd.n1196 vdd.n1195 681.178
R4020 vdd.n1196 vdd.n1189 681.178
R4021 vdd.n1202 vdd.n1189 681.178
R4022 vdd.n1203 vdd.n1202 681.178
R4023 vdd.n1205 vdd.n1203 681.178
R4024 vdd.n1218 vdd.n1217 681.178
R4025 vdd.n1217 vdd.n1216 681.178
R4026 vdd.n1216 vdd.n1180 681.178
R4027 vdd.n1211 vdd.n1180 681.178
R4028 vdd.n1211 vdd.n1210 681.178
R4029 vdd.n1210 vdd.n1209 681.178
R4030 vdd.n2275 vdd.n2268 681.178
R4031 vdd.n2284 vdd.n2268 681.178
R4032 vdd.n2284 vdd.n2266 681.178
R4033 vdd.n2290 vdd.n2266 681.178
R4034 vdd.n2291 vdd.n2290 681.178
R4035 vdd.n2293 vdd.n2291 681.178
R4036 vdd.n2282 vdd.n2281 681.178
R4037 vdd.n2283 vdd.n2282 681.178
R4038 vdd.n2283 vdd.n2262 681.178
R4039 vdd.n2299 vdd.n2262 681.178
R4040 vdd.n2299 vdd.n2298 681.178
R4041 vdd.n2298 vdd.n2297 681.178
R4042 vdd.n2320 vdd.n2313 681.178
R4043 vdd.n2329 vdd.n2313 681.178
R4044 vdd.n2329 vdd.n2311 681.178
R4045 vdd.n2335 vdd.n2311 681.178
R4046 vdd.n2336 vdd.n2335 681.178
R4047 vdd.n2338 vdd.n2336 681.178
R4048 vdd.n2327 vdd.n2326 681.178
R4049 vdd.n2328 vdd.n2327 681.178
R4050 vdd.n2328 vdd.n2307 681.178
R4051 vdd.n2344 vdd.n2307 681.178
R4052 vdd.n2344 vdd.n2343 681.178
R4053 vdd.n2343 vdd.n2342 681.178
R4054 vdd.n2370 vdd.n2363 681.178
R4055 vdd.n2379 vdd.n2363 681.178
R4056 vdd.n2379 vdd.n2361 681.178
R4057 vdd.n2385 vdd.n2361 681.178
R4058 vdd.n2386 vdd.n2385 681.178
R4059 vdd.n2388 vdd.n2386 681.178
R4060 vdd.n2377 vdd.n2376 681.178
R4061 vdd.n2378 vdd.n2377 681.178
R4062 vdd.n2378 vdd.n2357 681.178
R4063 vdd.n2394 vdd.n2357 681.178
R4064 vdd.n2394 vdd.n2393 681.178
R4065 vdd.n2393 vdd.n2392 681.178
R4066 vdd.n2416 vdd.n2409 681.178
R4067 vdd.n2425 vdd.n2409 681.178
R4068 vdd.n2425 vdd.n2407 681.178
R4069 vdd.n2431 vdd.n2407 681.178
R4070 vdd.n2432 vdd.n2431 681.178
R4071 vdd.n2434 vdd.n2432 681.178
R4072 vdd.n2423 vdd.n2422 681.178
R4073 vdd.n2424 vdd.n2423 681.178
R4074 vdd.n2424 vdd.n2403 681.178
R4075 vdd.n2440 vdd.n2403 681.178
R4076 vdd.n2440 vdd.n2439 681.178
R4077 vdd.n2439 vdd.n2438 681.178
R4078 vdd.n2464 vdd.n2457 681.178
R4079 vdd.n2473 vdd.n2457 681.178
R4080 vdd.n2473 vdd.n2455 681.178
R4081 vdd.n2479 vdd.n2455 681.178
R4082 vdd.n2480 vdd.n2479 681.178
R4083 vdd.n2482 vdd.n2480 681.178
R4084 vdd.n2471 vdd.n2470 681.178
R4085 vdd.n2472 vdd.n2471 681.178
R4086 vdd.n2472 vdd.n2451 681.178
R4087 vdd.n2488 vdd.n2451 681.178
R4088 vdd.n2488 vdd.n2487 681.178
R4089 vdd.n2487 vdd.n2486 681.178
R4090 vdd.n2610 vdd.n2609 681.178
R4091 vdd.n2611 vdd.n2610 681.178
R4092 vdd.n2611 vdd.n2589 681.178
R4093 vdd.n2626 vdd.n2589 681.178
R4094 vdd.n2626 vdd.n2590 681.178
R4095 vdd.n2618 vdd.n2590 681.178
R4096 vdd.n2603 vdd.n2596 681.178
R4097 vdd.n2612 vdd.n2596 681.178
R4098 vdd.n2612 vdd.n2598 681.178
R4099 vdd.n2598 vdd.n2592 681.178
R4100 vdd.n2623 vdd.n2592 681.178
R4101 vdd.n2623 vdd.n2622 681.178
R4102 vdd.n2564 vdd.n2563 681.178
R4103 vdd.n2565 vdd.n2564 681.178
R4104 vdd.n2565 vdd.n2543 681.178
R4105 vdd.n2580 vdd.n2543 681.178
R4106 vdd.n2580 vdd.n2544 681.178
R4107 vdd.n2572 vdd.n2544 681.178
R4108 vdd.n2557 vdd.n2550 681.178
R4109 vdd.n2566 vdd.n2550 681.178
R4110 vdd.n2566 vdd.n2552 681.178
R4111 vdd.n2552 vdd.n2546 681.178
R4112 vdd.n2577 vdd.n2546 681.178
R4113 vdd.n2577 vdd.n2576 681.178
R4114 vdd.n2657 vdd.n2656 681.178
R4115 vdd.n2658 vdd.n2657 681.178
R4116 vdd.n2658 vdd.n2636 681.178
R4117 vdd.n2673 vdd.n2636 681.178
R4118 vdd.n2673 vdd.n2637 681.178
R4119 vdd.n2665 vdd.n2637 681.178
R4120 vdd.n2650 vdd.n2643 681.178
R4121 vdd.n2659 vdd.n2643 681.178
R4122 vdd.n2659 vdd.n2645 681.178
R4123 vdd.n2645 vdd.n2639 681.178
R4124 vdd.n2670 vdd.n2639 681.178
R4125 vdd.n2670 vdd.n2669 681.178
R4126 vdd.n2705 vdd.n2704 681.178
R4127 vdd.n2706 vdd.n2705 681.178
R4128 vdd.n2706 vdd.n2684 681.178
R4129 vdd.n2721 vdd.n2684 681.178
R4130 vdd.n2721 vdd.n2685 681.178
R4131 vdd.n2713 vdd.n2685 681.178
R4132 vdd.n2698 vdd.n2691 681.178
R4133 vdd.n2707 vdd.n2691 681.178
R4134 vdd.n2707 vdd.n2693 681.178
R4135 vdd.n2693 vdd.n2687 681.178
R4136 vdd.n2718 vdd.n2687 681.178
R4137 vdd.n2718 vdd.n2717 681.178
R4138 vdd.n2751 vdd.n2750 681.178
R4139 vdd.n2752 vdd.n2751 681.178
R4140 vdd.n2752 vdd.n2730 681.178
R4141 vdd.n2767 vdd.n2730 681.178
R4142 vdd.n2767 vdd.n2731 681.178
R4143 vdd.n2759 vdd.n2731 681.178
R4144 vdd.n2744 vdd.n2737 681.178
R4145 vdd.n2753 vdd.n2737 681.178
R4146 vdd.n2753 vdd.n2739 681.178
R4147 vdd.n2739 vdd.n2733 681.178
R4148 vdd.n2764 vdd.n2733 681.178
R4149 vdd.n2764 vdd.n2763 681.178
R4150 vdd.n1005 vdd.n993 681.178
R4151 vdd.n1015 vdd.n993 681.178
R4152 vdd.n1015 vdd.n994 681.178
R4153 vdd.n994 vdd.n990 681.178
R4154 vdd.n1024 vdd.n990 681.178
R4155 vdd.n1025 vdd.n1024 681.178
R4156 vdd.n1007 vdd.n1003 681.178
R4157 vdd.n1003 vdd.n996 681.178
R4158 vdd.n998 vdd.n996 681.178
R4159 vdd.n1013 vdd.n998 681.178
R4160 vdd.n1013 vdd.n988 681.178
R4161 vdd.n1027 vdd.n988 681.178
R4162 vdd.n2893 vdd.n2892 681.178
R4163 vdd.n2894 vdd.n2893 681.178
R4164 vdd.n2894 vdd.n2872 681.178
R4165 vdd.n2909 vdd.n2872 681.178
R4166 vdd.n2909 vdd.n2873 681.178
R4167 vdd.n2901 vdd.n2873 681.178
R4168 vdd.n2886 vdd.n2879 681.178
R4169 vdd.n2895 vdd.n2879 681.178
R4170 vdd.n2895 vdd.n2881 681.178
R4171 vdd.n2881 vdd.n2875 681.178
R4172 vdd.n2906 vdd.n2875 681.178
R4173 vdd.n2906 vdd.n2905 681.178
R4174 vdd.n2846 vdd.n2845 681.178
R4175 vdd.n2847 vdd.n2846 681.178
R4176 vdd.n2847 vdd.n2825 681.178
R4177 vdd.n2862 vdd.n2825 681.178
R4178 vdd.n2862 vdd.n2826 681.178
R4179 vdd.n2854 vdd.n2826 681.178
R4180 vdd.n2839 vdd.n2832 681.178
R4181 vdd.n2848 vdd.n2832 681.178
R4182 vdd.n2848 vdd.n2834 681.178
R4183 vdd.n2834 vdd.n2828 681.178
R4184 vdd.n2859 vdd.n2828 681.178
R4185 vdd.n2859 vdd.n2858 681.178
R4186 vdd.n2800 vdd.n2799 681.178
R4187 vdd.n2801 vdd.n2800 681.178
R4188 vdd.n2801 vdd.n2779 681.178
R4189 vdd.n2816 vdd.n2779 681.178
R4190 vdd.n2816 vdd.n2780 681.178
R4191 vdd.n2808 vdd.n2780 681.178
R4192 vdd.n2793 vdd.n2786 681.178
R4193 vdd.n2802 vdd.n2786 681.178
R4194 vdd.n2802 vdd.n2788 681.178
R4195 vdd.n2788 vdd.n2782 681.178
R4196 vdd.n2813 vdd.n2782 681.178
R4197 vdd.n2813 vdd.n2812 681.178
R4198 vdd.n2940 vdd.n2939 681.178
R4199 vdd.n2941 vdd.n2940 681.178
R4200 vdd.n2941 vdd.n2919 681.178
R4201 vdd.n2956 vdd.n2919 681.178
R4202 vdd.n2956 vdd.n2920 681.178
R4203 vdd.n2948 vdd.n2920 681.178
R4204 vdd.n2933 vdd.n2926 681.178
R4205 vdd.n2942 vdd.n2926 681.178
R4206 vdd.n2942 vdd.n2928 681.178
R4207 vdd.n2928 vdd.n2922 681.178
R4208 vdd.n2953 vdd.n2922 681.178
R4209 vdd.n2953 vdd.n2952 681.178
R4210 vdd.n2988 vdd.n2987 681.178
R4211 vdd.n2989 vdd.n2988 681.178
R4212 vdd.n2989 vdd.n2967 681.178
R4213 vdd.n3004 vdd.n2967 681.178
R4214 vdd.n3004 vdd.n2968 681.178
R4215 vdd.n2996 vdd.n2968 681.178
R4216 vdd.n2981 vdd.n2974 681.178
R4217 vdd.n2990 vdd.n2974 681.178
R4218 vdd.n2990 vdd.n2976 681.178
R4219 vdd.n2976 vdd.n2970 681.178
R4220 vdd.n3001 vdd.n2970 681.178
R4221 vdd.n3001 vdd.n3000 681.178
R4222 vdd.n3034 vdd.n3033 681.178
R4223 vdd.n3035 vdd.n3034 681.178
R4224 vdd.n3035 vdd.n3013 681.178
R4225 vdd.n3050 vdd.n3013 681.178
R4226 vdd.n3050 vdd.n3014 681.178
R4227 vdd.n3042 vdd.n3014 681.178
R4228 vdd.n3027 vdd.n3020 681.178
R4229 vdd.n3036 vdd.n3020 681.178
R4230 vdd.n3036 vdd.n3022 681.178
R4231 vdd.n3022 vdd.n3016 681.178
R4232 vdd.n3047 vdd.n3016 681.178
R4233 vdd.n3047 vdd.n3046 681.178
R4234 vdd.n3128 vdd.n3127 681.178
R4235 vdd.n3129 vdd.n3128 681.178
R4236 vdd.n3129 vdd.n3107 681.178
R4237 vdd.n3144 vdd.n3107 681.178
R4238 vdd.n3144 vdd.n3108 681.178
R4239 vdd.n3136 vdd.n3108 681.178
R4240 vdd.n3121 vdd.n3114 681.178
R4241 vdd.n3130 vdd.n3114 681.178
R4242 vdd.n3130 vdd.n3116 681.178
R4243 vdd.n3116 vdd.n3110 681.178
R4244 vdd.n3141 vdd.n3110 681.178
R4245 vdd.n3141 vdd.n3140 681.178
R4246 vdd.n3082 vdd.n3081 681.178
R4247 vdd.n3083 vdd.n3082 681.178
R4248 vdd.n3083 vdd.n3061 681.178
R4249 vdd.n3098 vdd.n3061 681.178
R4250 vdd.n3098 vdd.n3062 681.178
R4251 vdd.n3090 vdd.n3062 681.178
R4252 vdd.n3075 vdd.n3068 681.178
R4253 vdd.n3084 vdd.n3068 681.178
R4254 vdd.n3084 vdd.n3070 681.178
R4255 vdd.n3070 vdd.n3064 681.178
R4256 vdd.n3095 vdd.n3064 681.178
R4257 vdd.n3095 vdd.n3094 681.178
R4258 vdd.n3175 vdd.n3174 681.178
R4259 vdd.n3176 vdd.n3175 681.178
R4260 vdd.n3176 vdd.n3154 681.178
R4261 vdd.n3191 vdd.n3154 681.178
R4262 vdd.n3191 vdd.n3155 681.178
R4263 vdd.n3183 vdd.n3155 681.178
R4264 vdd.n3168 vdd.n3161 681.178
R4265 vdd.n3177 vdd.n3161 681.178
R4266 vdd.n3177 vdd.n3163 681.178
R4267 vdd.n3163 vdd.n3157 681.178
R4268 vdd.n3188 vdd.n3157 681.178
R4269 vdd.n3188 vdd.n3187 681.178
R4270 vdd.n3223 vdd.n3222 681.178
R4271 vdd.n3224 vdd.n3223 681.178
R4272 vdd.n3224 vdd.n3202 681.178
R4273 vdd.n3239 vdd.n3202 681.178
R4274 vdd.n3239 vdd.n3203 681.178
R4275 vdd.n3231 vdd.n3203 681.178
R4276 vdd.n3216 vdd.n3209 681.178
R4277 vdd.n3225 vdd.n3209 681.178
R4278 vdd.n3225 vdd.n3211 681.178
R4279 vdd.n3211 vdd.n3205 681.178
R4280 vdd.n3236 vdd.n3205 681.178
R4281 vdd.n3236 vdd.n3235 681.178
R4282 vdd.n3269 vdd.n3268 681.178
R4283 vdd.n3270 vdd.n3269 681.178
R4284 vdd.n3270 vdd.n3248 681.178
R4285 vdd.n3285 vdd.n3248 681.178
R4286 vdd.n3285 vdd.n3249 681.178
R4287 vdd.n3277 vdd.n3249 681.178
R4288 vdd.n3262 vdd.n3255 681.178
R4289 vdd.n3271 vdd.n3255 681.178
R4290 vdd.n3271 vdd.n3257 681.178
R4291 vdd.n3257 vdd.n3251 681.178
R4292 vdd.n3282 vdd.n3251 681.178
R4293 vdd.n3282 vdd.n3281 681.178
R4294 vdd.n769 vdd.n757 681.178
R4295 vdd.n779 vdd.n757 681.178
R4296 vdd.n779 vdd.n758 681.178
R4297 vdd.n758 vdd.n754 681.178
R4298 vdd.n788 vdd.n754 681.178
R4299 vdd.n789 vdd.n788 681.178
R4300 vdd.n771 vdd.n767 681.178
R4301 vdd.n767 vdd.n760 681.178
R4302 vdd.n762 vdd.n760 681.178
R4303 vdd.n777 vdd.n762 681.178
R4304 vdd.n777 vdd.n752 681.178
R4305 vdd.n791 vdd.n752 681.178
R4306 vdd.n3364 vdd.n3363 681.178
R4307 vdd.n3365 vdd.n3364 681.178
R4308 vdd.n3365 vdd.n3343 681.178
R4309 vdd.n3380 vdd.n3343 681.178
R4310 vdd.n3380 vdd.n3344 681.178
R4311 vdd.n3372 vdd.n3344 681.178
R4312 vdd.n3357 vdd.n3350 681.178
R4313 vdd.n3366 vdd.n3350 681.178
R4314 vdd.n3366 vdd.n3352 681.178
R4315 vdd.n3352 vdd.n3346 681.178
R4316 vdd.n3377 vdd.n3346 681.178
R4317 vdd.n3377 vdd.n3376 681.178
R4318 vdd.n3318 vdd.n3317 681.178
R4319 vdd.n3319 vdd.n3318 681.178
R4320 vdd.n3319 vdd.n3297 681.178
R4321 vdd.n3334 vdd.n3297 681.178
R4322 vdd.n3334 vdd.n3298 681.178
R4323 vdd.n3326 vdd.n3298 681.178
R4324 vdd.n3311 vdd.n3304 681.178
R4325 vdd.n3320 vdd.n3304 681.178
R4326 vdd.n3320 vdd.n3306 681.178
R4327 vdd.n3306 vdd.n3300 681.178
R4328 vdd.n3331 vdd.n3300 681.178
R4329 vdd.n3331 vdd.n3330 681.178
R4330 vdd.n3411 vdd.n3410 681.178
R4331 vdd.n3412 vdd.n3411 681.178
R4332 vdd.n3412 vdd.n3390 681.178
R4333 vdd.n3427 vdd.n3390 681.178
R4334 vdd.n3427 vdd.n3391 681.178
R4335 vdd.n3419 vdd.n3391 681.178
R4336 vdd.n3404 vdd.n3397 681.178
R4337 vdd.n3413 vdd.n3397 681.178
R4338 vdd.n3413 vdd.n3399 681.178
R4339 vdd.n3399 vdd.n3393 681.178
R4340 vdd.n3424 vdd.n3393 681.178
R4341 vdd.n3424 vdd.n3423 681.178
R4342 vdd.n3459 vdd.n3458 681.178
R4343 vdd.n3460 vdd.n3459 681.178
R4344 vdd.n3460 vdd.n3438 681.178
R4345 vdd.n3475 vdd.n3438 681.178
R4346 vdd.n3475 vdd.n3439 681.178
R4347 vdd.n3467 vdd.n3439 681.178
R4348 vdd.n3452 vdd.n3445 681.178
R4349 vdd.n3461 vdd.n3445 681.178
R4350 vdd.n3461 vdd.n3447 681.178
R4351 vdd.n3447 vdd.n3441 681.178
R4352 vdd.n3472 vdd.n3441 681.178
R4353 vdd.n3472 vdd.n3471 681.178
R4354 vdd.n3505 vdd.n3504 681.178
R4355 vdd.n3506 vdd.n3505 681.178
R4356 vdd.n3506 vdd.n3484 681.178
R4357 vdd.n3521 vdd.n3484 681.178
R4358 vdd.n3521 vdd.n3485 681.178
R4359 vdd.n3513 vdd.n3485 681.178
R4360 vdd.n3498 vdd.n3491 681.178
R4361 vdd.n3507 vdd.n3491 681.178
R4362 vdd.n3507 vdd.n3493 681.178
R4363 vdd.n3493 vdd.n3487 681.178
R4364 vdd.n3518 vdd.n3487 681.178
R4365 vdd.n3518 vdd.n3517 681.178
R4366 vdd.n587 vdd.n586 681.178
R4367 vdd.n588 vdd.n587 681.178
R4368 vdd.n588 vdd.n566 681.178
R4369 vdd.n603 vdd.n566 681.178
R4370 vdd.n603 vdd.n567 681.178
R4371 vdd.n595 vdd.n567 681.178
R4372 vdd.n580 vdd.n573 681.178
R4373 vdd.n589 vdd.n573 681.178
R4374 vdd.n589 vdd.n575 681.178
R4375 vdd.n575 vdd.n569 681.178
R4376 vdd.n600 vdd.n569 681.178
R4377 vdd.n600 vdd.n599 681.178
R4378 vdd.n3600 vdd.n3599 681.178
R4379 vdd.n3601 vdd.n3600 681.178
R4380 vdd.n3601 vdd.n3579 681.178
R4381 vdd.n3616 vdd.n3579 681.178
R4382 vdd.n3616 vdd.n3580 681.178
R4383 vdd.n3608 vdd.n3580 681.178
R4384 vdd.n3593 vdd.n3586 681.178
R4385 vdd.n3602 vdd.n3586 681.178
R4386 vdd.n3602 vdd.n3588 681.178
R4387 vdd.n3588 vdd.n3582 681.178
R4388 vdd.n3613 vdd.n3582 681.178
R4389 vdd.n3613 vdd.n3612 681.178
R4390 vdd.n3554 vdd.n3553 681.178
R4391 vdd.n3555 vdd.n3554 681.178
R4392 vdd.n3555 vdd.n3533 681.178
R4393 vdd.n3570 vdd.n3533 681.178
R4394 vdd.n3570 vdd.n3534 681.178
R4395 vdd.n3562 vdd.n3534 681.178
R4396 vdd.n3547 vdd.n3540 681.178
R4397 vdd.n3556 vdd.n3540 681.178
R4398 vdd.n3556 vdd.n3542 681.178
R4399 vdd.n3542 vdd.n3536 681.178
R4400 vdd.n3567 vdd.n3536 681.178
R4401 vdd.n3567 vdd.n3566 681.178
R4402 vdd.n6614 vdd.n6613 681.178
R4403 vdd.n6615 vdd.n6614 681.178
R4404 vdd.n6615 vdd.n6593 681.178
R4405 vdd.n6630 vdd.n6593 681.178
R4406 vdd.n6630 vdd.n6594 681.178
R4407 vdd.n6622 vdd.n6594 681.178
R4408 vdd.n6607 vdd.n6600 681.178
R4409 vdd.n6616 vdd.n6600 681.178
R4410 vdd.n6616 vdd.n6602 681.178
R4411 vdd.n6602 vdd.n6596 681.178
R4412 vdd.n6627 vdd.n6596 681.178
R4413 vdd.n6627 vdd.n6626 681.178
R4414 vdd.n6568 vdd.n6567 681.178
R4415 vdd.n6569 vdd.n6568 681.178
R4416 vdd.n6569 vdd.n6547 681.178
R4417 vdd.n6584 vdd.n6547 681.178
R4418 vdd.n6584 vdd.n6548 681.178
R4419 vdd.n6576 vdd.n6548 681.178
R4420 vdd.n6561 vdd.n6554 681.178
R4421 vdd.n6570 vdd.n6554 681.178
R4422 vdd.n6570 vdd.n6556 681.178
R4423 vdd.n6556 vdd.n6550 681.178
R4424 vdd.n6581 vdd.n6550 681.178
R4425 vdd.n6581 vdd.n6580 681.178
R4426 vdd.n9628 vdd.n9627 681.178
R4427 vdd.n9629 vdd.n9628 681.178
R4428 vdd.n9629 vdd.n9607 681.178
R4429 vdd.n9644 vdd.n9607 681.178
R4430 vdd.n9644 vdd.n9608 681.178
R4431 vdd.n9636 vdd.n9608 681.178
R4432 vdd.n9621 vdd.n9614 681.178
R4433 vdd.n9630 vdd.n9614 681.178
R4434 vdd.n9630 vdd.n9616 681.178
R4435 vdd.n9616 vdd.n9610 681.178
R4436 vdd.n9641 vdd.n9610 681.178
R4437 vdd.n9641 vdd.n9640 681.178
R4438 vdd.n9582 vdd.n9581 681.178
R4439 vdd.n9583 vdd.n9582 681.178
R4440 vdd.n9583 vdd.n9561 681.178
R4441 vdd.n9598 vdd.n9561 681.178
R4442 vdd.n9598 vdd.n9562 681.178
R4443 vdd.n9590 vdd.n9562 681.178
R4444 vdd.n9575 vdd.n9568 681.178
R4445 vdd.n9584 vdd.n9568 681.178
R4446 vdd.n9584 vdd.n9570 681.178
R4447 vdd.n9570 vdd.n9564 681.178
R4448 vdd.n9595 vdd.n9564 681.178
R4449 vdd.n9595 vdd.n9594 681.178
R4450 vdd.n9674 vdd.n9673 681.178
R4451 vdd.n9675 vdd.n9674 681.178
R4452 vdd.n9675 vdd.n9653 681.178
R4453 vdd.n9690 vdd.n9653 681.178
R4454 vdd.n9690 vdd.n9654 681.178
R4455 vdd.n9682 vdd.n9654 681.178
R4456 vdd.n9667 vdd.n9660 681.178
R4457 vdd.n9676 vdd.n9660 681.178
R4458 vdd.n9676 vdd.n9662 681.178
R4459 vdd.n9662 vdd.n9656 681.178
R4460 vdd.n9687 vdd.n9656 681.178
R4461 vdd.n9687 vdd.n9686 681.178
R4462 vdd.n9720 vdd.n9719 681.178
R4463 vdd.n9721 vdd.n9720 681.178
R4464 vdd.n9721 vdd.n9699 681.178
R4465 vdd.n9736 vdd.n9699 681.178
R4466 vdd.n9736 vdd.n9700 681.178
R4467 vdd.n9728 vdd.n9700 681.178
R4468 vdd.n9713 vdd.n9706 681.178
R4469 vdd.n9722 vdd.n9706 681.178
R4470 vdd.n9722 vdd.n9708 681.178
R4471 vdd.n9708 vdd.n9702 681.178
R4472 vdd.n9733 vdd.n9702 681.178
R4473 vdd.n9733 vdd.n9732 681.178
R4474 vdd.n9818 vdd.n9817 681.178
R4475 vdd.n9819 vdd.n9818 681.178
R4476 vdd.n9819 vdd.n9797 681.178
R4477 vdd.n9834 vdd.n9797 681.178
R4478 vdd.n9834 vdd.n9798 681.178
R4479 vdd.n9826 vdd.n9798 681.178
R4480 vdd.n9811 vdd.n9804 681.178
R4481 vdd.n9820 vdd.n9804 681.178
R4482 vdd.n9820 vdd.n9806 681.178
R4483 vdd.n9806 vdd.n9800 681.178
R4484 vdd.n9831 vdd.n9800 681.178
R4485 vdd.n9831 vdd.n9830 681.178
R4486 vdd.n9864 vdd.n9863 681.178
R4487 vdd.n9865 vdd.n9864 681.178
R4488 vdd.n9865 vdd.n9843 681.178
R4489 vdd.n9880 vdd.n9843 681.178
R4490 vdd.n9880 vdd.n9844 681.178
R4491 vdd.n9872 vdd.n9844 681.178
R4492 vdd.n9857 vdd.n9850 681.178
R4493 vdd.n9866 vdd.n9850 681.178
R4494 vdd.n9866 vdd.n9852 681.178
R4495 vdd.n9852 vdd.n9846 681.178
R4496 vdd.n9877 vdd.n9846 681.178
R4497 vdd.n9877 vdd.n9876 681.178
R4498 vdd.n9910 vdd.n9909 681.178
R4499 vdd.n9911 vdd.n9910 681.178
R4500 vdd.n9911 vdd.n9889 681.178
R4501 vdd.n9926 vdd.n9889 681.178
R4502 vdd.n9926 vdd.n9890 681.178
R4503 vdd.n9918 vdd.n9890 681.178
R4504 vdd.n9903 vdd.n9896 681.178
R4505 vdd.n9912 vdd.n9896 681.178
R4506 vdd.n9912 vdd.n9898 681.178
R4507 vdd.n9898 vdd.n9892 681.178
R4508 vdd.n9923 vdd.n9892 681.178
R4509 vdd.n9923 vdd.n9922 681.178
R4510 vdd.n9956 vdd.n9955 681.178
R4511 vdd.n9957 vdd.n9956 681.178
R4512 vdd.n9957 vdd.n9935 681.178
R4513 vdd.n9972 vdd.n9935 681.178
R4514 vdd.n9972 vdd.n9936 681.178
R4515 vdd.n9964 vdd.n9936 681.178
R4516 vdd.n9949 vdd.n9942 681.178
R4517 vdd.n9958 vdd.n9942 681.178
R4518 vdd.n9958 vdd.n9944 681.178
R4519 vdd.n9944 vdd.n9938 681.178
R4520 vdd.n9969 vdd.n9938 681.178
R4521 vdd.n9969 vdd.n9968 681.178
R4522 vdd.n10054 vdd.n10053 681.178
R4523 vdd.n10055 vdd.n10054 681.178
R4524 vdd.n10055 vdd.n10033 681.178
R4525 vdd.n10070 vdd.n10033 681.178
R4526 vdd.n10070 vdd.n10034 681.178
R4527 vdd.n10062 vdd.n10034 681.178
R4528 vdd.n10047 vdd.n10040 681.178
R4529 vdd.n10056 vdd.n10040 681.178
R4530 vdd.n10056 vdd.n10042 681.178
R4531 vdd.n10042 vdd.n10036 681.178
R4532 vdd.n10067 vdd.n10036 681.178
R4533 vdd.n10067 vdd.n10066 681.178
R4534 vdd.n70 vdd.n69 681.178
R4535 vdd.n71 vdd.n70 681.178
R4536 vdd.n71 vdd.n49 681.178
R4537 vdd.n86 vdd.n49 681.178
R4538 vdd.n86 vdd.n50 681.178
R4539 vdd.n78 vdd.n50 681.178
R4540 vdd.n63 vdd.n56 681.178
R4541 vdd.n72 vdd.n56 681.178
R4542 vdd.n72 vdd.n58 681.178
R4543 vdd.n58 vdd.n52 681.178
R4544 vdd.n83 vdd.n52 681.178
R4545 vdd.n83 vdd.n82 681.178
R4546 vdd.n24 vdd.n23 681.178
R4547 vdd.n25 vdd.n24 681.178
R4548 vdd.n25 vdd.n3 681.178
R4549 vdd.n40 vdd.n3 681.178
R4550 vdd.n40 vdd.n4 681.178
R4551 vdd.n32 vdd.n4 681.178
R4552 vdd.n17 vdd.n10 681.178
R4553 vdd.n26 vdd.n10 681.178
R4554 vdd.n26 vdd.n12 681.178
R4555 vdd.n12 vdd.n6 681.178
R4556 vdd.n37 vdd.n6 681.178
R4557 vdd.n37 vdd.n36 681.178
R4558 vdd.n10100 vdd.n10099 681.178
R4559 vdd.n10101 vdd.n10100 681.178
R4560 vdd.n10101 vdd.n10079 681.178
R4561 vdd.n10116 vdd.n10079 681.178
R4562 vdd.n10116 vdd.n10080 681.178
R4563 vdd.n10108 vdd.n10080 681.178
R4564 vdd.n10093 vdd.n10086 681.178
R4565 vdd.n10102 vdd.n10086 681.178
R4566 vdd.n10102 vdd.n10088 681.178
R4567 vdd.n10088 vdd.n10082 681.178
R4568 vdd.n10113 vdd.n10082 681.178
R4569 vdd.n10113 vdd.n10112 681.178
R4570 vdd.n10148 vdd.n10147 681.178
R4571 vdd.n10149 vdd.n10148 681.178
R4572 vdd.n10149 vdd.n10127 681.178
R4573 vdd.n10164 vdd.n10127 681.178
R4574 vdd.n10164 vdd.n10128 681.178
R4575 vdd.n10156 vdd.n10128 681.178
R4576 vdd.n10141 vdd.n10134 681.178
R4577 vdd.n10150 vdd.n10134 681.178
R4578 vdd.n10150 vdd.n10136 681.178
R4579 vdd.n10136 vdd.n10130 681.178
R4580 vdd.n10161 vdd.n10130 681.178
R4581 vdd.n10161 vdd.n10160 681.178
R4582 vdd.n10194 vdd.n10193 681.178
R4583 vdd.n10195 vdd.n10194 681.178
R4584 vdd.n10195 vdd.n10173 681.178
R4585 vdd.n10210 vdd.n10173 681.178
R4586 vdd.n10210 vdd.n10174 681.178
R4587 vdd.n10202 vdd.n10174 681.178
R4588 vdd.n10187 vdd.n10180 681.178
R4589 vdd.n10196 vdd.n10180 681.178
R4590 vdd.n10196 vdd.n10182 681.178
R4591 vdd.n10182 vdd.n10176 681.178
R4592 vdd.n10207 vdd.n10176 681.178
R4593 vdd.n10207 vdd.n10206 681.178
R4594 vdd.n10000 vdd.n9988 681.178
R4595 vdd.n10010 vdd.n9988 681.178
R4596 vdd.n10010 vdd.n9989 681.178
R4597 vdd.n9989 vdd.n9985 681.178
R4598 vdd.n10019 vdd.n9985 681.178
R4599 vdd.n10020 vdd.n10019 681.178
R4600 vdd.n10002 vdd.n9998 681.178
R4601 vdd.n9998 vdd.n9991 681.178
R4602 vdd.n9993 vdd.n9991 681.178
R4603 vdd.n10008 vdd.n9993 681.178
R4604 vdd.n10008 vdd.n9983 681.178
R4605 vdd.n10022 vdd.n9983 681.178
R4606 vdd.n10336 vdd.n10335 681.178
R4607 vdd.n10337 vdd.n10336 681.178
R4608 vdd.n10337 vdd.n10315 681.178
R4609 vdd.n10352 vdd.n10315 681.178
R4610 vdd.n10352 vdd.n10316 681.178
R4611 vdd.n10344 vdd.n10316 681.178
R4612 vdd.n10329 vdd.n10322 681.178
R4613 vdd.n10338 vdd.n10322 681.178
R4614 vdd.n10338 vdd.n10324 681.178
R4615 vdd.n10324 vdd.n10318 681.178
R4616 vdd.n10349 vdd.n10318 681.178
R4617 vdd.n10349 vdd.n10348 681.178
R4618 vdd.n10289 vdd.n10288 681.178
R4619 vdd.n10290 vdd.n10289 681.178
R4620 vdd.n10290 vdd.n10268 681.178
R4621 vdd.n10305 vdd.n10268 681.178
R4622 vdd.n10305 vdd.n10269 681.178
R4623 vdd.n10297 vdd.n10269 681.178
R4624 vdd.n10282 vdd.n10275 681.178
R4625 vdd.n10291 vdd.n10275 681.178
R4626 vdd.n10291 vdd.n10277 681.178
R4627 vdd.n10277 vdd.n10271 681.178
R4628 vdd.n10302 vdd.n10271 681.178
R4629 vdd.n10302 vdd.n10301 681.178
R4630 vdd.n10243 vdd.n10242 681.178
R4631 vdd.n10244 vdd.n10243 681.178
R4632 vdd.n10244 vdd.n10222 681.178
R4633 vdd.n10259 vdd.n10222 681.178
R4634 vdd.n10259 vdd.n10223 681.178
R4635 vdd.n10251 vdd.n10223 681.178
R4636 vdd.n10236 vdd.n10229 681.178
R4637 vdd.n10245 vdd.n10229 681.178
R4638 vdd.n10245 vdd.n10231 681.178
R4639 vdd.n10231 vdd.n10225 681.178
R4640 vdd.n10256 vdd.n10225 681.178
R4641 vdd.n10256 vdd.n10255 681.178
R4642 vdd.n10383 vdd.n10382 681.178
R4643 vdd.n10384 vdd.n10383 681.178
R4644 vdd.n10384 vdd.n10362 681.178
R4645 vdd.n10399 vdd.n10362 681.178
R4646 vdd.n10399 vdd.n10363 681.178
R4647 vdd.n10391 vdd.n10363 681.178
R4648 vdd.n10376 vdd.n10369 681.178
R4649 vdd.n10385 vdd.n10369 681.178
R4650 vdd.n10385 vdd.n10371 681.178
R4651 vdd.n10371 vdd.n10365 681.178
R4652 vdd.n10396 vdd.n10365 681.178
R4653 vdd.n10396 vdd.n10395 681.178
R4654 vdd.n10431 vdd.n10430 681.178
R4655 vdd.n10432 vdd.n10431 681.178
R4656 vdd.n10432 vdd.n10410 681.178
R4657 vdd.n10447 vdd.n10410 681.178
R4658 vdd.n10447 vdd.n10411 681.178
R4659 vdd.n10439 vdd.n10411 681.178
R4660 vdd.n10424 vdd.n10417 681.178
R4661 vdd.n10433 vdd.n10417 681.178
R4662 vdd.n10433 vdd.n10419 681.178
R4663 vdd.n10419 vdd.n10413 681.178
R4664 vdd.n10444 vdd.n10413 681.178
R4665 vdd.n10444 vdd.n10443 681.178
R4666 vdd.n10477 vdd.n10476 681.178
R4667 vdd.n10478 vdd.n10477 681.178
R4668 vdd.n10478 vdd.n10456 681.178
R4669 vdd.n10493 vdd.n10456 681.178
R4670 vdd.n10493 vdd.n10457 681.178
R4671 vdd.n10485 vdd.n10457 681.178
R4672 vdd.n10470 vdd.n10463 681.178
R4673 vdd.n10479 vdd.n10463 681.178
R4674 vdd.n10479 vdd.n10465 681.178
R4675 vdd.n10465 vdd.n10459 681.178
R4676 vdd.n10490 vdd.n10459 681.178
R4677 vdd.n10490 vdd.n10489 681.178
R4678 vdd.n10571 vdd.n10570 681.178
R4679 vdd.n10572 vdd.n10571 681.178
R4680 vdd.n10572 vdd.n10550 681.178
R4681 vdd.n10587 vdd.n10550 681.178
R4682 vdd.n10587 vdd.n10551 681.178
R4683 vdd.n10579 vdd.n10551 681.178
R4684 vdd.n10564 vdd.n10557 681.178
R4685 vdd.n10573 vdd.n10557 681.178
R4686 vdd.n10573 vdd.n10559 681.178
R4687 vdd.n10559 vdd.n10553 681.178
R4688 vdd.n10584 vdd.n10553 681.178
R4689 vdd.n10584 vdd.n10583 681.178
R4690 vdd.n10525 vdd.n10524 681.178
R4691 vdd.n10526 vdd.n10525 681.178
R4692 vdd.n10526 vdd.n10504 681.178
R4693 vdd.n10541 vdd.n10504 681.178
R4694 vdd.n10541 vdd.n10505 681.178
R4695 vdd.n10533 vdd.n10505 681.178
R4696 vdd.n10518 vdd.n10511 681.178
R4697 vdd.n10527 vdd.n10511 681.178
R4698 vdd.n10527 vdd.n10513 681.178
R4699 vdd.n10513 vdd.n10507 681.178
R4700 vdd.n10538 vdd.n10507 681.178
R4701 vdd.n10538 vdd.n10537 681.178
R4702 vdd.n10618 vdd.n10617 681.178
R4703 vdd.n10619 vdd.n10618 681.178
R4704 vdd.n10619 vdd.n10597 681.178
R4705 vdd.n10634 vdd.n10597 681.178
R4706 vdd.n10634 vdd.n10598 681.178
R4707 vdd.n10626 vdd.n10598 681.178
R4708 vdd.n10611 vdd.n10604 681.178
R4709 vdd.n10620 vdd.n10604 681.178
R4710 vdd.n10620 vdd.n10606 681.178
R4711 vdd.n10606 vdd.n10600 681.178
R4712 vdd.n10631 vdd.n10600 681.178
R4713 vdd.n10631 vdd.n10630 681.178
R4714 vdd.n10666 vdd.n10665 681.178
R4715 vdd.n10667 vdd.n10666 681.178
R4716 vdd.n10667 vdd.n10645 681.178
R4717 vdd.n10682 vdd.n10645 681.178
R4718 vdd.n10682 vdd.n10646 681.178
R4719 vdd.n10674 vdd.n10646 681.178
R4720 vdd.n10659 vdd.n10652 681.178
R4721 vdd.n10668 vdd.n10652 681.178
R4722 vdd.n10668 vdd.n10654 681.178
R4723 vdd.n10654 vdd.n10648 681.178
R4724 vdd.n10679 vdd.n10648 681.178
R4725 vdd.n10679 vdd.n10678 681.178
R4726 vdd.n10712 vdd.n10711 681.178
R4727 vdd.n10713 vdd.n10712 681.178
R4728 vdd.n10713 vdd.n10691 681.178
R4729 vdd.n10728 vdd.n10691 681.178
R4730 vdd.n10728 vdd.n10692 681.178
R4731 vdd.n10720 vdd.n10692 681.178
R4732 vdd.n10705 vdd.n10698 681.178
R4733 vdd.n10714 vdd.n10698 681.178
R4734 vdd.n10714 vdd.n10700 681.178
R4735 vdd.n10700 vdd.n10694 681.178
R4736 vdd.n10725 vdd.n10694 681.178
R4737 vdd.n10725 vdd.n10724 681.178
R4738 vdd.n9764 vdd.n9752 681.178
R4739 vdd.n9774 vdd.n9752 681.178
R4740 vdd.n9774 vdd.n9753 681.178
R4741 vdd.n9753 vdd.n9749 681.178
R4742 vdd.n9783 vdd.n9749 681.178
R4743 vdd.n9784 vdd.n9783 681.178
R4744 vdd.n9766 vdd.n9762 681.178
R4745 vdd.n9762 vdd.n9755 681.178
R4746 vdd.n9757 vdd.n9755 681.178
R4747 vdd.n9772 vdd.n9757 681.178
R4748 vdd.n9772 vdd.n9747 681.178
R4749 vdd.n9786 vdd.n9747 681.178
R4750 vdd.n10807 vdd.n10806 681.178
R4751 vdd.n10808 vdd.n10807 681.178
R4752 vdd.n10808 vdd.n10786 681.178
R4753 vdd.n10823 vdd.n10786 681.178
R4754 vdd.n10823 vdd.n10787 681.178
R4755 vdd.n10815 vdd.n10787 681.178
R4756 vdd.n10800 vdd.n10793 681.178
R4757 vdd.n10809 vdd.n10793 681.178
R4758 vdd.n10809 vdd.n10795 681.178
R4759 vdd.n10795 vdd.n10789 681.178
R4760 vdd.n10820 vdd.n10789 681.178
R4761 vdd.n10820 vdd.n10819 681.178
R4762 vdd.n10761 vdd.n10760 681.178
R4763 vdd.n10762 vdd.n10761 681.178
R4764 vdd.n10762 vdd.n10740 681.178
R4765 vdd.n10777 vdd.n10740 681.178
R4766 vdd.n10777 vdd.n10741 681.178
R4767 vdd.n10769 vdd.n10741 681.178
R4768 vdd.n10754 vdd.n10747 681.178
R4769 vdd.n10763 vdd.n10747 681.178
R4770 vdd.n10763 vdd.n10749 681.178
R4771 vdd.n10749 vdd.n10743 681.178
R4772 vdd.n10774 vdd.n10743 681.178
R4773 vdd.n10774 vdd.n10773 681.178
R4774 vdd.n10854 vdd.n10853 681.178
R4775 vdd.n10855 vdd.n10854 681.178
R4776 vdd.n10855 vdd.n10833 681.178
R4777 vdd.n10870 vdd.n10833 681.178
R4778 vdd.n10870 vdd.n10834 681.178
R4779 vdd.n10862 vdd.n10834 681.178
R4780 vdd.n10847 vdd.n10840 681.178
R4781 vdd.n10856 vdd.n10840 681.178
R4782 vdd.n10856 vdd.n10842 681.178
R4783 vdd.n10842 vdd.n10836 681.178
R4784 vdd.n10867 vdd.n10836 681.178
R4785 vdd.n10867 vdd.n10866 681.178
R4786 vdd.n10902 vdd.n10901 681.178
R4787 vdd.n10903 vdd.n10902 681.178
R4788 vdd.n10903 vdd.n10881 681.178
R4789 vdd.n10918 vdd.n10881 681.178
R4790 vdd.n10918 vdd.n10882 681.178
R4791 vdd.n10910 vdd.n10882 681.178
R4792 vdd.n10895 vdd.n10888 681.178
R4793 vdd.n10904 vdd.n10888 681.178
R4794 vdd.n10904 vdd.n10890 681.178
R4795 vdd.n10890 vdd.n10884 681.178
R4796 vdd.n10915 vdd.n10884 681.178
R4797 vdd.n10915 vdd.n10914 681.178
R4798 vdd.n10948 vdd.n10947 681.178
R4799 vdd.n10949 vdd.n10948 681.178
R4800 vdd.n10949 vdd.n10927 681.178
R4801 vdd.n10964 vdd.n10927 681.178
R4802 vdd.n10964 vdd.n10928 681.178
R4803 vdd.n10956 vdd.n10928 681.178
R4804 vdd.n10941 vdd.n10934 681.178
R4805 vdd.n10950 vdd.n10934 681.178
R4806 vdd.n10950 vdd.n10936 681.178
R4807 vdd.n10936 vdd.n10930 681.178
R4808 vdd.n10961 vdd.n10930 681.178
R4809 vdd.n10961 vdd.n10960 681.178
R4810 vdd.n10989 vdd.n10982 681.178
R4811 vdd.n10998 vdd.n10982 681.178
R4812 vdd.n10998 vdd.n10980 681.178
R4813 vdd.n11004 vdd.n10980 681.178
R4814 vdd.n11005 vdd.n11004 681.178
R4815 vdd.n11007 vdd.n11005 681.178
R4816 vdd.n10996 vdd.n10995 681.178
R4817 vdd.n10997 vdd.n10996 681.178
R4818 vdd.n10997 vdd.n10976 681.178
R4819 vdd.n11013 vdd.n10976 681.178
R4820 vdd.n11013 vdd.n11012 681.178
R4821 vdd.n11012 vdd.n11011 681.178
R4822 vdd.n11034 vdd.n11027 681.178
R4823 vdd.n11043 vdd.n11027 681.178
R4824 vdd.n11043 vdd.n11025 681.178
R4825 vdd.n11049 vdd.n11025 681.178
R4826 vdd.n11050 vdd.n11049 681.178
R4827 vdd.n11052 vdd.n11050 681.178
R4828 vdd.n11041 vdd.n11040 681.178
R4829 vdd.n11042 vdd.n11041 681.178
R4830 vdd.n11042 vdd.n11021 681.178
R4831 vdd.n11058 vdd.n11021 681.178
R4832 vdd.n11058 vdd.n11057 681.178
R4833 vdd.n11057 vdd.n11056 681.178
R4834 vdd.n11084 vdd.n11077 681.178
R4835 vdd.n11093 vdd.n11077 681.178
R4836 vdd.n11093 vdd.n11075 681.178
R4837 vdd.n11099 vdd.n11075 681.178
R4838 vdd.n11100 vdd.n11099 681.178
R4839 vdd.n11102 vdd.n11100 681.178
R4840 vdd.n11091 vdd.n11090 681.178
R4841 vdd.n11092 vdd.n11091 681.178
R4842 vdd.n11092 vdd.n11071 681.178
R4843 vdd.n11108 vdd.n11071 681.178
R4844 vdd.n11108 vdd.n11107 681.178
R4845 vdd.n11107 vdd.n11106 681.178
R4846 vdd.n11130 vdd.n11123 681.178
R4847 vdd.n11139 vdd.n11123 681.178
R4848 vdd.n11139 vdd.n11121 681.178
R4849 vdd.n11145 vdd.n11121 681.178
R4850 vdd.n11146 vdd.n11145 681.178
R4851 vdd.n11148 vdd.n11146 681.178
R4852 vdd.n11137 vdd.n11136 681.178
R4853 vdd.n11138 vdd.n11137 681.178
R4854 vdd.n11138 vdd.n11117 681.178
R4855 vdd.n11154 vdd.n11117 681.178
R4856 vdd.n11154 vdd.n11153 681.178
R4857 vdd.n11153 vdd.n11152 681.178
R4858 vdd.n11178 vdd.n11171 681.178
R4859 vdd.n11187 vdd.n11171 681.178
R4860 vdd.n11187 vdd.n11169 681.178
R4861 vdd.n11193 vdd.n11169 681.178
R4862 vdd.n11194 vdd.n11193 681.178
R4863 vdd.n11196 vdd.n11194 681.178
R4864 vdd.n11185 vdd.n11184 681.178
R4865 vdd.n11186 vdd.n11185 681.178
R4866 vdd.n11186 vdd.n11165 681.178
R4867 vdd.n11202 vdd.n11165 681.178
R4868 vdd.n11202 vdd.n11201 681.178
R4869 vdd.n11201 vdd.n11200 681.178
R4870 vdd.n442 vdd.n441 681.178
R4871 vdd.n443 vdd.n442 681.178
R4872 vdd.n443 vdd.n436 681.178
R4873 vdd.n449 vdd.n436 681.178
R4874 vdd.n450 vdd.n449 681.178
R4875 vdd.n452 vdd.n450 681.178
R4876 vdd.n465 vdd.n464 681.178
R4877 vdd.n464 vdd.n463 681.178
R4878 vdd.n463 vdd.n427 681.178
R4879 vdd.n458 vdd.n427 681.178
R4880 vdd.n458 vdd.n457 681.178
R4881 vdd.n457 vdd.n456 681.178
R4882 vdd.n11225 vdd.n11218 681.178
R4883 vdd.n11234 vdd.n11218 681.178
R4884 vdd.n11234 vdd.n11216 681.178
R4885 vdd.n11240 vdd.n11216 681.178
R4886 vdd.n11241 vdd.n11240 681.178
R4887 vdd.n11243 vdd.n11241 681.178
R4888 vdd.n11232 vdd.n11231 681.178
R4889 vdd.n11233 vdd.n11232 681.178
R4890 vdd.n11233 vdd.n11212 681.178
R4891 vdd.n11249 vdd.n11212 681.178
R4892 vdd.n11249 vdd.n11248 681.178
R4893 vdd.n11248 vdd.n11247 681.178
R4894 vdd.n11270 vdd.n11263 681.178
R4895 vdd.n11279 vdd.n11263 681.178
R4896 vdd.n11279 vdd.n11261 681.178
R4897 vdd.n11285 vdd.n11261 681.178
R4898 vdd.n11286 vdd.n11285 681.178
R4899 vdd.n11288 vdd.n11286 681.178
R4900 vdd.n11277 vdd.n11276 681.178
R4901 vdd.n11278 vdd.n11277 681.178
R4902 vdd.n11278 vdd.n11257 681.178
R4903 vdd.n11294 vdd.n11257 681.178
R4904 vdd.n11294 vdd.n11293 681.178
R4905 vdd.n11293 vdd.n11292 681.178
R4906 vdd.n11316 vdd.n11309 681.178
R4907 vdd.n11325 vdd.n11309 681.178
R4908 vdd.n11325 vdd.n11307 681.178
R4909 vdd.n11331 vdd.n11307 681.178
R4910 vdd.n11332 vdd.n11331 681.178
R4911 vdd.n11334 vdd.n11332 681.178
R4912 vdd.n11323 vdd.n11322 681.178
R4913 vdd.n11324 vdd.n11323 681.178
R4914 vdd.n11324 vdd.n11303 681.178
R4915 vdd.n11340 vdd.n11303 681.178
R4916 vdd.n11340 vdd.n11339 681.178
R4917 vdd.n11339 vdd.n11338 681.178
R4918 vdd.n11367 vdd.n11360 681.178
R4919 vdd.n11376 vdd.n11360 681.178
R4920 vdd.n11376 vdd.n11358 681.178
R4921 vdd.n11382 vdd.n11358 681.178
R4922 vdd.n11383 vdd.n11382 681.178
R4923 vdd.n11385 vdd.n11383 681.178
R4924 vdd.n11374 vdd.n11373 681.178
R4925 vdd.n11375 vdd.n11374 681.178
R4926 vdd.n11375 vdd.n11354 681.178
R4927 vdd.n11391 vdd.n11354 681.178
R4928 vdd.n11391 vdd.n11390 681.178
R4929 vdd.n11390 vdd.n11389 681.178
R4930 vdd.n11413 vdd.n11406 681.178
R4931 vdd.n11422 vdd.n11406 681.178
R4932 vdd.n11422 vdd.n11404 681.178
R4933 vdd.n11428 vdd.n11404 681.178
R4934 vdd.n11429 vdd.n11428 681.178
R4935 vdd.n11431 vdd.n11429 681.178
R4936 vdd.n11420 vdd.n11419 681.178
R4937 vdd.n11421 vdd.n11420 681.178
R4938 vdd.n11421 vdd.n11400 681.178
R4939 vdd.n11437 vdd.n11400 681.178
R4940 vdd.n11437 vdd.n11436 681.178
R4941 vdd.n11436 vdd.n11435 681.178
R4942 vdd.n11461 vdd.n11454 681.178
R4943 vdd.n11470 vdd.n11454 681.178
R4944 vdd.n11470 vdd.n11452 681.178
R4945 vdd.n11476 vdd.n11452 681.178
R4946 vdd.n11477 vdd.n11476 681.178
R4947 vdd.n11479 vdd.n11477 681.178
R4948 vdd.n11468 vdd.n11467 681.178
R4949 vdd.n11469 vdd.n11468 681.178
R4950 vdd.n11469 vdd.n11448 681.178
R4951 vdd.n11485 vdd.n11448 681.178
R4952 vdd.n11485 vdd.n11484 681.178
R4953 vdd.n11484 vdd.n11483 681.178
R4954 vdd.n11507 vdd.n11500 681.178
R4955 vdd.n11516 vdd.n11500 681.178
R4956 vdd.n11516 vdd.n11498 681.178
R4957 vdd.n11522 vdd.n11498 681.178
R4958 vdd.n11523 vdd.n11522 681.178
R4959 vdd.n11525 vdd.n11523 681.178
R4960 vdd.n11514 vdd.n11513 681.178
R4961 vdd.n11515 vdd.n11514 681.178
R4962 vdd.n11515 vdd.n11494 681.178
R4963 vdd.n11531 vdd.n11494 681.178
R4964 vdd.n11531 vdd.n11530 681.178
R4965 vdd.n11530 vdd.n11529 681.178
R4966 vdd.n11552 vdd.n11545 681.178
R4967 vdd.n11561 vdd.n11545 681.178
R4968 vdd.n11561 vdd.n11543 681.178
R4969 vdd.n11567 vdd.n11543 681.178
R4970 vdd.n11568 vdd.n11567 681.178
R4971 vdd.n11570 vdd.n11568 681.178
R4972 vdd.n11559 vdd.n11558 681.178
R4973 vdd.n11560 vdd.n11559 681.178
R4974 vdd.n11560 vdd.n11539 681.178
R4975 vdd.n11576 vdd.n11539 681.178
R4976 vdd.n11576 vdd.n11575 681.178
R4977 vdd.n11575 vdd.n11574 681.178
R4978 vdd.n11602 vdd.n11595 681.178
R4979 vdd.n11611 vdd.n11595 681.178
R4980 vdd.n11611 vdd.n11593 681.178
R4981 vdd.n11617 vdd.n11593 681.178
R4982 vdd.n11618 vdd.n11617 681.178
R4983 vdd.n11620 vdd.n11618 681.178
R4984 vdd.n11609 vdd.n11608 681.178
R4985 vdd.n11610 vdd.n11609 681.178
R4986 vdd.n11610 vdd.n11589 681.178
R4987 vdd.n11626 vdd.n11589 681.178
R4988 vdd.n11626 vdd.n11625 681.178
R4989 vdd.n11625 vdd.n11624 681.178
R4990 vdd.n11648 vdd.n11641 681.178
R4991 vdd.n11657 vdd.n11641 681.178
R4992 vdd.n11657 vdd.n11639 681.178
R4993 vdd.n11663 vdd.n11639 681.178
R4994 vdd.n11664 vdd.n11663 681.178
R4995 vdd.n11666 vdd.n11664 681.178
R4996 vdd.n11655 vdd.n11654 681.178
R4997 vdd.n11656 vdd.n11655 681.178
R4998 vdd.n11656 vdd.n11635 681.178
R4999 vdd.n11672 vdd.n11635 681.178
R5000 vdd.n11672 vdd.n11671 681.178
R5001 vdd.n11671 vdd.n11670 681.178
R5002 vdd.n11696 vdd.n11689 681.178
R5003 vdd.n11705 vdd.n11689 681.178
R5004 vdd.n11705 vdd.n11687 681.178
R5005 vdd.n11711 vdd.n11687 681.178
R5006 vdd.n11712 vdd.n11711 681.178
R5007 vdd.n11714 vdd.n11712 681.178
R5008 vdd.n11703 vdd.n11702 681.178
R5009 vdd.n11704 vdd.n11703 681.178
R5010 vdd.n11704 vdd.n11683 681.178
R5011 vdd.n11720 vdd.n11683 681.178
R5012 vdd.n11720 vdd.n11719 681.178
R5013 vdd.n11719 vdd.n11718 681.178
R5014 vdd.n207 vdd.n206 681.178
R5015 vdd.n208 vdd.n207 681.178
R5016 vdd.n208 vdd.n201 681.178
R5017 vdd.n214 vdd.n201 681.178
R5018 vdd.n215 vdd.n214 681.178
R5019 vdd.n217 vdd.n215 681.178
R5020 vdd.n230 vdd.n229 681.178
R5021 vdd.n229 vdd.n228 681.178
R5022 vdd.n228 vdd.n192 681.178
R5023 vdd.n223 vdd.n192 681.178
R5024 vdd.n223 vdd.n222 681.178
R5025 vdd.n222 vdd.n221 681.178
R5026 vdd.n11743 vdd.n11736 681.178
R5027 vdd.n11752 vdd.n11736 681.178
R5028 vdd.n11752 vdd.n11734 681.178
R5029 vdd.n11758 vdd.n11734 681.178
R5030 vdd.n11759 vdd.n11758 681.178
R5031 vdd.n11761 vdd.n11759 681.178
R5032 vdd.n11750 vdd.n11749 681.178
R5033 vdd.n11751 vdd.n11750 681.178
R5034 vdd.n11751 vdd.n11730 681.178
R5035 vdd.n11767 vdd.n11730 681.178
R5036 vdd.n11767 vdd.n11766 681.178
R5037 vdd.n11766 vdd.n11765 681.178
R5038 vdd.n11788 vdd.n11781 681.178
R5039 vdd.n11797 vdd.n11781 681.178
R5040 vdd.n11797 vdd.n11779 681.178
R5041 vdd.n11803 vdd.n11779 681.178
R5042 vdd.n11804 vdd.n11803 681.178
R5043 vdd.n11806 vdd.n11804 681.178
R5044 vdd.n11795 vdd.n11794 681.178
R5045 vdd.n11796 vdd.n11795 681.178
R5046 vdd.n11796 vdd.n11775 681.178
R5047 vdd.n11812 vdd.n11775 681.178
R5048 vdd.n11812 vdd.n11811 681.178
R5049 vdd.n11811 vdd.n11810 681.178
R5050 vdd.n11838 vdd.n11831 681.178
R5051 vdd.n11847 vdd.n11831 681.178
R5052 vdd.n11847 vdd.n11829 681.178
R5053 vdd.n11853 vdd.n11829 681.178
R5054 vdd.n11854 vdd.n11853 681.178
R5055 vdd.n11856 vdd.n11854 681.178
R5056 vdd.n11845 vdd.n11844 681.178
R5057 vdd.n11846 vdd.n11845 681.178
R5058 vdd.n11846 vdd.n11825 681.178
R5059 vdd.n11862 vdd.n11825 681.178
R5060 vdd.n11862 vdd.n11861 681.178
R5061 vdd.n11861 vdd.n11860 681.178
R5062 vdd.n11884 vdd.n11877 681.178
R5063 vdd.n11893 vdd.n11877 681.178
R5064 vdd.n11893 vdd.n11875 681.178
R5065 vdd.n11899 vdd.n11875 681.178
R5066 vdd.n11900 vdd.n11899 681.178
R5067 vdd.n11902 vdd.n11900 681.178
R5068 vdd.n11891 vdd.n11890 681.178
R5069 vdd.n11892 vdd.n11891 681.178
R5070 vdd.n11892 vdd.n11871 681.178
R5071 vdd.n11908 vdd.n11871 681.178
R5072 vdd.n11908 vdd.n11907 681.178
R5073 vdd.n11907 vdd.n11906 681.178
R5074 vdd.n11932 vdd.n11925 681.178
R5075 vdd.n11941 vdd.n11925 681.178
R5076 vdd.n11941 vdd.n11923 681.178
R5077 vdd.n11947 vdd.n11923 681.178
R5078 vdd.n11948 vdd.n11947 681.178
R5079 vdd.n11950 vdd.n11948 681.178
R5080 vdd.n11939 vdd.n11938 681.178
R5081 vdd.n11940 vdd.n11939 681.178
R5082 vdd.n11940 vdd.n11919 681.178
R5083 vdd.n11956 vdd.n11919 681.178
R5084 vdd.n11956 vdd.n11955 681.178
R5085 vdd.n11955 vdd.n11954 681.178
R5086 vdd.t1047 vdd.n105 287.382
R5087 vdd.t507 vdd.n105 287.382
R5088 vdd.t507 vdd.n107 287.382
R5089 vdd.n107 vdd.t509 287.382
R5090 vdd.n128 vdd.t509 287.382
R5091 vdd.t1182 vdd.n128 287.382
R5092 vdd.t7 vdd.n151 287.382
R5093 vdd.t913 vdd.n151 287.382
R5094 vdd.t913 vdd.n153 287.382
R5095 vdd.n153 vdd.t915 287.382
R5096 vdd.n174 vdd.t915 287.382
R5097 vdd.t977 vdd.n174 287.382
R5098 vdd.t1475 vdd.n248 287.382
R5099 vdd.t736 vdd.n248 287.382
R5100 vdd.t736 vdd.n250 287.382
R5101 vdd.n250 vdd.t738 287.382
R5102 vdd.n271 vdd.t738 287.382
R5103 vdd.t527 vdd.n271 287.382
R5104 vdd.t562 vdd.n294 287.382
R5105 vdd.t161 vdd.n294 287.382
R5106 vdd.t161 vdd.n296 287.382
R5107 vdd.n296 vdd.t163 287.382
R5108 vdd.n317 vdd.t163 287.382
R5109 vdd.t1238 vdd.n317 287.382
R5110 vdd.t1298 vdd.n340 287.382
R5111 vdd.t572 vdd.n340 287.382
R5112 vdd.t572 vdd.n342 287.382
R5113 vdd.n342 vdd.t574 287.382
R5114 vdd.n363 vdd.t574 287.382
R5115 vdd.t156 vdd.n363 287.382
R5116 vdd.t1485 vdd.n386 287.382
R5117 vdd.t1413 vdd.n386 287.382
R5118 vdd.t1413 vdd.n388 287.382
R5119 vdd.n388 vdd.t1415 287.382
R5120 vdd.n409 vdd.t1415 287.382
R5121 vdd.t959 vdd.n409 287.382
R5122 vdd.t209 vdd.n483 287.382
R5123 vdd.t925 vdd.n483 287.382
R5124 vdd.t925 vdd.n485 287.382
R5125 vdd.n485 vdd.t927 287.382
R5126 vdd.n506 vdd.t927 287.382
R5127 vdd.t336 vdd.n506 287.382
R5128 vdd.t375 vdd.n529 287.382
R5129 vdd.t127 vdd.n529 287.382
R5130 vdd.t127 vdd.n531 287.382
R5131 vdd.n531 vdd.t126 287.382
R5132 vdd.n552 vdd.t126 287.382
R5133 vdd.t122 vdd.n552 287.382
R5134 vdd.t728 vdd.n6696 287.382
R5135 vdd.t362 vdd.n6696 287.382
R5136 vdd.t362 vdd.n6688 287.382
R5137 vdd.t363 vdd.n6688 287.382
R5138 vdd.t363 vdd.n6722 287.382
R5139 vdd.n6722 vdd.t1288 287.382
R5140 vdd.t235 vdd.n6742 287.382
R5141 vdd.t624 vdd.n6742 287.382
R5142 vdd.t624 vdd.n6734 287.382
R5143 vdd.t625 vdd.n6734 287.382
R5144 vdd.t625 vdd.n6768 287.382
R5145 vdd.n6768 vdd.t207 287.382
R5146 vdd.t155 vdd.n6840 287.382
R5147 vdd.t152 vdd.n6840 287.382
R5148 vdd.t152 vdd.n6832 287.382
R5149 vdd.t153 vdd.n6832 287.382
R5150 vdd.t153 vdd.n6866 287.382
R5151 vdd.n6866 vdd.t1318 287.382
R5152 vdd.t413 vdd.n6886 287.382
R5153 vdd.t217 vdd.n6886 287.382
R5154 vdd.t217 vdd.n6878 287.382
R5155 vdd.t218 vdd.n6878 287.382
R5156 vdd.t218 vdd.n6912 287.382
R5157 vdd.n6912 vdd.t205 287.382
R5158 vdd.t983 vdd.n6932 287.382
R5159 vdd.t980 vdd.n6932 287.382
R5160 vdd.t980 vdd.n6924 287.382
R5161 vdd.t981 vdd.n6924 287.382
R5162 vdd.t981 vdd.n6958 287.382
R5163 vdd.n6958 vdd.t558 287.382
R5164 vdd.t1107 vdd.n6978 287.382
R5165 vdd.t806 vdd.n6978 287.382
R5166 vdd.t806 vdd.n6970 287.382
R5167 vdd.t807 vdd.n6970 287.382
R5168 vdd.t807 vdd.n7004 287.382
R5169 vdd.n7004 vdd.t377 287.382
R5170 vdd.t353 vdd.n7076 287.382
R5171 vdd.t302 vdd.n7076 287.382
R5172 vdd.t302 vdd.n7068 287.382
R5173 vdd.t303 vdd.n7068 287.382
R5174 vdd.t303 vdd.n7102 287.382
R5175 vdd.n7102 vdd.t587 287.382
R5176 vdd.t634 vdd.n8534 287.382
R5177 vdd.t1451 vdd.n8534 287.382
R5178 vdd.t1451 vdd.n8526 287.382
R5179 vdd.t1452 vdd.n8526 287.382
R5180 vdd.t1452 vdd.n8560 287.382
R5181 vdd.n8560 vdd.t482 287.382
R5182 vdd.t1463 vdd.n7121 287.382
R5183 vdd.t521 vdd.n7121 287.382
R5184 vdd.t521 vdd.n7123 287.382
R5185 vdd.n7123 vdd.t520 287.382
R5186 vdd.n7144 vdd.t520 287.382
R5187 vdd.t1025 vdd.n7144 287.382
R5188 vdd.t1310 vdd.n7167 287.382
R5189 vdd.t183 vdd.n7167 287.382
R5190 vdd.t183 vdd.n7169 287.382
R5191 vdd.n7169 vdd.t182 287.382
R5192 vdd.n7190 vdd.t182 287.382
R5193 vdd.t979 vdd.n7190 287.382
R5194 vdd.t1049 vdd.n7264 287.382
R5195 vdd.t883 vdd.n7264 287.382
R5196 vdd.t883 vdd.n7266 287.382
R5197 vdd.n7266 vdd.t882 287.382
R5198 vdd.n7287 vdd.t882 287.382
R5199 vdd.t1285 vdd.n7287 287.382
R5200 vdd.t1360 vdd.n7310 287.382
R5201 vdd.t532 vdd.n7310 287.382
R5202 vdd.t532 vdd.n7312 287.382
R5203 vdd.n7312 vdd.t534 287.382
R5204 vdd.n7333 vdd.t534 287.382
R5205 vdd.t536 vdd.n7333 287.382
R5206 vdd.t593 vdd.n7356 287.382
R5207 vdd.t1092 vdd.n7356 287.382
R5208 vdd.t1092 vdd.n7358 287.382
R5209 vdd.n7358 vdd.t1091 287.382
R5210 vdd.n7379 vdd.t1091 287.382
R5211 vdd.t1094 vdd.n7379 287.382
R5212 vdd.t379 vdd.n7402 287.382
R5213 vdd.t1253 vdd.n7402 287.382
R5214 vdd.t1253 vdd.n7404 287.382
R5215 vdd.n7404 vdd.t1252 287.382
R5216 vdd.n7425 vdd.t1252 287.382
R5217 vdd.t1255 vdd.n7425 287.382
R5218 vdd.t1326 vdd.n7499 287.382
R5219 vdd.t931 vdd.n7499 287.382
R5220 vdd.t931 vdd.n7501 287.382
R5221 vdd.n7501 vdd.t930 287.382
R5222 vdd.n7522 vdd.t930 287.382
R5223 vdd.t143 vdd.n7522 287.382
R5224 vdd.t484 vdd.n6648 287.382
R5225 vdd.t704 vdd.n6648 287.382
R5226 vdd.t704 vdd.n6650 287.382
R5227 vdd.n6650 vdd.t703 287.382
R5228 vdd.n6671 vdd.t703 287.382
R5229 vdd.t1088 vdd.n6671 287.382
R5230 vdd.t898 vdd.n7543 287.382
R5231 vdd.t1273 vdd.n7543 287.382
R5232 vdd.t1273 vdd.n7545 287.382
R5233 vdd.n7545 vdd.t1272 287.382
R5234 vdd.n7566 vdd.t1272 287.382
R5235 vdd.t1263 vdd.n7566 287.382
R5236 vdd.t166 vdd.n7588 287.382
R5237 vdd.t886 vdd.n7588 287.382
R5238 vdd.t886 vdd.n7590 287.382
R5239 vdd.n7590 vdd.t885 287.382
R5240 vdd.n7611 vdd.t885 287.382
R5241 vdd.t809 vdd.n7611 287.382
R5242 vdd.t589 vdd.n7638 287.382
R5243 vdd.t223 vdd.n7638 287.382
R5244 vdd.t223 vdd.n7640 287.382
R5245 vdd.n7640 vdd.t225 287.382
R5246 vdd.n7661 vdd.t225 287.382
R5247 vdd.t1226 vdd.n7661 287.382
R5248 vdd.t862 vdd.n7684 287.382
R5249 vdd.t251 vdd.n7684 287.382
R5250 vdd.t251 vdd.n7686 287.382
R5251 vdd.n7686 vdd.t250 287.382
R5252 vdd.n7707 vdd.t250 287.382
R5253 vdd.t874 vdd.n7707 287.382
R5254 vdd.t1342 vdd.n7732 287.382
R5255 vdd.t1265 vdd.n7732 287.382
R5256 vdd.t1265 vdd.n7734 287.382
R5257 vdd.n7734 vdd.t1264 287.382
R5258 vdd.n7755 vdd.t1264 287.382
R5259 vdd.t1078 vdd.n7755 287.382
R5260 vdd.n7442 vdd.t1154 287.382
R5261 vdd.t443 vdd.n7442 287.382
R5262 vdd.n7450 vdd.t443 287.382
R5263 vdd.n7450 vdd.t442 287.382
R5264 vdd.n7467 vdd.t442 287.382
R5265 vdd.t892 vdd.n7467 287.382
R5266 vdd.t896 vdd.n7779 287.382
R5267 vdd.t518 vdd.n7779 287.382
R5268 vdd.t518 vdd.n7781 287.382
R5269 vdd.n7781 vdd.t517 287.382
R5270 vdd.n7802 vdd.t517 287.382
R5271 vdd.t1506 vdd.n7802 287.382
R5272 vdd.t837 vdd.n7824 287.382
R5273 vdd.t239 vdd.n7824 287.382
R5274 vdd.t239 vdd.n7826 287.382
R5275 vdd.n7826 vdd.t238 287.382
R5276 vdd.n7847 vdd.t238 287.382
R5277 vdd.t241 vdd.n7847 287.382
R5278 vdd.t1375 vdd.n7870 287.382
R5279 vdd.t541 vdd.n7870 287.382
R5280 vdd.t541 vdd.n7872 287.382
R5281 vdd.n7872 vdd.t540 287.382
R5282 vdd.n7893 vdd.t540 287.382
R5283 vdd.t543 vdd.n7893 287.382
R5284 vdd.t486 vdd.n7921 287.382
R5285 vdd.t68 vdd.n7921 287.382
R5286 vdd.t68 vdd.n7923 287.382
R5287 vdd.n7923 vdd.t67 287.382
R5288 vdd.n7944 vdd.t67 287.382
R5289 vdd.t306 vdd.n7944 287.382
R5290 vdd.t872 vdd.n7967 287.382
R5291 vdd.t319 vdd.n7967 287.382
R5292 vdd.t319 vdd.n7969 287.382
R5293 vdd.n7969 vdd.t318 287.382
R5294 vdd.n7990 vdd.t318 287.382
R5295 vdd.t620 vdd.n7990 287.382
R5296 vdd.t1330 vdd.n8015 287.382
R5297 vdd.t962 vdd.n8015 287.382
R5298 vdd.t962 vdd.n8017 287.382
R5299 vdd.n8017 vdd.t961 287.382
R5300 vdd.n8038 vdd.t961 287.382
R5301 vdd.t978 vdd.n8038 287.382
R5302 vdd.t36 vdd.n8061 287.382
R5303 vdd.t643 vdd.n8061 287.382
R5304 vdd.t643 vdd.n8063 287.382
R5305 vdd.n8063 vdd.t642 287.382
R5306 vdd.n8084 vdd.t642 287.382
R5307 vdd.t22 vdd.n8084 287.382
R5308 vdd.t835 vdd.n8106 287.382
R5309 vdd.t130 vdd.n8106 287.382
R5310 vdd.t130 vdd.n8108 287.382
R5311 vdd.n8108 vdd.t129 287.382
R5312 vdd.n8129 vdd.t129 287.382
R5313 vdd.t335 vdd.n8129 287.382
R5314 vdd.t201 vdd.n8156 287.382
R5315 vdd.t325 vdd.n8156 287.382
R5316 vdd.t325 vdd.n8158 287.382
R5317 vdd.n8158 vdd.t324 287.382
R5318 vdd.n8179 vdd.t324 287.382
R5319 vdd.t70 vdd.n8179 287.382
R5320 vdd.t973 vdd.n8202 287.382
R5321 vdd.t248 vdd.n8202 287.382
R5322 vdd.t248 vdd.n8204 287.382
R5323 vdd.n8204 vdd.t247 287.382
R5324 vdd.n8225 vdd.t247 287.382
R5325 vdd.t1442 vdd.n8225 287.382
R5326 vdd.t1346 vdd.n8250 287.382
R5327 vdd.t1448 vdd.n8250 287.382
R5328 vdd.t1448 vdd.n8252 287.382
R5329 vdd.n8252 vdd.t1450 287.382
R5330 vdd.n8273 vdd.t1450 287.382
R5331 vdd.t743 vdd.n8273 287.382
R5332 vdd.n7207 vdd.t1459 287.382
R5333 vdd.t1394 vdd.n7207 287.382
R5334 vdd.n7215 vdd.t1394 287.382
R5335 vdd.n7215 vdd.t1393 287.382
R5336 vdd.n7232 vdd.t1393 287.382
R5337 vdd.t277 vdd.n7232 287.382
R5338 vdd.t854 vdd.n8297 287.382
R5339 vdd.t1176 vdd.n8297 287.382
R5340 vdd.t1176 vdd.n8299 287.382
R5341 vdd.n8299 vdd.t1175 287.382
R5342 vdd.n8320 vdd.t1175 287.382
R5343 vdd.t1112 vdd.n8320 287.382
R5344 vdd.t56 vdd.n8342 287.382
R5345 vdd.t450 vdd.n8342 287.382
R5346 vdd.t450 vdd.n8344 287.382
R5347 vdd.n8344 vdd.t449 287.382
R5348 vdd.n8365 vdd.t449 287.382
R5349 vdd.t343 vdd.n8365 287.382
R5350 vdd.t9 vdd.n8392 287.382
R5351 vdd.t879 vdd.n8392 287.382
R5352 vdd.t879 vdd.n8394 287.382
R5353 vdd.n8394 vdd.t878 287.382
R5354 vdd.n8415 vdd.t878 287.382
R5355 vdd.t881 vdd.n8415 287.382
R5356 vdd.t40 vdd.n8438 287.382
R5357 vdd.t1420 vdd.n8438 287.382
R5358 vdd.t1420 vdd.n8440 287.382
R5359 vdd.n8440 vdd.t1419 287.382
R5360 vdd.n8461 vdd.t1419 287.382
R5361 vdd.t1149 vdd.n8461 287.382
R5362 vdd.t211 vdd.n8486 287.382
R5363 vdd.t1064 vdd.n8486 287.382
R5364 vdd.t1064 vdd.n8488 287.382
R5365 vdd.n8488 vdd.t1063 287.382
R5366 vdd.n8509 vdd.t1063 287.382
R5367 vdd.t1066 vdd.n8509 287.382
R5368 vdd.t284 vdd.n8627 287.382
R5369 vdd.t1079 vdd.n8627 287.382
R5370 vdd.t1079 vdd.n8619 287.382
R5371 vdd.t1080 vdd.n8619 287.382
R5372 vdd.t1080 vdd.n8653 287.382
R5373 vdd.n8653 vdd.t848 287.382
R5374 vdd.t412 vdd.n8581 287.382
R5375 vdd.t764 vdd.n8581 287.382
R5376 vdd.t764 vdd.n8573 287.382
R5377 vdd.t762 vdd.n8573 287.382
R5378 vdd.t762 vdd.n8607 287.382
R5379 vdd.n8607 vdd.t773 287.382
R5380 vdd.t1143 vdd.n8674 287.382
R5381 vdd.t254 vdd.n8674 287.382
R5382 vdd.t254 vdd.n8666 287.382
R5383 vdd.t255 vdd.n8666 287.382
R5384 vdd.t255 vdd.n8700 287.382
R5385 vdd.n8700 vdd.t1314 287.382
R5386 vdd.t658 vdd.n8722 287.382
R5387 vdd.t933 vdd.n8722 287.382
R5388 vdd.t933 vdd.n8714 287.382
R5389 vdd.t934 vdd.n8714 287.382
R5390 vdd.t934 vdd.n8748 287.382
R5391 vdd.n8748 vdd.t856 287.382
R5392 vdd.t1507 vdd.n8768 287.382
R5393 vdd.t190 vdd.n8768 287.382
R5394 vdd.t190 vdd.n8760 287.382
R5395 vdd.t188 vdd.n8760 287.382
R5396 vdd.t188 vdd.n8794 287.382
R5397 vdd.n8794 vdd.t1467 287.382
R5398 vdd.t1089 vdd.n7023 287.382
R5399 vdd.t82 vdd.n7023 287.382
R5400 vdd.t82 vdd.n7042 287.382
R5401 vdd.n7042 vdd.t80 287.382
R5402 vdd.t80 vdd.n7017 287.382
R5403 vdd.t97 vdd.n7017 287.382
R5404 vdd.t66 vdd.n8910 287.382
R5405 vdd.t139 vdd.n8910 287.382
R5406 vdd.t139 vdd.n8902 287.382
R5407 vdd.t137 vdd.n8902 287.382
R5408 vdd.t137 vdd.n8936 287.382
R5409 vdd.n8936 vdd.t825 287.382
R5410 vdd.t1195 vdd.n8863 287.382
R5411 vdd.t584 vdd.n8863 287.382
R5412 vdd.t584 vdd.n8855 287.382
R5413 vdd.t585 vdd.n8855 287.382
R5414 vdd.t585 vdd.n8889 287.382
R5415 vdd.n8889 vdd.t765 287.382
R5416 vdd.t264 vdd.n8817 287.382
R5417 vdd.t1201 vdd.n8817 287.382
R5418 vdd.t1201 vdd.n8809 287.382
R5419 vdd.t1199 vdd.n8809 287.382
R5420 vdd.t1199 vdd.n8843 287.382
R5421 vdd.n8843 vdd.t1129 287.382
R5422 vdd.t758 vdd.n8957 287.382
R5423 vdd.t755 vdd.n8957 287.382
R5424 vdd.t755 vdd.n8949 287.382
R5425 vdd.t756 vdd.n8949 287.382
R5426 vdd.t756 vdd.n8983 287.382
R5427 vdd.n8983 vdd.t458 287.382
R5428 vdd.t1062 vdd.n9005 287.382
R5429 vdd.t640 vdd.n9005 287.382
R5430 vdd.t640 vdd.n8997 287.382
R5431 vdd.t638 vdd.n8997 287.382
R5432 vdd.t638 vdd.n9031 287.382
R5433 vdd.n9031 vdd.t864 287.382
R5434 vdd.t1108 vdd.n9051 287.382
R5435 vdd.t1526 vdd.n9051 287.382
R5436 vdd.t1526 vdd.n9043 287.382
R5437 vdd.t1524 vdd.n9043 287.382
R5438 vdd.t1524 vdd.n9077 287.382
R5439 vdd.n9077 vdd.t1477 287.382
R5440 vdd.t64 vdd.n9145 287.382
R5441 vdd.t77 vdd.n9145 287.382
R5442 vdd.t77 vdd.n9137 287.382
R5443 vdd.t78 vdd.n9137 287.382
R5444 vdd.t78 vdd.n9171 287.382
R5445 vdd.n9171 vdd.t1006 287.382
R5446 vdd.t1024 vdd.n9099 287.382
R5447 vdd.t785 vdd.n9099 287.382
R5448 vdd.t785 vdd.n9091 287.382
R5449 vdd.t783 vdd.n9091 287.382
R5450 vdd.t783 vdd.n9125 287.382
R5451 vdd.n9125 vdd.t430 287.382
R5452 vdd.t1270 vdd.n9192 287.382
R5453 vdd.t1267 vdd.n9192 287.382
R5454 vdd.t1267 vdd.n9184 287.382
R5455 vdd.t1268 vdd.n9184 287.382
R5456 vdd.t1268 vdd.n9218 287.382
R5457 vdd.n9218 vdd.t566 287.382
R5458 vdd.t675 vdd.n9240 287.382
R5459 vdd.t744 vdd.n9240 287.382
R5460 vdd.t744 vdd.n9232 287.382
R5461 vdd.t745 vdd.n9232 287.382
R5462 vdd.t745 vdd.n9266 287.382
R5463 vdd.n9266 vdd.t42 287.382
R5464 vdd.t547 vdd.n9286 287.382
R5465 vdd.t401 vdd.n9286 287.382
R5466 vdd.t401 vdd.n9278 287.382
R5467 vdd.t399 vdd.n9278 287.382
R5468 vdd.t399 vdd.n9312 287.382
R5469 vdd.n9312 vdd.t1302 287.382
R5470 vdd.t1362 vdd.n6787 287.382
R5471 vdd.t693 vdd.n6787 287.382
R5472 vdd.t693 vdd.n6806 287.382
R5473 vdd.n6806 vdd.t691 287.382
R5474 vdd.t691 vdd.n6781 287.382
R5475 vdd.t89 vdd.n6781 287.382
R5476 vdd.t523 vdd.n9381 287.382
R5477 vdd.t176 vdd.n9381 287.382
R5478 vdd.t176 vdd.n9373 287.382
R5479 vdd.t177 vdd.n9373 287.382
R5480 vdd.t177 vdd.n9407 287.382
R5481 vdd.n9407 vdd.t988 287.382
R5482 vdd.t1031 vdd.n9335 287.382
R5483 vdd.t1028 vdd.n9335 287.382
R5484 vdd.t1028 vdd.n9327 287.382
R5485 vdd.t1029 vdd.n9327 287.382
R5486 vdd.t1029 vdd.n9361 287.382
R5487 vdd.n9361 vdd.t627 287.382
R5488 vdd.t428 vdd.n9428 287.382
R5489 vdd.t546 vdd.n9428 287.382
R5490 vdd.t546 vdd.n9420 287.382
R5491 vdd.t544 vdd.n9420 287.382
R5492 vdd.t544 vdd.n9454 287.382
R5493 vdd.n9454 vdd.t601 287.382
R5494 vdd.t1191 vdd.n9476 287.382
R5495 vdd.t661 vdd.n9476 287.382
R5496 vdd.t661 vdd.n9468 287.382
R5497 vdd.t662 vdd.n9468 287.382
R5498 vdd.t662 vdd.n9502 287.382
R5499 vdd.n9502 vdd.t860 287.382
R5500 vdd.t76 vdd.n9522 287.382
R5501 vdd.t1518 vdd.n9522 287.382
R5502 vdd.t1518 vdd.n9514 287.382
R5503 vdd.t1519 vdd.n9514 287.382
R5504 vdd.t1519 vdd.n9548 287.382
R5505 vdd.n9548 vdd.t1041 287.382
R5506 vdd.t441 vdd.n3682 287.382
R5507 vdd.t474 vdd.n3682 287.382
R5508 vdd.t474 vdd.n3674 287.382
R5509 vdd.t475 vdd.n3674 287.382
R5510 vdd.t475 vdd.n3708 287.382
R5511 vdd.n3708 vdd.t1483 287.382
R5512 vdd.t234 vdd.n3728 287.382
R5513 vdd.t680 vdd.n3728 287.382
R5514 vdd.t680 vdd.n3720 287.382
R5515 vdd.t681 vdd.n3720 287.382
R5516 vdd.t681 vdd.n3754 287.382
R5517 vdd.n3754 vdd.t464 287.382
R5518 vdd.t503 vdd.n3826 287.382
R5519 vdd.t192 vdd.n3826 287.382
R5520 vdd.t192 vdd.n3818 287.382
R5521 vdd.t193 vdd.n3818 287.382
R5522 vdd.t193 vdd.n3852 287.382
R5523 vdd.n3852 vdd.t599 287.382
R5524 vdd.t136 vdd.n3872 287.382
R5525 vdd.t1279 vdd.n3872 287.382
R5526 vdd.t1279 vdd.n3864 287.382
R5527 vdd.t1280 vdd.n3864 287.382
R5528 vdd.t1280 vdd.n3898 287.382
R5529 vdd.n3898 vdd.t460 287.382
R5530 vdd.t611 vdd.n3918 287.382
R5531 vdd.t1132 vdd.n3918 287.382
R5532 vdd.t1132 vdd.n3910 287.382
R5533 vdd.t1133 vdd.n3910 287.382
R5534 vdd.t1133 vdd.n3944 287.382
R5535 vdd.n3944 vdd.t1057 287.382
R5536 vdd.t802 vdd.n3964 287.382
R5537 vdd.t1207 vdd.n3964 287.382
R5538 vdd.t1207 vdd.n3956 287.382
R5539 vdd.t1208 vdd.n3956 287.382
R5540 vdd.t1208 vdd.n3990 287.382
R5541 vdd.n3990 vdd.t603 287.382
R5542 vdd.t473 vdd.n4062 287.382
R5543 vdd.t1407 vdd.n4062 287.382
R5544 vdd.t1407 vdd.n4054 287.382
R5545 vdd.t1408 vdd.n4054 287.382
R5546 vdd.t1408 vdd.n4088 287.382
R5547 vdd.n4088 vdd.t468 287.382
R5548 vdd.t327 vdd.n5520 287.382
R5549 vdd.t759 vdd.n5520 287.382
R5550 vdd.t759 vdd.n5512 287.382
R5551 vdd.t760 vdd.n5512 287.382
R5552 vdd.t760 vdd.n5546 287.382
R5553 vdd.n5546 vdd.t556 287.382
R5554 vdd.t203 vdd.n4107 287.382
R5555 vdd.t394 vdd.n4107 287.382
R5556 vdd.t394 vdd.n4109 287.382
R5557 vdd.n4109 vdd.t393 287.382
R5558 vdd.n4130 vdd.t393 287.382
R5559 vdd.t440 vdd.n4130 287.382
R5560 vdd.t554 vdd.n4153 287.382
R5561 vdd.t621 vdd.n4153 287.382
R5562 vdd.t621 vdd.n4155 287.382
R5563 vdd.n4155 vdd.t623 287.382
R5564 vdd.n4176 vdd.t623 287.382
R5565 vdd.t477 vdd.n4176 287.382
R5566 vdd.t1290 vdd.n4250 287.382
R5567 vdd.t1183 vdd.n4250 287.382
R5568 vdd.t1183 vdd.n4252 287.382
R5569 vdd.n4252 vdd.t1185 287.382
R5570 vdd.n4273 vdd.t1185 287.382
R5571 vdd.t114 vdd.n4273 287.382
R5572 vdd.t1316 vdd.n4296 287.382
R5573 vdd.t419 vdd.n4296 287.382
R5574 vdd.t419 vdd.n4298 287.382
R5575 vdd.n4298 vdd.t421 287.382
R5576 vdd.n4319 vdd.t421 287.382
R5577 vdd.t810 vdd.n4319 287.382
R5578 vdd.t1055 vdd.n4342 287.382
R5579 vdd.t1424 vdd.n4342 287.382
R5580 vdd.t1424 vdd.n4344 287.382
R5581 vdd.n4344 vdd.t1426 287.382
R5582 vdd.n4365 vdd.t1426 287.382
R5583 vdd.t1427 vdd.n4365 287.382
R5584 vdd.t570 vdd.n4388 287.382
R5585 vdd.t1435 vdd.n4388 287.382
R5586 vdd.t1435 vdd.n4390 287.382
R5587 vdd.n4390 vdd.t1437 287.382
R5588 vdd.n4411 vdd.t1437 287.382
R5589 vdd.t1225 vdd.n4411 287.382
R5590 vdd.t1045 vdd.n4485 287.382
R5591 vdd.t1231 vdd.n4485 287.382
R5592 vdd.t1231 vdd.n4487 287.382
R5593 vdd.n4487 vdd.t1233 287.382
R5594 vdd.n4508 vdd.t1233 287.382
R5595 vdd.t951 vdd.n4508 287.382
R5596 vdd.t560 vdd.n3634 287.382
R5597 vdd.t1034 vdd.n3634 287.382
R5598 vdd.t1034 vdd.n3636 287.382
R5599 vdd.n3636 vdd.t1036 287.382
R5600 vdd.n3657 vdd.t1036 287.382
R5601 vdd.t230 vdd.n3657 287.382
R5602 vdd.t1000 vdd.n4529 287.382
R5603 vdd.t696 vdd.n4529 287.382
R5604 vdd.t696 vdd.n4531 287.382
R5605 vdd.n4531 vdd.t698 287.382
R5606 vdd.n4552 vdd.t698 287.382
R5607 vdd.t1148 vdd.n4552 287.382
R5608 vdd.t174 vdd.n4574 287.382
R5609 vdd.t447 vdd.n4574 287.382
R5610 vdd.t447 vdd.n4576 287.382
R5611 vdd.n4576 vdd.t446 287.382
R5612 vdd.n4597 vdd.t446 287.382
R5613 vdd.t145 vdd.n4597 287.382
R5614 vdd.t197 vdd.n4624 287.382
R5615 vdd.t149 vdd.n4624 287.382
R5616 vdd.t149 vdd.n4626 287.382
R5617 vdd.n4626 vdd.t151 287.382
R5618 vdd.n4647 vdd.t151 287.382
R5619 vdd.t1178 vdd.n4647 287.382
R5620 vdd.t34 vdd.n4670 287.382
R5621 vdd.t668 vdd.n4670 287.382
R5622 vdd.t668 vdd.n4672 287.382
R5623 vdd.n4672 vdd.t667 287.382
R5624 vdd.n4693 vdd.t667 287.382
R5625 vdd.t670 vdd.n4693 287.382
R5626 vdd.t1473 vdd.n4718 287.382
R5627 vdd.t470 vdd.n4718 287.382
R5628 vdd.t470 vdd.n4720 287.382
R5629 vdd.n4720 vdd.t472 287.382
R5630 vdd.n4741 vdd.t472 287.382
R5631 vdd.t1032 vdd.n4741 287.382
R5632 vdd.n4428 vdd.t1457 287.382
R5633 vdd.t1239 vdd.n4428 287.382
R5634 vdd.n4436 vdd.t1239 287.382
R5635 vdd.n4436 vdd.t1241 287.382
R5636 vdd.n4453 vdd.t1241 287.382
R5637 vdd.t455 vdd.n4453 287.382
R5638 vdd.t827 vdd.n4765 287.382
R5639 vdd.t227 vdd.n4765 287.382
R5640 vdd.t227 vdd.n4767 287.382
R5641 vdd.n4767 vdd.t229 287.382
R5642 vdd.n4788 vdd.t229 287.382
R5643 vdd.t72 vdd.n4788 287.382
R5644 vdd.t52 vdd.n4810 287.382
R5645 vdd.t365 vdd.n4810 287.382
R5646 vdd.t365 vdd.n4812 287.382
R5647 vdd.n4812 vdd.t367 287.382
R5648 vdd.n4833 vdd.t367 287.382
R5649 vdd.t1256 vdd.n4833 287.382
R5650 vdd.t1371 vdd.n4856 287.382
R5651 vdd.t414 vdd.n4856 287.382
R5652 vdd.t414 vdd.n4858 287.382
R5653 vdd.n4858 vdd.t416 287.382
R5654 vdd.n4879 vdd.t416 287.382
R5655 vdd.t411 vdd.n4879 287.382
R5656 vdd.t1487 vdd.n4907 287.382
R5657 vdd.t1227 vdd.n4907 287.382
R5658 vdd.t1227 vdd.n4909 287.382
R5659 vdd.n4909 vdd.t1229 287.382
R5660 vdd.n4930 vdd.t1229 287.382
R5661 vdd.t1090 vdd.n4930 287.382
R5662 vdd.t858 vdd.n4953 287.382
R5663 vdd.t510 vdd.n4953 287.382
R5664 vdd.t510 vdd.n4955 287.382
R5665 vdd.n4955 vdd.t512 287.382
R5666 vdd.n4976 vdd.t512 287.382
R5667 vdd.t1165 vdd.n4976 287.382
R5668 vdd.t1300 vdd.n5001 287.382
R5669 vdd.t1099 vdd.n5001 287.382
R5670 vdd.t1099 vdd.n5003 287.382
R5671 vdd.n5003 vdd.t1101 287.382
R5672 vdd.n5024 vdd.t1101 287.382
R5673 vdd.t308 vdd.n5024 287.382
R5674 vdd.t1010 vdd.n5047 287.382
R5675 vdd.t1167 vdd.n5047 287.382
R5676 vdd.t1167 vdd.n5049 287.382
R5677 vdd.n5049 vdd.t1166 287.382
R5678 vdd.n5070 vdd.t1166 287.382
R5679 vdd.t1412 vdd.n5070 287.382
R5680 vdd.t50 vdd.n5092 287.382
R5681 vdd.t107 vdd.n5092 287.382
R5682 vdd.t107 vdd.n5094 287.382
R5683 vdd.n5094 vdd.t109 287.382
R5684 vdd.n5115 vdd.t109 287.382
R5685 vdd.t607 vdd.n5115 287.382
R5686 vdd.t1043 vdd.n5142 287.382
R5687 vdd.t344 vdd.n5142 287.382
R5688 vdd.t344 vdd.n5144 287.382
R5689 vdd.n5144 vdd.t346 287.382
R5690 vdd.n5165 vdd.t346 287.382
R5691 vdd.t191 vdd.n5165 287.382
R5692 vdd.t942 vdd.n5188 287.382
R5693 vdd.t322 vdd.n5188 287.382
R5694 vdd.t322 vdd.n5190 287.382
R5695 vdd.n5190 vdd.t321 287.382
R5696 vdd.n5211 vdd.t321 287.382
R5697 vdd.t1278 vdd.n5211 287.382
R5698 vdd.t1304 vdd.n5236 287.382
R5699 vdd.t700 vdd.n5236 287.382
R5700 vdd.t700 vdd.n5238 287.382
R5701 vdd.n5238 vdd.t699 287.382
R5702 vdd.n5259 vdd.t699 287.382
R5703 vdd.t537 vdd.n5259 287.382
R5704 vdd.n4193 vdd.t1455 287.382
R5705 vdd.t710 vdd.n4193 287.382
R5706 vdd.n4201 vdd.t710 287.382
R5707 vdd.n4201 vdd.t712 287.382
R5708 vdd.n4218 vdd.t712 287.382
R5709 vdd.t1067 vdd.n4218 287.382
R5710 vdd.t844 vdd.n5283 287.382
R5711 vdd.t1109 vdd.n5283 287.382
R5712 vdd.t1109 vdd.n5285 287.382
R5713 vdd.n5285 vdd.t1111 287.382
R5714 vdd.n5306 vdd.t1111 287.382
R5715 vdd.t888 vdd.n5306 287.382
R5716 vdd.t172 vdd.n5328 287.382
R5717 vdd.t1503 vdd.n5328 287.382
R5718 vdd.t1503 vdd.n5330 287.382
R5719 vdd.n5330 vdd.t1505 287.382
R5720 vdd.n5351 vdd.t1505 287.382
R5721 vdd.t660 vdd.n5351 287.382
R5722 vdd.t456 vdd.n5378 287.382
R5723 vdd.t719 vdd.n5378 287.382
R5724 vdd.t719 vdd.n5380 287.382
R5725 vdd.n5380 vdd.t718 287.382
R5726 vdd.n5401 vdd.t718 287.382
R5727 vdd.t63 vdd.n5401 287.382
R5728 vdd.t1012 vdd.n5424 287.382
R5729 vdd.t500 vdd.n5424 287.382
R5730 vdd.t500 vdd.n5426 287.382
R5731 vdd.n5426 vdd.t499 287.382
R5732 vdd.n5447 vdd.t499 287.382
R5733 vdd.t1411 vdd.n5447 287.382
R5734 vdd.t1051 vdd.n5472 287.382
R5735 vdd.t504 vdd.n5472 287.382
R5736 vdd.t504 vdd.n5474 287.382
R5737 vdd.n5474 vdd.t506 287.382
R5738 vdd.n5495 vdd.t506 287.382
R5739 vdd.t269 vdd.n5495 287.382
R5740 vdd.t716 vdd.n5613 287.382
R5741 vdd.t713 vdd.n5613 287.382
R5742 vdd.t713 vdd.n5605 287.382
R5743 vdd.t714 vdd.n5605 287.382
R5744 vdd.t714 vdd.n5639 287.382
R5745 vdd.n5639 vdd.t906 287.382
R5746 vdd.t1237 vdd.n5567 287.382
R5747 vdd.t185 vdd.n5567 287.382
R5748 vdd.t185 vdd.n5559 287.382
R5749 vdd.t186 vdd.n5559 287.382
R5750 vdd.t186 vdd.n5593 287.382
R5751 vdd.n5593 vdd.t164 287.382
R5752 vdd.t144 vdd.n5660 287.382
R5753 vdd.t396 vdd.n5660 287.382
R5754 vdd.t396 vdd.n5652 287.382
R5755 vdd.t397 vdd.n5652 287.382
R5756 vdd.t397 vdd.n5686 287.382
R5757 vdd.n5686 vdd.t595 287.382
R5758 vdd.t924 vdd.n5708 287.382
R5759 vdd.t1214 vdd.n5708 287.382
R5760 vdd.t1214 vdd.n5700 287.382
R5761 vdd.t1215 vdd.n5700 287.382
R5762 vdd.t1215 vdd.n5734 287.382
R5763 vdd.n5734 vdd.t990 287.382
R5764 vdd.t424 vdd.n5754 287.382
R5765 vdd.t583 vdd.n5754 287.382
R5766 vdd.t583 vdd.n5746 287.382
R5767 vdd.t581 vdd.n5746 287.382
R5768 vdd.t581 vdd.n5780 287.382
R5769 vdd.n5780 vdd.t13 287.382
R5770 vdd.t1422 vdd.n4009 287.382
R5771 vdd.t1517 vdd.n4009 287.382
R5772 vdd.t1517 vdd.n4028 287.382
R5773 vdd.n4028 vdd.t1515 287.382
R5774 vdd.t1515 vdd.n4003 287.382
R5775 vdd.t99 vdd.n4003 287.382
R5776 vdd.t23 vdd.n5896 287.382
R5777 vdd.t330 vdd.n5896 287.382
R5778 vdd.t330 vdd.n5888 287.382
R5779 vdd.t328 vdd.n5888 287.382
R5780 vdd.t328 vdd.n5922 287.382
R5781 vdd.n5922 vdd.t866 287.382
R5782 vdd.t786 vdd.n5849 287.382
R5783 vdd.t1527 vdd.n5849 287.382
R5784 vdd.t1527 vdd.n5841 287.382
R5785 vdd.t1528 vdd.n5841 287.382
R5786 vdd.t1528 vdd.n5875 287.382
R5787 vdd.n5875 vdd.t767 287.382
R5788 vdd.t928 vdd.n5803 287.382
R5789 vdd.t777 vdd.n5803 287.382
R5790 vdd.t777 vdd.n5795 287.382
R5791 vdd.t778 vdd.n5795 287.382
R5792 vdd.t778 vdd.n5829 287.382
R5793 vdd.n5829 vdd.t1373 287.382
R5794 vdd.t679 vdd.n5943 287.382
R5795 vdd.t676 vdd.n5943 287.382
R5796 vdd.t676 vdd.n5935 287.382
R5797 vdd.t677 vdd.n5935 287.382
R5798 vdd.t677 vdd.n5969 287.382
R5799 vdd.n5969 vdd.t1479 287.382
R5800 vdd.t1258 vdd.n5991 287.382
R5801 vdd.t1192 vdd.n5991 287.382
R5802 vdd.t1192 vdd.n5983 287.382
R5803 vdd.t1193 vdd.n5983 287.382
R5804 vdd.t1193 vdd.n6017 287.382
R5805 vdd.n6017 vdd.t1002 287.382
R5806 vdd.t429 vdd.n6037 287.382
R5807 vdd.t2 vdd.n6037 287.382
R5808 vdd.t2 vdd.n6029 287.382
R5809 vdd.t0 vdd.n6029 287.382
R5810 vdd.t0 vdd.n6063 287.382
R5811 vdd.n6063 vdd.t1489 287.382
R5812 vdd.t305 vdd.n6131 287.382
R5813 vdd.t631 vdd.n6131 287.382
R5814 vdd.t631 vdd.n6123 287.382
R5815 vdd.t632 vdd.n6123 287.382
R5816 vdd.t632 vdd.n6157 287.382
R5817 vdd.n6157 vdd.t969 287.382
R5818 vdd.t671 vdd.n6085 287.382
R5819 vdd.t1206 vdd.n6085 287.382
R5820 vdd.t1206 vdd.n6077 287.382
R5821 vdd.t1204 vdd.n6077 287.382
R5822 vdd.t1204 vdd.n6111 287.382
R5823 vdd.n6111 vdd.t434 287.382
R5824 vdd.t387 vdd.n6178 287.382
R5825 vdd.t1157 vdd.n6178 287.382
R5826 vdd.t1157 vdd.n6170 287.382
R5827 vdd.t1158 vdd.n6170 287.382
R5828 vdd.t1158 vdd.n6204 287.382
R5829 vdd.n6204 vdd.t1336 287.382
R5830 vdd.t246 vdd.n6226 287.382
R5831 vdd.t1403 vdd.n6226 287.382
R5832 vdd.t1403 vdd.n6218 287.382
R5833 vdd.t1404 vdd.n6218 287.382
R5834 vdd.t1404 vdd.n6252 287.382
R5835 vdd.n6252 vdd.t32 287.382
R5836 vdd.t1026 vdd.n6272 287.382
R5837 vdd.t944 vdd.n6272 287.382
R5838 vdd.t944 vdd.n6264 287.382
R5839 vdd.t945 vdd.n6264 287.382
R5840 vdd.t945 vdd.n6298 287.382
R5841 vdd.n6298 vdd.t496 287.382
R5842 vdd.t724 vdd.n3773 287.382
R5843 vdd.t721 vdd.n3773 287.382
R5844 vdd.t721 vdd.n3792 287.382
R5845 vdd.n3792 vdd.t722 287.382
R5846 vdd.t722 vdd.n3767 287.382
R5847 vdd.t93 vdd.n3767 287.382
R5848 vdd.t20 vdd.n6367 287.382
R5849 vdd.t17 vdd.n6367 287.382
R5850 vdd.t17 vdd.n6359 287.382
R5851 vdd.t18 vdd.n6359 287.382
R5852 vdd.t18 vdd.n6393 287.382
R5853 vdd.n6393 vdd.t868 287.382
R5854 vdd.t331 vdd.n6321 287.382
R5855 vdd.t749 vdd.n6321 287.382
R5856 vdd.t749 vdd.n6313 287.382
R5857 vdd.t750 vdd.n6313 287.382
R5858 vdd.t750 vdd.n6347 287.382
R5859 vdd.n6347 vdd.t432 287.382
R5860 vdd.t615 vdd.n6414 287.382
R5861 vdd.t686 vdd.n6414 287.382
R5862 vdd.t686 vdd.n6406 287.382
R5863 vdd.t684 vdd.n6406 287.382
R5864 vdd.t684 vdd.n6440 287.382
R5865 vdd.n6440 vdd.t1053 287.382
R5866 vdd.t1367 vdd.n6462 287.382
R5867 vdd.t1169 vdd.n6462 287.382
R5868 vdd.t1169 vdd.n6454 287.382
R5869 vdd.t1170 vdd.n6454 287.382
R5870 vdd.t1170 vdd.n6488 287.382
R5871 vdd.n6488 vdd.t894 287.382
R5872 vdd.t314 vdd.n6508 287.382
R5873 vdd.t121 vdd.n6508 287.382
R5874 vdd.t121 vdd.n6500 287.382
R5875 vdd.t119 vdd.n6500 287.382
R5876 vdd.t119 vdd.n6534 287.382
R5877 vdd.n6534 vdd.t564 287.382
R5878 vdd.t695 vdd.n668 287.382
R5879 vdd.t46 vdd.n668 287.382
R5880 vdd.t46 vdd.n660 287.382
R5881 vdd.t47 vdd.n660 287.382
R5882 vdd.t47 vdd.n694 287.382
R5883 vdd.n694 vdd.t1465 287.382
R5884 vdd.t1406 vdd.n714 287.382
R5885 vdd.t123 vdd.n714 287.382
R5886 vdd.t123 vdd.n706 287.382
R5887 vdd.t124 vdd.n706 287.382
R5888 vdd.t124 vdd.n740 287.382
R5889 vdd.n740 vdd.t1501 287.382
R5890 vdd.t1202 vdd.n812 287.382
R5891 vdd.t291 vdd.n812 287.382
R5892 vdd.t291 vdd.n804 287.382
R5893 vdd.t289 vdd.n804 287.382
R5894 vdd.t289 vdd.n838 287.382
R5895 vdd.n838 vdd.t1358 287.382
R5896 vdd.t1383 vdd.n858 287.382
R5897 vdd.t427 vdd.n858 287.382
R5898 vdd.t427 vdd.n850 287.382
R5899 vdd.t425 vdd.n850 287.382
R5900 vdd.t425 vdd.n884 287.382
R5901 vdd.n884 vdd.t1497 287.382
R5902 vdd.t361 vdd.n904 287.382
R5903 vdd.t215 vdd.n904 287.382
R5904 vdd.t215 vdd.n896 287.382
R5905 vdd.t213 vdd.n896 287.382
R5906 vdd.t213 vdd.n930 287.382
R5907 vdd.n930 vdd.t1312 287.382
R5908 vdd.t236 vdd.n950 287.382
R5909 vdd.t923 vdd.n950 287.382
R5910 vdd.t923 vdd.n942 287.382
R5911 vdd.t921 vdd.n942 287.382
R5912 vdd.t921 vdd.n976 287.382
R5913 vdd.n976 vdd.t462 287.382
R5914 vdd.t1259 vdd.n1048 287.382
R5915 vdd.t957 vdd.n1048 287.382
R5916 vdd.t957 vdd.n1040 287.382
R5917 vdd.t955 vdd.n1040 287.382
R5918 vdd.t955 vdd.n1074 287.382
R5919 vdd.n1074 vdd.t1469 287.382
R5920 vdd.t1213 vdd.n2506 287.382
R5921 vdd.t181 vdd.n2506 287.382
R5922 vdd.t181 vdd.n2498 287.382
R5923 vdd.t179 vdd.n2498 287.382
R5924 vdd.t179 vdd.n2532 287.382
R5925 vdd.n2532 vdd.t381 287.382
R5926 vdd.t3 vdd.n1093 287.382
R5927 vdd.t111 vdd.n1093 287.382
R5928 vdd.t111 vdd.n1095 287.382
R5929 vdd.n1095 vdd.t113 287.382
R5930 vdd.n1116 vdd.t113 287.382
R5931 vdd.t947 vdd.n1116 287.382
R5932 vdd.t195 vdd.n1139 287.382
R5933 vdd.t731 vdd.n1139 287.382
R5934 vdd.t731 vdd.n1141 287.382
R5935 vdd.n1141 vdd.t730 287.382
R5936 vdd.n1162 vdd.t730 287.382
R5937 vdd.t747 vdd.n1162 287.382
R5938 vdd.t1308 vdd.n1236 287.382
R5939 vdd.t1368 vdd.n1236 287.382
R5940 vdd.t1368 vdd.n1238 287.382
R5941 vdd.n1238 vdd.t1370 287.382
R5942 vdd.n1259 vdd.t1370 287.382
R5943 vdd.t86 vdd.n1259 287.382
R5944 vdd.t1495 vdd.n1282 287.382
R5945 vdd.t1103 vdd.n1282 287.382
R5946 vdd.t1103 vdd.n1284 287.382
R5947 vdd.n1284 vdd.t1105 287.382
R5948 vdd.n1305 vdd.t1105 287.382
R5949 vdd.t157 vdd.n1305 287.382
R5950 vdd.t1356 vdd.n1328 287.382
R5951 vdd.t311 vdd.n1328 287.382
R5952 vdd.t311 vdd.n1330 287.382
R5953 vdd.n1330 vdd.t313 287.382
R5954 vdd.n1351 vdd.t313 287.382
R5955 vdd.t65 vdd.n1351 287.382
R5956 vdd.t591 vdd.n1374 287.382
R5957 vdd.t918 vdd.n1374 287.382
R5958 vdd.t918 vdd.n1376 287.382
R5959 vdd.n1376 vdd.t917 287.382
R5960 vdd.n1397 vdd.t917 287.382
R5961 vdd.t920 vdd.n1397 287.382
R5962 vdd.t385 vdd.n1471 287.382
R5963 vdd.t409 vdd.n1471 287.382
R5964 vdd.t409 vdd.n1473 287.382
R5965 vdd.n1473 vdd.t408 287.382
R5966 vdd.n1494 vdd.t408 287.382
R5967 vdd.t1447 vdd.n1494 287.382
R5968 vdd.t552 vdd.n620 287.382
R5969 vdd.t348 vdd.n620 287.382
R5970 vdd.t348 vdd.n622 287.382
R5971 vdd.n622 vdd.t347 287.382
R5972 vdd.n643 vdd.t347 287.382
R5973 vdd.t893 vdd.n643 287.382
R5974 vdd.t823 vdd.n1515 287.382
R5975 vdd.t1222 vdd.n1515 287.382
R5976 vdd.t1222 vdd.n1517 287.382
R5977 vdd.n1517 vdd.t1224 287.382
R5978 vdd.n1538 vdd.t1224 287.382
R5979 vdd.t1142 vdd.n1538 287.382
R5980 vdd.t833 vdd.n1560 287.382
R5981 vdd.t1188 vdd.n1560 287.382
R5982 vdd.t1188 vdd.n1562 287.382
R5983 vdd.n1562 vdd.t1190 287.382
R5984 vdd.n1583 vdd.t1190 287.382
R5985 vdd.t1121 vdd.n1583 287.382
R5986 vdd.t466 vdd.n1610 287.382
R5987 vdd.t1068 vdd.n1610 287.382
R5988 vdd.t1068 vdd.n1612 287.382
R5989 vdd.n1612 vdd.t1070 287.382
R5990 vdd.n1633 vdd.t1070 287.382
R5991 vdd.t1033 vdd.n1633 287.382
R5992 vdd.t998 vdd.n1656 287.382
R5993 vdd.t953 vdd.n1656 287.382
R5994 vdd.t953 vdd.n1658 287.382
R5995 vdd.n1658 vdd.t952 287.382
R5996 vdd.n1679 vdd.t952 287.382
R5997 vdd.t309 vdd.n1679 287.382
R5998 vdd.t1493 vdd.n1704 287.382
R5999 vdd.t83 vdd.n1704 287.382
R6000 vdd.t83 vdd.n1706 287.382
R6001 vdd.n1706 vdd.t85 287.382
R6002 vdd.n1727 vdd.t85 287.382
R6003 vdd.t1018 vdd.n1727 287.382
R6004 vdd.n1414 vdd.t101 287.382
R6005 vdd.t1072 vdd.n1414 287.382
R6006 vdd.n1422 vdd.t1072 287.382
R6007 vdd.n1422 vdd.t1074 287.382
R6008 vdd.n1439 vdd.t1074 287.382
R6009 vdd.t1443 vdd.n1439 287.382
R6010 vdd.t870 vdd.n1751 287.382
R6011 vdd.t664 vdd.n1751 287.382
R6012 vdd.t664 vdd.n1753 287.382
R6013 vdd.n1753 vdd.t666 287.382
R6014 vdd.n1774 vdd.t666 287.382
R6015 vdd.t683 vdd.n1774 287.382
R6016 vdd.t170 vdd.n1796 287.382
R6017 vdd.t368 vdd.n1796 287.382
R6018 vdd.t368 vdd.n1798 287.382
R6019 vdd.n1798 vdd.t370 287.382
R6020 vdd.n1819 vdd.t370 287.382
R6021 vdd.t132 vdd.n1819 287.382
R6022 vdd.t1127 vdd.n1842 287.382
R6023 vdd.t654 vdd.n1842 287.382
R6024 vdd.t654 vdd.n1844 287.382
R6025 vdd.n1844 vdd.t656 287.382
R6026 vdd.n1865 vdd.t656 287.382
R6027 vdd.t657 vdd.n1865 287.382
R6028 vdd.t1324 vdd.n1893 287.382
R6029 vdd.t787 vdd.n1893 287.382
R6030 vdd.t787 vdd.n1895 287.382
R6031 vdd.n1895 vdd.t789 287.382
R6032 vdd.n1916 vdd.t789 287.382
R6033 vdd.t1283 vdd.n1916 287.382
R6034 vdd.t992 vdd.n1939 287.382
R6035 vdd.t388 vdd.n1939 287.382
R6036 vdd.t388 vdd.n1941 287.382
R6037 vdd.n1941 vdd.t390 287.382
R6038 vdd.n1962 vdd.t390 287.382
R6039 vdd.t391 vdd.n1962 287.382
R6040 vdd.t371 vdd.n1987 287.382
R6041 vdd.t158 vdd.n1987 287.382
R6042 vdd.t158 vdd.n1989 287.382
R6043 vdd.n1989 vdd.t160 287.382
R6044 vdd.n2010 vdd.t160 287.382
R6045 vdd.t268 vdd.n2010 287.382
R6046 vdd.t971 vdd.n2033 287.382
R6047 vdd.t1218 vdd.n2033 287.382
R6048 vdd.t1218 vdd.n2035 287.382
R6049 vdd.n2035 vdd.t1217 287.382
R6050 vdd.n2056 vdd.t1217 287.382
R6051 vdd.t1220 vdd.n2056 287.382
R6052 vdd.t168 vdd.n2078 287.382
R6053 vdd.t841 vdd.n2078 287.382
R6054 vdd.t841 vdd.n2080 287.382
R6055 vdd.n2080 vdd.t843 287.382
R6056 vdd.n2101 vdd.t843 287.382
R6057 vdd.t226 vdd.n2101 287.382
R6058 vdd.t1344 vdd.n2128 287.382
R6059 vdd.t635 vdd.n2128 287.382
R6060 vdd.t635 vdd.n2130 287.382
R6061 vdd.n2130 vdd.t637 287.382
R6062 vdd.n2151 vdd.t637 287.382
R6063 vdd.t110 vdd.n2151 287.382
R6064 vdd.t940 vdd.n2174 287.382
R6065 vdd.t232 vdd.n2174 287.382
R6066 vdd.t232 vdd.n2176 287.382
R6067 vdd.n2176 vdd.t231 287.382
R6068 vdd.n2197 vdd.t231 287.382
R6069 vdd.t1131 vdd.n2197 287.382
R6070 vdd.t1481 vdd.n2222 287.382
R6071 vdd.t1116 vdd.n2222 287.382
R6072 vdd.t1116 vdd.n2224 287.382
R6073 vdd.n2224 vdd.t1118 287.382
R6074 vdd.n2245 vdd.t1118 287.382
R6075 vdd.t1119 vdd.n2245 287.382
R6076 vdd.n1179 vdd.t95 287.382
R6077 vdd.t672 vdd.n1179 287.382
R6078 vdd.n1187 vdd.t672 287.382
R6079 vdd.n1187 vdd.t674 287.382
R6080 vdd.n1204 vdd.t674 287.382
R6081 vdd.t1163 vdd.n1204 287.382
R6082 vdd.t900 vdd.n2269 287.382
R6083 vdd.t296 vdd.n2269 287.382
R6084 vdd.t296 vdd.n2271 287.382
R6085 vdd.n2271 vdd.t298 287.382
R6086 vdd.n2292 vdd.t298 287.382
R6087 vdd.t929 vdd.n2292 287.382
R6088 vdd.t771 vdd.n2314 287.382
R6089 vdd.t116 vdd.n2314 287.382
R6090 vdd.t116 vdd.n2316 287.382
R6091 vdd.n2316 vdd.t118 287.382
R6092 vdd.n2337 vdd.t118 287.382
R6093 vdd.t516 vdd.n2337 287.382
R6094 vdd.t492 vdd.n2364 287.382
R6095 vdd.t1038 vdd.n2364 287.382
R6096 vdd.t1038 vdd.n2366 287.382
R6097 vdd.n2366 vdd.t1040 287.382
R6098 vdd.n2387 vdd.t1040 287.382
R6099 vdd.t103 vdd.n2387 287.382
R6100 vdd.t975 vdd.n2410 287.382
R6101 vdd.t875 vdd.n2410 287.382
R6102 vdd.t875 vdd.n2412 287.382
R6103 vdd.n2412 vdd.t877 287.382
R6104 vdd.n2433 vdd.t877 287.382
R6105 vdd.t606 vdd.n2433 287.382
R6106 vdd.t1348 vdd.n2458 287.382
R6107 vdd.t1444 vdd.n2458 287.382
R6108 vdd.t1444 vdd.n2460 287.382
R6109 vdd.n2460 vdd.t1446 287.382
R6110 vdd.n2481 vdd.t1446 287.382
R6111 vdd.t1423 vdd.n2481 287.382
R6112 vdd.t423 vdd.n2599 287.382
R6113 vdd.t526 vdd.n2599 287.382
R6114 vdd.t526 vdd.n2591 287.382
R6115 vdd.t524 vdd.n2591 287.382
R6116 vdd.t524 vdd.n2625 287.382
R6117 vdd.n2625 vdd.t815 287.382
R6118 vdd.t1027 vdd.n2553 287.382
R6119 vdd.t334 vdd.n2553 287.382
R6120 vdd.t334 vdd.n2545 287.382
R6121 vdd.t332 vdd.n2545 287.382
R6122 vdd.t332 vdd.n2579 287.382
R6123 vdd.n2579 vdd.t769 287.382
R6124 vdd.t916 vdd.n2646 287.382
R6125 vdd.t618 vdd.n2646 287.382
R6126 vdd.t618 vdd.n2638 287.382
R6127 vdd.t616 vdd.n2638 287.382
R6128 vdd.t616 vdd.n2672 287.382
R6129 vdd.n2672 vdd.t1350 287.382
R6130 vdd.t717 vdd.n2694 287.382
R6131 vdd.t1098 vdd.n2694 287.382
R6132 vdd.t1098 vdd.n2686 287.382
R6133 vdd.t1096 vdd.n2686 287.382
R6134 vdd.t1096 vdd.n2720 287.382
R6135 vdd.n2720 vdd.t1016 287.382
R6136 vdd.t392 vdd.n2740 287.382
R6137 vdd.t1141 vdd.n2740 287.382
R6138 vdd.t1141 vdd.n2732 287.382
R6139 vdd.t1139 vdd.n2732 287.382
R6140 vdd.t1139 vdd.n2766 287.382
R6141 vdd.n2766 vdd.t494 287.382
R6142 vdd.t1230 vdd.n995 287.382
R6143 vdd.t404 vdd.n995 287.382
R6144 vdd.t404 vdd.n1014 287.382
R6145 vdd.n1014 vdd.t402 287.382
R6146 vdd.t402 vdd.n989 287.382
R6147 vdd.t91 vdd.n989 287.382
R6148 vdd.t445 vdd.n2882 287.382
R6149 vdd.t75 vdd.n2882 287.382
R6150 vdd.t75 vdd.n2874 287.382
R6151 vdd.t73 vdd.n2874 287.382
R6152 vdd.t73 vdd.n2908 287.382
R6153 vdd.n2908 vdd.t44 287.382
R6154 vdd.t1106 vdd.n2835 287.382
R6155 vdd.t133 vdd.n2835 287.382
R6156 vdd.t133 vdd.n2827 287.382
R6157 vdd.t134 vdd.n2827 287.382
R6158 vdd.t134 vdd.n2861 287.382
R6159 vdd.n2861 vdd.t438 287.382
R6160 vdd.t729 vdd.n2789 287.382
R6161 vdd.t614 vdd.n2789 287.382
R6162 vdd.t614 vdd.n2781 287.382
R6163 vdd.t612 vdd.n2781 287.382
R6164 vdd.t612 vdd.n2815 287.382
R6165 vdd.n2815 vdd.t1125 287.382
R6166 vdd.t605 vdd.n2929 287.382
R6167 vdd.t222 vdd.n2929 287.382
R6168 vdd.t222 vdd.n2921 287.382
R6169 vdd.t220 vdd.n2921 287.382
R6170 vdd.t220 vdd.n2955 287.382
R6171 vdd.n2955 vdd.t11 287.382
R6172 vdd.t1221 vdd.n2977 287.382
R6173 vdd.t1386 vdd.n2977 287.382
R6174 vdd.t1386 vdd.n2969 287.382
R6175 vdd.t1384 vdd.n2969 287.382
R6176 vdd.t1384 vdd.n3003 287.382
R6177 vdd.n3003 vdd.t38 287.382
R6178 vdd.t1434 vdd.n3023 287.382
R6179 vdd.t454 vdd.n3023 287.382
R6180 vdd.t454 vdd.n3015 287.382
R6181 vdd.t452 vdd.n3015 287.382
R6182 vdd.t452 vdd.n3049 287.382
R6183 vdd.n3049 vdd.t1296 287.382
R6184 vdd.t1156 vdd.n3117 287.382
R6185 vdd.t801 vdd.n3117 287.382
R6186 vdd.t801 vdd.n3109 287.382
R6187 vdd.t799 vdd.n3109 287.382
R6188 vdd.t799 vdd.n3143 287.382
R6189 vdd.n3143 vdd.t852 287.382
R6190 vdd.t21 vdd.n3071 287.382
R6191 vdd.t276 vdd.n3071 287.382
R6192 vdd.t276 vdd.n3063 287.382
R6193 vdd.t274 vdd.n3063 287.382
R6194 vdd.t274 vdd.n3097 287.382
R6195 vdd.n3097 vdd.t790 287.382
R6196 vdd.t245 vdd.n3164 287.382
R6197 vdd.t280 vdd.n3164 287.382
R6198 vdd.t280 vdd.n3156 287.382
R6199 vdd.t278 vdd.n3156 287.382
R6200 vdd.t278 vdd.n3190 287.382
R6201 vdd.n3190 vdd.t373 287.382
R6202 vdd.t1282 vdd.n3212 287.382
R6203 vdd.t1212 vdd.n3212 287.382
R6204 vdd.t1212 vdd.n3204 287.382
R6205 vdd.t1210 vdd.n3204 287.382
R6206 vdd.t1210 vdd.n3238 287.382
R6207 vdd.n3238 vdd.t967 287.382
R6208 vdd.t798 vdd.n3258 287.382
R6209 vdd.t1277 vdd.n3258 287.382
R6210 vdd.t1277 vdd.n3250 287.382
R6211 vdd.t1275 vdd.n3250 287.382
R6212 vdd.t1275 vdd.n3284 287.382
R6213 vdd.n3284 vdd.t1328 287.382
R6214 vdd.t1410 vdd.n759 287.382
R6215 vdd.t1433 vdd.n759 287.382
R6216 vdd.t1433 vdd.n778 287.382
R6217 vdd.n778 vdd.t1431 287.382
R6218 vdd.t1431 vdd.n753 287.382
R6219 vdd.t87 vdd.n753 287.382
R6220 vdd.t1203 vdd.n3353 287.382
R6221 vdd.t265 vdd.n3353 287.382
R6222 vdd.t265 vdd.n3345 287.382
R6223 vdd.t266 vdd.n3345 287.382
R6224 vdd.t266 vdd.n3379 287.382
R6225 vdd.n3379 vdd.t819 287.382
R6226 vdd.t310 vdd.n3307 287.382
R6227 vdd.t1508 vdd.n3307 287.382
R6228 vdd.t1508 vdd.n3299 287.382
R6229 vdd.t1509 vdd.n3299 287.382
R6230 vdd.t1509 vdd.n3333 287.382
R6231 vdd.n3333 vdd.t436 287.382
R6232 vdd.t1124 vdd.n3400 287.382
R6233 vdd.t1137 vdd.n3400 287.382
R6234 vdd.t1137 vdd.n3392 287.382
R6235 vdd.t1135 vdd.n3392 287.382
R6236 vdd.t1135 vdd.n3426 287.382
R6237 vdd.n3426 vdd.t1332 287.382
R6238 vdd.t1061 vdd.n3448 287.382
R6239 vdd.t648 vdd.n3448 287.382
R6240 vdd.t648 vdd.n3440 287.382
R6241 vdd.t649 vdd.n3440 287.382
R6242 vdd.t649 vdd.n3474 287.382
R6243 vdd.n3474 vdd.t904 287.382
R6244 vdd.t1123 vdd.n3494 287.382
R6245 vdd.t830 vdd.n3494 287.382
R6246 vdd.t830 vdd.n3486 287.382
R6247 vdd.t831 vdd.n3486 287.382
R6248 vdd.t831 vdd.n3520 287.382
R6249 vdd.n3520 vdd.t488 287.382
R6250 vdd.t748 vdd.n576 287.382
R6251 vdd.t1153 vdd.n576 287.382
R6252 vdd.t1153 vdd.n568 287.382
R6253 vdd.t1151 vdd.n568 287.382
R6254 vdd.t1151 vdd.n602 287.382
R6255 vdd.n602 vdd.t30 287.382
R6256 vdd.t1382 vdd.n3589 287.382
R6257 vdd.t1428 vdd.n3589 287.382
R6258 vdd.t1428 vdd.n3581 287.382
R6259 vdd.t1429 vdd.n3581 287.382
R6260 vdd.t1429 vdd.n3615 287.382
R6261 vdd.n3615 vdd.t24 287.382
R6262 vdd.t1150 vdd.n3543 287.382
R6263 vdd.t1172 vdd.n3543 287.382
R6264 vdd.t1172 vdd.n3535 287.382
R6265 vdd.t1173 vdd.n3535 287.382
R6266 vdd.t1173 vdd.n3569 287.382
R6267 vdd.n3569 vdd.t986 287.382
R6268 vdd.t1095 vdd.n6603 287.382
R6269 vdd.t709 vdd.n6603 287.382
R6270 vdd.t709 vdd.n6595 287.382
R6271 vdd.t707 vdd.n6595 287.382
R6272 vdd.t707 vdd.n6629 287.382
R6273 vdd.n6629 vdd.t28 287.382
R6274 vdd.t1243 vdd.n6557 287.382
R6275 vdd.t549 vdd.n6557 287.382
R6276 vdd.t549 vdd.n6549 287.382
R6277 vdd.t550 vdd.n6549 287.382
R6278 vdd.t550 vdd.n6583 287.382
R6279 vdd.n6583 vdd.t1186 287.382
R6280 vdd.t706 vdd.n9617 287.382
R6281 vdd.t912 vdd.n9617 287.382
R6282 vdd.t912 vdd.n9609 287.382
R6283 vdd.t910 vdd.n9609 287.382
R6284 vdd.t910 vdd.n9643 287.382
R6285 vdd.n9643 vdd.t26 287.382
R6286 vdd.t237 vdd.n9571 287.382
R6287 vdd.t1113 vdd.n9571 287.382
R6288 vdd.t1113 vdd.n9563 287.382
R6289 vdd.t1114 vdd.n9563 287.382
R6290 vdd.t1114 vdd.n9597 287.382
R6291 vdd.n9597 vdd.t984 287.382
R6292 vdd.t1514 vdd.n9663 287.382
R6293 vdd.t1511 vdd.n9663 287.382
R6294 vdd.t1511 vdd.n9655 287.382
R6295 vdd.t1512 vdd.n9655 287.382
R6296 vdd.t1512 vdd.n9689 287.382
R6297 vdd.n9689 vdd.t1354 287.382
R6298 vdd.t71 vdd.n9709 287.382
R6299 vdd.t1387 vdd.n9709 287.382
R6300 vdd.t1387 vdd.n9701 287.382
R6301 vdd.t1388 vdd.n9701 287.382
R6302 vdd.t1388 vdd.n9735 287.382
R6303 vdd.n9735 vdd.t1322 287.382
R6304 vdd.t360 vdd.n9807 287.382
R6305 vdd.t727 vdd.n9807 287.382
R6306 vdd.t727 vdd.n9799 287.382
R6307 vdd.t725 vdd.n9799 287.382
R6308 vdd.t725 vdd.n9833 287.382
R6309 vdd.n9833 vdd.t478 287.382
R6310 vdd.t1284 vdd.n9853 287.382
R6311 vdd.t1179 vdd.n9853 287.382
R6312 vdd.t1179 vdd.n9845 287.382
R6313 vdd.t1180 vdd.n9845 287.382
R6314 vdd.t1180 vdd.n9879 287.382
R6315 vdd.n9879 vdd.t1059 287.382
R6316 vdd.t1023 vdd.n9899 287.382
R6317 vdd.t259 vdd.n9899 287.382
R6318 vdd.t259 vdd.n9891 287.382
R6319 vdd.t257 vdd.n9891 287.382
R6320 vdd.t257 vdd.n9925 287.382
R6321 vdd.n9925 vdd.t15 287.382
R6322 vdd.t960 vdd.n9945 287.382
R6323 vdd.t62 vdd.n9945 287.382
R6324 vdd.t62 vdd.n9937 287.382
R6325 vdd.t60 vdd.n9937 287.382
R6326 vdd.t60 vdd.n9971 287.382
R6327 vdd.n9971 vdd.t490 287.382
R6328 vdd.t548 vdd.n10043 287.382
R6329 vdd.t337 vdd.n10043 287.382
R6330 vdd.t337 vdd.n10035 287.382
R6331 vdd.t338 vdd.n10035 287.382
R6332 vdd.t338 vdd.n10069 287.382
R6333 vdd.n10069 vdd.t1334 287.382
R6334 vdd.t422 vdd.n59 287.382
R6335 vdd.t242 vdd.n59 287.382
R6336 vdd.t242 vdd.n51 287.382
R6337 vdd.t243 vdd.n51 287.382
R6338 vdd.t243 vdd.n85 287.382
R6339 vdd.n85 vdd.t1008 287.382
R6340 vdd.t260 vdd.n13 287.382
R6341 vdd.t653 vdd.n13 287.382
R6342 vdd.t653 vdd.n5 287.382
R6343 vdd.t651 vdd.n5 287.382
R6344 vdd.t651 vdd.n39 287.382
R6345 vdd.n39 vdd.t839 287.382
R6346 vdd.t1164 vdd.n10089 287.382
R6347 vdd.t1087 vdd.n10089 287.382
R6348 vdd.t1087 vdd.n10081 287.382
R6349 vdd.t1085 vdd.n10081 287.382
R6350 vdd.t1085 vdd.n10115 287.382
R6351 vdd.n10115 vdd.t568 287.382
R6352 vdd.t1438 vdd.n10137 287.382
R6353 vdd.t780 vdd.n10137 287.382
R6354 vdd.t780 vdd.n10129 287.382
R6355 vdd.t781 vdd.n10129 287.382
R6356 vdd.t781 vdd.n10163 287.382
R6357 vdd.n10163 vdd.t908 287.382
R6358 vdd.t418 vdd.n10183 287.382
R6359 vdd.t1020 vdd.n10183 287.382
R6360 vdd.t1020 vdd.n10175 287.382
R6361 vdd.t1021 vdd.n10175 287.382
R6362 vdd.t1021 vdd.n10209 287.382
R6363 vdd.n10209 vdd.t597 287.382
R6364 vdd.t694 vdd.n9990 287.382
R6365 vdd.t1397 vdd.n9990 287.382
R6366 vdd.t1397 vdd.n10009 287.382
R6367 vdd.n10009 vdd.t1398 287.382
R6368 vdd.t1398 vdd.n9984 287.382
R6369 vdd.t575 vdd.n9984 287.382
R6370 vdd.t702 vdd.n10325 287.382
R6371 vdd.t687 vdd.n10325 287.382
R6372 vdd.t687 vdd.n10317 287.382
R6373 vdd.t688 vdd.n10317 287.382
R6374 vdd.t688 vdd.n10351 287.382
R6375 vdd.n10351 vdd.t938 287.382
R6376 vdd.t502 vdd.n10278 287.382
R6377 vdd.t299 vdd.n10278 287.382
R6378 vdd.t299 vdd.n10270 287.382
R6379 vdd.t300 vdd.n10270 287.382
R6380 vdd.t300 vdd.n10304 287.382
R6381 vdd.n10304 vdd.t54 287.382
R6382 vdd.t659 vdd.n10232 287.382
R6383 vdd.t1416 vdd.n10232 287.382
R6384 vdd.t1416 vdd.n10224 287.382
R6385 vdd.t1417 vdd.n10224 287.382
R6386 vdd.t1417 vdd.n10258 287.382
R6387 vdd.n10258 vdd.t1379 287.382
R6388 vdd.t1138 vdd.n10372 287.382
R6389 vdd.t354 vdd.n10372 287.382
R6390 vdd.t354 vdd.n10364 287.382
R6391 vdd.t355 vdd.n10364 287.382
R6392 vdd.t355 vdd.n10398 287.382
R6393 vdd.n10398 vdd.t383 287.382
R6394 vdd.t1454 vdd.n10420 287.382
R6395 vdd.t1400 vdd.n10420 287.382
R6396 vdd.t1400 vdd.n10412 287.382
R6397 vdd.t1401 vdd.n10412 287.382
R6398 vdd.t1401 vdd.n10446 287.382
R6399 vdd.n10446 vdd.t846 287.382
R6400 vdd.t1257 vdd.n10466 287.382
R6401 vdd.t803 vdd.n10466 287.382
R6402 vdd.t803 vdd.n10458 287.382
R6403 vdd.t804 vdd.n10458 287.382
R6404 vdd.t804 vdd.n10492 287.382
R6405 vdd.n10492 vdd.t1306 287.382
R6406 vdd.t1366 vdd.n10560 287.382
R6407 vdd.t1260 vdd.n10560 287.382
R6408 vdd.t1260 vdd.n10552 287.382
R6409 vdd.t1261 vdd.n10552 287.382
R6410 vdd.t1261 vdd.n10586 287.382
R6411 vdd.n10586 vdd.t1004 287.382
R6412 vdd.t1102 vdd.n10514 287.382
R6413 vdd.t261 vdd.n10514 287.382
R6414 vdd.t261 vdd.n10506 287.382
R6415 vdd.t262 vdd.n10506 287.382
R6416 vdd.t262 vdd.n10540 287.382
R6417 vdd.n10540 vdd.t775 287.382
R6418 vdd.t1019 vdd.n10607 287.382
R6419 vdd.t1077 vdd.n10607 287.382
R6420 vdd.t1077 vdd.n10599 287.382
R6421 vdd.t1075 vdd.n10599 287.382
R6422 vdd.t1075 vdd.n10633 287.382
R6423 vdd.n10633 vdd.t1491 287.382
R6424 vdd.t253 vdd.n10655 287.382
R6425 vdd.t610 vdd.n10655 287.382
R6426 vdd.t610 vdd.n10647 287.382
R6427 vdd.t608 vdd.n10647 287.382
R6428 vdd.t608 vdd.n10681 287.382
R6429 vdd.n10681 vdd.t817 287.382
R6430 vdd.t292 vdd.n10701 287.382
R6431 vdd.t146 vdd.n10701 287.382
R6432 vdd.t146 vdd.n10693 287.382
R6433 vdd.t147 vdd.n10693 287.382
R6434 vdd.t147 vdd.n10727 287.382
R6435 vdd.n10727 vdd.t1352 287.382
R6436 vdd.t964 vdd.n9754 287.382
R6437 vdd.t1363 vdd.n9754 287.382
R6438 vdd.t1363 vdd.n9773 287.382
R6439 vdd.n9773 vdd.t1364 287.382
R6440 vdd.t1364 vdd.n9748 287.382
R6441 vdd.t1461 vdd.n9748 287.382
R6442 vdd.t742 vdd.n10796 287.382
R6443 vdd.t1234 vdd.n10796 287.382
R6444 vdd.t1234 vdd.n10788 287.382
R6445 vdd.t1235 vdd.n10788 287.382
R6446 vdd.t1235 vdd.n10822 287.382
R6447 vdd.n10822 vdd.t902 287.382
R6448 vdd.t1247 vdd.n10750 287.382
R6449 vdd.t1244 vdd.n10750 287.382
R6450 vdd.t1244 vdd.n10742 287.382
R6451 vdd.t1245 vdd.n10742 287.382
R6452 vdd.t1245 vdd.n10776 287.382
R6453 vdd.n10776 vdd.t629 287.382
R6454 vdd.t417 vdd.n10843 287.382
R6455 vdd.t1162 vdd.n10843 287.382
R6456 vdd.t1162 vdd.n10835 287.382
R6457 vdd.t1160 vdd.n10835 287.382
R6458 vdd.t1160 vdd.n10869 287.382
R6459 vdd.n10869 vdd.t480 287.382
R6460 vdd.t285 vdd.n10891 287.382
R6461 vdd.t948 vdd.n10891 287.382
R6462 vdd.t948 vdd.n10883 287.382
R6463 vdd.t949 vdd.n10883 287.382
R6464 vdd.t949 vdd.n10917 287.382
R6465 vdd.n10917 vdd.t936 287.382
R6466 vdd.t690 vdd.n10937 287.382
R6467 vdd.t1196 vdd.n10937 287.382
R6468 vdd.t1196 vdd.n10929 287.382
R6469 vdd.t1197 vdd.n10929 287.382
R6470 vdd.t1197 vdd.n10963 287.382
R6471 vdd.n10963 vdd.t5 287.382
R6472 vdd.t821 vdd.n10983 287.382
R6473 vdd.t286 vdd.n10983 287.382
R6474 vdd.t286 vdd.n10985 287.382
R6475 vdd.n10985 vdd.t288 287.382
R6476 vdd.n11006 vdd.t288 287.382
R6477 vdd.t498 vdd.n11006 287.382
R6478 vdd.t58 vdd.n11028 287.382
R6479 vdd.t645 vdd.n11028 287.382
R6480 vdd.t645 vdd.n11030 287.382
R6481 vdd.n11030 vdd.t647 287.382
R6482 vdd.n11051 vdd.t647 287.382
R6483 vdd.t1251 vdd.n11051 287.382
R6484 vdd.t1499 vdd.n11078 287.382
R6485 vdd.t733 vdd.n11078 287.382
R6486 vdd.t733 vdd.n11080 287.382
R6487 vdd.n11080 vdd.t735 287.382
R6488 vdd.n11101 vdd.t735 287.382
R6489 vdd.t538 vdd.n11101 287.382
R6490 vdd.t996 vdd.n11124 287.382
R6491 vdd.t294 vdd.n11124 287.382
R6492 vdd.t294 vdd.n11126 287.382
R6493 vdd.n11126 vdd.t293 287.382
R6494 vdd.n11147 vdd.t293 287.382
R6495 vdd.t539 vdd.n11147 287.382
R6496 vdd.t1294 vdd.n11172 287.382
R6497 vdd.t350 vdd.n11172 287.382
R6498 vdd.t350 vdd.n11174 287.382
R6499 vdd.n11174 vdd.t352 287.382
R6500 vdd.n11195 vdd.t352 287.382
R6501 vdd.t216 vdd.n11195 287.382
R6502 vdd.n426 vdd.t579 287.382
R6503 vdd.t740 vdd.n426 287.382
R6504 vdd.n434 vdd.t740 287.382
R6505 vdd.n434 vdd.t739 287.382
R6506 vdd.n451 vdd.t739 287.382
R6507 vdd.t1122 vdd.n451 287.382
R6508 vdd.t965 vdd.n11219 287.382
R6509 vdd.t514 vdd.n11219 287.382
R6510 vdd.t514 vdd.n11221 287.382
R6511 vdd.n11221 vdd.t513 287.382
R6512 vdd.n11242 vdd.t513 287.382
R6513 vdd.t115 vdd.n11242 287.382
R6514 vdd.t796 vdd.n11264 287.382
R6515 vdd.t889 vdd.n11264 287.382
R6516 vdd.t889 vdd.n11266 287.382
R6517 vdd.n11266 vdd.t891 287.382
R6518 vdd.n11287 vdd.t891 287.382
R6519 vdd.t531 vdd.n11287 287.382
R6520 vdd.t1377 vdd.n11310 287.382
R6521 vdd.t405 vdd.n11310 287.382
R6522 vdd.t405 vdd.n11312 287.382
R6523 vdd.n11312 vdd.t407 287.382
R6524 vdd.n11333 vdd.t407 287.382
R6525 vdd.t1037 vdd.n11333 287.382
R6526 vdd.t199 vdd.n11361 287.382
R6527 vdd.t1145 vdd.n11361 287.382
R6528 vdd.t1145 vdd.n11363 287.382
R6529 vdd.n11363 vdd.t1144 287.382
R6530 vdd.n11384 vdd.t1144 287.382
R6531 vdd.t1147 vdd.n11384 287.382
R6532 vdd.t850 vdd.n11407 287.382
R6533 vdd.t282 vdd.n11407 287.382
R6534 vdd.t282 vdd.n11409 287.382
R6535 vdd.n11409 vdd.t281 287.382
R6536 vdd.n11430 vdd.t281 287.382
R6537 vdd.t958 vdd.n11430 287.382
R6538 vdd.t1340 vdd.n11455 287.382
R6539 vdd.t1521 vdd.n11455 287.382
R6540 vdd.t1521 vdd.n11457 287.382
R6541 vdd.n11457 vdd.t1523 287.382
R6542 vdd.n11478 vdd.t1523 287.382
R6543 vdd.t1242 vdd.n11478 287.382
R6544 vdd.t811 vdd.n11501 287.382
R6545 vdd.t270 vdd.n11501 287.382
R6546 vdd.t270 vdd.n11503 287.382
R6547 vdd.n11503 vdd.t272 287.382
R6548 vdd.n11524 vdd.t272 287.382
R6549 vdd.t273 vdd.n11524 287.382
R6550 vdd.t794 vdd.n11546 287.382
R6551 vdd.t1439 vdd.n11546 287.382
R6552 vdd.t1439 vdd.n11548 287.382
R6553 vdd.n11548 vdd.t1441 287.382
R6554 vdd.n11569 vdd.t1441 287.382
R6555 vdd.t307 vdd.n11569 287.382
R6556 vdd.t1286 vdd.n11596 287.382
R6557 vdd.t1390 vdd.n11596 287.382
R6558 vdd.t1390 vdd.n11598 287.382
R6559 vdd.n11598 vdd.t1392 287.382
R6560 vdd.n11619 vdd.t1392 287.382
R6561 vdd.t535 vdd.n11619 287.382
R6562 vdd.t994 vdd.n11642 287.382
R6563 vdd.t1248 vdd.n11642 287.382
R6564 vdd.t1248 vdd.n11644 287.382
R6565 vdd.n11644 vdd.t1250 287.382
R6566 vdd.n11665 vdd.t1250 287.382
R6567 vdd.t641 vdd.n11665 287.382
R6568 vdd.t1338 vdd.n11690 287.382
R6569 vdd.t528 vdd.n11690 287.382
R6570 vdd.t528 vdd.n11692 287.382
R6571 vdd.n11692 vdd.t530 287.382
R6572 vdd.n11713 vdd.t530 287.382
R6573 vdd.t1120 vdd.n11713 287.382
R6574 vdd.n191 vdd.t577 287.382
R6575 vdd.t141 vdd.n191 287.382
R6576 vdd.n199 vdd.t141 287.382
R6577 vdd.n199 vdd.t140 287.382
R6578 vdd.n216 vdd.t140 287.382
R6579 vdd.t1381 vdd.n216 287.382
R6580 vdd.t1014 vdd.n11737 287.382
R6581 vdd.t357 vdd.n11737 287.382
R6582 vdd.t357 vdd.n11739 287.382
R6583 vdd.n11739 vdd.t359 287.382
R6584 vdd.n11760 vdd.t359 287.382
R6585 vdd.t49 vdd.n11760 287.382
R6586 vdd.t792 vdd.n11782 287.382
R6587 vdd.t104 vdd.n11782 287.382
R6588 vdd.t104 vdd.n11784 287.382
R6589 vdd.n11784 vdd.t106 287.382
R6590 vdd.n11805 vdd.t106 287.382
R6591 vdd.t1396 vdd.n11805 287.382
R6592 vdd.t1320 vdd.n11832 287.382
R6593 vdd.t316 vdd.n11832 287.382
R6594 vdd.t316 vdd.n11834 287.382
R6595 vdd.n11834 vdd.t315 287.382
R6596 vdd.n11855 vdd.t315 287.382
R6597 vdd.t1271 vdd.n11855 287.382
R6598 vdd.t813 vdd.n11878 287.382
R6599 vdd.t752 vdd.n11878 287.382
R6600 vdd.t752 vdd.n11880 287.382
R6601 vdd.n11880 vdd.t754 287.382
R6602 vdd.n11901 vdd.t754 287.382
R6603 vdd.t619 vdd.n11901 287.382
R6604 vdd.t1292 vdd.n11926 287.382
R6605 vdd.t340 vdd.n11926 287.382
R6606 vdd.t340 vdd.n11928 287.382
R6607 vdd.n11928 vdd.t342 287.382
R6608 vdd.n11949 vdd.t342 287.382
R6609 vdd.t1071 vdd.n11949 287.382
R6610 vdd.n110 vdd.n109 242.685
R6611 vdd.n156 vdd.n155 242.685
R6612 vdd.n253 vdd.n252 242.685
R6613 vdd.n299 vdd.n298 242.685
R6614 vdd.n345 vdd.n344 242.685
R6615 vdd.n391 vdd.n390 242.685
R6616 vdd.n488 vdd.n487 242.685
R6617 vdd.n534 vdd.n533 242.685
R6618 vdd.n7126 vdd.n7125 242.685
R6619 vdd.n7172 vdd.n7171 242.685
R6620 vdd.n7269 vdd.n7268 242.685
R6621 vdd.n7315 vdd.n7314 242.685
R6622 vdd.n7361 vdd.n7360 242.685
R6623 vdd.n7407 vdd.n7406 242.685
R6624 vdd.n7504 vdd.n7503 242.685
R6625 vdd.n6653 vdd.n6652 242.685
R6626 vdd.n7548 vdd.n7547 242.685
R6627 vdd.n7593 vdd.n7592 242.685
R6628 vdd.n7643 vdd.n7642 242.685
R6629 vdd.n7689 vdd.n7688 242.685
R6630 vdd.n7737 vdd.n7736 242.685
R6631 vdd.n7455 vdd.n7440 242.685
R6632 vdd.n7784 vdd.n7783 242.685
R6633 vdd.n7829 vdd.n7828 242.685
R6634 vdd.n7875 vdd.n7874 242.685
R6635 vdd.n7926 vdd.n7925 242.685
R6636 vdd.n7972 vdd.n7971 242.685
R6637 vdd.n8020 vdd.n8019 242.685
R6638 vdd.n8066 vdd.n8065 242.685
R6639 vdd.n8111 vdd.n8110 242.685
R6640 vdd.n8161 vdd.n8160 242.685
R6641 vdd.n8207 vdd.n8206 242.685
R6642 vdd.n8255 vdd.n8254 242.685
R6643 vdd.n7220 vdd.n7205 242.685
R6644 vdd.n8302 vdd.n8301 242.685
R6645 vdd.n8347 vdd.n8346 242.685
R6646 vdd.n8397 vdd.n8396 242.685
R6647 vdd.n8443 vdd.n8442 242.685
R6648 vdd.n8491 vdd.n8490 242.685
R6649 vdd.n4112 vdd.n4111 242.685
R6650 vdd.n4158 vdd.n4157 242.685
R6651 vdd.n4255 vdd.n4254 242.685
R6652 vdd.n4301 vdd.n4300 242.685
R6653 vdd.n4347 vdd.n4346 242.685
R6654 vdd.n4393 vdd.n4392 242.685
R6655 vdd.n4490 vdd.n4489 242.685
R6656 vdd.n3639 vdd.n3638 242.685
R6657 vdd.n4534 vdd.n4533 242.685
R6658 vdd.n4579 vdd.n4578 242.685
R6659 vdd.n4629 vdd.n4628 242.685
R6660 vdd.n4675 vdd.n4674 242.685
R6661 vdd.n4723 vdd.n4722 242.685
R6662 vdd.n4441 vdd.n4426 242.685
R6663 vdd.n4770 vdd.n4769 242.685
R6664 vdd.n4815 vdd.n4814 242.685
R6665 vdd.n4861 vdd.n4860 242.685
R6666 vdd.n4912 vdd.n4911 242.685
R6667 vdd.n4958 vdd.n4957 242.685
R6668 vdd.n5006 vdd.n5005 242.685
R6669 vdd.n5052 vdd.n5051 242.685
R6670 vdd.n5097 vdd.n5096 242.685
R6671 vdd.n5147 vdd.n5146 242.685
R6672 vdd.n5193 vdd.n5192 242.685
R6673 vdd.n5241 vdd.n5240 242.685
R6674 vdd.n4206 vdd.n4191 242.685
R6675 vdd.n5288 vdd.n5287 242.685
R6676 vdd.n5333 vdd.n5332 242.685
R6677 vdd.n5383 vdd.n5382 242.685
R6678 vdd.n5429 vdd.n5428 242.685
R6679 vdd.n5477 vdd.n5476 242.685
R6680 vdd.n1098 vdd.n1097 242.685
R6681 vdd.n1144 vdd.n1143 242.685
R6682 vdd.n1241 vdd.n1240 242.685
R6683 vdd.n1287 vdd.n1286 242.685
R6684 vdd.n1333 vdd.n1332 242.685
R6685 vdd.n1379 vdd.n1378 242.685
R6686 vdd.n1476 vdd.n1475 242.685
R6687 vdd.n625 vdd.n624 242.685
R6688 vdd.n1520 vdd.n1519 242.685
R6689 vdd.n1565 vdd.n1564 242.685
R6690 vdd.n1615 vdd.n1614 242.685
R6691 vdd.n1661 vdd.n1660 242.685
R6692 vdd.n1709 vdd.n1708 242.685
R6693 vdd.n1427 vdd.n1412 242.685
R6694 vdd.n1756 vdd.n1755 242.685
R6695 vdd.n1801 vdd.n1800 242.685
R6696 vdd.n1847 vdd.n1846 242.685
R6697 vdd.n1898 vdd.n1897 242.685
R6698 vdd.n1944 vdd.n1943 242.685
R6699 vdd.n1992 vdd.n1991 242.685
R6700 vdd.n2038 vdd.n2037 242.685
R6701 vdd.n2083 vdd.n2082 242.685
R6702 vdd.n2133 vdd.n2132 242.685
R6703 vdd.n2179 vdd.n2178 242.685
R6704 vdd.n2227 vdd.n2226 242.685
R6705 vdd.n1192 vdd.n1177 242.685
R6706 vdd.n2274 vdd.n2273 242.685
R6707 vdd.n2319 vdd.n2318 242.685
R6708 vdd.n2369 vdd.n2368 242.685
R6709 vdd.n2415 vdd.n2414 242.685
R6710 vdd.n2463 vdd.n2462 242.685
R6711 vdd.n10988 vdd.n10987 242.685
R6712 vdd.n11033 vdd.n11032 242.685
R6713 vdd.n11083 vdd.n11082 242.685
R6714 vdd.n11129 vdd.n11128 242.685
R6715 vdd.n11177 vdd.n11176 242.685
R6716 vdd.n439 vdd.n424 242.685
R6717 vdd.n11224 vdd.n11223 242.685
R6718 vdd.n11269 vdd.n11268 242.685
R6719 vdd.n11315 vdd.n11314 242.685
R6720 vdd.n11366 vdd.n11365 242.685
R6721 vdd.n11412 vdd.n11411 242.685
R6722 vdd.n11460 vdd.n11459 242.685
R6723 vdd.n11506 vdd.n11505 242.685
R6724 vdd.n11551 vdd.n11550 242.685
R6725 vdd.n11601 vdd.n11600 242.685
R6726 vdd.n11647 vdd.n11646 242.685
R6727 vdd.n11695 vdd.n11694 242.685
R6728 vdd.n204 vdd.n189 242.685
R6729 vdd.n11742 vdd.n11741 242.685
R6730 vdd.n11787 vdd.n11786 242.685
R6731 vdd.n11837 vdd.n11836 242.685
R6732 vdd.n11883 vdd.n11882 242.685
R6733 vdd.n11931 vdd.n11930 242.685
R6734 vdd.n130 vdd.n100 242.684
R6735 vdd.n176 vdd.n146 242.684
R6736 vdd.n273 vdd.n243 242.684
R6737 vdd.n319 vdd.n289 242.684
R6738 vdd.n365 vdd.n335 242.684
R6739 vdd.n411 vdd.n381 242.684
R6740 vdd.n508 vdd.n478 242.684
R6741 vdd.n554 vdd.n524 242.684
R6742 vdd.n6701 vdd.n6698 242.684
R6743 vdd.n6716 vdd.n6691 242.684
R6744 vdd.n6747 vdd.n6744 242.684
R6745 vdd.n6762 vdd.n6737 242.684
R6746 vdd.n6845 vdd.n6842 242.684
R6747 vdd.n6860 vdd.n6835 242.684
R6748 vdd.n6891 vdd.n6888 242.684
R6749 vdd.n6906 vdd.n6881 242.684
R6750 vdd.n6937 vdd.n6934 242.684
R6751 vdd.n6952 vdd.n6927 242.684
R6752 vdd.n6983 vdd.n6980 242.684
R6753 vdd.n6998 vdd.n6973 242.684
R6754 vdd.n7081 vdd.n7078 242.684
R6755 vdd.n7096 vdd.n7071 242.684
R6756 vdd.n8539 vdd.n8536 242.684
R6757 vdd.n8554 vdd.n8529 242.684
R6758 vdd.n7146 vdd.n7116 242.684
R6759 vdd.n7192 vdd.n7162 242.684
R6760 vdd.n7289 vdd.n7259 242.684
R6761 vdd.n7335 vdd.n7305 242.684
R6762 vdd.n7381 vdd.n7351 242.684
R6763 vdd.n7427 vdd.n7397 242.684
R6764 vdd.n7524 vdd.n7494 242.684
R6765 vdd.n6673 vdd.n6643 242.684
R6766 vdd.n7568 vdd.n7538 242.684
R6767 vdd.n7613 vdd.n7583 242.684
R6768 vdd.n7663 vdd.n7633 242.684
R6769 vdd.n7709 vdd.n7679 242.684
R6770 vdd.n7757 vdd.n7727 242.684
R6771 vdd.n7469 vdd.n7448 242.684
R6772 vdd.n7804 vdd.n7774 242.684
R6773 vdd.n7849 vdd.n7819 242.684
R6774 vdd.n7895 vdd.n7865 242.684
R6775 vdd.n7946 vdd.n7916 242.684
R6776 vdd.n7992 vdd.n7962 242.684
R6777 vdd.n8040 vdd.n8010 242.684
R6778 vdd.n8086 vdd.n8056 242.684
R6779 vdd.n8131 vdd.n8101 242.684
R6780 vdd.n8181 vdd.n8151 242.684
R6781 vdd.n8227 vdd.n8197 242.684
R6782 vdd.n8275 vdd.n8245 242.684
R6783 vdd.n7234 vdd.n7213 242.684
R6784 vdd.n8322 vdd.n8292 242.684
R6785 vdd.n8367 vdd.n8337 242.684
R6786 vdd.n8417 vdd.n8387 242.684
R6787 vdd.n8463 vdd.n8433 242.684
R6788 vdd.n8511 vdd.n8481 242.684
R6789 vdd.n8632 vdd.n8629 242.684
R6790 vdd.n8647 vdd.n8622 242.684
R6791 vdd.n8586 vdd.n8583 242.684
R6792 vdd.n8601 vdd.n8576 242.684
R6793 vdd.n8679 vdd.n8676 242.684
R6794 vdd.n8694 vdd.n8669 242.684
R6795 vdd.n8727 vdd.n8724 242.684
R6796 vdd.n8742 vdd.n8717 242.684
R6797 vdd.n8773 vdd.n8770 242.684
R6798 vdd.n8788 vdd.n8763 242.684
R6799 vdd.n7034 vdd.n7029 242.684
R6800 vdd.n7054 vdd.n7014 242.684
R6801 vdd.n8915 vdd.n8912 242.684
R6802 vdd.n8930 vdd.n8905 242.684
R6803 vdd.n8868 vdd.n8865 242.684
R6804 vdd.n8883 vdd.n8858 242.684
R6805 vdd.n8822 vdd.n8819 242.684
R6806 vdd.n8837 vdd.n8812 242.684
R6807 vdd.n8962 vdd.n8959 242.684
R6808 vdd.n8977 vdd.n8952 242.684
R6809 vdd.n9010 vdd.n9007 242.684
R6810 vdd.n9025 vdd.n9000 242.684
R6811 vdd.n9056 vdd.n9053 242.684
R6812 vdd.n9071 vdd.n9046 242.684
R6813 vdd.n9150 vdd.n9147 242.684
R6814 vdd.n9165 vdd.n9140 242.684
R6815 vdd.n9104 vdd.n9101 242.684
R6816 vdd.n9119 vdd.n9094 242.684
R6817 vdd.n9197 vdd.n9194 242.684
R6818 vdd.n9212 vdd.n9187 242.684
R6819 vdd.n9245 vdd.n9242 242.684
R6820 vdd.n9260 vdd.n9235 242.684
R6821 vdd.n9291 vdd.n9288 242.684
R6822 vdd.n9306 vdd.n9281 242.684
R6823 vdd.n6798 vdd.n6793 242.684
R6824 vdd.n6818 vdd.n6778 242.684
R6825 vdd.n9386 vdd.n9383 242.684
R6826 vdd.n9401 vdd.n9376 242.684
R6827 vdd.n9340 vdd.n9337 242.684
R6828 vdd.n9355 vdd.n9330 242.684
R6829 vdd.n9433 vdd.n9430 242.684
R6830 vdd.n9448 vdd.n9423 242.684
R6831 vdd.n9481 vdd.n9478 242.684
R6832 vdd.n9496 vdd.n9471 242.684
R6833 vdd.n9527 vdd.n9524 242.684
R6834 vdd.n9542 vdd.n9517 242.684
R6835 vdd.n3687 vdd.n3684 242.684
R6836 vdd.n3702 vdd.n3677 242.684
R6837 vdd.n3733 vdd.n3730 242.684
R6838 vdd.n3748 vdd.n3723 242.684
R6839 vdd.n3831 vdd.n3828 242.684
R6840 vdd.n3846 vdd.n3821 242.684
R6841 vdd.n3877 vdd.n3874 242.684
R6842 vdd.n3892 vdd.n3867 242.684
R6843 vdd.n3923 vdd.n3920 242.684
R6844 vdd.n3938 vdd.n3913 242.684
R6845 vdd.n3969 vdd.n3966 242.684
R6846 vdd.n3984 vdd.n3959 242.684
R6847 vdd.n4067 vdd.n4064 242.684
R6848 vdd.n4082 vdd.n4057 242.684
R6849 vdd.n5525 vdd.n5522 242.684
R6850 vdd.n5540 vdd.n5515 242.684
R6851 vdd.n4132 vdd.n4102 242.684
R6852 vdd.n4178 vdd.n4148 242.684
R6853 vdd.n4275 vdd.n4245 242.684
R6854 vdd.n4321 vdd.n4291 242.684
R6855 vdd.n4367 vdd.n4337 242.684
R6856 vdd.n4413 vdd.n4383 242.684
R6857 vdd.n4510 vdd.n4480 242.684
R6858 vdd.n3659 vdd.n3629 242.684
R6859 vdd.n4554 vdd.n4524 242.684
R6860 vdd.n4599 vdd.n4569 242.684
R6861 vdd.n4649 vdd.n4619 242.684
R6862 vdd.n4695 vdd.n4665 242.684
R6863 vdd.n4743 vdd.n4713 242.684
R6864 vdd.n4455 vdd.n4434 242.684
R6865 vdd.n4790 vdd.n4760 242.684
R6866 vdd.n4835 vdd.n4805 242.684
R6867 vdd.n4881 vdd.n4851 242.684
R6868 vdd.n4932 vdd.n4902 242.684
R6869 vdd.n4978 vdd.n4948 242.684
R6870 vdd.n5026 vdd.n4996 242.684
R6871 vdd.n5072 vdd.n5042 242.684
R6872 vdd.n5117 vdd.n5087 242.684
R6873 vdd.n5167 vdd.n5137 242.684
R6874 vdd.n5213 vdd.n5183 242.684
R6875 vdd.n5261 vdd.n5231 242.684
R6876 vdd.n4220 vdd.n4199 242.684
R6877 vdd.n5308 vdd.n5278 242.684
R6878 vdd.n5353 vdd.n5323 242.684
R6879 vdd.n5403 vdd.n5373 242.684
R6880 vdd.n5449 vdd.n5419 242.684
R6881 vdd.n5497 vdd.n5467 242.684
R6882 vdd.n5618 vdd.n5615 242.684
R6883 vdd.n5633 vdd.n5608 242.684
R6884 vdd.n5572 vdd.n5569 242.684
R6885 vdd.n5587 vdd.n5562 242.684
R6886 vdd.n5665 vdd.n5662 242.684
R6887 vdd.n5680 vdd.n5655 242.684
R6888 vdd.n5713 vdd.n5710 242.684
R6889 vdd.n5728 vdd.n5703 242.684
R6890 vdd.n5759 vdd.n5756 242.684
R6891 vdd.n5774 vdd.n5749 242.684
R6892 vdd.n4020 vdd.n4015 242.684
R6893 vdd.n4040 vdd.n4000 242.684
R6894 vdd.n5901 vdd.n5898 242.684
R6895 vdd.n5916 vdd.n5891 242.684
R6896 vdd.n5854 vdd.n5851 242.684
R6897 vdd.n5869 vdd.n5844 242.684
R6898 vdd.n5808 vdd.n5805 242.684
R6899 vdd.n5823 vdd.n5798 242.684
R6900 vdd.n5948 vdd.n5945 242.684
R6901 vdd.n5963 vdd.n5938 242.684
R6902 vdd.n5996 vdd.n5993 242.684
R6903 vdd.n6011 vdd.n5986 242.684
R6904 vdd.n6042 vdd.n6039 242.684
R6905 vdd.n6057 vdd.n6032 242.684
R6906 vdd.n6136 vdd.n6133 242.684
R6907 vdd.n6151 vdd.n6126 242.684
R6908 vdd.n6090 vdd.n6087 242.684
R6909 vdd.n6105 vdd.n6080 242.684
R6910 vdd.n6183 vdd.n6180 242.684
R6911 vdd.n6198 vdd.n6173 242.684
R6912 vdd.n6231 vdd.n6228 242.684
R6913 vdd.n6246 vdd.n6221 242.684
R6914 vdd.n6277 vdd.n6274 242.684
R6915 vdd.n6292 vdd.n6267 242.684
R6916 vdd.n3784 vdd.n3779 242.684
R6917 vdd.n3804 vdd.n3764 242.684
R6918 vdd.n6372 vdd.n6369 242.684
R6919 vdd.n6387 vdd.n6362 242.684
R6920 vdd.n6326 vdd.n6323 242.684
R6921 vdd.n6341 vdd.n6316 242.684
R6922 vdd.n6419 vdd.n6416 242.684
R6923 vdd.n6434 vdd.n6409 242.684
R6924 vdd.n6467 vdd.n6464 242.684
R6925 vdd.n6482 vdd.n6457 242.684
R6926 vdd.n6513 vdd.n6510 242.684
R6927 vdd.n6528 vdd.n6503 242.684
R6928 vdd.n673 vdd.n670 242.684
R6929 vdd.n688 vdd.n663 242.684
R6930 vdd.n719 vdd.n716 242.684
R6931 vdd.n734 vdd.n709 242.684
R6932 vdd.n817 vdd.n814 242.684
R6933 vdd.n832 vdd.n807 242.684
R6934 vdd.n863 vdd.n860 242.684
R6935 vdd.n878 vdd.n853 242.684
R6936 vdd.n909 vdd.n906 242.684
R6937 vdd.n924 vdd.n899 242.684
R6938 vdd.n955 vdd.n952 242.684
R6939 vdd.n970 vdd.n945 242.684
R6940 vdd.n1053 vdd.n1050 242.684
R6941 vdd.n1068 vdd.n1043 242.684
R6942 vdd.n2511 vdd.n2508 242.684
R6943 vdd.n2526 vdd.n2501 242.684
R6944 vdd.n1118 vdd.n1088 242.684
R6945 vdd.n1164 vdd.n1134 242.684
R6946 vdd.n1261 vdd.n1231 242.684
R6947 vdd.n1307 vdd.n1277 242.684
R6948 vdd.n1353 vdd.n1323 242.684
R6949 vdd.n1399 vdd.n1369 242.684
R6950 vdd.n1496 vdd.n1466 242.684
R6951 vdd.n645 vdd.n615 242.684
R6952 vdd.n1540 vdd.n1510 242.684
R6953 vdd.n1585 vdd.n1555 242.684
R6954 vdd.n1635 vdd.n1605 242.684
R6955 vdd.n1681 vdd.n1651 242.684
R6956 vdd.n1729 vdd.n1699 242.684
R6957 vdd.n1441 vdd.n1420 242.684
R6958 vdd.n1776 vdd.n1746 242.684
R6959 vdd.n1821 vdd.n1791 242.684
R6960 vdd.n1867 vdd.n1837 242.684
R6961 vdd.n1918 vdd.n1888 242.684
R6962 vdd.n1964 vdd.n1934 242.684
R6963 vdd.n2012 vdd.n1982 242.684
R6964 vdd.n2058 vdd.n2028 242.684
R6965 vdd.n2103 vdd.n2073 242.684
R6966 vdd.n2153 vdd.n2123 242.684
R6967 vdd.n2199 vdd.n2169 242.684
R6968 vdd.n2247 vdd.n2217 242.684
R6969 vdd.n1206 vdd.n1185 242.684
R6970 vdd.n2294 vdd.n2264 242.684
R6971 vdd.n2339 vdd.n2309 242.684
R6972 vdd.n2389 vdd.n2359 242.684
R6973 vdd.n2435 vdd.n2405 242.684
R6974 vdd.n2483 vdd.n2453 242.684
R6975 vdd.n2604 vdd.n2601 242.684
R6976 vdd.n2619 vdd.n2594 242.684
R6977 vdd.n2558 vdd.n2555 242.684
R6978 vdd.n2573 vdd.n2548 242.684
R6979 vdd.n2651 vdd.n2648 242.684
R6980 vdd.n2666 vdd.n2641 242.684
R6981 vdd.n2699 vdd.n2696 242.684
R6982 vdd.n2714 vdd.n2689 242.684
R6983 vdd.n2745 vdd.n2742 242.684
R6984 vdd.n2760 vdd.n2735 242.684
R6985 vdd.n1006 vdd.n1001 242.684
R6986 vdd.n1026 vdd.n986 242.684
R6987 vdd.n2887 vdd.n2884 242.684
R6988 vdd.n2902 vdd.n2877 242.684
R6989 vdd.n2840 vdd.n2837 242.684
R6990 vdd.n2855 vdd.n2830 242.684
R6991 vdd.n2794 vdd.n2791 242.684
R6992 vdd.n2809 vdd.n2784 242.684
R6993 vdd.n2934 vdd.n2931 242.684
R6994 vdd.n2949 vdd.n2924 242.684
R6995 vdd.n2982 vdd.n2979 242.684
R6996 vdd.n2997 vdd.n2972 242.684
R6997 vdd.n3028 vdd.n3025 242.684
R6998 vdd.n3043 vdd.n3018 242.684
R6999 vdd.n3122 vdd.n3119 242.684
R7000 vdd.n3137 vdd.n3112 242.684
R7001 vdd.n3076 vdd.n3073 242.684
R7002 vdd.n3091 vdd.n3066 242.684
R7003 vdd.n3169 vdd.n3166 242.684
R7004 vdd.n3184 vdd.n3159 242.684
R7005 vdd.n3217 vdd.n3214 242.684
R7006 vdd.n3232 vdd.n3207 242.684
R7007 vdd.n3263 vdd.n3260 242.684
R7008 vdd.n3278 vdd.n3253 242.684
R7009 vdd.n770 vdd.n765 242.684
R7010 vdd.n790 vdd.n750 242.684
R7011 vdd.n3358 vdd.n3355 242.684
R7012 vdd.n3373 vdd.n3348 242.684
R7013 vdd.n3312 vdd.n3309 242.684
R7014 vdd.n3327 vdd.n3302 242.684
R7015 vdd.n3405 vdd.n3402 242.684
R7016 vdd.n3420 vdd.n3395 242.684
R7017 vdd.n3453 vdd.n3450 242.684
R7018 vdd.n3468 vdd.n3443 242.684
R7019 vdd.n3499 vdd.n3496 242.684
R7020 vdd.n3514 vdd.n3489 242.684
R7021 vdd.n581 vdd.n578 242.684
R7022 vdd.n596 vdd.n571 242.684
R7023 vdd.n3594 vdd.n3591 242.684
R7024 vdd.n3609 vdd.n3584 242.684
R7025 vdd.n3548 vdd.n3545 242.684
R7026 vdd.n3563 vdd.n3538 242.684
R7027 vdd.n6608 vdd.n6605 242.684
R7028 vdd.n6623 vdd.n6598 242.684
R7029 vdd.n6562 vdd.n6559 242.684
R7030 vdd.n6577 vdd.n6552 242.684
R7031 vdd.n9622 vdd.n9619 242.684
R7032 vdd.n9637 vdd.n9612 242.684
R7033 vdd.n9576 vdd.n9573 242.684
R7034 vdd.n9591 vdd.n9566 242.684
R7035 vdd.n9668 vdd.n9665 242.684
R7036 vdd.n9683 vdd.n9658 242.684
R7037 vdd.n9714 vdd.n9711 242.684
R7038 vdd.n9729 vdd.n9704 242.684
R7039 vdd.n9812 vdd.n9809 242.684
R7040 vdd.n9827 vdd.n9802 242.684
R7041 vdd.n9858 vdd.n9855 242.684
R7042 vdd.n9873 vdd.n9848 242.684
R7043 vdd.n9904 vdd.n9901 242.684
R7044 vdd.n9919 vdd.n9894 242.684
R7045 vdd.n9950 vdd.n9947 242.684
R7046 vdd.n9965 vdd.n9940 242.684
R7047 vdd.n10048 vdd.n10045 242.684
R7048 vdd.n10063 vdd.n10038 242.684
R7049 vdd.n64 vdd.n61 242.684
R7050 vdd.n79 vdd.n54 242.684
R7051 vdd.n18 vdd.n15 242.684
R7052 vdd.n33 vdd.n8 242.684
R7053 vdd.n10094 vdd.n10091 242.684
R7054 vdd.n10109 vdd.n10084 242.684
R7055 vdd.n10142 vdd.n10139 242.684
R7056 vdd.n10157 vdd.n10132 242.684
R7057 vdd.n10188 vdd.n10185 242.684
R7058 vdd.n10203 vdd.n10178 242.684
R7059 vdd.n10001 vdd.n9996 242.684
R7060 vdd.n10021 vdd.n9981 242.684
R7061 vdd.n10330 vdd.n10327 242.684
R7062 vdd.n10345 vdd.n10320 242.684
R7063 vdd.n10283 vdd.n10280 242.684
R7064 vdd.n10298 vdd.n10273 242.684
R7065 vdd.n10237 vdd.n10234 242.684
R7066 vdd.n10252 vdd.n10227 242.684
R7067 vdd.n10377 vdd.n10374 242.684
R7068 vdd.n10392 vdd.n10367 242.684
R7069 vdd.n10425 vdd.n10422 242.684
R7070 vdd.n10440 vdd.n10415 242.684
R7071 vdd.n10471 vdd.n10468 242.684
R7072 vdd.n10486 vdd.n10461 242.684
R7073 vdd.n10565 vdd.n10562 242.684
R7074 vdd.n10580 vdd.n10555 242.684
R7075 vdd.n10519 vdd.n10516 242.684
R7076 vdd.n10534 vdd.n10509 242.684
R7077 vdd.n10612 vdd.n10609 242.684
R7078 vdd.n10627 vdd.n10602 242.684
R7079 vdd.n10660 vdd.n10657 242.684
R7080 vdd.n10675 vdd.n10650 242.684
R7081 vdd.n10706 vdd.n10703 242.684
R7082 vdd.n10721 vdd.n10696 242.684
R7083 vdd.n9765 vdd.n9760 242.684
R7084 vdd.n9785 vdd.n9745 242.684
R7085 vdd.n10801 vdd.n10798 242.684
R7086 vdd.n10816 vdd.n10791 242.684
R7087 vdd.n10755 vdd.n10752 242.684
R7088 vdd.n10770 vdd.n10745 242.684
R7089 vdd.n10848 vdd.n10845 242.684
R7090 vdd.n10863 vdd.n10838 242.684
R7091 vdd.n10896 vdd.n10893 242.684
R7092 vdd.n10911 vdd.n10886 242.684
R7093 vdd.n10942 vdd.n10939 242.684
R7094 vdd.n10957 vdd.n10932 242.684
R7095 vdd.n11008 vdd.n10978 242.684
R7096 vdd.n11053 vdd.n11023 242.684
R7097 vdd.n11103 vdd.n11073 242.684
R7098 vdd.n11149 vdd.n11119 242.684
R7099 vdd.n11197 vdd.n11167 242.684
R7100 vdd.n453 vdd.n432 242.684
R7101 vdd.n11244 vdd.n11214 242.684
R7102 vdd.n11289 vdd.n11259 242.684
R7103 vdd.n11335 vdd.n11305 242.684
R7104 vdd.n11386 vdd.n11356 242.684
R7105 vdd.n11432 vdd.n11402 242.684
R7106 vdd.n11480 vdd.n11450 242.684
R7107 vdd.n11526 vdd.n11496 242.684
R7108 vdd.n11571 vdd.n11541 242.684
R7109 vdd.n11621 vdd.n11591 242.684
R7110 vdd.n11667 vdd.n11637 242.684
R7111 vdd.n11715 vdd.n11685 242.684
R7112 vdd.n218 vdd.n197 242.684
R7113 vdd.n11762 vdd.n11732 242.684
R7114 vdd.n11807 vdd.n11777 242.684
R7115 vdd.n11857 vdd.n11827 242.684
R7116 vdd.n11903 vdd.n11873 242.684
R7117 vdd.n11951 vdd.n11921 242.684
R7118 vdd.n11994 vdd.n11986 93.7417
R7119 vdd.n12004 vdd.n11964 93.7417
R7120 vdd.n11975 vdd.n11967 93.7417
R7121 vdd.n124 vdd.n123 93.7417
R7122 vdd.n123 vdd.n97 93.7417
R7123 vdd.n122 vdd.n95 93.7417
R7124 vdd.n137 vdd.n95 93.7417
R7125 vdd.n114 vdd.n103 93.7417
R7126 vdd.n115 vdd.n114 93.7417
R7127 vdd.n170 vdd.n169 93.7417
R7128 vdd.n169 vdd.n143 93.7417
R7129 vdd.n168 vdd.n141 93.7417
R7130 vdd.n183 vdd.n141 93.7417
R7131 vdd.n160 vdd.n149 93.7417
R7132 vdd.n161 vdd.n160 93.7417
R7133 vdd.n267 vdd.n266 93.7417
R7134 vdd.n266 vdd.n240 93.7417
R7135 vdd.n265 vdd.n238 93.7417
R7136 vdd.n280 vdd.n238 93.7417
R7137 vdd.n257 vdd.n246 93.7417
R7138 vdd.n258 vdd.n257 93.7417
R7139 vdd.n313 vdd.n312 93.7417
R7140 vdd.n312 vdd.n286 93.7417
R7141 vdd.n311 vdd.n284 93.7417
R7142 vdd.n326 vdd.n284 93.7417
R7143 vdd.n303 vdd.n292 93.7417
R7144 vdd.n304 vdd.n303 93.7417
R7145 vdd.n359 vdd.n358 93.7417
R7146 vdd.n358 vdd.n332 93.7417
R7147 vdd.n357 vdd.n330 93.7417
R7148 vdd.n372 vdd.n330 93.7417
R7149 vdd.n349 vdd.n338 93.7417
R7150 vdd.n350 vdd.n349 93.7417
R7151 vdd.n405 vdd.n404 93.7417
R7152 vdd.n404 vdd.n378 93.7417
R7153 vdd.n403 vdd.n376 93.7417
R7154 vdd.n418 vdd.n376 93.7417
R7155 vdd.n395 vdd.n384 93.7417
R7156 vdd.n396 vdd.n395 93.7417
R7157 vdd.n502 vdd.n501 93.7417
R7158 vdd.n501 vdd.n475 93.7417
R7159 vdd.n500 vdd.n473 93.7417
R7160 vdd.n515 vdd.n473 93.7417
R7161 vdd.n492 vdd.n481 93.7417
R7162 vdd.n493 vdd.n492 93.7417
R7163 vdd.n548 vdd.n547 93.7417
R7164 vdd.n547 vdd.n521 93.7417
R7165 vdd.n546 vdd.n519 93.7417
R7166 vdd.n561 vdd.n519 93.7417
R7167 vdd.n538 vdd.n527 93.7417
R7168 vdd.n539 vdd.n538 93.7417
R7169 vdd.n6690 vdd.n6685 93.7417
R7170 vdd.n6713 vdd.n6690 93.7417
R7171 vdd.n6725 vdd.n6683 93.7417
R7172 vdd.n6711 vdd.n6683 93.7417
R7173 vdd.n6704 vdd.n6703 93.7417
R7174 vdd.n6703 vdd.n6692 93.7417
R7175 vdd.n6736 vdd.n6731 93.7417
R7176 vdd.n6759 vdd.n6736 93.7417
R7177 vdd.n6771 vdd.n6729 93.7417
R7178 vdd.n6757 vdd.n6729 93.7417
R7179 vdd.n6750 vdd.n6749 93.7417
R7180 vdd.n6749 vdd.n6738 93.7417
R7181 vdd.n6834 vdd.n6829 93.7417
R7182 vdd.n6857 vdd.n6834 93.7417
R7183 vdd.n6869 vdd.n6827 93.7417
R7184 vdd.n6855 vdd.n6827 93.7417
R7185 vdd.n6848 vdd.n6847 93.7417
R7186 vdd.n6847 vdd.n6836 93.7417
R7187 vdd.n6880 vdd.n6875 93.7417
R7188 vdd.n6903 vdd.n6880 93.7417
R7189 vdd.n6915 vdd.n6873 93.7417
R7190 vdd.n6901 vdd.n6873 93.7417
R7191 vdd.n6894 vdd.n6893 93.7417
R7192 vdd.n6893 vdd.n6882 93.7417
R7193 vdd.n6926 vdd.n6921 93.7417
R7194 vdd.n6949 vdd.n6926 93.7417
R7195 vdd.n6961 vdd.n6919 93.7417
R7196 vdd.n6947 vdd.n6919 93.7417
R7197 vdd.n6940 vdd.n6939 93.7417
R7198 vdd.n6939 vdd.n6928 93.7417
R7199 vdd.n6972 vdd.n6967 93.7417
R7200 vdd.n6995 vdd.n6972 93.7417
R7201 vdd.n7007 vdd.n6965 93.7417
R7202 vdd.n6993 vdd.n6965 93.7417
R7203 vdd.n6986 vdd.n6985 93.7417
R7204 vdd.n6985 vdd.n6974 93.7417
R7205 vdd.n7070 vdd.n7065 93.7417
R7206 vdd.n7093 vdd.n7070 93.7417
R7207 vdd.n7105 vdd.n7063 93.7417
R7208 vdd.n7091 vdd.n7063 93.7417
R7209 vdd.n7084 vdd.n7083 93.7417
R7210 vdd.n7083 vdd.n7072 93.7417
R7211 vdd.n8528 vdd.n8523 93.7417
R7212 vdd.n8551 vdd.n8528 93.7417
R7213 vdd.n8563 vdd.n8521 93.7417
R7214 vdd.n8549 vdd.n8521 93.7417
R7215 vdd.n8542 vdd.n8541 93.7417
R7216 vdd.n8541 vdd.n8530 93.7417
R7217 vdd.n7140 vdd.n7139 93.7417
R7218 vdd.n7139 vdd.n7113 93.7417
R7219 vdd.n7138 vdd.n7111 93.7417
R7220 vdd.n7153 vdd.n7111 93.7417
R7221 vdd.n7130 vdd.n7119 93.7417
R7222 vdd.n7131 vdd.n7130 93.7417
R7223 vdd.n7186 vdd.n7185 93.7417
R7224 vdd.n7185 vdd.n7159 93.7417
R7225 vdd.n7184 vdd.n7157 93.7417
R7226 vdd.n7199 vdd.n7157 93.7417
R7227 vdd.n7176 vdd.n7165 93.7417
R7228 vdd.n7177 vdd.n7176 93.7417
R7229 vdd.n7283 vdd.n7282 93.7417
R7230 vdd.n7282 vdd.n7256 93.7417
R7231 vdd.n7281 vdd.n7254 93.7417
R7232 vdd.n7296 vdd.n7254 93.7417
R7233 vdd.n7273 vdd.n7262 93.7417
R7234 vdd.n7274 vdd.n7273 93.7417
R7235 vdd.n7329 vdd.n7328 93.7417
R7236 vdd.n7328 vdd.n7302 93.7417
R7237 vdd.n7327 vdd.n7300 93.7417
R7238 vdd.n7342 vdd.n7300 93.7417
R7239 vdd.n7319 vdd.n7308 93.7417
R7240 vdd.n7320 vdd.n7319 93.7417
R7241 vdd.n7375 vdd.n7374 93.7417
R7242 vdd.n7374 vdd.n7348 93.7417
R7243 vdd.n7373 vdd.n7346 93.7417
R7244 vdd.n7388 vdd.n7346 93.7417
R7245 vdd.n7365 vdd.n7354 93.7417
R7246 vdd.n7366 vdd.n7365 93.7417
R7247 vdd.n7421 vdd.n7420 93.7417
R7248 vdd.n7420 vdd.n7394 93.7417
R7249 vdd.n7419 vdd.n7392 93.7417
R7250 vdd.n7434 vdd.n7392 93.7417
R7251 vdd.n7411 vdd.n7400 93.7417
R7252 vdd.n7412 vdd.n7411 93.7417
R7253 vdd.n7518 vdd.n7517 93.7417
R7254 vdd.n7517 vdd.n7491 93.7417
R7255 vdd.n7516 vdd.n7489 93.7417
R7256 vdd.n7531 vdd.n7489 93.7417
R7257 vdd.n7508 vdd.n7497 93.7417
R7258 vdd.n7509 vdd.n7508 93.7417
R7259 vdd.n6667 vdd.n6666 93.7417
R7260 vdd.n6666 vdd.n6640 93.7417
R7261 vdd.n6665 vdd.n6638 93.7417
R7262 vdd.n6680 vdd.n6638 93.7417
R7263 vdd.n6657 vdd.n6646 93.7417
R7264 vdd.n6658 vdd.n6657 93.7417
R7265 vdd.n7562 vdd.n7561 93.7417
R7266 vdd.n7561 vdd.n7535 93.7417
R7267 vdd.n7560 vdd.n7533 93.7417
R7268 vdd.n7575 vdd.n7533 93.7417
R7269 vdd.n7552 vdd.n7541 93.7417
R7270 vdd.n7553 vdd.n7552 93.7417
R7271 vdd.n7607 vdd.n7606 93.7417
R7272 vdd.n7606 vdd.n7580 93.7417
R7273 vdd.n7605 vdd.n7578 93.7417
R7274 vdd.n7620 vdd.n7578 93.7417
R7275 vdd.n7597 vdd.n7586 93.7417
R7276 vdd.n7598 vdd.n7597 93.7417
R7277 vdd.n7657 vdd.n7656 93.7417
R7278 vdd.n7656 vdd.n7630 93.7417
R7279 vdd.n7655 vdd.n7628 93.7417
R7280 vdd.n7670 vdd.n7628 93.7417
R7281 vdd.n7647 vdd.n7636 93.7417
R7282 vdd.n7648 vdd.n7647 93.7417
R7283 vdd.n7703 vdd.n7702 93.7417
R7284 vdd.n7702 vdd.n7676 93.7417
R7285 vdd.n7701 vdd.n7674 93.7417
R7286 vdd.n7716 vdd.n7674 93.7417
R7287 vdd.n7693 vdd.n7682 93.7417
R7288 vdd.n7694 vdd.n7693 93.7417
R7289 vdd.n7751 vdd.n7750 93.7417
R7290 vdd.n7750 vdd.n7724 93.7417
R7291 vdd.n7749 vdd.n7722 93.7417
R7292 vdd.n7764 vdd.n7722 93.7417
R7293 vdd.n7741 vdd.n7730 93.7417
R7294 vdd.n7742 vdd.n7741 93.7417
R7295 vdd.n7463 vdd.n7462 93.7417
R7296 vdd.n7462 vdd.n7446 93.7417
R7297 vdd.n7461 vdd.n7444 93.7417
R7298 vdd.n7477 vdd.n7444 93.7417
R7299 vdd.n7454 vdd.n7453 93.7417
R7300 vdd.n7453 vdd.n7439 93.7417
R7301 vdd.n7798 vdd.n7797 93.7417
R7302 vdd.n7797 vdd.n7771 93.7417
R7303 vdd.n7796 vdd.n7769 93.7417
R7304 vdd.n7811 vdd.n7769 93.7417
R7305 vdd.n7788 vdd.n7777 93.7417
R7306 vdd.n7789 vdd.n7788 93.7417
R7307 vdd.n7843 vdd.n7842 93.7417
R7308 vdd.n7842 vdd.n7816 93.7417
R7309 vdd.n7841 vdd.n7814 93.7417
R7310 vdd.n7856 vdd.n7814 93.7417
R7311 vdd.n7833 vdd.n7822 93.7417
R7312 vdd.n7834 vdd.n7833 93.7417
R7313 vdd.n7889 vdd.n7888 93.7417
R7314 vdd.n7888 vdd.n7862 93.7417
R7315 vdd.n7887 vdd.n7860 93.7417
R7316 vdd.n7902 vdd.n7860 93.7417
R7317 vdd.n7879 vdd.n7868 93.7417
R7318 vdd.n7880 vdd.n7879 93.7417
R7319 vdd.n7940 vdd.n7939 93.7417
R7320 vdd.n7939 vdd.n7913 93.7417
R7321 vdd.n7938 vdd.n7911 93.7417
R7322 vdd.n7953 vdd.n7911 93.7417
R7323 vdd.n7930 vdd.n7919 93.7417
R7324 vdd.n7931 vdd.n7930 93.7417
R7325 vdd.n7986 vdd.n7985 93.7417
R7326 vdd.n7985 vdd.n7959 93.7417
R7327 vdd.n7984 vdd.n7957 93.7417
R7328 vdd.n7999 vdd.n7957 93.7417
R7329 vdd.n7976 vdd.n7965 93.7417
R7330 vdd.n7977 vdd.n7976 93.7417
R7331 vdd.n8034 vdd.n8033 93.7417
R7332 vdd.n8033 vdd.n8007 93.7417
R7333 vdd.n8032 vdd.n8005 93.7417
R7334 vdd.n8047 vdd.n8005 93.7417
R7335 vdd.n8024 vdd.n8013 93.7417
R7336 vdd.n8025 vdd.n8024 93.7417
R7337 vdd.n8080 vdd.n8079 93.7417
R7338 vdd.n8079 vdd.n8053 93.7417
R7339 vdd.n8078 vdd.n8051 93.7417
R7340 vdd.n8093 vdd.n8051 93.7417
R7341 vdd.n8070 vdd.n8059 93.7417
R7342 vdd.n8071 vdd.n8070 93.7417
R7343 vdd.n8125 vdd.n8124 93.7417
R7344 vdd.n8124 vdd.n8098 93.7417
R7345 vdd.n8123 vdd.n8096 93.7417
R7346 vdd.n8138 vdd.n8096 93.7417
R7347 vdd.n8115 vdd.n8104 93.7417
R7348 vdd.n8116 vdd.n8115 93.7417
R7349 vdd.n8175 vdd.n8174 93.7417
R7350 vdd.n8174 vdd.n8148 93.7417
R7351 vdd.n8173 vdd.n8146 93.7417
R7352 vdd.n8188 vdd.n8146 93.7417
R7353 vdd.n8165 vdd.n8154 93.7417
R7354 vdd.n8166 vdd.n8165 93.7417
R7355 vdd.n8221 vdd.n8220 93.7417
R7356 vdd.n8220 vdd.n8194 93.7417
R7357 vdd.n8219 vdd.n8192 93.7417
R7358 vdd.n8234 vdd.n8192 93.7417
R7359 vdd.n8211 vdd.n8200 93.7417
R7360 vdd.n8212 vdd.n8211 93.7417
R7361 vdd.n8269 vdd.n8268 93.7417
R7362 vdd.n8268 vdd.n8242 93.7417
R7363 vdd.n8267 vdd.n8240 93.7417
R7364 vdd.n8282 vdd.n8240 93.7417
R7365 vdd.n8259 vdd.n8248 93.7417
R7366 vdd.n8260 vdd.n8259 93.7417
R7367 vdd.n7228 vdd.n7227 93.7417
R7368 vdd.n7227 vdd.n7211 93.7417
R7369 vdd.n7226 vdd.n7209 93.7417
R7370 vdd.n7242 vdd.n7209 93.7417
R7371 vdd.n7219 vdd.n7218 93.7417
R7372 vdd.n7218 vdd.n7204 93.7417
R7373 vdd.n8316 vdd.n8315 93.7417
R7374 vdd.n8315 vdd.n8289 93.7417
R7375 vdd.n8314 vdd.n8287 93.7417
R7376 vdd.n8329 vdd.n8287 93.7417
R7377 vdd.n8306 vdd.n8295 93.7417
R7378 vdd.n8307 vdd.n8306 93.7417
R7379 vdd.n8361 vdd.n8360 93.7417
R7380 vdd.n8360 vdd.n8334 93.7417
R7381 vdd.n8359 vdd.n8332 93.7417
R7382 vdd.n8374 vdd.n8332 93.7417
R7383 vdd.n8351 vdd.n8340 93.7417
R7384 vdd.n8352 vdd.n8351 93.7417
R7385 vdd.n8411 vdd.n8410 93.7417
R7386 vdd.n8410 vdd.n8384 93.7417
R7387 vdd.n8409 vdd.n8382 93.7417
R7388 vdd.n8424 vdd.n8382 93.7417
R7389 vdd.n8401 vdd.n8390 93.7417
R7390 vdd.n8402 vdd.n8401 93.7417
R7391 vdd.n8457 vdd.n8456 93.7417
R7392 vdd.n8456 vdd.n8430 93.7417
R7393 vdd.n8455 vdd.n8428 93.7417
R7394 vdd.n8470 vdd.n8428 93.7417
R7395 vdd.n8447 vdd.n8436 93.7417
R7396 vdd.n8448 vdd.n8447 93.7417
R7397 vdd.n8505 vdd.n8504 93.7417
R7398 vdd.n8504 vdd.n8478 93.7417
R7399 vdd.n8503 vdd.n8476 93.7417
R7400 vdd.n8518 vdd.n8476 93.7417
R7401 vdd.n8495 vdd.n8484 93.7417
R7402 vdd.n8496 vdd.n8495 93.7417
R7403 vdd.n8621 vdd.n8616 93.7417
R7404 vdd.n8644 vdd.n8621 93.7417
R7405 vdd.n8656 vdd.n8614 93.7417
R7406 vdd.n8642 vdd.n8614 93.7417
R7407 vdd.n8635 vdd.n8634 93.7417
R7408 vdd.n8634 vdd.n8623 93.7417
R7409 vdd.n8575 vdd.n8570 93.7417
R7410 vdd.n8598 vdd.n8575 93.7417
R7411 vdd.n8610 vdd.n8568 93.7417
R7412 vdd.n8596 vdd.n8568 93.7417
R7413 vdd.n8589 vdd.n8588 93.7417
R7414 vdd.n8588 vdd.n8577 93.7417
R7415 vdd.n8668 vdd.n8663 93.7417
R7416 vdd.n8691 vdd.n8668 93.7417
R7417 vdd.n8703 vdd.n8661 93.7417
R7418 vdd.n8689 vdd.n8661 93.7417
R7419 vdd.n8682 vdd.n8681 93.7417
R7420 vdd.n8681 vdd.n8670 93.7417
R7421 vdd.n8716 vdd.n8711 93.7417
R7422 vdd.n8739 vdd.n8716 93.7417
R7423 vdd.n8751 vdd.n8709 93.7417
R7424 vdd.n8737 vdd.n8709 93.7417
R7425 vdd.n8730 vdd.n8729 93.7417
R7426 vdd.n8729 vdd.n8718 93.7417
R7427 vdd.n8762 vdd.n8757 93.7417
R7428 vdd.n8785 vdd.n8762 93.7417
R7429 vdd.n8797 vdd.n8755 93.7417
R7430 vdd.n8783 vdd.n8755 93.7417
R7431 vdd.n8776 vdd.n8775 93.7417
R7432 vdd.n8775 vdd.n8764 93.7417
R7433 vdd.n7050 vdd.n7049 93.7417
R7434 vdd.n7050 vdd.n7015 93.7417
R7435 vdd.n7047 vdd.n7019 93.7417
R7436 vdd.n7039 vdd.n7019 93.7417
R7437 vdd.n7027 vdd.n7020 93.7417
R7438 vdd.n7037 vdd.n7027 93.7417
R7439 vdd.n8904 vdd.n8899 93.7417
R7440 vdd.n8927 vdd.n8904 93.7417
R7441 vdd.n8939 vdd.n8897 93.7417
R7442 vdd.n8925 vdd.n8897 93.7417
R7443 vdd.n8918 vdd.n8917 93.7417
R7444 vdd.n8917 vdd.n8906 93.7417
R7445 vdd.n8857 vdd.n8852 93.7417
R7446 vdd.n8880 vdd.n8857 93.7417
R7447 vdd.n8892 vdd.n8850 93.7417
R7448 vdd.n8878 vdd.n8850 93.7417
R7449 vdd.n8871 vdd.n8870 93.7417
R7450 vdd.n8870 vdd.n8859 93.7417
R7451 vdd.n8811 vdd.n8806 93.7417
R7452 vdd.n8834 vdd.n8811 93.7417
R7453 vdd.n8846 vdd.n8804 93.7417
R7454 vdd.n8832 vdd.n8804 93.7417
R7455 vdd.n8825 vdd.n8824 93.7417
R7456 vdd.n8824 vdd.n8813 93.7417
R7457 vdd.n8951 vdd.n8946 93.7417
R7458 vdd.n8974 vdd.n8951 93.7417
R7459 vdd.n8986 vdd.n8944 93.7417
R7460 vdd.n8972 vdd.n8944 93.7417
R7461 vdd.n8965 vdd.n8964 93.7417
R7462 vdd.n8964 vdd.n8953 93.7417
R7463 vdd.n8999 vdd.n8994 93.7417
R7464 vdd.n9022 vdd.n8999 93.7417
R7465 vdd.n9034 vdd.n8992 93.7417
R7466 vdd.n9020 vdd.n8992 93.7417
R7467 vdd.n9013 vdd.n9012 93.7417
R7468 vdd.n9012 vdd.n9001 93.7417
R7469 vdd.n9045 vdd.n9040 93.7417
R7470 vdd.n9068 vdd.n9045 93.7417
R7471 vdd.n9080 vdd.n9038 93.7417
R7472 vdd.n9066 vdd.n9038 93.7417
R7473 vdd.n9059 vdd.n9058 93.7417
R7474 vdd.n9058 vdd.n9047 93.7417
R7475 vdd.n9139 vdd.n9134 93.7417
R7476 vdd.n9162 vdd.n9139 93.7417
R7477 vdd.n9174 vdd.n9132 93.7417
R7478 vdd.n9160 vdd.n9132 93.7417
R7479 vdd.n9153 vdd.n9152 93.7417
R7480 vdd.n9152 vdd.n9141 93.7417
R7481 vdd.n9093 vdd.n9088 93.7417
R7482 vdd.n9116 vdd.n9093 93.7417
R7483 vdd.n9128 vdd.n9086 93.7417
R7484 vdd.n9114 vdd.n9086 93.7417
R7485 vdd.n9107 vdd.n9106 93.7417
R7486 vdd.n9106 vdd.n9095 93.7417
R7487 vdd.n9186 vdd.n9181 93.7417
R7488 vdd.n9209 vdd.n9186 93.7417
R7489 vdd.n9221 vdd.n9179 93.7417
R7490 vdd.n9207 vdd.n9179 93.7417
R7491 vdd.n9200 vdd.n9199 93.7417
R7492 vdd.n9199 vdd.n9188 93.7417
R7493 vdd.n9234 vdd.n9229 93.7417
R7494 vdd.n9257 vdd.n9234 93.7417
R7495 vdd.n9269 vdd.n9227 93.7417
R7496 vdd.n9255 vdd.n9227 93.7417
R7497 vdd.n9248 vdd.n9247 93.7417
R7498 vdd.n9247 vdd.n9236 93.7417
R7499 vdd.n9280 vdd.n9275 93.7417
R7500 vdd.n9303 vdd.n9280 93.7417
R7501 vdd.n9315 vdd.n9273 93.7417
R7502 vdd.n9301 vdd.n9273 93.7417
R7503 vdd.n9294 vdd.n9293 93.7417
R7504 vdd.n9293 vdd.n9282 93.7417
R7505 vdd.n6814 vdd.n6813 93.7417
R7506 vdd.n6814 vdd.n6779 93.7417
R7507 vdd.n6811 vdd.n6783 93.7417
R7508 vdd.n6803 vdd.n6783 93.7417
R7509 vdd.n6791 vdd.n6784 93.7417
R7510 vdd.n6801 vdd.n6791 93.7417
R7511 vdd.n9375 vdd.n9370 93.7417
R7512 vdd.n9398 vdd.n9375 93.7417
R7513 vdd.n9410 vdd.n9368 93.7417
R7514 vdd.n9396 vdd.n9368 93.7417
R7515 vdd.n9389 vdd.n9388 93.7417
R7516 vdd.n9388 vdd.n9377 93.7417
R7517 vdd.n9329 vdd.n9324 93.7417
R7518 vdd.n9352 vdd.n9329 93.7417
R7519 vdd.n9364 vdd.n9322 93.7417
R7520 vdd.n9350 vdd.n9322 93.7417
R7521 vdd.n9343 vdd.n9342 93.7417
R7522 vdd.n9342 vdd.n9331 93.7417
R7523 vdd.n9422 vdd.n9417 93.7417
R7524 vdd.n9445 vdd.n9422 93.7417
R7525 vdd.n9457 vdd.n9415 93.7417
R7526 vdd.n9443 vdd.n9415 93.7417
R7527 vdd.n9436 vdd.n9435 93.7417
R7528 vdd.n9435 vdd.n9424 93.7417
R7529 vdd.n9470 vdd.n9465 93.7417
R7530 vdd.n9493 vdd.n9470 93.7417
R7531 vdd.n9505 vdd.n9463 93.7417
R7532 vdd.n9491 vdd.n9463 93.7417
R7533 vdd.n9484 vdd.n9483 93.7417
R7534 vdd.n9483 vdd.n9472 93.7417
R7535 vdd.n9516 vdd.n9511 93.7417
R7536 vdd.n9539 vdd.n9516 93.7417
R7537 vdd.n9551 vdd.n9509 93.7417
R7538 vdd.n9537 vdd.n9509 93.7417
R7539 vdd.n9530 vdd.n9529 93.7417
R7540 vdd.n9529 vdd.n9518 93.7417
R7541 vdd.n3676 vdd.n3671 93.7417
R7542 vdd.n3699 vdd.n3676 93.7417
R7543 vdd.n3711 vdd.n3669 93.7417
R7544 vdd.n3697 vdd.n3669 93.7417
R7545 vdd.n3690 vdd.n3689 93.7417
R7546 vdd.n3689 vdd.n3678 93.7417
R7547 vdd.n3722 vdd.n3717 93.7417
R7548 vdd.n3745 vdd.n3722 93.7417
R7549 vdd.n3757 vdd.n3715 93.7417
R7550 vdd.n3743 vdd.n3715 93.7417
R7551 vdd.n3736 vdd.n3735 93.7417
R7552 vdd.n3735 vdd.n3724 93.7417
R7553 vdd.n3820 vdd.n3815 93.7417
R7554 vdd.n3843 vdd.n3820 93.7417
R7555 vdd.n3855 vdd.n3813 93.7417
R7556 vdd.n3841 vdd.n3813 93.7417
R7557 vdd.n3834 vdd.n3833 93.7417
R7558 vdd.n3833 vdd.n3822 93.7417
R7559 vdd.n3866 vdd.n3861 93.7417
R7560 vdd.n3889 vdd.n3866 93.7417
R7561 vdd.n3901 vdd.n3859 93.7417
R7562 vdd.n3887 vdd.n3859 93.7417
R7563 vdd.n3880 vdd.n3879 93.7417
R7564 vdd.n3879 vdd.n3868 93.7417
R7565 vdd.n3912 vdd.n3907 93.7417
R7566 vdd.n3935 vdd.n3912 93.7417
R7567 vdd.n3947 vdd.n3905 93.7417
R7568 vdd.n3933 vdd.n3905 93.7417
R7569 vdd.n3926 vdd.n3925 93.7417
R7570 vdd.n3925 vdd.n3914 93.7417
R7571 vdd.n3958 vdd.n3953 93.7417
R7572 vdd.n3981 vdd.n3958 93.7417
R7573 vdd.n3993 vdd.n3951 93.7417
R7574 vdd.n3979 vdd.n3951 93.7417
R7575 vdd.n3972 vdd.n3971 93.7417
R7576 vdd.n3971 vdd.n3960 93.7417
R7577 vdd.n4056 vdd.n4051 93.7417
R7578 vdd.n4079 vdd.n4056 93.7417
R7579 vdd.n4091 vdd.n4049 93.7417
R7580 vdd.n4077 vdd.n4049 93.7417
R7581 vdd.n4070 vdd.n4069 93.7417
R7582 vdd.n4069 vdd.n4058 93.7417
R7583 vdd.n5514 vdd.n5509 93.7417
R7584 vdd.n5537 vdd.n5514 93.7417
R7585 vdd.n5549 vdd.n5507 93.7417
R7586 vdd.n5535 vdd.n5507 93.7417
R7587 vdd.n5528 vdd.n5527 93.7417
R7588 vdd.n5527 vdd.n5516 93.7417
R7589 vdd.n4126 vdd.n4125 93.7417
R7590 vdd.n4125 vdd.n4099 93.7417
R7591 vdd.n4124 vdd.n4097 93.7417
R7592 vdd.n4139 vdd.n4097 93.7417
R7593 vdd.n4116 vdd.n4105 93.7417
R7594 vdd.n4117 vdd.n4116 93.7417
R7595 vdd.n4172 vdd.n4171 93.7417
R7596 vdd.n4171 vdd.n4145 93.7417
R7597 vdd.n4170 vdd.n4143 93.7417
R7598 vdd.n4185 vdd.n4143 93.7417
R7599 vdd.n4162 vdd.n4151 93.7417
R7600 vdd.n4163 vdd.n4162 93.7417
R7601 vdd.n4269 vdd.n4268 93.7417
R7602 vdd.n4268 vdd.n4242 93.7417
R7603 vdd.n4267 vdd.n4240 93.7417
R7604 vdd.n4282 vdd.n4240 93.7417
R7605 vdd.n4259 vdd.n4248 93.7417
R7606 vdd.n4260 vdd.n4259 93.7417
R7607 vdd.n4315 vdd.n4314 93.7417
R7608 vdd.n4314 vdd.n4288 93.7417
R7609 vdd.n4313 vdd.n4286 93.7417
R7610 vdd.n4328 vdd.n4286 93.7417
R7611 vdd.n4305 vdd.n4294 93.7417
R7612 vdd.n4306 vdd.n4305 93.7417
R7613 vdd.n4361 vdd.n4360 93.7417
R7614 vdd.n4360 vdd.n4334 93.7417
R7615 vdd.n4359 vdd.n4332 93.7417
R7616 vdd.n4374 vdd.n4332 93.7417
R7617 vdd.n4351 vdd.n4340 93.7417
R7618 vdd.n4352 vdd.n4351 93.7417
R7619 vdd.n4407 vdd.n4406 93.7417
R7620 vdd.n4406 vdd.n4380 93.7417
R7621 vdd.n4405 vdd.n4378 93.7417
R7622 vdd.n4420 vdd.n4378 93.7417
R7623 vdd.n4397 vdd.n4386 93.7417
R7624 vdd.n4398 vdd.n4397 93.7417
R7625 vdd.n4504 vdd.n4503 93.7417
R7626 vdd.n4503 vdd.n4477 93.7417
R7627 vdd.n4502 vdd.n4475 93.7417
R7628 vdd.n4517 vdd.n4475 93.7417
R7629 vdd.n4494 vdd.n4483 93.7417
R7630 vdd.n4495 vdd.n4494 93.7417
R7631 vdd.n3653 vdd.n3652 93.7417
R7632 vdd.n3652 vdd.n3626 93.7417
R7633 vdd.n3651 vdd.n3624 93.7417
R7634 vdd.n3666 vdd.n3624 93.7417
R7635 vdd.n3643 vdd.n3632 93.7417
R7636 vdd.n3644 vdd.n3643 93.7417
R7637 vdd.n4548 vdd.n4547 93.7417
R7638 vdd.n4547 vdd.n4521 93.7417
R7639 vdd.n4546 vdd.n4519 93.7417
R7640 vdd.n4561 vdd.n4519 93.7417
R7641 vdd.n4538 vdd.n4527 93.7417
R7642 vdd.n4539 vdd.n4538 93.7417
R7643 vdd.n4593 vdd.n4592 93.7417
R7644 vdd.n4592 vdd.n4566 93.7417
R7645 vdd.n4591 vdd.n4564 93.7417
R7646 vdd.n4606 vdd.n4564 93.7417
R7647 vdd.n4583 vdd.n4572 93.7417
R7648 vdd.n4584 vdd.n4583 93.7417
R7649 vdd.n4643 vdd.n4642 93.7417
R7650 vdd.n4642 vdd.n4616 93.7417
R7651 vdd.n4641 vdd.n4614 93.7417
R7652 vdd.n4656 vdd.n4614 93.7417
R7653 vdd.n4633 vdd.n4622 93.7417
R7654 vdd.n4634 vdd.n4633 93.7417
R7655 vdd.n4689 vdd.n4688 93.7417
R7656 vdd.n4688 vdd.n4662 93.7417
R7657 vdd.n4687 vdd.n4660 93.7417
R7658 vdd.n4702 vdd.n4660 93.7417
R7659 vdd.n4679 vdd.n4668 93.7417
R7660 vdd.n4680 vdd.n4679 93.7417
R7661 vdd.n4737 vdd.n4736 93.7417
R7662 vdd.n4736 vdd.n4710 93.7417
R7663 vdd.n4735 vdd.n4708 93.7417
R7664 vdd.n4750 vdd.n4708 93.7417
R7665 vdd.n4727 vdd.n4716 93.7417
R7666 vdd.n4728 vdd.n4727 93.7417
R7667 vdd.n4449 vdd.n4448 93.7417
R7668 vdd.n4448 vdd.n4432 93.7417
R7669 vdd.n4447 vdd.n4430 93.7417
R7670 vdd.n4463 vdd.n4430 93.7417
R7671 vdd.n4440 vdd.n4439 93.7417
R7672 vdd.n4439 vdd.n4425 93.7417
R7673 vdd.n4784 vdd.n4783 93.7417
R7674 vdd.n4783 vdd.n4757 93.7417
R7675 vdd.n4782 vdd.n4755 93.7417
R7676 vdd.n4797 vdd.n4755 93.7417
R7677 vdd.n4774 vdd.n4763 93.7417
R7678 vdd.n4775 vdd.n4774 93.7417
R7679 vdd.n4829 vdd.n4828 93.7417
R7680 vdd.n4828 vdd.n4802 93.7417
R7681 vdd.n4827 vdd.n4800 93.7417
R7682 vdd.n4842 vdd.n4800 93.7417
R7683 vdd.n4819 vdd.n4808 93.7417
R7684 vdd.n4820 vdd.n4819 93.7417
R7685 vdd.n4875 vdd.n4874 93.7417
R7686 vdd.n4874 vdd.n4848 93.7417
R7687 vdd.n4873 vdd.n4846 93.7417
R7688 vdd.n4888 vdd.n4846 93.7417
R7689 vdd.n4865 vdd.n4854 93.7417
R7690 vdd.n4866 vdd.n4865 93.7417
R7691 vdd.n4926 vdd.n4925 93.7417
R7692 vdd.n4925 vdd.n4899 93.7417
R7693 vdd.n4924 vdd.n4897 93.7417
R7694 vdd.n4939 vdd.n4897 93.7417
R7695 vdd.n4916 vdd.n4905 93.7417
R7696 vdd.n4917 vdd.n4916 93.7417
R7697 vdd.n4972 vdd.n4971 93.7417
R7698 vdd.n4971 vdd.n4945 93.7417
R7699 vdd.n4970 vdd.n4943 93.7417
R7700 vdd.n4985 vdd.n4943 93.7417
R7701 vdd.n4962 vdd.n4951 93.7417
R7702 vdd.n4963 vdd.n4962 93.7417
R7703 vdd.n5020 vdd.n5019 93.7417
R7704 vdd.n5019 vdd.n4993 93.7417
R7705 vdd.n5018 vdd.n4991 93.7417
R7706 vdd.n5033 vdd.n4991 93.7417
R7707 vdd.n5010 vdd.n4999 93.7417
R7708 vdd.n5011 vdd.n5010 93.7417
R7709 vdd.n5066 vdd.n5065 93.7417
R7710 vdd.n5065 vdd.n5039 93.7417
R7711 vdd.n5064 vdd.n5037 93.7417
R7712 vdd.n5079 vdd.n5037 93.7417
R7713 vdd.n5056 vdd.n5045 93.7417
R7714 vdd.n5057 vdd.n5056 93.7417
R7715 vdd.n5111 vdd.n5110 93.7417
R7716 vdd.n5110 vdd.n5084 93.7417
R7717 vdd.n5109 vdd.n5082 93.7417
R7718 vdd.n5124 vdd.n5082 93.7417
R7719 vdd.n5101 vdd.n5090 93.7417
R7720 vdd.n5102 vdd.n5101 93.7417
R7721 vdd.n5161 vdd.n5160 93.7417
R7722 vdd.n5160 vdd.n5134 93.7417
R7723 vdd.n5159 vdd.n5132 93.7417
R7724 vdd.n5174 vdd.n5132 93.7417
R7725 vdd.n5151 vdd.n5140 93.7417
R7726 vdd.n5152 vdd.n5151 93.7417
R7727 vdd.n5207 vdd.n5206 93.7417
R7728 vdd.n5206 vdd.n5180 93.7417
R7729 vdd.n5205 vdd.n5178 93.7417
R7730 vdd.n5220 vdd.n5178 93.7417
R7731 vdd.n5197 vdd.n5186 93.7417
R7732 vdd.n5198 vdd.n5197 93.7417
R7733 vdd.n5255 vdd.n5254 93.7417
R7734 vdd.n5254 vdd.n5228 93.7417
R7735 vdd.n5253 vdd.n5226 93.7417
R7736 vdd.n5268 vdd.n5226 93.7417
R7737 vdd.n5245 vdd.n5234 93.7417
R7738 vdd.n5246 vdd.n5245 93.7417
R7739 vdd.n4214 vdd.n4213 93.7417
R7740 vdd.n4213 vdd.n4197 93.7417
R7741 vdd.n4212 vdd.n4195 93.7417
R7742 vdd.n4228 vdd.n4195 93.7417
R7743 vdd.n4205 vdd.n4204 93.7417
R7744 vdd.n4204 vdd.n4190 93.7417
R7745 vdd.n5302 vdd.n5301 93.7417
R7746 vdd.n5301 vdd.n5275 93.7417
R7747 vdd.n5300 vdd.n5273 93.7417
R7748 vdd.n5315 vdd.n5273 93.7417
R7749 vdd.n5292 vdd.n5281 93.7417
R7750 vdd.n5293 vdd.n5292 93.7417
R7751 vdd.n5347 vdd.n5346 93.7417
R7752 vdd.n5346 vdd.n5320 93.7417
R7753 vdd.n5345 vdd.n5318 93.7417
R7754 vdd.n5360 vdd.n5318 93.7417
R7755 vdd.n5337 vdd.n5326 93.7417
R7756 vdd.n5338 vdd.n5337 93.7417
R7757 vdd.n5397 vdd.n5396 93.7417
R7758 vdd.n5396 vdd.n5370 93.7417
R7759 vdd.n5395 vdd.n5368 93.7417
R7760 vdd.n5410 vdd.n5368 93.7417
R7761 vdd.n5387 vdd.n5376 93.7417
R7762 vdd.n5388 vdd.n5387 93.7417
R7763 vdd.n5443 vdd.n5442 93.7417
R7764 vdd.n5442 vdd.n5416 93.7417
R7765 vdd.n5441 vdd.n5414 93.7417
R7766 vdd.n5456 vdd.n5414 93.7417
R7767 vdd.n5433 vdd.n5422 93.7417
R7768 vdd.n5434 vdd.n5433 93.7417
R7769 vdd.n5491 vdd.n5490 93.7417
R7770 vdd.n5490 vdd.n5464 93.7417
R7771 vdd.n5489 vdd.n5462 93.7417
R7772 vdd.n5504 vdd.n5462 93.7417
R7773 vdd.n5481 vdd.n5470 93.7417
R7774 vdd.n5482 vdd.n5481 93.7417
R7775 vdd.n5607 vdd.n5602 93.7417
R7776 vdd.n5630 vdd.n5607 93.7417
R7777 vdd.n5642 vdd.n5600 93.7417
R7778 vdd.n5628 vdd.n5600 93.7417
R7779 vdd.n5621 vdd.n5620 93.7417
R7780 vdd.n5620 vdd.n5609 93.7417
R7781 vdd.n5561 vdd.n5556 93.7417
R7782 vdd.n5584 vdd.n5561 93.7417
R7783 vdd.n5596 vdd.n5554 93.7417
R7784 vdd.n5582 vdd.n5554 93.7417
R7785 vdd.n5575 vdd.n5574 93.7417
R7786 vdd.n5574 vdd.n5563 93.7417
R7787 vdd.n5654 vdd.n5649 93.7417
R7788 vdd.n5677 vdd.n5654 93.7417
R7789 vdd.n5689 vdd.n5647 93.7417
R7790 vdd.n5675 vdd.n5647 93.7417
R7791 vdd.n5668 vdd.n5667 93.7417
R7792 vdd.n5667 vdd.n5656 93.7417
R7793 vdd.n5702 vdd.n5697 93.7417
R7794 vdd.n5725 vdd.n5702 93.7417
R7795 vdd.n5737 vdd.n5695 93.7417
R7796 vdd.n5723 vdd.n5695 93.7417
R7797 vdd.n5716 vdd.n5715 93.7417
R7798 vdd.n5715 vdd.n5704 93.7417
R7799 vdd.n5748 vdd.n5743 93.7417
R7800 vdd.n5771 vdd.n5748 93.7417
R7801 vdd.n5783 vdd.n5741 93.7417
R7802 vdd.n5769 vdd.n5741 93.7417
R7803 vdd.n5762 vdd.n5761 93.7417
R7804 vdd.n5761 vdd.n5750 93.7417
R7805 vdd.n4036 vdd.n4035 93.7417
R7806 vdd.n4036 vdd.n4001 93.7417
R7807 vdd.n4033 vdd.n4005 93.7417
R7808 vdd.n4025 vdd.n4005 93.7417
R7809 vdd.n4013 vdd.n4006 93.7417
R7810 vdd.n4023 vdd.n4013 93.7417
R7811 vdd.n5890 vdd.n5885 93.7417
R7812 vdd.n5913 vdd.n5890 93.7417
R7813 vdd.n5925 vdd.n5883 93.7417
R7814 vdd.n5911 vdd.n5883 93.7417
R7815 vdd.n5904 vdd.n5903 93.7417
R7816 vdd.n5903 vdd.n5892 93.7417
R7817 vdd.n5843 vdd.n5838 93.7417
R7818 vdd.n5866 vdd.n5843 93.7417
R7819 vdd.n5878 vdd.n5836 93.7417
R7820 vdd.n5864 vdd.n5836 93.7417
R7821 vdd.n5857 vdd.n5856 93.7417
R7822 vdd.n5856 vdd.n5845 93.7417
R7823 vdd.n5797 vdd.n5792 93.7417
R7824 vdd.n5820 vdd.n5797 93.7417
R7825 vdd.n5832 vdd.n5790 93.7417
R7826 vdd.n5818 vdd.n5790 93.7417
R7827 vdd.n5811 vdd.n5810 93.7417
R7828 vdd.n5810 vdd.n5799 93.7417
R7829 vdd.n5937 vdd.n5932 93.7417
R7830 vdd.n5960 vdd.n5937 93.7417
R7831 vdd.n5972 vdd.n5930 93.7417
R7832 vdd.n5958 vdd.n5930 93.7417
R7833 vdd.n5951 vdd.n5950 93.7417
R7834 vdd.n5950 vdd.n5939 93.7417
R7835 vdd.n5985 vdd.n5980 93.7417
R7836 vdd.n6008 vdd.n5985 93.7417
R7837 vdd.n6020 vdd.n5978 93.7417
R7838 vdd.n6006 vdd.n5978 93.7417
R7839 vdd.n5999 vdd.n5998 93.7417
R7840 vdd.n5998 vdd.n5987 93.7417
R7841 vdd.n6031 vdd.n6026 93.7417
R7842 vdd.n6054 vdd.n6031 93.7417
R7843 vdd.n6066 vdd.n6024 93.7417
R7844 vdd.n6052 vdd.n6024 93.7417
R7845 vdd.n6045 vdd.n6044 93.7417
R7846 vdd.n6044 vdd.n6033 93.7417
R7847 vdd.n6125 vdd.n6120 93.7417
R7848 vdd.n6148 vdd.n6125 93.7417
R7849 vdd.n6160 vdd.n6118 93.7417
R7850 vdd.n6146 vdd.n6118 93.7417
R7851 vdd.n6139 vdd.n6138 93.7417
R7852 vdd.n6138 vdd.n6127 93.7417
R7853 vdd.n6079 vdd.n6074 93.7417
R7854 vdd.n6102 vdd.n6079 93.7417
R7855 vdd.n6114 vdd.n6072 93.7417
R7856 vdd.n6100 vdd.n6072 93.7417
R7857 vdd.n6093 vdd.n6092 93.7417
R7858 vdd.n6092 vdd.n6081 93.7417
R7859 vdd.n6172 vdd.n6167 93.7417
R7860 vdd.n6195 vdd.n6172 93.7417
R7861 vdd.n6207 vdd.n6165 93.7417
R7862 vdd.n6193 vdd.n6165 93.7417
R7863 vdd.n6186 vdd.n6185 93.7417
R7864 vdd.n6185 vdd.n6174 93.7417
R7865 vdd.n6220 vdd.n6215 93.7417
R7866 vdd.n6243 vdd.n6220 93.7417
R7867 vdd.n6255 vdd.n6213 93.7417
R7868 vdd.n6241 vdd.n6213 93.7417
R7869 vdd.n6234 vdd.n6233 93.7417
R7870 vdd.n6233 vdd.n6222 93.7417
R7871 vdd.n6266 vdd.n6261 93.7417
R7872 vdd.n6289 vdd.n6266 93.7417
R7873 vdd.n6301 vdd.n6259 93.7417
R7874 vdd.n6287 vdd.n6259 93.7417
R7875 vdd.n6280 vdd.n6279 93.7417
R7876 vdd.n6279 vdd.n6268 93.7417
R7877 vdd.n3800 vdd.n3799 93.7417
R7878 vdd.n3800 vdd.n3765 93.7417
R7879 vdd.n3797 vdd.n3769 93.7417
R7880 vdd.n3789 vdd.n3769 93.7417
R7881 vdd.n3777 vdd.n3770 93.7417
R7882 vdd.n3787 vdd.n3777 93.7417
R7883 vdd.n6361 vdd.n6356 93.7417
R7884 vdd.n6384 vdd.n6361 93.7417
R7885 vdd.n6396 vdd.n6354 93.7417
R7886 vdd.n6382 vdd.n6354 93.7417
R7887 vdd.n6375 vdd.n6374 93.7417
R7888 vdd.n6374 vdd.n6363 93.7417
R7889 vdd.n6315 vdd.n6310 93.7417
R7890 vdd.n6338 vdd.n6315 93.7417
R7891 vdd.n6350 vdd.n6308 93.7417
R7892 vdd.n6336 vdd.n6308 93.7417
R7893 vdd.n6329 vdd.n6328 93.7417
R7894 vdd.n6328 vdd.n6317 93.7417
R7895 vdd.n6408 vdd.n6403 93.7417
R7896 vdd.n6431 vdd.n6408 93.7417
R7897 vdd.n6443 vdd.n6401 93.7417
R7898 vdd.n6429 vdd.n6401 93.7417
R7899 vdd.n6422 vdd.n6421 93.7417
R7900 vdd.n6421 vdd.n6410 93.7417
R7901 vdd.n6456 vdd.n6451 93.7417
R7902 vdd.n6479 vdd.n6456 93.7417
R7903 vdd.n6491 vdd.n6449 93.7417
R7904 vdd.n6477 vdd.n6449 93.7417
R7905 vdd.n6470 vdd.n6469 93.7417
R7906 vdd.n6469 vdd.n6458 93.7417
R7907 vdd.n6502 vdd.n6497 93.7417
R7908 vdd.n6525 vdd.n6502 93.7417
R7909 vdd.n6537 vdd.n6495 93.7417
R7910 vdd.n6523 vdd.n6495 93.7417
R7911 vdd.n6516 vdd.n6515 93.7417
R7912 vdd.n6515 vdd.n6504 93.7417
R7913 vdd.n662 vdd.n657 93.7417
R7914 vdd.n685 vdd.n662 93.7417
R7915 vdd.n697 vdd.n655 93.7417
R7916 vdd.n683 vdd.n655 93.7417
R7917 vdd.n676 vdd.n675 93.7417
R7918 vdd.n675 vdd.n664 93.7417
R7919 vdd.n708 vdd.n703 93.7417
R7920 vdd.n731 vdd.n708 93.7417
R7921 vdd.n743 vdd.n701 93.7417
R7922 vdd.n729 vdd.n701 93.7417
R7923 vdd.n722 vdd.n721 93.7417
R7924 vdd.n721 vdd.n710 93.7417
R7925 vdd.n806 vdd.n801 93.7417
R7926 vdd.n829 vdd.n806 93.7417
R7927 vdd.n841 vdd.n799 93.7417
R7928 vdd.n827 vdd.n799 93.7417
R7929 vdd.n820 vdd.n819 93.7417
R7930 vdd.n819 vdd.n808 93.7417
R7931 vdd.n852 vdd.n847 93.7417
R7932 vdd.n875 vdd.n852 93.7417
R7933 vdd.n887 vdd.n845 93.7417
R7934 vdd.n873 vdd.n845 93.7417
R7935 vdd.n866 vdd.n865 93.7417
R7936 vdd.n865 vdd.n854 93.7417
R7937 vdd.n898 vdd.n893 93.7417
R7938 vdd.n921 vdd.n898 93.7417
R7939 vdd.n933 vdd.n891 93.7417
R7940 vdd.n919 vdd.n891 93.7417
R7941 vdd.n912 vdd.n911 93.7417
R7942 vdd.n911 vdd.n900 93.7417
R7943 vdd.n944 vdd.n939 93.7417
R7944 vdd.n967 vdd.n944 93.7417
R7945 vdd.n979 vdd.n937 93.7417
R7946 vdd.n965 vdd.n937 93.7417
R7947 vdd.n958 vdd.n957 93.7417
R7948 vdd.n957 vdd.n946 93.7417
R7949 vdd.n1042 vdd.n1037 93.7417
R7950 vdd.n1065 vdd.n1042 93.7417
R7951 vdd.n1077 vdd.n1035 93.7417
R7952 vdd.n1063 vdd.n1035 93.7417
R7953 vdd.n1056 vdd.n1055 93.7417
R7954 vdd.n1055 vdd.n1044 93.7417
R7955 vdd.n2500 vdd.n2495 93.7417
R7956 vdd.n2523 vdd.n2500 93.7417
R7957 vdd.n2535 vdd.n2493 93.7417
R7958 vdd.n2521 vdd.n2493 93.7417
R7959 vdd.n2514 vdd.n2513 93.7417
R7960 vdd.n2513 vdd.n2502 93.7417
R7961 vdd.n1112 vdd.n1111 93.7417
R7962 vdd.n1111 vdd.n1085 93.7417
R7963 vdd.n1110 vdd.n1083 93.7417
R7964 vdd.n1125 vdd.n1083 93.7417
R7965 vdd.n1102 vdd.n1091 93.7417
R7966 vdd.n1103 vdd.n1102 93.7417
R7967 vdd.n1158 vdd.n1157 93.7417
R7968 vdd.n1157 vdd.n1131 93.7417
R7969 vdd.n1156 vdd.n1129 93.7417
R7970 vdd.n1171 vdd.n1129 93.7417
R7971 vdd.n1148 vdd.n1137 93.7417
R7972 vdd.n1149 vdd.n1148 93.7417
R7973 vdd.n1255 vdd.n1254 93.7417
R7974 vdd.n1254 vdd.n1228 93.7417
R7975 vdd.n1253 vdd.n1226 93.7417
R7976 vdd.n1268 vdd.n1226 93.7417
R7977 vdd.n1245 vdd.n1234 93.7417
R7978 vdd.n1246 vdd.n1245 93.7417
R7979 vdd.n1301 vdd.n1300 93.7417
R7980 vdd.n1300 vdd.n1274 93.7417
R7981 vdd.n1299 vdd.n1272 93.7417
R7982 vdd.n1314 vdd.n1272 93.7417
R7983 vdd.n1291 vdd.n1280 93.7417
R7984 vdd.n1292 vdd.n1291 93.7417
R7985 vdd.n1347 vdd.n1346 93.7417
R7986 vdd.n1346 vdd.n1320 93.7417
R7987 vdd.n1345 vdd.n1318 93.7417
R7988 vdd.n1360 vdd.n1318 93.7417
R7989 vdd.n1337 vdd.n1326 93.7417
R7990 vdd.n1338 vdd.n1337 93.7417
R7991 vdd.n1393 vdd.n1392 93.7417
R7992 vdd.n1392 vdd.n1366 93.7417
R7993 vdd.n1391 vdd.n1364 93.7417
R7994 vdd.n1406 vdd.n1364 93.7417
R7995 vdd.n1383 vdd.n1372 93.7417
R7996 vdd.n1384 vdd.n1383 93.7417
R7997 vdd.n1490 vdd.n1489 93.7417
R7998 vdd.n1489 vdd.n1463 93.7417
R7999 vdd.n1488 vdd.n1461 93.7417
R8000 vdd.n1503 vdd.n1461 93.7417
R8001 vdd.n1480 vdd.n1469 93.7417
R8002 vdd.n1481 vdd.n1480 93.7417
R8003 vdd.n639 vdd.n638 93.7417
R8004 vdd.n638 vdd.n612 93.7417
R8005 vdd.n637 vdd.n610 93.7417
R8006 vdd.n652 vdd.n610 93.7417
R8007 vdd.n629 vdd.n618 93.7417
R8008 vdd.n630 vdd.n629 93.7417
R8009 vdd.n1534 vdd.n1533 93.7417
R8010 vdd.n1533 vdd.n1507 93.7417
R8011 vdd.n1532 vdd.n1505 93.7417
R8012 vdd.n1547 vdd.n1505 93.7417
R8013 vdd.n1524 vdd.n1513 93.7417
R8014 vdd.n1525 vdd.n1524 93.7417
R8015 vdd.n1579 vdd.n1578 93.7417
R8016 vdd.n1578 vdd.n1552 93.7417
R8017 vdd.n1577 vdd.n1550 93.7417
R8018 vdd.n1592 vdd.n1550 93.7417
R8019 vdd.n1569 vdd.n1558 93.7417
R8020 vdd.n1570 vdd.n1569 93.7417
R8021 vdd.n1629 vdd.n1628 93.7417
R8022 vdd.n1628 vdd.n1602 93.7417
R8023 vdd.n1627 vdd.n1600 93.7417
R8024 vdd.n1642 vdd.n1600 93.7417
R8025 vdd.n1619 vdd.n1608 93.7417
R8026 vdd.n1620 vdd.n1619 93.7417
R8027 vdd.n1675 vdd.n1674 93.7417
R8028 vdd.n1674 vdd.n1648 93.7417
R8029 vdd.n1673 vdd.n1646 93.7417
R8030 vdd.n1688 vdd.n1646 93.7417
R8031 vdd.n1665 vdd.n1654 93.7417
R8032 vdd.n1666 vdd.n1665 93.7417
R8033 vdd.n1723 vdd.n1722 93.7417
R8034 vdd.n1722 vdd.n1696 93.7417
R8035 vdd.n1721 vdd.n1694 93.7417
R8036 vdd.n1736 vdd.n1694 93.7417
R8037 vdd.n1713 vdd.n1702 93.7417
R8038 vdd.n1714 vdd.n1713 93.7417
R8039 vdd.n1435 vdd.n1434 93.7417
R8040 vdd.n1434 vdd.n1418 93.7417
R8041 vdd.n1433 vdd.n1416 93.7417
R8042 vdd.n1449 vdd.n1416 93.7417
R8043 vdd.n1426 vdd.n1425 93.7417
R8044 vdd.n1425 vdd.n1411 93.7417
R8045 vdd.n1770 vdd.n1769 93.7417
R8046 vdd.n1769 vdd.n1743 93.7417
R8047 vdd.n1768 vdd.n1741 93.7417
R8048 vdd.n1783 vdd.n1741 93.7417
R8049 vdd.n1760 vdd.n1749 93.7417
R8050 vdd.n1761 vdd.n1760 93.7417
R8051 vdd.n1815 vdd.n1814 93.7417
R8052 vdd.n1814 vdd.n1788 93.7417
R8053 vdd.n1813 vdd.n1786 93.7417
R8054 vdd.n1828 vdd.n1786 93.7417
R8055 vdd.n1805 vdd.n1794 93.7417
R8056 vdd.n1806 vdd.n1805 93.7417
R8057 vdd.n1861 vdd.n1860 93.7417
R8058 vdd.n1860 vdd.n1834 93.7417
R8059 vdd.n1859 vdd.n1832 93.7417
R8060 vdd.n1874 vdd.n1832 93.7417
R8061 vdd.n1851 vdd.n1840 93.7417
R8062 vdd.n1852 vdd.n1851 93.7417
R8063 vdd.n1912 vdd.n1911 93.7417
R8064 vdd.n1911 vdd.n1885 93.7417
R8065 vdd.n1910 vdd.n1883 93.7417
R8066 vdd.n1925 vdd.n1883 93.7417
R8067 vdd.n1902 vdd.n1891 93.7417
R8068 vdd.n1903 vdd.n1902 93.7417
R8069 vdd.n1958 vdd.n1957 93.7417
R8070 vdd.n1957 vdd.n1931 93.7417
R8071 vdd.n1956 vdd.n1929 93.7417
R8072 vdd.n1971 vdd.n1929 93.7417
R8073 vdd.n1948 vdd.n1937 93.7417
R8074 vdd.n1949 vdd.n1948 93.7417
R8075 vdd.n2006 vdd.n2005 93.7417
R8076 vdd.n2005 vdd.n1979 93.7417
R8077 vdd.n2004 vdd.n1977 93.7417
R8078 vdd.n2019 vdd.n1977 93.7417
R8079 vdd.n1996 vdd.n1985 93.7417
R8080 vdd.n1997 vdd.n1996 93.7417
R8081 vdd.n2052 vdd.n2051 93.7417
R8082 vdd.n2051 vdd.n2025 93.7417
R8083 vdd.n2050 vdd.n2023 93.7417
R8084 vdd.n2065 vdd.n2023 93.7417
R8085 vdd.n2042 vdd.n2031 93.7417
R8086 vdd.n2043 vdd.n2042 93.7417
R8087 vdd.n2097 vdd.n2096 93.7417
R8088 vdd.n2096 vdd.n2070 93.7417
R8089 vdd.n2095 vdd.n2068 93.7417
R8090 vdd.n2110 vdd.n2068 93.7417
R8091 vdd.n2087 vdd.n2076 93.7417
R8092 vdd.n2088 vdd.n2087 93.7417
R8093 vdd.n2147 vdd.n2146 93.7417
R8094 vdd.n2146 vdd.n2120 93.7417
R8095 vdd.n2145 vdd.n2118 93.7417
R8096 vdd.n2160 vdd.n2118 93.7417
R8097 vdd.n2137 vdd.n2126 93.7417
R8098 vdd.n2138 vdd.n2137 93.7417
R8099 vdd.n2193 vdd.n2192 93.7417
R8100 vdd.n2192 vdd.n2166 93.7417
R8101 vdd.n2191 vdd.n2164 93.7417
R8102 vdd.n2206 vdd.n2164 93.7417
R8103 vdd.n2183 vdd.n2172 93.7417
R8104 vdd.n2184 vdd.n2183 93.7417
R8105 vdd.n2241 vdd.n2240 93.7417
R8106 vdd.n2240 vdd.n2214 93.7417
R8107 vdd.n2239 vdd.n2212 93.7417
R8108 vdd.n2254 vdd.n2212 93.7417
R8109 vdd.n2231 vdd.n2220 93.7417
R8110 vdd.n2232 vdd.n2231 93.7417
R8111 vdd.n1200 vdd.n1199 93.7417
R8112 vdd.n1199 vdd.n1183 93.7417
R8113 vdd.n1198 vdd.n1181 93.7417
R8114 vdd.n1214 vdd.n1181 93.7417
R8115 vdd.n1191 vdd.n1190 93.7417
R8116 vdd.n1190 vdd.n1176 93.7417
R8117 vdd.n2288 vdd.n2287 93.7417
R8118 vdd.n2287 vdd.n2261 93.7417
R8119 vdd.n2286 vdd.n2259 93.7417
R8120 vdd.n2301 vdd.n2259 93.7417
R8121 vdd.n2278 vdd.n2267 93.7417
R8122 vdd.n2279 vdd.n2278 93.7417
R8123 vdd.n2333 vdd.n2332 93.7417
R8124 vdd.n2332 vdd.n2306 93.7417
R8125 vdd.n2331 vdd.n2304 93.7417
R8126 vdd.n2346 vdd.n2304 93.7417
R8127 vdd.n2323 vdd.n2312 93.7417
R8128 vdd.n2324 vdd.n2323 93.7417
R8129 vdd.n2383 vdd.n2382 93.7417
R8130 vdd.n2382 vdd.n2356 93.7417
R8131 vdd.n2381 vdd.n2354 93.7417
R8132 vdd.n2396 vdd.n2354 93.7417
R8133 vdd.n2373 vdd.n2362 93.7417
R8134 vdd.n2374 vdd.n2373 93.7417
R8135 vdd.n2429 vdd.n2428 93.7417
R8136 vdd.n2428 vdd.n2402 93.7417
R8137 vdd.n2427 vdd.n2400 93.7417
R8138 vdd.n2442 vdd.n2400 93.7417
R8139 vdd.n2419 vdd.n2408 93.7417
R8140 vdd.n2420 vdd.n2419 93.7417
R8141 vdd.n2477 vdd.n2476 93.7417
R8142 vdd.n2476 vdd.n2450 93.7417
R8143 vdd.n2475 vdd.n2448 93.7417
R8144 vdd.n2490 vdd.n2448 93.7417
R8145 vdd.n2467 vdd.n2456 93.7417
R8146 vdd.n2468 vdd.n2467 93.7417
R8147 vdd.n2593 vdd.n2588 93.7417
R8148 vdd.n2616 vdd.n2593 93.7417
R8149 vdd.n2628 vdd.n2586 93.7417
R8150 vdd.n2614 vdd.n2586 93.7417
R8151 vdd.n2607 vdd.n2606 93.7417
R8152 vdd.n2606 vdd.n2595 93.7417
R8153 vdd.n2547 vdd.n2542 93.7417
R8154 vdd.n2570 vdd.n2547 93.7417
R8155 vdd.n2582 vdd.n2540 93.7417
R8156 vdd.n2568 vdd.n2540 93.7417
R8157 vdd.n2561 vdd.n2560 93.7417
R8158 vdd.n2560 vdd.n2549 93.7417
R8159 vdd.n2640 vdd.n2635 93.7417
R8160 vdd.n2663 vdd.n2640 93.7417
R8161 vdd.n2675 vdd.n2633 93.7417
R8162 vdd.n2661 vdd.n2633 93.7417
R8163 vdd.n2654 vdd.n2653 93.7417
R8164 vdd.n2653 vdd.n2642 93.7417
R8165 vdd.n2688 vdd.n2683 93.7417
R8166 vdd.n2711 vdd.n2688 93.7417
R8167 vdd.n2723 vdd.n2681 93.7417
R8168 vdd.n2709 vdd.n2681 93.7417
R8169 vdd.n2702 vdd.n2701 93.7417
R8170 vdd.n2701 vdd.n2690 93.7417
R8171 vdd.n2734 vdd.n2729 93.7417
R8172 vdd.n2757 vdd.n2734 93.7417
R8173 vdd.n2769 vdd.n2727 93.7417
R8174 vdd.n2755 vdd.n2727 93.7417
R8175 vdd.n2748 vdd.n2747 93.7417
R8176 vdd.n2747 vdd.n2736 93.7417
R8177 vdd.n1022 vdd.n1021 93.7417
R8178 vdd.n1022 vdd.n987 93.7417
R8179 vdd.n1019 vdd.n991 93.7417
R8180 vdd.n1011 vdd.n991 93.7417
R8181 vdd.n999 vdd.n992 93.7417
R8182 vdd.n1009 vdd.n999 93.7417
R8183 vdd.n2876 vdd.n2871 93.7417
R8184 vdd.n2899 vdd.n2876 93.7417
R8185 vdd.n2911 vdd.n2869 93.7417
R8186 vdd.n2897 vdd.n2869 93.7417
R8187 vdd.n2890 vdd.n2889 93.7417
R8188 vdd.n2889 vdd.n2878 93.7417
R8189 vdd.n2829 vdd.n2824 93.7417
R8190 vdd.n2852 vdd.n2829 93.7417
R8191 vdd.n2864 vdd.n2822 93.7417
R8192 vdd.n2850 vdd.n2822 93.7417
R8193 vdd.n2843 vdd.n2842 93.7417
R8194 vdd.n2842 vdd.n2831 93.7417
R8195 vdd.n2783 vdd.n2778 93.7417
R8196 vdd.n2806 vdd.n2783 93.7417
R8197 vdd.n2818 vdd.n2776 93.7417
R8198 vdd.n2804 vdd.n2776 93.7417
R8199 vdd.n2797 vdd.n2796 93.7417
R8200 vdd.n2796 vdd.n2785 93.7417
R8201 vdd.n2923 vdd.n2918 93.7417
R8202 vdd.n2946 vdd.n2923 93.7417
R8203 vdd.n2958 vdd.n2916 93.7417
R8204 vdd.n2944 vdd.n2916 93.7417
R8205 vdd.n2937 vdd.n2936 93.7417
R8206 vdd.n2936 vdd.n2925 93.7417
R8207 vdd.n2971 vdd.n2966 93.7417
R8208 vdd.n2994 vdd.n2971 93.7417
R8209 vdd.n3006 vdd.n2964 93.7417
R8210 vdd.n2992 vdd.n2964 93.7417
R8211 vdd.n2985 vdd.n2984 93.7417
R8212 vdd.n2984 vdd.n2973 93.7417
R8213 vdd.n3017 vdd.n3012 93.7417
R8214 vdd.n3040 vdd.n3017 93.7417
R8215 vdd.n3052 vdd.n3010 93.7417
R8216 vdd.n3038 vdd.n3010 93.7417
R8217 vdd.n3031 vdd.n3030 93.7417
R8218 vdd.n3030 vdd.n3019 93.7417
R8219 vdd.n3111 vdd.n3106 93.7417
R8220 vdd.n3134 vdd.n3111 93.7417
R8221 vdd.n3146 vdd.n3104 93.7417
R8222 vdd.n3132 vdd.n3104 93.7417
R8223 vdd.n3125 vdd.n3124 93.7417
R8224 vdd.n3124 vdd.n3113 93.7417
R8225 vdd.n3065 vdd.n3060 93.7417
R8226 vdd.n3088 vdd.n3065 93.7417
R8227 vdd.n3100 vdd.n3058 93.7417
R8228 vdd.n3086 vdd.n3058 93.7417
R8229 vdd.n3079 vdd.n3078 93.7417
R8230 vdd.n3078 vdd.n3067 93.7417
R8231 vdd.n3158 vdd.n3153 93.7417
R8232 vdd.n3181 vdd.n3158 93.7417
R8233 vdd.n3193 vdd.n3151 93.7417
R8234 vdd.n3179 vdd.n3151 93.7417
R8235 vdd.n3172 vdd.n3171 93.7417
R8236 vdd.n3171 vdd.n3160 93.7417
R8237 vdd.n3206 vdd.n3201 93.7417
R8238 vdd.n3229 vdd.n3206 93.7417
R8239 vdd.n3241 vdd.n3199 93.7417
R8240 vdd.n3227 vdd.n3199 93.7417
R8241 vdd.n3220 vdd.n3219 93.7417
R8242 vdd.n3219 vdd.n3208 93.7417
R8243 vdd.n3252 vdd.n3247 93.7417
R8244 vdd.n3275 vdd.n3252 93.7417
R8245 vdd.n3287 vdd.n3245 93.7417
R8246 vdd.n3273 vdd.n3245 93.7417
R8247 vdd.n3266 vdd.n3265 93.7417
R8248 vdd.n3265 vdd.n3254 93.7417
R8249 vdd.n786 vdd.n785 93.7417
R8250 vdd.n786 vdd.n751 93.7417
R8251 vdd.n783 vdd.n755 93.7417
R8252 vdd.n775 vdd.n755 93.7417
R8253 vdd.n763 vdd.n756 93.7417
R8254 vdd.n773 vdd.n763 93.7417
R8255 vdd.n3347 vdd.n3342 93.7417
R8256 vdd.n3370 vdd.n3347 93.7417
R8257 vdd.n3382 vdd.n3340 93.7417
R8258 vdd.n3368 vdd.n3340 93.7417
R8259 vdd.n3361 vdd.n3360 93.7417
R8260 vdd.n3360 vdd.n3349 93.7417
R8261 vdd.n3301 vdd.n3296 93.7417
R8262 vdd.n3324 vdd.n3301 93.7417
R8263 vdd.n3336 vdd.n3294 93.7417
R8264 vdd.n3322 vdd.n3294 93.7417
R8265 vdd.n3315 vdd.n3314 93.7417
R8266 vdd.n3314 vdd.n3303 93.7417
R8267 vdd.n3394 vdd.n3389 93.7417
R8268 vdd.n3417 vdd.n3394 93.7417
R8269 vdd.n3429 vdd.n3387 93.7417
R8270 vdd.n3415 vdd.n3387 93.7417
R8271 vdd.n3408 vdd.n3407 93.7417
R8272 vdd.n3407 vdd.n3396 93.7417
R8273 vdd.n3442 vdd.n3437 93.7417
R8274 vdd.n3465 vdd.n3442 93.7417
R8275 vdd.n3477 vdd.n3435 93.7417
R8276 vdd.n3463 vdd.n3435 93.7417
R8277 vdd.n3456 vdd.n3455 93.7417
R8278 vdd.n3455 vdd.n3444 93.7417
R8279 vdd.n3488 vdd.n3483 93.7417
R8280 vdd.n3511 vdd.n3488 93.7417
R8281 vdd.n3523 vdd.n3481 93.7417
R8282 vdd.n3509 vdd.n3481 93.7417
R8283 vdd.n3502 vdd.n3501 93.7417
R8284 vdd.n3501 vdd.n3490 93.7417
R8285 vdd.n570 vdd.n565 93.7417
R8286 vdd.n593 vdd.n570 93.7417
R8287 vdd.n605 vdd.n563 93.7417
R8288 vdd.n591 vdd.n563 93.7417
R8289 vdd.n584 vdd.n583 93.7417
R8290 vdd.n583 vdd.n572 93.7417
R8291 vdd.n3583 vdd.n3578 93.7417
R8292 vdd.n3606 vdd.n3583 93.7417
R8293 vdd.n3618 vdd.n3576 93.7417
R8294 vdd.n3604 vdd.n3576 93.7417
R8295 vdd.n3597 vdd.n3596 93.7417
R8296 vdd.n3596 vdd.n3585 93.7417
R8297 vdd.n3537 vdd.n3532 93.7417
R8298 vdd.n3560 vdd.n3537 93.7417
R8299 vdd.n3572 vdd.n3530 93.7417
R8300 vdd.n3558 vdd.n3530 93.7417
R8301 vdd.n3551 vdd.n3550 93.7417
R8302 vdd.n3550 vdd.n3539 93.7417
R8303 vdd.n6597 vdd.n6592 93.7417
R8304 vdd.n6620 vdd.n6597 93.7417
R8305 vdd.n6632 vdd.n6590 93.7417
R8306 vdd.n6618 vdd.n6590 93.7417
R8307 vdd.n6611 vdd.n6610 93.7417
R8308 vdd.n6610 vdd.n6599 93.7417
R8309 vdd.n6551 vdd.n6546 93.7417
R8310 vdd.n6574 vdd.n6551 93.7417
R8311 vdd.n6586 vdd.n6544 93.7417
R8312 vdd.n6572 vdd.n6544 93.7417
R8313 vdd.n6565 vdd.n6564 93.7417
R8314 vdd.n6564 vdd.n6553 93.7417
R8315 vdd.n9611 vdd.n9606 93.7417
R8316 vdd.n9634 vdd.n9611 93.7417
R8317 vdd.n9646 vdd.n9604 93.7417
R8318 vdd.n9632 vdd.n9604 93.7417
R8319 vdd.n9625 vdd.n9624 93.7417
R8320 vdd.n9624 vdd.n9613 93.7417
R8321 vdd.n9565 vdd.n9560 93.7417
R8322 vdd.n9588 vdd.n9565 93.7417
R8323 vdd.n9600 vdd.n9558 93.7417
R8324 vdd.n9586 vdd.n9558 93.7417
R8325 vdd.n9579 vdd.n9578 93.7417
R8326 vdd.n9578 vdd.n9567 93.7417
R8327 vdd.n9657 vdd.n9652 93.7417
R8328 vdd.n9680 vdd.n9657 93.7417
R8329 vdd.n9692 vdd.n9650 93.7417
R8330 vdd.n9678 vdd.n9650 93.7417
R8331 vdd.n9671 vdd.n9670 93.7417
R8332 vdd.n9670 vdd.n9659 93.7417
R8333 vdd.n9703 vdd.n9698 93.7417
R8334 vdd.n9726 vdd.n9703 93.7417
R8335 vdd.n9738 vdd.n9696 93.7417
R8336 vdd.n9724 vdd.n9696 93.7417
R8337 vdd.n9717 vdd.n9716 93.7417
R8338 vdd.n9716 vdd.n9705 93.7417
R8339 vdd.n9801 vdd.n9796 93.7417
R8340 vdd.n9824 vdd.n9801 93.7417
R8341 vdd.n9836 vdd.n9794 93.7417
R8342 vdd.n9822 vdd.n9794 93.7417
R8343 vdd.n9815 vdd.n9814 93.7417
R8344 vdd.n9814 vdd.n9803 93.7417
R8345 vdd.n9847 vdd.n9842 93.7417
R8346 vdd.n9870 vdd.n9847 93.7417
R8347 vdd.n9882 vdd.n9840 93.7417
R8348 vdd.n9868 vdd.n9840 93.7417
R8349 vdd.n9861 vdd.n9860 93.7417
R8350 vdd.n9860 vdd.n9849 93.7417
R8351 vdd.n9893 vdd.n9888 93.7417
R8352 vdd.n9916 vdd.n9893 93.7417
R8353 vdd.n9928 vdd.n9886 93.7417
R8354 vdd.n9914 vdd.n9886 93.7417
R8355 vdd.n9907 vdd.n9906 93.7417
R8356 vdd.n9906 vdd.n9895 93.7417
R8357 vdd.n9939 vdd.n9934 93.7417
R8358 vdd.n9962 vdd.n9939 93.7417
R8359 vdd.n9974 vdd.n9932 93.7417
R8360 vdd.n9960 vdd.n9932 93.7417
R8361 vdd.n9953 vdd.n9952 93.7417
R8362 vdd.n9952 vdd.n9941 93.7417
R8363 vdd.n10037 vdd.n10032 93.7417
R8364 vdd.n10060 vdd.n10037 93.7417
R8365 vdd.n10072 vdd.n10030 93.7417
R8366 vdd.n10058 vdd.n10030 93.7417
R8367 vdd.n10051 vdd.n10050 93.7417
R8368 vdd.n10050 vdd.n10039 93.7417
R8369 vdd.n53 vdd.n48 93.7417
R8370 vdd.n76 vdd.n53 93.7417
R8371 vdd.n88 vdd.n46 93.7417
R8372 vdd.n74 vdd.n46 93.7417
R8373 vdd.n67 vdd.n66 93.7417
R8374 vdd.n66 vdd.n55 93.7417
R8375 vdd.n7 vdd.n2 93.7417
R8376 vdd.n30 vdd.n7 93.7417
R8377 vdd.n42 vdd.n0 93.7417
R8378 vdd.n28 vdd.n0 93.7417
R8379 vdd.n21 vdd.n20 93.7417
R8380 vdd.n20 vdd.n9 93.7417
R8381 vdd.n10083 vdd.n10078 93.7417
R8382 vdd.n10106 vdd.n10083 93.7417
R8383 vdd.n10118 vdd.n10076 93.7417
R8384 vdd.n10104 vdd.n10076 93.7417
R8385 vdd.n10097 vdd.n10096 93.7417
R8386 vdd.n10096 vdd.n10085 93.7417
R8387 vdd.n10131 vdd.n10126 93.7417
R8388 vdd.n10154 vdd.n10131 93.7417
R8389 vdd.n10166 vdd.n10124 93.7417
R8390 vdd.n10152 vdd.n10124 93.7417
R8391 vdd.n10145 vdd.n10144 93.7417
R8392 vdd.n10144 vdd.n10133 93.7417
R8393 vdd.n10177 vdd.n10172 93.7417
R8394 vdd.n10200 vdd.n10177 93.7417
R8395 vdd.n10212 vdd.n10170 93.7417
R8396 vdd.n10198 vdd.n10170 93.7417
R8397 vdd.n10191 vdd.n10190 93.7417
R8398 vdd.n10190 vdd.n10179 93.7417
R8399 vdd.n10017 vdd.n10016 93.7417
R8400 vdd.n10017 vdd.n9982 93.7417
R8401 vdd.n10014 vdd.n9986 93.7417
R8402 vdd.n10006 vdd.n9986 93.7417
R8403 vdd.n9994 vdd.n9987 93.7417
R8404 vdd.n10004 vdd.n9994 93.7417
R8405 vdd.n10319 vdd.n10314 93.7417
R8406 vdd.n10342 vdd.n10319 93.7417
R8407 vdd.n10354 vdd.n10312 93.7417
R8408 vdd.n10340 vdd.n10312 93.7417
R8409 vdd.n10333 vdd.n10332 93.7417
R8410 vdd.n10332 vdd.n10321 93.7417
R8411 vdd.n10272 vdd.n10267 93.7417
R8412 vdd.n10295 vdd.n10272 93.7417
R8413 vdd.n10307 vdd.n10265 93.7417
R8414 vdd.n10293 vdd.n10265 93.7417
R8415 vdd.n10286 vdd.n10285 93.7417
R8416 vdd.n10285 vdd.n10274 93.7417
R8417 vdd.n10226 vdd.n10221 93.7417
R8418 vdd.n10249 vdd.n10226 93.7417
R8419 vdd.n10261 vdd.n10219 93.7417
R8420 vdd.n10247 vdd.n10219 93.7417
R8421 vdd.n10240 vdd.n10239 93.7417
R8422 vdd.n10239 vdd.n10228 93.7417
R8423 vdd.n10366 vdd.n10361 93.7417
R8424 vdd.n10389 vdd.n10366 93.7417
R8425 vdd.n10401 vdd.n10359 93.7417
R8426 vdd.n10387 vdd.n10359 93.7417
R8427 vdd.n10380 vdd.n10379 93.7417
R8428 vdd.n10379 vdd.n10368 93.7417
R8429 vdd.n10414 vdd.n10409 93.7417
R8430 vdd.n10437 vdd.n10414 93.7417
R8431 vdd.n10449 vdd.n10407 93.7417
R8432 vdd.n10435 vdd.n10407 93.7417
R8433 vdd.n10428 vdd.n10427 93.7417
R8434 vdd.n10427 vdd.n10416 93.7417
R8435 vdd.n10460 vdd.n10455 93.7417
R8436 vdd.n10483 vdd.n10460 93.7417
R8437 vdd.n10495 vdd.n10453 93.7417
R8438 vdd.n10481 vdd.n10453 93.7417
R8439 vdd.n10474 vdd.n10473 93.7417
R8440 vdd.n10473 vdd.n10462 93.7417
R8441 vdd.n10554 vdd.n10549 93.7417
R8442 vdd.n10577 vdd.n10554 93.7417
R8443 vdd.n10589 vdd.n10547 93.7417
R8444 vdd.n10575 vdd.n10547 93.7417
R8445 vdd.n10568 vdd.n10567 93.7417
R8446 vdd.n10567 vdd.n10556 93.7417
R8447 vdd.n10508 vdd.n10503 93.7417
R8448 vdd.n10531 vdd.n10508 93.7417
R8449 vdd.n10543 vdd.n10501 93.7417
R8450 vdd.n10529 vdd.n10501 93.7417
R8451 vdd.n10522 vdd.n10521 93.7417
R8452 vdd.n10521 vdd.n10510 93.7417
R8453 vdd.n10601 vdd.n10596 93.7417
R8454 vdd.n10624 vdd.n10601 93.7417
R8455 vdd.n10636 vdd.n10594 93.7417
R8456 vdd.n10622 vdd.n10594 93.7417
R8457 vdd.n10615 vdd.n10614 93.7417
R8458 vdd.n10614 vdd.n10603 93.7417
R8459 vdd.n10649 vdd.n10644 93.7417
R8460 vdd.n10672 vdd.n10649 93.7417
R8461 vdd.n10684 vdd.n10642 93.7417
R8462 vdd.n10670 vdd.n10642 93.7417
R8463 vdd.n10663 vdd.n10662 93.7417
R8464 vdd.n10662 vdd.n10651 93.7417
R8465 vdd.n10695 vdd.n10690 93.7417
R8466 vdd.n10718 vdd.n10695 93.7417
R8467 vdd.n10730 vdd.n10688 93.7417
R8468 vdd.n10716 vdd.n10688 93.7417
R8469 vdd.n10709 vdd.n10708 93.7417
R8470 vdd.n10708 vdd.n10697 93.7417
R8471 vdd.n9781 vdd.n9780 93.7417
R8472 vdd.n9781 vdd.n9746 93.7417
R8473 vdd.n9778 vdd.n9750 93.7417
R8474 vdd.n9770 vdd.n9750 93.7417
R8475 vdd.n9758 vdd.n9751 93.7417
R8476 vdd.n9768 vdd.n9758 93.7417
R8477 vdd.n10790 vdd.n10785 93.7417
R8478 vdd.n10813 vdd.n10790 93.7417
R8479 vdd.n10825 vdd.n10783 93.7417
R8480 vdd.n10811 vdd.n10783 93.7417
R8481 vdd.n10804 vdd.n10803 93.7417
R8482 vdd.n10803 vdd.n10792 93.7417
R8483 vdd.n10744 vdd.n10739 93.7417
R8484 vdd.n10767 vdd.n10744 93.7417
R8485 vdd.n10779 vdd.n10737 93.7417
R8486 vdd.n10765 vdd.n10737 93.7417
R8487 vdd.n10758 vdd.n10757 93.7417
R8488 vdd.n10757 vdd.n10746 93.7417
R8489 vdd.n10837 vdd.n10832 93.7417
R8490 vdd.n10860 vdd.n10837 93.7417
R8491 vdd.n10872 vdd.n10830 93.7417
R8492 vdd.n10858 vdd.n10830 93.7417
R8493 vdd.n10851 vdd.n10850 93.7417
R8494 vdd.n10850 vdd.n10839 93.7417
R8495 vdd.n10885 vdd.n10880 93.7417
R8496 vdd.n10908 vdd.n10885 93.7417
R8497 vdd.n10920 vdd.n10878 93.7417
R8498 vdd.n10906 vdd.n10878 93.7417
R8499 vdd.n10899 vdd.n10898 93.7417
R8500 vdd.n10898 vdd.n10887 93.7417
R8501 vdd.n10931 vdd.n10926 93.7417
R8502 vdd.n10954 vdd.n10931 93.7417
R8503 vdd.n10966 vdd.n10924 93.7417
R8504 vdd.n10952 vdd.n10924 93.7417
R8505 vdd.n10945 vdd.n10944 93.7417
R8506 vdd.n10944 vdd.n10933 93.7417
R8507 vdd.n11002 vdd.n11001 93.7417
R8508 vdd.n11001 vdd.n10975 93.7417
R8509 vdd.n11000 vdd.n10973 93.7417
R8510 vdd.n11015 vdd.n10973 93.7417
R8511 vdd.n10992 vdd.n10981 93.7417
R8512 vdd.n10993 vdd.n10992 93.7417
R8513 vdd.n11047 vdd.n11046 93.7417
R8514 vdd.n11046 vdd.n11020 93.7417
R8515 vdd.n11045 vdd.n11018 93.7417
R8516 vdd.n11060 vdd.n11018 93.7417
R8517 vdd.n11037 vdd.n11026 93.7417
R8518 vdd.n11038 vdd.n11037 93.7417
R8519 vdd.n11097 vdd.n11096 93.7417
R8520 vdd.n11096 vdd.n11070 93.7417
R8521 vdd.n11095 vdd.n11068 93.7417
R8522 vdd.n11110 vdd.n11068 93.7417
R8523 vdd.n11087 vdd.n11076 93.7417
R8524 vdd.n11088 vdd.n11087 93.7417
R8525 vdd.n11143 vdd.n11142 93.7417
R8526 vdd.n11142 vdd.n11116 93.7417
R8527 vdd.n11141 vdd.n11114 93.7417
R8528 vdd.n11156 vdd.n11114 93.7417
R8529 vdd.n11133 vdd.n11122 93.7417
R8530 vdd.n11134 vdd.n11133 93.7417
R8531 vdd.n11191 vdd.n11190 93.7417
R8532 vdd.n11190 vdd.n11164 93.7417
R8533 vdd.n11189 vdd.n11162 93.7417
R8534 vdd.n11204 vdd.n11162 93.7417
R8535 vdd.n11181 vdd.n11170 93.7417
R8536 vdd.n11182 vdd.n11181 93.7417
R8537 vdd.n447 vdd.n446 93.7417
R8538 vdd.n446 vdd.n430 93.7417
R8539 vdd.n445 vdd.n428 93.7417
R8540 vdd.n461 vdd.n428 93.7417
R8541 vdd.n438 vdd.n437 93.7417
R8542 vdd.n437 vdd.n423 93.7417
R8543 vdd.n11238 vdd.n11237 93.7417
R8544 vdd.n11237 vdd.n11211 93.7417
R8545 vdd.n11236 vdd.n11209 93.7417
R8546 vdd.n11251 vdd.n11209 93.7417
R8547 vdd.n11228 vdd.n11217 93.7417
R8548 vdd.n11229 vdd.n11228 93.7417
R8549 vdd.n11283 vdd.n11282 93.7417
R8550 vdd.n11282 vdd.n11256 93.7417
R8551 vdd.n11281 vdd.n11254 93.7417
R8552 vdd.n11296 vdd.n11254 93.7417
R8553 vdd.n11273 vdd.n11262 93.7417
R8554 vdd.n11274 vdd.n11273 93.7417
R8555 vdd.n11329 vdd.n11328 93.7417
R8556 vdd.n11328 vdd.n11302 93.7417
R8557 vdd.n11327 vdd.n11300 93.7417
R8558 vdd.n11342 vdd.n11300 93.7417
R8559 vdd.n11319 vdd.n11308 93.7417
R8560 vdd.n11320 vdd.n11319 93.7417
R8561 vdd.n11380 vdd.n11379 93.7417
R8562 vdd.n11379 vdd.n11353 93.7417
R8563 vdd.n11378 vdd.n11351 93.7417
R8564 vdd.n11393 vdd.n11351 93.7417
R8565 vdd.n11370 vdd.n11359 93.7417
R8566 vdd.n11371 vdd.n11370 93.7417
R8567 vdd.n11426 vdd.n11425 93.7417
R8568 vdd.n11425 vdd.n11399 93.7417
R8569 vdd.n11424 vdd.n11397 93.7417
R8570 vdd.n11439 vdd.n11397 93.7417
R8571 vdd.n11416 vdd.n11405 93.7417
R8572 vdd.n11417 vdd.n11416 93.7417
R8573 vdd.n11474 vdd.n11473 93.7417
R8574 vdd.n11473 vdd.n11447 93.7417
R8575 vdd.n11472 vdd.n11445 93.7417
R8576 vdd.n11487 vdd.n11445 93.7417
R8577 vdd.n11464 vdd.n11453 93.7417
R8578 vdd.n11465 vdd.n11464 93.7417
R8579 vdd.n11520 vdd.n11519 93.7417
R8580 vdd.n11519 vdd.n11493 93.7417
R8581 vdd.n11518 vdd.n11491 93.7417
R8582 vdd.n11533 vdd.n11491 93.7417
R8583 vdd.n11510 vdd.n11499 93.7417
R8584 vdd.n11511 vdd.n11510 93.7417
R8585 vdd.n11565 vdd.n11564 93.7417
R8586 vdd.n11564 vdd.n11538 93.7417
R8587 vdd.n11563 vdd.n11536 93.7417
R8588 vdd.n11578 vdd.n11536 93.7417
R8589 vdd.n11555 vdd.n11544 93.7417
R8590 vdd.n11556 vdd.n11555 93.7417
R8591 vdd.n11615 vdd.n11614 93.7417
R8592 vdd.n11614 vdd.n11588 93.7417
R8593 vdd.n11613 vdd.n11586 93.7417
R8594 vdd.n11628 vdd.n11586 93.7417
R8595 vdd.n11605 vdd.n11594 93.7417
R8596 vdd.n11606 vdd.n11605 93.7417
R8597 vdd.n11661 vdd.n11660 93.7417
R8598 vdd.n11660 vdd.n11634 93.7417
R8599 vdd.n11659 vdd.n11632 93.7417
R8600 vdd.n11674 vdd.n11632 93.7417
R8601 vdd.n11651 vdd.n11640 93.7417
R8602 vdd.n11652 vdd.n11651 93.7417
R8603 vdd.n11709 vdd.n11708 93.7417
R8604 vdd.n11708 vdd.n11682 93.7417
R8605 vdd.n11707 vdd.n11680 93.7417
R8606 vdd.n11722 vdd.n11680 93.7417
R8607 vdd.n11699 vdd.n11688 93.7417
R8608 vdd.n11700 vdd.n11699 93.7417
R8609 vdd.n212 vdd.n211 93.7417
R8610 vdd.n211 vdd.n195 93.7417
R8611 vdd.n210 vdd.n193 93.7417
R8612 vdd.n226 vdd.n193 93.7417
R8613 vdd.n203 vdd.n202 93.7417
R8614 vdd.n202 vdd.n188 93.7417
R8615 vdd.n11756 vdd.n11755 93.7417
R8616 vdd.n11755 vdd.n11729 93.7417
R8617 vdd.n11754 vdd.n11727 93.7417
R8618 vdd.n11769 vdd.n11727 93.7417
R8619 vdd.n11746 vdd.n11735 93.7417
R8620 vdd.n11747 vdd.n11746 93.7417
R8621 vdd.n11801 vdd.n11800 93.7417
R8622 vdd.n11800 vdd.n11774 93.7417
R8623 vdd.n11799 vdd.n11772 93.7417
R8624 vdd.n11814 vdd.n11772 93.7417
R8625 vdd.n11791 vdd.n11780 93.7417
R8626 vdd.n11792 vdd.n11791 93.7417
R8627 vdd.n11851 vdd.n11850 93.7417
R8628 vdd.n11850 vdd.n11824 93.7417
R8629 vdd.n11849 vdd.n11822 93.7417
R8630 vdd.n11864 vdd.n11822 93.7417
R8631 vdd.n11841 vdd.n11830 93.7417
R8632 vdd.n11842 vdd.n11841 93.7417
R8633 vdd.n11897 vdd.n11896 93.7417
R8634 vdd.n11896 vdd.n11870 93.7417
R8635 vdd.n11895 vdd.n11868 93.7417
R8636 vdd.n11910 vdd.n11868 93.7417
R8637 vdd.n11887 vdd.n11876 93.7417
R8638 vdd.n11888 vdd.n11887 93.7417
R8639 vdd.n11945 vdd.n11944 93.7417
R8640 vdd.n11944 vdd.n11918 93.7417
R8641 vdd.n11943 vdd.n11916 93.7417
R8642 vdd.n11958 vdd.n11916 93.7417
R8643 vdd.n11935 vdd.n11924 93.7417
R8644 vdd.n11936 vdd.n11935 93.7417
R8645 vdd.n113 vdd.n112 84.1148
R8646 vdd.n131 vdd.n101 84.1148
R8647 vdd.n159 vdd.n158 84.1148
R8648 vdd.n177 vdd.n147 84.1148
R8649 vdd.n256 vdd.n255 84.1148
R8650 vdd.n274 vdd.n244 84.1148
R8651 vdd.n302 vdd.n301 84.1148
R8652 vdd.n320 vdd.n290 84.1148
R8653 vdd.n348 vdd.n347 84.1148
R8654 vdd.n366 vdd.n336 84.1148
R8655 vdd.n394 vdd.n393 84.1148
R8656 vdd.n412 vdd.n382 84.1148
R8657 vdd.n491 vdd.n490 84.1148
R8658 vdd.n509 vdd.n479 84.1148
R8659 vdd.n537 vdd.n536 84.1148
R8660 vdd.n555 vdd.n525 84.1148
R8661 vdd.n6718 vdd.n6717 84.1148
R8662 vdd.n6702 vdd.n6699 84.1148
R8663 vdd.n6764 vdd.n6763 84.1148
R8664 vdd.n6748 vdd.n6745 84.1148
R8665 vdd.n6862 vdd.n6861 84.1148
R8666 vdd.n6846 vdd.n6843 84.1148
R8667 vdd.n6908 vdd.n6907 84.1148
R8668 vdd.n6892 vdd.n6889 84.1148
R8669 vdd.n6954 vdd.n6953 84.1148
R8670 vdd.n6938 vdd.n6935 84.1148
R8671 vdd.n7000 vdd.n6999 84.1148
R8672 vdd.n6984 vdd.n6981 84.1148
R8673 vdd.n7098 vdd.n7097 84.1148
R8674 vdd.n7082 vdd.n7079 84.1148
R8675 vdd.n8556 vdd.n8555 84.1148
R8676 vdd.n8540 vdd.n8537 84.1148
R8677 vdd.n7129 vdd.n7128 84.1148
R8678 vdd.n7147 vdd.n7117 84.1148
R8679 vdd.n7175 vdd.n7174 84.1148
R8680 vdd.n7193 vdd.n7163 84.1148
R8681 vdd.n7272 vdd.n7271 84.1148
R8682 vdd.n7290 vdd.n7260 84.1148
R8683 vdd.n7318 vdd.n7317 84.1148
R8684 vdd.n7336 vdd.n7306 84.1148
R8685 vdd.n7364 vdd.n7363 84.1148
R8686 vdd.n7382 vdd.n7352 84.1148
R8687 vdd.n7410 vdd.n7409 84.1148
R8688 vdd.n7428 vdd.n7398 84.1148
R8689 vdd.n7507 vdd.n7506 84.1148
R8690 vdd.n7525 vdd.n7495 84.1148
R8691 vdd.n6656 vdd.n6655 84.1148
R8692 vdd.n6674 vdd.n6644 84.1148
R8693 vdd.n7551 vdd.n7550 84.1148
R8694 vdd.n7569 vdd.n7539 84.1148
R8695 vdd.n7596 vdd.n7595 84.1148
R8696 vdd.n7614 vdd.n7584 84.1148
R8697 vdd.n7646 vdd.n7645 84.1148
R8698 vdd.n7664 vdd.n7634 84.1148
R8699 vdd.n7692 vdd.n7691 84.1148
R8700 vdd.n7710 vdd.n7680 84.1148
R8701 vdd.n7740 vdd.n7739 84.1148
R8702 vdd.n7758 vdd.n7728 84.1148
R8703 vdd.n7456 vdd.n7438 84.1148
R8704 vdd.n7470 vdd.n7449 84.1148
R8705 vdd.n7787 vdd.n7786 84.1148
R8706 vdd.n7805 vdd.n7775 84.1148
R8707 vdd.n7832 vdd.n7831 84.1148
R8708 vdd.n7850 vdd.n7820 84.1148
R8709 vdd.n7878 vdd.n7877 84.1148
R8710 vdd.n7896 vdd.n7866 84.1148
R8711 vdd.n7929 vdd.n7928 84.1148
R8712 vdd.n7947 vdd.n7917 84.1148
R8713 vdd.n7975 vdd.n7974 84.1148
R8714 vdd.n7993 vdd.n7963 84.1148
R8715 vdd.n8023 vdd.n8022 84.1148
R8716 vdd.n8041 vdd.n8011 84.1148
R8717 vdd.n8069 vdd.n8068 84.1148
R8718 vdd.n8087 vdd.n8057 84.1148
R8719 vdd.n8114 vdd.n8113 84.1148
R8720 vdd.n8132 vdd.n8102 84.1148
R8721 vdd.n8164 vdd.n8163 84.1148
R8722 vdd.n8182 vdd.n8152 84.1148
R8723 vdd.n8210 vdd.n8209 84.1148
R8724 vdd.n8228 vdd.n8198 84.1148
R8725 vdd.n8258 vdd.n8257 84.1148
R8726 vdd.n8276 vdd.n8246 84.1148
R8727 vdd.n7221 vdd.n7203 84.1148
R8728 vdd.n7235 vdd.n7214 84.1148
R8729 vdd.n8305 vdd.n8304 84.1148
R8730 vdd.n8323 vdd.n8293 84.1148
R8731 vdd.n8350 vdd.n8349 84.1148
R8732 vdd.n8368 vdd.n8338 84.1148
R8733 vdd.n8400 vdd.n8399 84.1148
R8734 vdd.n8418 vdd.n8388 84.1148
R8735 vdd.n8446 vdd.n8445 84.1148
R8736 vdd.n8464 vdd.n8434 84.1148
R8737 vdd.n8494 vdd.n8493 84.1148
R8738 vdd.n8512 vdd.n8482 84.1148
R8739 vdd.n8649 vdd.n8648 84.1148
R8740 vdd.n8633 vdd.n8630 84.1148
R8741 vdd.n8603 vdd.n8602 84.1148
R8742 vdd.n8587 vdd.n8584 84.1148
R8743 vdd.n8696 vdd.n8695 84.1148
R8744 vdd.n8680 vdd.n8677 84.1148
R8745 vdd.n8744 vdd.n8743 84.1148
R8746 vdd.n8728 vdd.n8725 84.1148
R8747 vdd.n8790 vdd.n8789 84.1148
R8748 vdd.n8774 vdd.n8771 84.1148
R8749 vdd.n7057 vdd.n7056 84.1148
R8750 vdd.n7036 vdd.n7028 84.1148
R8751 vdd.n8932 vdd.n8931 84.1148
R8752 vdd.n8916 vdd.n8913 84.1148
R8753 vdd.n8885 vdd.n8884 84.1148
R8754 vdd.n8869 vdd.n8866 84.1148
R8755 vdd.n8839 vdd.n8838 84.1148
R8756 vdd.n8823 vdd.n8820 84.1148
R8757 vdd.n8979 vdd.n8978 84.1148
R8758 vdd.n8963 vdd.n8960 84.1148
R8759 vdd.n9027 vdd.n9026 84.1148
R8760 vdd.n9011 vdd.n9008 84.1148
R8761 vdd.n9073 vdd.n9072 84.1148
R8762 vdd.n9057 vdd.n9054 84.1148
R8763 vdd.n9167 vdd.n9166 84.1148
R8764 vdd.n9151 vdd.n9148 84.1148
R8765 vdd.n9121 vdd.n9120 84.1148
R8766 vdd.n9105 vdd.n9102 84.1148
R8767 vdd.n9214 vdd.n9213 84.1148
R8768 vdd.n9198 vdd.n9195 84.1148
R8769 vdd.n9262 vdd.n9261 84.1148
R8770 vdd.n9246 vdd.n9243 84.1148
R8771 vdd.n9308 vdd.n9307 84.1148
R8772 vdd.n9292 vdd.n9289 84.1148
R8773 vdd.n6821 vdd.n6820 84.1148
R8774 vdd.n6800 vdd.n6792 84.1148
R8775 vdd.n9403 vdd.n9402 84.1148
R8776 vdd.n9387 vdd.n9384 84.1148
R8777 vdd.n9357 vdd.n9356 84.1148
R8778 vdd.n9341 vdd.n9338 84.1148
R8779 vdd.n9450 vdd.n9449 84.1148
R8780 vdd.n9434 vdd.n9431 84.1148
R8781 vdd.n9498 vdd.n9497 84.1148
R8782 vdd.n9482 vdd.n9479 84.1148
R8783 vdd.n9544 vdd.n9543 84.1148
R8784 vdd.n9528 vdd.n9525 84.1148
R8785 vdd.n3704 vdd.n3703 84.1148
R8786 vdd.n3688 vdd.n3685 84.1148
R8787 vdd.n3750 vdd.n3749 84.1148
R8788 vdd.n3734 vdd.n3731 84.1148
R8789 vdd.n3848 vdd.n3847 84.1148
R8790 vdd.n3832 vdd.n3829 84.1148
R8791 vdd.n3894 vdd.n3893 84.1148
R8792 vdd.n3878 vdd.n3875 84.1148
R8793 vdd.n3940 vdd.n3939 84.1148
R8794 vdd.n3924 vdd.n3921 84.1148
R8795 vdd.n3986 vdd.n3985 84.1148
R8796 vdd.n3970 vdd.n3967 84.1148
R8797 vdd.n4084 vdd.n4083 84.1148
R8798 vdd.n4068 vdd.n4065 84.1148
R8799 vdd.n5542 vdd.n5541 84.1148
R8800 vdd.n5526 vdd.n5523 84.1148
R8801 vdd.n4115 vdd.n4114 84.1148
R8802 vdd.n4133 vdd.n4103 84.1148
R8803 vdd.n4161 vdd.n4160 84.1148
R8804 vdd.n4179 vdd.n4149 84.1148
R8805 vdd.n4258 vdd.n4257 84.1148
R8806 vdd.n4276 vdd.n4246 84.1148
R8807 vdd.n4304 vdd.n4303 84.1148
R8808 vdd.n4322 vdd.n4292 84.1148
R8809 vdd.n4350 vdd.n4349 84.1148
R8810 vdd.n4368 vdd.n4338 84.1148
R8811 vdd.n4396 vdd.n4395 84.1148
R8812 vdd.n4414 vdd.n4384 84.1148
R8813 vdd.n4493 vdd.n4492 84.1148
R8814 vdd.n4511 vdd.n4481 84.1148
R8815 vdd.n3642 vdd.n3641 84.1148
R8816 vdd.n3660 vdd.n3630 84.1148
R8817 vdd.n4537 vdd.n4536 84.1148
R8818 vdd.n4555 vdd.n4525 84.1148
R8819 vdd.n4582 vdd.n4581 84.1148
R8820 vdd.n4600 vdd.n4570 84.1148
R8821 vdd.n4632 vdd.n4631 84.1148
R8822 vdd.n4650 vdd.n4620 84.1148
R8823 vdd.n4678 vdd.n4677 84.1148
R8824 vdd.n4696 vdd.n4666 84.1148
R8825 vdd.n4726 vdd.n4725 84.1148
R8826 vdd.n4744 vdd.n4714 84.1148
R8827 vdd.n4442 vdd.n4424 84.1148
R8828 vdd.n4456 vdd.n4435 84.1148
R8829 vdd.n4773 vdd.n4772 84.1148
R8830 vdd.n4791 vdd.n4761 84.1148
R8831 vdd.n4818 vdd.n4817 84.1148
R8832 vdd.n4836 vdd.n4806 84.1148
R8833 vdd.n4864 vdd.n4863 84.1148
R8834 vdd.n4882 vdd.n4852 84.1148
R8835 vdd.n4915 vdd.n4914 84.1148
R8836 vdd.n4933 vdd.n4903 84.1148
R8837 vdd.n4961 vdd.n4960 84.1148
R8838 vdd.n4979 vdd.n4949 84.1148
R8839 vdd.n5009 vdd.n5008 84.1148
R8840 vdd.n5027 vdd.n4997 84.1148
R8841 vdd.n5055 vdd.n5054 84.1148
R8842 vdd.n5073 vdd.n5043 84.1148
R8843 vdd.n5100 vdd.n5099 84.1148
R8844 vdd.n5118 vdd.n5088 84.1148
R8845 vdd.n5150 vdd.n5149 84.1148
R8846 vdd.n5168 vdd.n5138 84.1148
R8847 vdd.n5196 vdd.n5195 84.1148
R8848 vdd.n5214 vdd.n5184 84.1148
R8849 vdd.n5244 vdd.n5243 84.1148
R8850 vdd.n5262 vdd.n5232 84.1148
R8851 vdd.n4207 vdd.n4189 84.1148
R8852 vdd.n4221 vdd.n4200 84.1148
R8853 vdd.n5291 vdd.n5290 84.1148
R8854 vdd.n5309 vdd.n5279 84.1148
R8855 vdd.n5336 vdd.n5335 84.1148
R8856 vdd.n5354 vdd.n5324 84.1148
R8857 vdd.n5386 vdd.n5385 84.1148
R8858 vdd.n5404 vdd.n5374 84.1148
R8859 vdd.n5432 vdd.n5431 84.1148
R8860 vdd.n5450 vdd.n5420 84.1148
R8861 vdd.n5480 vdd.n5479 84.1148
R8862 vdd.n5498 vdd.n5468 84.1148
R8863 vdd.n5635 vdd.n5634 84.1148
R8864 vdd.n5619 vdd.n5616 84.1148
R8865 vdd.n5589 vdd.n5588 84.1148
R8866 vdd.n5573 vdd.n5570 84.1148
R8867 vdd.n5682 vdd.n5681 84.1148
R8868 vdd.n5666 vdd.n5663 84.1148
R8869 vdd.n5730 vdd.n5729 84.1148
R8870 vdd.n5714 vdd.n5711 84.1148
R8871 vdd.n5776 vdd.n5775 84.1148
R8872 vdd.n5760 vdd.n5757 84.1148
R8873 vdd.n4043 vdd.n4042 84.1148
R8874 vdd.n4022 vdd.n4014 84.1148
R8875 vdd.n5918 vdd.n5917 84.1148
R8876 vdd.n5902 vdd.n5899 84.1148
R8877 vdd.n5871 vdd.n5870 84.1148
R8878 vdd.n5855 vdd.n5852 84.1148
R8879 vdd.n5825 vdd.n5824 84.1148
R8880 vdd.n5809 vdd.n5806 84.1148
R8881 vdd.n5965 vdd.n5964 84.1148
R8882 vdd.n5949 vdd.n5946 84.1148
R8883 vdd.n6013 vdd.n6012 84.1148
R8884 vdd.n5997 vdd.n5994 84.1148
R8885 vdd.n6059 vdd.n6058 84.1148
R8886 vdd.n6043 vdd.n6040 84.1148
R8887 vdd.n6153 vdd.n6152 84.1148
R8888 vdd.n6137 vdd.n6134 84.1148
R8889 vdd.n6107 vdd.n6106 84.1148
R8890 vdd.n6091 vdd.n6088 84.1148
R8891 vdd.n6200 vdd.n6199 84.1148
R8892 vdd.n6184 vdd.n6181 84.1148
R8893 vdd.n6248 vdd.n6247 84.1148
R8894 vdd.n6232 vdd.n6229 84.1148
R8895 vdd.n6294 vdd.n6293 84.1148
R8896 vdd.n6278 vdd.n6275 84.1148
R8897 vdd.n3807 vdd.n3806 84.1148
R8898 vdd.n3786 vdd.n3778 84.1148
R8899 vdd.n6389 vdd.n6388 84.1148
R8900 vdd.n6373 vdd.n6370 84.1148
R8901 vdd.n6343 vdd.n6342 84.1148
R8902 vdd.n6327 vdd.n6324 84.1148
R8903 vdd.n6436 vdd.n6435 84.1148
R8904 vdd.n6420 vdd.n6417 84.1148
R8905 vdd.n6484 vdd.n6483 84.1148
R8906 vdd.n6468 vdd.n6465 84.1148
R8907 vdd.n6530 vdd.n6529 84.1148
R8908 vdd.n6514 vdd.n6511 84.1148
R8909 vdd.n690 vdd.n689 84.1148
R8910 vdd.n674 vdd.n671 84.1148
R8911 vdd.n736 vdd.n735 84.1148
R8912 vdd.n720 vdd.n717 84.1148
R8913 vdd.n834 vdd.n833 84.1148
R8914 vdd.n818 vdd.n815 84.1148
R8915 vdd.n880 vdd.n879 84.1148
R8916 vdd.n864 vdd.n861 84.1148
R8917 vdd.n926 vdd.n925 84.1148
R8918 vdd.n910 vdd.n907 84.1148
R8919 vdd.n972 vdd.n971 84.1148
R8920 vdd.n956 vdd.n953 84.1148
R8921 vdd.n1070 vdd.n1069 84.1148
R8922 vdd.n1054 vdd.n1051 84.1148
R8923 vdd.n2528 vdd.n2527 84.1148
R8924 vdd.n2512 vdd.n2509 84.1148
R8925 vdd.n1101 vdd.n1100 84.1148
R8926 vdd.n1119 vdd.n1089 84.1148
R8927 vdd.n1147 vdd.n1146 84.1148
R8928 vdd.n1165 vdd.n1135 84.1148
R8929 vdd.n1244 vdd.n1243 84.1148
R8930 vdd.n1262 vdd.n1232 84.1148
R8931 vdd.n1290 vdd.n1289 84.1148
R8932 vdd.n1308 vdd.n1278 84.1148
R8933 vdd.n1336 vdd.n1335 84.1148
R8934 vdd.n1354 vdd.n1324 84.1148
R8935 vdd.n1382 vdd.n1381 84.1148
R8936 vdd.n1400 vdd.n1370 84.1148
R8937 vdd.n1479 vdd.n1478 84.1148
R8938 vdd.n1497 vdd.n1467 84.1148
R8939 vdd.n628 vdd.n627 84.1148
R8940 vdd.n646 vdd.n616 84.1148
R8941 vdd.n1523 vdd.n1522 84.1148
R8942 vdd.n1541 vdd.n1511 84.1148
R8943 vdd.n1568 vdd.n1567 84.1148
R8944 vdd.n1586 vdd.n1556 84.1148
R8945 vdd.n1618 vdd.n1617 84.1148
R8946 vdd.n1636 vdd.n1606 84.1148
R8947 vdd.n1664 vdd.n1663 84.1148
R8948 vdd.n1682 vdd.n1652 84.1148
R8949 vdd.n1712 vdd.n1711 84.1148
R8950 vdd.n1730 vdd.n1700 84.1148
R8951 vdd.n1428 vdd.n1410 84.1148
R8952 vdd.n1442 vdd.n1421 84.1148
R8953 vdd.n1759 vdd.n1758 84.1148
R8954 vdd.n1777 vdd.n1747 84.1148
R8955 vdd.n1804 vdd.n1803 84.1148
R8956 vdd.n1822 vdd.n1792 84.1148
R8957 vdd.n1850 vdd.n1849 84.1148
R8958 vdd.n1868 vdd.n1838 84.1148
R8959 vdd.n1901 vdd.n1900 84.1148
R8960 vdd.n1919 vdd.n1889 84.1148
R8961 vdd.n1947 vdd.n1946 84.1148
R8962 vdd.n1965 vdd.n1935 84.1148
R8963 vdd.n1995 vdd.n1994 84.1148
R8964 vdd.n2013 vdd.n1983 84.1148
R8965 vdd.n2041 vdd.n2040 84.1148
R8966 vdd.n2059 vdd.n2029 84.1148
R8967 vdd.n2086 vdd.n2085 84.1148
R8968 vdd.n2104 vdd.n2074 84.1148
R8969 vdd.n2136 vdd.n2135 84.1148
R8970 vdd.n2154 vdd.n2124 84.1148
R8971 vdd.n2182 vdd.n2181 84.1148
R8972 vdd.n2200 vdd.n2170 84.1148
R8973 vdd.n2230 vdd.n2229 84.1148
R8974 vdd.n2248 vdd.n2218 84.1148
R8975 vdd.n1193 vdd.n1175 84.1148
R8976 vdd.n1207 vdd.n1186 84.1148
R8977 vdd.n2277 vdd.n2276 84.1148
R8978 vdd.n2295 vdd.n2265 84.1148
R8979 vdd.n2322 vdd.n2321 84.1148
R8980 vdd.n2340 vdd.n2310 84.1148
R8981 vdd.n2372 vdd.n2371 84.1148
R8982 vdd.n2390 vdd.n2360 84.1148
R8983 vdd.n2418 vdd.n2417 84.1148
R8984 vdd.n2436 vdd.n2406 84.1148
R8985 vdd.n2466 vdd.n2465 84.1148
R8986 vdd.n2484 vdd.n2454 84.1148
R8987 vdd.n2621 vdd.n2620 84.1148
R8988 vdd.n2605 vdd.n2602 84.1148
R8989 vdd.n2575 vdd.n2574 84.1148
R8990 vdd.n2559 vdd.n2556 84.1148
R8991 vdd.n2668 vdd.n2667 84.1148
R8992 vdd.n2652 vdd.n2649 84.1148
R8993 vdd.n2716 vdd.n2715 84.1148
R8994 vdd.n2700 vdd.n2697 84.1148
R8995 vdd.n2762 vdd.n2761 84.1148
R8996 vdd.n2746 vdd.n2743 84.1148
R8997 vdd.n1029 vdd.n1028 84.1148
R8998 vdd.n1008 vdd.n1000 84.1148
R8999 vdd.n2904 vdd.n2903 84.1148
R9000 vdd.n2888 vdd.n2885 84.1148
R9001 vdd.n2857 vdd.n2856 84.1148
R9002 vdd.n2841 vdd.n2838 84.1148
R9003 vdd.n2811 vdd.n2810 84.1148
R9004 vdd.n2795 vdd.n2792 84.1148
R9005 vdd.n2951 vdd.n2950 84.1148
R9006 vdd.n2935 vdd.n2932 84.1148
R9007 vdd.n2999 vdd.n2998 84.1148
R9008 vdd.n2983 vdd.n2980 84.1148
R9009 vdd.n3045 vdd.n3044 84.1148
R9010 vdd.n3029 vdd.n3026 84.1148
R9011 vdd.n3139 vdd.n3138 84.1148
R9012 vdd.n3123 vdd.n3120 84.1148
R9013 vdd.n3093 vdd.n3092 84.1148
R9014 vdd.n3077 vdd.n3074 84.1148
R9015 vdd.n3186 vdd.n3185 84.1148
R9016 vdd.n3170 vdd.n3167 84.1148
R9017 vdd.n3234 vdd.n3233 84.1148
R9018 vdd.n3218 vdd.n3215 84.1148
R9019 vdd.n3280 vdd.n3279 84.1148
R9020 vdd.n3264 vdd.n3261 84.1148
R9021 vdd.n793 vdd.n792 84.1148
R9022 vdd.n772 vdd.n764 84.1148
R9023 vdd.n3375 vdd.n3374 84.1148
R9024 vdd.n3359 vdd.n3356 84.1148
R9025 vdd.n3329 vdd.n3328 84.1148
R9026 vdd.n3313 vdd.n3310 84.1148
R9027 vdd.n3422 vdd.n3421 84.1148
R9028 vdd.n3406 vdd.n3403 84.1148
R9029 vdd.n3470 vdd.n3469 84.1148
R9030 vdd.n3454 vdd.n3451 84.1148
R9031 vdd.n3516 vdd.n3515 84.1148
R9032 vdd.n3500 vdd.n3497 84.1148
R9033 vdd.n598 vdd.n597 84.1148
R9034 vdd.n582 vdd.n579 84.1148
R9035 vdd.n3611 vdd.n3610 84.1148
R9036 vdd.n3595 vdd.n3592 84.1148
R9037 vdd.n3565 vdd.n3564 84.1148
R9038 vdd.n3549 vdd.n3546 84.1148
R9039 vdd.n6625 vdd.n6624 84.1148
R9040 vdd.n6609 vdd.n6606 84.1148
R9041 vdd.n6579 vdd.n6578 84.1148
R9042 vdd.n6563 vdd.n6560 84.1148
R9043 vdd.n9639 vdd.n9638 84.1148
R9044 vdd.n9623 vdd.n9620 84.1148
R9045 vdd.n9593 vdd.n9592 84.1148
R9046 vdd.n9577 vdd.n9574 84.1148
R9047 vdd.n9685 vdd.n9684 84.1148
R9048 vdd.n9669 vdd.n9666 84.1148
R9049 vdd.n9731 vdd.n9730 84.1148
R9050 vdd.n9715 vdd.n9712 84.1148
R9051 vdd.n9829 vdd.n9828 84.1148
R9052 vdd.n9813 vdd.n9810 84.1148
R9053 vdd.n9875 vdd.n9874 84.1148
R9054 vdd.n9859 vdd.n9856 84.1148
R9055 vdd.n9921 vdd.n9920 84.1148
R9056 vdd.n9905 vdd.n9902 84.1148
R9057 vdd.n9967 vdd.n9966 84.1148
R9058 vdd.n9951 vdd.n9948 84.1148
R9059 vdd.n10065 vdd.n10064 84.1148
R9060 vdd.n10049 vdd.n10046 84.1148
R9061 vdd.n81 vdd.n80 84.1148
R9062 vdd.n65 vdd.n62 84.1148
R9063 vdd.n35 vdd.n34 84.1148
R9064 vdd.n19 vdd.n16 84.1148
R9065 vdd.n10111 vdd.n10110 84.1148
R9066 vdd.n10095 vdd.n10092 84.1148
R9067 vdd.n10159 vdd.n10158 84.1148
R9068 vdd.n10143 vdd.n10140 84.1148
R9069 vdd.n10205 vdd.n10204 84.1148
R9070 vdd.n10189 vdd.n10186 84.1148
R9071 vdd.n10024 vdd.n10023 84.1148
R9072 vdd.n10003 vdd.n9995 84.1148
R9073 vdd.n10347 vdd.n10346 84.1148
R9074 vdd.n10331 vdd.n10328 84.1148
R9075 vdd.n10300 vdd.n10299 84.1148
R9076 vdd.n10284 vdd.n10281 84.1148
R9077 vdd.n10254 vdd.n10253 84.1148
R9078 vdd.n10238 vdd.n10235 84.1148
R9079 vdd.n10394 vdd.n10393 84.1148
R9080 vdd.n10378 vdd.n10375 84.1148
R9081 vdd.n10442 vdd.n10441 84.1148
R9082 vdd.n10426 vdd.n10423 84.1148
R9083 vdd.n10488 vdd.n10487 84.1148
R9084 vdd.n10472 vdd.n10469 84.1148
R9085 vdd.n10582 vdd.n10581 84.1148
R9086 vdd.n10566 vdd.n10563 84.1148
R9087 vdd.n10536 vdd.n10535 84.1148
R9088 vdd.n10520 vdd.n10517 84.1148
R9089 vdd.n10629 vdd.n10628 84.1148
R9090 vdd.n10613 vdd.n10610 84.1148
R9091 vdd.n10677 vdd.n10676 84.1148
R9092 vdd.n10661 vdd.n10658 84.1148
R9093 vdd.n10723 vdd.n10722 84.1148
R9094 vdd.n10707 vdd.n10704 84.1148
R9095 vdd.n9788 vdd.n9787 84.1148
R9096 vdd.n9767 vdd.n9759 84.1148
R9097 vdd.n10818 vdd.n10817 84.1148
R9098 vdd.n10802 vdd.n10799 84.1148
R9099 vdd.n10772 vdd.n10771 84.1148
R9100 vdd.n10756 vdd.n10753 84.1148
R9101 vdd.n10865 vdd.n10864 84.1148
R9102 vdd.n10849 vdd.n10846 84.1148
R9103 vdd.n10913 vdd.n10912 84.1148
R9104 vdd.n10897 vdd.n10894 84.1148
R9105 vdd.n10959 vdd.n10958 84.1148
R9106 vdd.n10943 vdd.n10940 84.1148
R9107 vdd.n10991 vdd.n10990 84.1148
R9108 vdd.n11009 vdd.n10979 84.1148
R9109 vdd.n11036 vdd.n11035 84.1148
R9110 vdd.n11054 vdd.n11024 84.1148
R9111 vdd.n11086 vdd.n11085 84.1148
R9112 vdd.n11104 vdd.n11074 84.1148
R9113 vdd.n11132 vdd.n11131 84.1148
R9114 vdd.n11150 vdd.n11120 84.1148
R9115 vdd.n11180 vdd.n11179 84.1148
R9116 vdd.n11198 vdd.n11168 84.1148
R9117 vdd.n440 vdd.n422 84.1148
R9118 vdd.n454 vdd.n433 84.1148
R9119 vdd.n11227 vdd.n11226 84.1148
R9120 vdd.n11245 vdd.n11215 84.1148
R9121 vdd.n11272 vdd.n11271 84.1148
R9122 vdd.n11290 vdd.n11260 84.1148
R9123 vdd.n11318 vdd.n11317 84.1148
R9124 vdd.n11336 vdd.n11306 84.1148
R9125 vdd.n11369 vdd.n11368 84.1148
R9126 vdd.n11387 vdd.n11357 84.1148
R9127 vdd.n11415 vdd.n11414 84.1148
R9128 vdd.n11433 vdd.n11403 84.1148
R9129 vdd.n11463 vdd.n11462 84.1148
R9130 vdd.n11481 vdd.n11451 84.1148
R9131 vdd.n11509 vdd.n11508 84.1148
R9132 vdd.n11527 vdd.n11497 84.1148
R9133 vdd.n11554 vdd.n11553 84.1148
R9134 vdd.n11572 vdd.n11542 84.1148
R9135 vdd.n11604 vdd.n11603 84.1148
R9136 vdd.n11622 vdd.n11592 84.1148
R9137 vdd.n11650 vdd.n11649 84.1148
R9138 vdd.n11668 vdd.n11638 84.1148
R9139 vdd.n11698 vdd.n11697 84.1148
R9140 vdd.n11716 vdd.n11686 84.1148
R9141 vdd.n205 vdd.n187 84.1148
R9142 vdd.n219 vdd.n198 84.1148
R9143 vdd.n11745 vdd.n11744 84.1148
R9144 vdd.n11763 vdd.n11733 84.1148
R9145 vdd.n11790 vdd.n11789 84.1148
R9146 vdd.n11808 vdd.n11778 84.1148
R9147 vdd.n11840 vdd.n11839 84.1148
R9148 vdd.n11858 vdd.n11828 84.1148
R9149 vdd.n11886 vdd.n11885 84.1148
R9150 vdd.n11904 vdd.n11874 84.1148
R9151 vdd.n11934 vdd.n11933 84.1148
R9152 vdd.n11952 vdd.n11922 84.1148
R9153 vdd.n11993 vdd.n11988 63.3004
R9154 vdd.n11974 vdd.n11969 63.3004
R9155 vdd.n116 vdd.n113 63.3004
R9156 vdd.n132 vdd.n131 63.3004
R9157 vdd.n162 vdd.n159 63.3004
R9158 vdd.n178 vdd.n177 63.3004
R9159 vdd.n259 vdd.n256 63.3004
R9160 vdd.n275 vdd.n274 63.3004
R9161 vdd.n305 vdd.n302 63.3004
R9162 vdd.n321 vdd.n320 63.3004
R9163 vdd.n351 vdd.n348 63.3004
R9164 vdd.n367 vdd.n366 63.3004
R9165 vdd.n397 vdd.n394 63.3004
R9166 vdd.n413 vdd.n412 63.3004
R9167 vdd.n494 vdd.n491 63.3004
R9168 vdd.n510 vdd.n509 63.3004
R9169 vdd.n540 vdd.n537 63.3004
R9170 vdd.n556 vdd.n555 63.3004
R9171 vdd.n6717 vdd.n6714 63.3004
R9172 vdd.n6705 vdd.n6702 63.3004
R9173 vdd.n6763 vdd.n6760 63.3004
R9174 vdd.n6751 vdd.n6748 63.3004
R9175 vdd.n6861 vdd.n6858 63.3004
R9176 vdd.n6849 vdd.n6846 63.3004
R9177 vdd.n6907 vdd.n6904 63.3004
R9178 vdd.n6895 vdd.n6892 63.3004
R9179 vdd.n6953 vdd.n6950 63.3004
R9180 vdd.n6941 vdd.n6938 63.3004
R9181 vdd.n6999 vdd.n6996 63.3004
R9182 vdd.n6987 vdd.n6984 63.3004
R9183 vdd.n7097 vdd.n7094 63.3004
R9184 vdd.n7085 vdd.n7082 63.3004
R9185 vdd.n8555 vdd.n8552 63.3004
R9186 vdd.n8543 vdd.n8540 63.3004
R9187 vdd.n7132 vdd.n7129 63.3004
R9188 vdd.n7148 vdd.n7147 63.3004
R9189 vdd.n7178 vdd.n7175 63.3004
R9190 vdd.n7194 vdd.n7193 63.3004
R9191 vdd.n7275 vdd.n7272 63.3004
R9192 vdd.n7291 vdd.n7290 63.3004
R9193 vdd.n7321 vdd.n7318 63.3004
R9194 vdd.n7337 vdd.n7336 63.3004
R9195 vdd.n7367 vdd.n7364 63.3004
R9196 vdd.n7383 vdd.n7382 63.3004
R9197 vdd.n7413 vdd.n7410 63.3004
R9198 vdd.n7429 vdd.n7428 63.3004
R9199 vdd.n7510 vdd.n7507 63.3004
R9200 vdd.n7526 vdd.n7525 63.3004
R9201 vdd.n6659 vdd.n6656 63.3004
R9202 vdd.n6675 vdd.n6674 63.3004
R9203 vdd.n7554 vdd.n7551 63.3004
R9204 vdd.n7570 vdd.n7569 63.3004
R9205 vdd.n7599 vdd.n7596 63.3004
R9206 vdd.n7615 vdd.n7614 63.3004
R9207 vdd.n7649 vdd.n7646 63.3004
R9208 vdd.n7665 vdd.n7664 63.3004
R9209 vdd.n7695 vdd.n7692 63.3004
R9210 vdd.n7711 vdd.n7710 63.3004
R9211 vdd.n7743 vdd.n7740 63.3004
R9212 vdd.n7759 vdd.n7758 63.3004
R9213 vdd.n7471 vdd.n7470 63.3004
R9214 vdd.n7790 vdd.n7787 63.3004
R9215 vdd.n7806 vdd.n7805 63.3004
R9216 vdd.n7835 vdd.n7832 63.3004
R9217 vdd.n7851 vdd.n7850 63.3004
R9218 vdd.n7881 vdd.n7878 63.3004
R9219 vdd.n7897 vdd.n7896 63.3004
R9220 vdd.n7932 vdd.n7929 63.3004
R9221 vdd.n7948 vdd.n7947 63.3004
R9222 vdd.n7978 vdd.n7975 63.3004
R9223 vdd.n7994 vdd.n7993 63.3004
R9224 vdd.n8026 vdd.n8023 63.3004
R9225 vdd.n8042 vdd.n8041 63.3004
R9226 vdd.n8072 vdd.n8069 63.3004
R9227 vdd.n8088 vdd.n8087 63.3004
R9228 vdd.n8117 vdd.n8114 63.3004
R9229 vdd.n8133 vdd.n8132 63.3004
R9230 vdd.n8167 vdd.n8164 63.3004
R9231 vdd.n8183 vdd.n8182 63.3004
R9232 vdd.n8213 vdd.n8210 63.3004
R9233 vdd.n8229 vdd.n8228 63.3004
R9234 vdd.n8261 vdd.n8258 63.3004
R9235 vdd.n8277 vdd.n8276 63.3004
R9236 vdd.n7236 vdd.n7235 63.3004
R9237 vdd.n8308 vdd.n8305 63.3004
R9238 vdd.n8324 vdd.n8323 63.3004
R9239 vdd.n8353 vdd.n8350 63.3004
R9240 vdd.n8369 vdd.n8368 63.3004
R9241 vdd.n8403 vdd.n8400 63.3004
R9242 vdd.n8419 vdd.n8418 63.3004
R9243 vdd.n8449 vdd.n8446 63.3004
R9244 vdd.n8465 vdd.n8464 63.3004
R9245 vdd.n8497 vdd.n8494 63.3004
R9246 vdd.n8513 vdd.n8512 63.3004
R9247 vdd.n8648 vdd.n8645 63.3004
R9248 vdd.n8636 vdd.n8633 63.3004
R9249 vdd.n8602 vdd.n8599 63.3004
R9250 vdd.n8590 vdd.n8587 63.3004
R9251 vdd.n8695 vdd.n8692 63.3004
R9252 vdd.n8683 vdd.n8680 63.3004
R9253 vdd.n8743 vdd.n8740 63.3004
R9254 vdd.n8731 vdd.n8728 63.3004
R9255 vdd.n8789 vdd.n8786 63.3004
R9256 vdd.n8777 vdd.n8774 63.3004
R9257 vdd.n7032 vdd.n7028 63.3004
R9258 vdd.n8931 vdd.n8928 63.3004
R9259 vdd.n8919 vdd.n8916 63.3004
R9260 vdd.n8884 vdd.n8881 63.3004
R9261 vdd.n8872 vdd.n8869 63.3004
R9262 vdd.n8838 vdd.n8835 63.3004
R9263 vdd.n8826 vdd.n8823 63.3004
R9264 vdd.n8978 vdd.n8975 63.3004
R9265 vdd.n8966 vdd.n8963 63.3004
R9266 vdd.n9026 vdd.n9023 63.3004
R9267 vdd.n9014 vdd.n9011 63.3004
R9268 vdd.n9072 vdd.n9069 63.3004
R9269 vdd.n9060 vdd.n9057 63.3004
R9270 vdd.n9166 vdd.n9163 63.3004
R9271 vdd.n9154 vdd.n9151 63.3004
R9272 vdd.n9120 vdd.n9117 63.3004
R9273 vdd.n9108 vdd.n9105 63.3004
R9274 vdd.n9213 vdd.n9210 63.3004
R9275 vdd.n9201 vdd.n9198 63.3004
R9276 vdd.n9261 vdd.n9258 63.3004
R9277 vdd.n9249 vdd.n9246 63.3004
R9278 vdd.n9307 vdd.n9304 63.3004
R9279 vdd.n9295 vdd.n9292 63.3004
R9280 vdd.n6796 vdd.n6792 63.3004
R9281 vdd.n9402 vdd.n9399 63.3004
R9282 vdd.n9390 vdd.n9387 63.3004
R9283 vdd.n9356 vdd.n9353 63.3004
R9284 vdd.n9344 vdd.n9341 63.3004
R9285 vdd.n9449 vdd.n9446 63.3004
R9286 vdd.n9437 vdd.n9434 63.3004
R9287 vdd.n9497 vdd.n9494 63.3004
R9288 vdd.n9485 vdd.n9482 63.3004
R9289 vdd.n9543 vdd.n9540 63.3004
R9290 vdd.n9531 vdd.n9528 63.3004
R9291 vdd.n3703 vdd.n3700 63.3004
R9292 vdd.n3691 vdd.n3688 63.3004
R9293 vdd.n3749 vdd.n3746 63.3004
R9294 vdd.n3737 vdd.n3734 63.3004
R9295 vdd.n3847 vdd.n3844 63.3004
R9296 vdd.n3835 vdd.n3832 63.3004
R9297 vdd.n3893 vdd.n3890 63.3004
R9298 vdd.n3881 vdd.n3878 63.3004
R9299 vdd.n3939 vdd.n3936 63.3004
R9300 vdd.n3927 vdd.n3924 63.3004
R9301 vdd.n3985 vdd.n3982 63.3004
R9302 vdd.n3973 vdd.n3970 63.3004
R9303 vdd.n4083 vdd.n4080 63.3004
R9304 vdd.n4071 vdd.n4068 63.3004
R9305 vdd.n5541 vdd.n5538 63.3004
R9306 vdd.n5529 vdd.n5526 63.3004
R9307 vdd.n4118 vdd.n4115 63.3004
R9308 vdd.n4134 vdd.n4133 63.3004
R9309 vdd.n4164 vdd.n4161 63.3004
R9310 vdd.n4180 vdd.n4179 63.3004
R9311 vdd.n4261 vdd.n4258 63.3004
R9312 vdd.n4277 vdd.n4276 63.3004
R9313 vdd.n4307 vdd.n4304 63.3004
R9314 vdd.n4323 vdd.n4322 63.3004
R9315 vdd.n4353 vdd.n4350 63.3004
R9316 vdd.n4369 vdd.n4368 63.3004
R9317 vdd.n4399 vdd.n4396 63.3004
R9318 vdd.n4415 vdd.n4414 63.3004
R9319 vdd.n4496 vdd.n4493 63.3004
R9320 vdd.n4512 vdd.n4511 63.3004
R9321 vdd.n3645 vdd.n3642 63.3004
R9322 vdd.n3661 vdd.n3660 63.3004
R9323 vdd.n4540 vdd.n4537 63.3004
R9324 vdd.n4556 vdd.n4555 63.3004
R9325 vdd.n4585 vdd.n4582 63.3004
R9326 vdd.n4601 vdd.n4600 63.3004
R9327 vdd.n4635 vdd.n4632 63.3004
R9328 vdd.n4651 vdd.n4650 63.3004
R9329 vdd.n4681 vdd.n4678 63.3004
R9330 vdd.n4697 vdd.n4696 63.3004
R9331 vdd.n4729 vdd.n4726 63.3004
R9332 vdd.n4745 vdd.n4744 63.3004
R9333 vdd.n4457 vdd.n4456 63.3004
R9334 vdd.n4776 vdd.n4773 63.3004
R9335 vdd.n4792 vdd.n4791 63.3004
R9336 vdd.n4821 vdd.n4818 63.3004
R9337 vdd.n4837 vdd.n4836 63.3004
R9338 vdd.n4867 vdd.n4864 63.3004
R9339 vdd.n4883 vdd.n4882 63.3004
R9340 vdd.n4918 vdd.n4915 63.3004
R9341 vdd.n4934 vdd.n4933 63.3004
R9342 vdd.n4964 vdd.n4961 63.3004
R9343 vdd.n4980 vdd.n4979 63.3004
R9344 vdd.n5012 vdd.n5009 63.3004
R9345 vdd.n5028 vdd.n5027 63.3004
R9346 vdd.n5058 vdd.n5055 63.3004
R9347 vdd.n5074 vdd.n5073 63.3004
R9348 vdd.n5103 vdd.n5100 63.3004
R9349 vdd.n5119 vdd.n5118 63.3004
R9350 vdd.n5153 vdd.n5150 63.3004
R9351 vdd.n5169 vdd.n5168 63.3004
R9352 vdd.n5199 vdd.n5196 63.3004
R9353 vdd.n5215 vdd.n5214 63.3004
R9354 vdd.n5247 vdd.n5244 63.3004
R9355 vdd.n5263 vdd.n5262 63.3004
R9356 vdd.n4222 vdd.n4221 63.3004
R9357 vdd.n5294 vdd.n5291 63.3004
R9358 vdd.n5310 vdd.n5309 63.3004
R9359 vdd.n5339 vdd.n5336 63.3004
R9360 vdd.n5355 vdd.n5354 63.3004
R9361 vdd.n5389 vdd.n5386 63.3004
R9362 vdd.n5405 vdd.n5404 63.3004
R9363 vdd.n5435 vdd.n5432 63.3004
R9364 vdd.n5451 vdd.n5450 63.3004
R9365 vdd.n5483 vdd.n5480 63.3004
R9366 vdd.n5499 vdd.n5498 63.3004
R9367 vdd.n5634 vdd.n5631 63.3004
R9368 vdd.n5622 vdd.n5619 63.3004
R9369 vdd.n5588 vdd.n5585 63.3004
R9370 vdd.n5576 vdd.n5573 63.3004
R9371 vdd.n5681 vdd.n5678 63.3004
R9372 vdd.n5669 vdd.n5666 63.3004
R9373 vdd.n5729 vdd.n5726 63.3004
R9374 vdd.n5717 vdd.n5714 63.3004
R9375 vdd.n5775 vdd.n5772 63.3004
R9376 vdd.n5763 vdd.n5760 63.3004
R9377 vdd.n4018 vdd.n4014 63.3004
R9378 vdd.n5917 vdd.n5914 63.3004
R9379 vdd.n5905 vdd.n5902 63.3004
R9380 vdd.n5870 vdd.n5867 63.3004
R9381 vdd.n5858 vdd.n5855 63.3004
R9382 vdd.n5824 vdd.n5821 63.3004
R9383 vdd.n5812 vdd.n5809 63.3004
R9384 vdd.n5964 vdd.n5961 63.3004
R9385 vdd.n5952 vdd.n5949 63.3004
R9386 vdd.n6012 vdd.n6009 63.3004
R9387 vdd.n6000 vdd.n5997 63.3004
R9388 vdd.n6058 vdd.n6055 63.3004
R9389 vdd.n6046 vdd.n6043 63.3004
R9390 vdd.n6152 vdd.n6149 63.3004
R9391 vdd.n6140 vdd.n6137 63.3004
R9392 vdd.n6106 vdd.n6103 63.3004
R9393 vdd.n6094 vdd.n6091 63.3004
R9394 vdd.n6199 vdd.n6196 63.3004
R9395 vdd.n6187 vdd.n6184 63.3004
R9396 vdd.n6247 vdd.n6244 63.3004
R9397 vdd.n6235 vdd.n6232 63.3004
R9398 vdd.n6293 vdd.n6290 63.3004
R9399 vdd.n6281 vdd.n6278 63.3004
R9400 vdd.n3782 vdd.n3778 63.3004
R9401 vdd.n6388 vdd.n6385 63.3004
R9402 vdd.n6376 vdd.n6373 63.3004
R9403 vdd.n6342 vdd.n6339 63.3004
R9404 vdd.n6330 vdd.n6327 63.3004
R9405 vdd.n6435 vdd.n6432 63.3004
R9406 vdd.n6423 vdd.n6420 63.3004
R9407 vdd.n6483 vdd.n6480 63.3004
R9408 vdd.n6471 vdd.n6468 63.3004
R9409 vdd.n6529 vdd.n6526 63.3004
R9410 vdd.n6517 vdd.n6514 63.3004
R9411 vdd.n689 vdd.n686 63.3004
R9412 vdd.n677 vdd.n674 63.3004
R9413 vdd.n735 vdd.n732 63.3004
R9414 vdd.n723 vdd.n720 63.3004
R9415 vdd.n833 vdd.n830 63.3004
R9416 vdd.n821 vdd.n818 63.3004
R9417 vdd.n879 vdd.n876 63.3004
R9418 vdd.n867 vdd.n864 63.3004
R9419 vdd.n925 vdd.n922 63.3004
R9420 vdd.n913 vdd.n910 63.3004
R9421 vdd.n971 vdd.n968 63.3004
R9422 vdd.n959 vdd.n956 63.3004
R9423 vdd.n1069 vdd.n1066 63.3004
R9424 vdd.n1057 vdd.n1054 63.3004
R9425 vdd.n2527 vdd.n2524 63.3004
R9426 vdd.n2515 vdd.n2512 63.3004
R9427 vdd.n1104 vdd.n1101 63.3004
R9428 vdd.n1120 vdd.n1119 63.3004
R9429 vdd.n1150 vdd.n1147 63.3004
R9430 vdd.n1166 vdd.n1165 63.3004
R9431 vdd.n1247 vdd.n1244 63.3004
R9432 vdd.n1263 vdd.n1262 63.3004
R9433 vdd.n1293 vdd.n1290 63.3004
R9434 vdd.n1309 vdd.n1308 63.3004
R9435 vdd.n1339 vdd.n1336 63.3004
R9436 vdd.n1355 vdd.n1354 63.3004
R9437 vdd.n1385 vdd.n1382 63.3004
R9438 vdd.n1401 vdd.n1400 63.3004
R9439 vdd.n1482 vdd.n1479 63.3004
R9440 vdd.n1498 vdd.n1497 63.3004
R9441 vdd.n631 vdd.n628 63.3004
R9442 vdd.n647 vdd.n646 63.3004
R9443 vdd.n1526 vdd.n1523 63.3004
R9444 vdd.n1542 vdd.n1541 63.3004
R9445 vdd.n1571 vdd.n1568 63.3004
R9446 vdd.n1587 vdd.n1586 63.3004
R9447 vdd.n1621 vdd.n1618 63.3004
R9448 vdd.n1637 vdd.n1636 63.3004
R9449 vdd.n1667 vdd.n1664 63.3004
R9450 vdd.n1683 vdd.n1682 63.3004
R9451 vdd.n1715 vdd.n1712 63.3004
R9452 vdd.n1731 vdd.n1730 63.3004
R9453 vdd.n1443 vdd.n1442 63.3004
R9454 vdd.n1762 vdd.n1759 63.3004
R9455 vdd.n1778 vdd.n1777 63.3004
R9456 vdd.n1807 vdd.n1804 63.3004
R9457 vdd.n1823 vdd.n1822 63.3004
R9458 vdd.n1853 vdd.n1850 63.3004
R9459 vdd.n1869 vdd.n1868 63.3004
R9460 vdd.n1904 vdd.n1901 63.3004
R9461 vdd.n1920 vdd.n1919 63.3004
R9462 vdd.n1950 vdd.n1947 63.3004
R9463 vdd.n1966 vdd.n1965 63.3004
R9464 vdd.n1998 vdd.n1995 63.3004
R9465 vdd.n2014 vdd.n2013 63.3004
R9466 vdd.n2044 vdd.n2041 63.3004
R9467 vdd.n2060 vdd.n2059 63.3004
R9468 vdd.n2089 vdd.n2086 63.3004
R9469 vdd.n2105 vdd.n2104 63.3004
R9470 vdd.n2139 vdd.n2136 63.3004
R9471 vdd.n2155 vdd.n2154 63.3004
R9472 vdd.n2185 vdd.n2182 63.3004
R9473 vdd.n2201 vdd.n2200 63.3004
R9474 vdd.n2233 vdd.n2230 63.3004
R9475 vdd.n2249 vdd.n2248 63.3004
R9476 vdd.n1208 vdd.n1207 63.3004
R9477 vdd.n2280 vdd.n2277 63.3004
R9478 vdd.n2296 vdd.n2295 63.3004
R9479 vdd.n2325 vdd.n2322 63.3004
R9480 vdd.n2341 vdd.n2340 63.3004
R9481 vdd.n2375 vdd.n2372 63.3004
R9482 vdd.n2391 vdd.n2390 63.3004
R9483 vdd.n2421 vdd.n2418 63.3004
R9484 vdd.n2437 vdd.n2436 63.3004
R9485 vdd.n2469 vdd.n2466 63.3004
R9486 vdd.n2485 vdd.n2484 63.3004
R9487 vdd.n2620 vdd.n2617 63.3004
R9488 vdd.n2608 vdd.n2605 63.3004
R9489 vdd.n2574 vdd.n2571 63.3004
R9490 vdd.n2562 vdd.n2559 63.3004
R9491 vdd.n2667 vdd.n2664 63.3004
R9492 vdd.n2655 vdd.n2652 63.3004
R9493 vdd.n2715 vdd.n2712 63.3004
R9494 vdd.n2703 vdd.n2700 63.3004
R9495 vdd.n2761 vdd.n2758 63.3004
R9496 vdd.n2749 vdd.n2746 63.3004
R9497 vdd.n1004 vdd.n1000 63.3004
R9498 vdd.n2903 vdd.n2900 63.3004
R9499 vdd.n2891 vdd.n2888 63.3004
R9500 vdd.n2856 vdd.n2853 63.3004
R9501 vdd.n2844 vdd.n2841 63.3004
R9502 vdd.n2810 vdd.n2807 63.3004
R9503 vdd.n2798 vdd.n2795 63.3004
R9504 vdd.n2950 vdd.n2947 63.3004
R9505 vdd.n2938 vdd.n2935 63.3004
R9506 vdd.n2998 vdd.n2995 63.3004
R9507 vdd.n2986 vdd.n2983 63.3004
R9508 vdd.n3044 vdd.n3041 63.3004
R9509 vdd.n3032 vdd.n3029 63.3004
R9510 vdd.n3138 vdd.n3135 63.3004
R9511 vdd.n3126 vdd.n3123 63.3004
R9512 vdd.n3092 vdd.n3089 63.3004
R9513 vdd.n3080 vdd.n3077 63.3004
R9514 vdd.n3185 vdd.n3182 63.3004
R9515 vdd.n3173 vdd.n3170 63.3004
R9516 vdd.n3233 vdd.n3230 63.3004
R9517 vdd.n3221 vdd.n3218 63.3004
R9518 vdd.n3279 vdd.n3276 63.3004
R9519 vdd.n3267 vdd.n3264 63.3004
R9520 vdd.n768 vdd.n764 63.3004
R9521 vdd.n3374 vdd.n3371 63.3004
R9522 vdd.n3362 vdd.n3359 63.3004
R9523 vdd.n3328 vdd.n3325 63.3004
R9524 vdd.n3316 vdd.n3313 63.3004
R9525 vdd.n3421 vdd.n3418 63.3004
R9526 vdd.n3409 vdd.n3406 63.3004
R9527 vdd.n3469 vdd.n3466 63.3004
R9528 vdd.n3457 vdd.n3454 63.3004
R9529 vdd.n3515 vdd.n3512 63.3004
R9530 vdd.n3503 vdd.n3500 63.3004
R9531 vdd.n597 vdd.n594 63.3004
R9532 vdd.n585 vdd.n582 63.3004
R9533 vdd.n3610 vdd.n3607 63.3004
R9534 vdd.n3598 vdd.n3595 63.3004
R9535 vdd.n3564 vdd.n3561 63.3004
R9536 vdd.n3552 vdd.n3549 63.3004
R9537 vdd.n6624 vdd.n6621 63.3004
R9538 vdd.n6612 vdd.n6609 63.3004
R9539 vdd.n6578 vdd.n6575 63.3004
R9540 vdd.n6566 vdd.n6563 63.3004
R9541 vdd.n9638 vdd.n9635 63.3004
R9542 vdd.n9626 vdd.n9623 63.3004
R9543 vdd.n9592 vdd.n9589 63.3004
R9544 vdd.n9580 vdd.n9577 63.3004
R9545 vdd.n9684 vdd.n9681 63.3004
R9546 vdd.n9672 vdd.n9669 63.3004
R9547 vdd.n9730 vdd.n9727 63.3004
R9548 vdd.n9718 vdd.n9715 63.3004
R9549 vdd.n9828 vdd.n9825 63.3004
R9550 vdd.n9816 vdd.n9813 63.3004
R9551 vdd.n9874 vdd.n9871 63.3004
R9552 vdd.n9862 vdd.n9859 63.3004
R9553 vdd.n9920 vdd.n9917 63.3004
R9554 vdd.n9908 vdd.n9905 63.3004
R9555 vdd.n9966 vdd.n9963 63.3004
R9556 vdd.n9954 vdd.n9951 63.3004
R9557 vdd.n10064 vdd.n10061 63.3004
R9558 vdd.n10052 vdd.n10049 63.3004
R9559 vdd.n80 vdd.n77 63.3004
R9560 vdd.n68 vdd.n65 63.3004
R9561 vdd.n34 vdd.n31 63.3004
R9562 vdd.n22 vdd.n19 63.3004
R9563 vdd.n10110 vdd.n10107 63.3004
R9564 vdd.n10098 vdd.n10095 63.3004
R9565 vdd.n10158 vdd.n10155 63.3004
R9566 vdd.n10146 vdd.n10143 63.3004
R9567 vdd.n10204 vdd.n10201 63.3004
R9568 vdd.n10192 vdd.n10189 63.3004
R9569 vdd.n9999 vdd.n9995 63.3004
R9570 vdd.n10346 vdd.n10343 63.3004
R9571 vdd.n10334 vdd.n10331 63.3004
R9572 vdd.n10299 vdd.n10296 63.3004
R9573 vdd.n10287 vdd.n10284 63.3004
R9574 vdd.n10253 vdd.n10250 63.3004
R9575 vdd.n10241 vdd.n10238 63.3004
R9576 vdd.n10393 vdd.n10390 63.3004
R9577 vdd.n10381 vdd.n10378 63.3004
R9578 vdd.n10441 vdd.n10438 63.3004
R9579 vdd.n10429 vdd.n10426 63.3004
R9580 vdd.n10487 vdd.n10484 63.3004
R9581 vdd.n10475 vdd.n10472 63.3004
R9582 vdd.n10581 vdd.n10578 63.3004
R9583 vdd.n10569 vdd.n10566 63.3004
R9584 vdd.n10535 vdd.n10532 63.3004
R9585 vdd.n10523 vdd.n10520 63.3004
R9586 vdd.n10628 vdd.n10625 63.3004
R9587 vdd.n10616 vdd.n10613 63.3004
R9588 vdd.n10676 vdd.n10673 63.3004
R9589 vdd.n10664 vdd.n10661 63.3004
R9590 vdd.n10722 vdd.n10719 63.3004
R9591 vdd.n10710 vdd.n10707 63.3004
R9592 vdd.n9763 vdd.n9759 63.3004
R9593 vdd.n10817 vdd.n10814 63.3004
R9594 vdd.n10805 vdd.n10802 63.3004
R9595 vdd.n10771 vdd.n10768 63.3004
R9596 vdd.n10759 vdd.n10756 63.3004
R9597 vdd.n10864 vdd.n10861 63.3004
R9598 vdd.n10852 vdd.n10849 63.3004
R9599 vdd.n10912 vdd.n10909 63.3004
R9600 vdd.n10900 vdd.n10897 63.3004
R9601 vdd.n10958 vdd.n10955 63.3004
R9602 vdd.n10946 vdd.n10943 63.3004
R9603 vdd.n10994 vdd.n10991 63.3004
R9604 vdd.n11010 vdd.n11009 63.3004
R9605 vdd.n11039 vdd.n11036 63.3004
R9606 vdd.n11055 vdd.n11054 63.3004
R9607 vdd.n11089 vdd.n11086 63.3004
R9608 vdd.n11105 vdd.n11104 63.3004
R9609 vdd.n11135 vdd.n11132 63.3004
R9610 vdd.n11151 vdd.n11150 63.3004
R9611 vdd.n11183 vdd.n11180 63.3004
R9612 vdd.n11199 vdd.n11198 63.3004
R9613 vdd.n455 vdd.n454 63.3004
R9614 vdd.n11230 vdd.n11227 63.3004
R9615 vdd.n11246 vdd.n11245 63.3004
R9616 vdd.n11275 vdd.n11272 63.3004
R9617 vdd.n11291 vdd.n11290 63.3004
R9618 vdd.n11321 vdd.n11318 63.3004
R9619 vdd.n11337 vdd.n11336 63.3004
R9620 vdd.n11372 vdd.n11369 63.3004
R9621 vdd.n11388 vdd.n11387 63.3004
R9622 vdd.n11418 vdd.n11415 63.3004
R9623 vdd.n11434 vdd.n11433 63.3004
R9624 vdd.n11466 vdd.n11463 63.3004
R9625 vdd.n11482 vdd.n11481 63.3004
R9626 vdd.n11512 vdd.n11509 63.3004
R9627 vdd.n11528 vdd.n11527 63.3004
R9628 vdd.n11557 vdd.n11554 63.3004
R9629 vdd.n11573 vdd.n11572 63.3004
R9630 vdd.n11607 vdd.n11604 63.3004
R9631 vdd.n11623 vdd.n11622 63.3004
R9632 vdd.n11653 vdd.n11650 63.3004
R9633 vdd.n11669 vdd.n11668 63.3004
R9634 vdd.n11701 vdd.n11698 63.3004
R9635 vdd.n11717 vdd.n11716 63.3004
R9636 vdd.n220 vdd.n219 63.3004
R9637 vdd.n11748 vdd.n11745 63.3004
R9638 vdd.n11764 vdd.n11763 63.3004
R9639 vdd.n11793 vdd.n11790 63.3004
R9640 vdd.n11809 vdd.n11808 63.3004
R9641 vdd.n11843 vdd.n11840 63.3004
R9642 vdd.n11859 vdd.n11858 63.3004
R9643 vdd.n11889 vdd.n11886 63.3004
R9644 vdd.n11905 vdd.n11904 63.3004
R9645 vdd.n11937 vdd.n11934 63.3004
R9646 vdd.n11953 vdd.n11952 63.3004
R9647 vdd.n7483 vdd.n7438 50.8372
R9648 vdd.n7248 vdd.n7203 50.8372
R9649 vdd.n7058 vdd.n7057 50.8372
R9650 vdd.n6822 vdd.n6821 50.8372
R9651 vdd.n4469 vdd.n4424 50.8372
R9652 vdd.n4234 vdd.n4189 50.8372
R9653 vdd.n4044 vdd.n4043 50.8372
R9654 vdd.n3808 vdd.n3807 50.8372
R9655 vdd.n1455 vdd.n1410 50.8372
R9656 vdd.n1220 vdd.n1175 50.8372
R9657 vdd.n1030 vdd.n1029 50.8372
R9658 vdd.n794 vdd.n793 50.8372
R9659 vdd.n10025 vdd.n10024 50.8372
R9660 vdd.n9789 vdd.n9788 50.8372
R9661 vdd.n467 vdd.n422 50.8372
R9662 vdd.n232 vdd.n187 50.8372
R9663 vdd.n11980 vdd.n11979 35.2919
R9664 vdd.n12000 vdd.n11998 35.2919
R9665 vdd.n12000 vdd.n11999 35.2919
R9666 vdd.n112 vdd.n103 35.2919
R9667 vdd.n121 vdd.n103 35.2919
R9668 vdd.n122 vdd.n121 35.2919
R9669 vdd.n125 vdd.n122 35.2919
R9670 vdd.n125 vdd.n124 35.2919
R9671 vdd.n124 vdd.n101 35.2919
R9672 vdd.n158 vdd.n149 35.2919
R9673 vdd.n167 vdd.n149 35.2919
R9674 vdd.n168 vdd.n167 35.2919
R9675 vdd.n171 vdd.n168 35.2919
R9676 vdd.n171 vdd.n170 35.2919
R9677 vdd.n170 vdd.n147 35.2919
R9678 vdd.n255 vdd.n246 35.2919
R9679 vdd.n264 vdd.n246 35.2919
R9680 vdd.n265 vdd.n264 35.2919
R9681 vdd.n268 vdd.n265 35.2919
R9682 vdd.n268 vdd.n267 35.2919
R9683 vdd.n267 vdd.n244 35.2919
R9684 vdd.n301 vdd.n292 35.2919
R9685 vdd.n310 vdd.n292 35.2919
R9686 vdd.n311 vdd.n310 35.2919
R9687 vdd.n314 vdd.n311 35.2919
R9688 vdd.n314 vdd.n313 35.2919
R9689 vdd.n313 vdd.n290 35.2919
R9690 vdd.n347 vdd.n338 35.2919
R9691 vdd.n356 vdd.n338 35.2919
R9692 vdd.n357 vdd.n356 35.2919
R9693 vdd.n360 vdd.n357 35.2919
R9694 vdd.n360 vdd.n359 35.2919
R9695 vdd.n359 vdd.n336 35.2919
R9696 vdd.n393 vdd.n384 35.2919
R9697 vdd.n402 vdd.n384 35.2919
R9698 vdd.n403 vdd.n402 35.2919
R9699 vdd.n406 vdd.n403 35.2919
R9700 vdd.n406 vdd.n405 35.2919
R9701 vdd.n405 vdd.n382 35.2919
R9702 vdd.n490 vdd.n481 35.2919
R9703 vdd.n499 vdd.n481 35.2919
R9704 vdd.n500 vdd.n499 35.2919
R9705 vdd.n503 vdd.n500 35.2919
R9706 vdd.n503 vdd.n502 35.2919
R9707 vdd.n502 vdd.n479 35.2919
R9708 vdd.n536 vdd.n527 35.2919
R9709 vdd.n545 vdd.n527 35.2919
R9710 vdd.n546 vdd.n545 35.2919
R9711 vdd.n549 vdd.n546 35.2919
R9712 vdd.n549 vdd.n548 35.2919
R9713 vdd.n548 vdd.n525 35.2919
R9714 vdd.n6699 vdd.n6692 35.2919
R9715 vdd.n6710 vdd.n6692 35.2919
R9716 vdd.n6711 vdd.n6710 35.2919
R9717 vdd.n6712 vdd.n6711 35.2919
R9718 vdd.n6713 vdd.n6712 35.2919
R9719 vdd.n6718 vdd.n6713 35.2919
R9720 vdd.n6745 vdd.n6738 35.2919
R9721 vdd.n6756 vdd.n6738 35.2919
R9722 vdd.n6757 vdd.n6756 35.2919
R9723 vdd.n6758 vdd.n6757 35.2919
R9724 vdd.n6759 vdd.n6758 35.2919
R9725 vdd.n6764 vdd.n6759 35.2919
R9726 vdd.n6843 vdd.n6836 35.2919
R9727 vdd.n6854 vdd.n6836 35.2919
R9728 vdd.n6855 vdd.n6854 35.2919
R9729 vdd.n6856 vdd.n6855 35.2919
R9730 vdd.n6857 vdd.n6856 35.2919
R9731 vdd.n6862 vdd.n6857 35.2919
R9732 vdd.n6889 vdd.n6882 35.2919
R9733 vdd.n6900 vdd.n6882 35.2919
R9734 vdd.n6901 vdd.n6900 35.2919
R9735 vdd.n6902 vdd.n6901 35.2919
R9736 vdd.n6903 vdd.n6902 35.2919
R9737 vdd.n6908 vdd.n6903 35.2919
R9738 vdd.n6935 vdd.n6928 35.2919
R9739 vdd.n6946 vdd.n6928 35.2919
R9740 vdd.n6947 vdd.n6946 35.2919
R9741 vdd.n6948 vdd.n6947 35.2919
R9742 vdd.n6949 vdd.n6948 35.2919
R9743 vdd.n6954 vdd.n6949 35.2919
R9744 vdd.n6981 vdd.n6974 35.2919
R9745 vdd.n6992 vdd.n6974 35.2919
R9746 vdd.n6993 vdd.n6992 35.2919
R9747 vdd.n6994 vdd.n6993 35.2919
R9748 vdd.n6995 vdd.n6994 35.2919
R9749 vdd.n7000 vdd.n6995 35.2919
R9750 vdd.n7079 vdd.n7072 35.2919
R9751 vdd.n7090 vdd.n7072 35.2919
R9752 vdd.n7091 vdd.n7090 35.2919
R9753 vdd.n7092 vdd.n7091 35.2919
R9754 vdd.n7093 vdd.n7092 35.2919
R9755 vdd.n7098 vdd.n7093 35.2919
R9756 vdd.n8537 vdd.n8530 35.2919
R9757 vdd.n8548 vdd.n8530 35.2919
R9758 vdd.n8549 vdd.n8548 35.2919
R9759 vdd.n8550 vdd.n8549 35.2919
R9760 vdd.n8551 vdd.n8550 35.2919
R9761 vdd.n8556 vdd.n8551 35.2919
R9762 vdd.n7128 vdd.n7119 35.2919
R9763 vdd.n7137 vdd.n7119 35.2919
R9764 vdd.n7138 vdd.n7137 35.2919
R9765 vdd.n7141 vdd.n7138 35.2919
R9766 vdd.n7141 vdd.n7140 35.2919
R9767 vdd.n7140 vdd.n7117 35.2919
R9768 vdd.n7174 vdd.n7165 35.2919
R9769 vdd.n7183 vdd.n7165 35.2919
R9770 vdd.n7184 vdd.n7183 35.2919
R9771 vdd.n7187 vdd.n7184 35.2919
R9772 vdd.n7187 vdd.n7186 35.2919
R9773 vdd.n7186 vdd.n7163 35.2919
R9774 vdd.n7271 vdd.n7262 35.2919
R9775 vdd.n7280 vdd.n7262 35.2919
R9776 vdd.n7281 vdd.n7280 35.2919
R9777 vdd.n7284 vdd.n7281 35.2919
R9778 vdd.n7284 vdd.n7283 35.2919
R9779 vdd.n7283 vdd.n7260 35.2919
R9780 vdd.n7317 vdd.n7308 35.2919
R9781 vdd.n7326 vdd.n7308 35.2919
R9782 vdd.n7327 vdd.n7326 35.2919
R9783 vdd.n7330 vdd.n7327 35.2919
R9784 vdd.n7330 vdd.n7329 35.2919
R9785 vdd.n7329 vdd.n7306 35.2919
R9786 vdd.n7363 vdd.n7354 35.2919
R9787 vdd.n7372 vdd.n7354 35.2919
R9788 vdd.n7373 vdd.n7372 35.2919
R9789 vdd.n7376 vdd.n7373 35.2919
R9790 vdd.n7376 vdd.n7375 35.2919
R9791 vdd.n7375 vdd.n7352 35.2919
R9792 vdd.n7409 vdd.n7400 35.2919
R9793 vdd.n7418 vdd.n7400 35.2919
R9794 vdd.n7419 vdd.n7418 35.2919
R9795 vdd.n7422 vdd.n7419 35.2919
R9796 vdd.n7422 vdd.n7421 35.2919
R9797 vdd.n7421 vdd.n7398 35.2919
R9798 vdd.n7506 vdd.n7497 35.2919
R9799 vdd.n7515 vdd.n7497 35.2919
R9800 vdd.n7516 vdd.n7515 35.2919
R9801 vdd.n7519 vdd.n7516 35.2919
R9802 vdd.n7519 vdd.n7518 35.2919
R9803 vdd.n7518 vdd.n7495 35.2919
R9804 vdd.n6655 vdd.n6646 35.2919
R9805 vdd.n6664 vdd.n6646 35.2919
R9806 vdd.n6665 vdd.n6664 35.2919
R9807 vdd.n6668 vdd.n6665 35.2919
R9808 vdd.n6668 vdd.n6667 35.2919
R9809 vdd.n6667 vdd.n6644 35.2919
R9810 vdd.n7550 vdd.n7541 35.2919
R9811 vdd.n7559 vdd.n7541 35.2919
R9812 vdd.n7560 vdd.n7559 35.2919
R9813 vdd.n7563 vdd.n7560 35.2919
R9814 vdd.n7563 vdd.n7562 35.2919
R9815 vdd.n7562 vdd.n7539 35.2919
R9816 vdd.n7595 vdd.n7586 35.2919
R9817 vdd.n7604 vdd.n7586 35.2919
R9818 vdd.n7605 vdd.n7604 35.2919
R9819 vdd.n7608 vdd.n7605 35.2919
R9820 vdd.n7608 vdd.n7607 35.2919
R9821 vdd.n7607 vdd.n7584 35.2919
R9822 vdd.n7645 vdd.n7636 35.2919
R9823 vdd.n7654 vdd.n7636 35.2919
R9824 vdd.n7655 vdd.n7654 35.2919
R9825 vdd.n7658 vdd.n7655 35.2919
R9826 vdd.n7658 vdd.n7657 35.2919
R9827 vdd.n7657 vdd.n7634 35.2919
R9828 vdd.n7691 vdd.n7682 35.2919
R9829 vdd.n7700 vdd.n7682 35.2919
R9830 vdd.n7701 vdd.n7700 35.2919
R9831 vdd.n7704 vdd.n7701 35.2919
R9832 vdd.n7704 vdd.n7703 35.2919
R9833 vdd.n7703 vdd.n7680 35.2919
R9834 vdd.n7739 vdd.n7730 35.2919
R9835 vdd.n7748 vdd.n7730 35.2919
R9836 vdd.n7749 vdd.n7748 35.2919
R9837 vdd.n7752 vdd.n7749 35.2919
R9838 vdd.n7752 vdd.n7751 35.2919
R9839 vdd.n7751 vdd.n7728 35.2919
R9840 vdd.n7456 vdd.n7454 35.2919
R9841 vdd.n7460 vdd.n7454 35.2919
R9842 vdd.n7461 vdd.n7460 35.2919
R9843 vdd.n7464 vdd.n7461 35.2919
R9844 vdd.n7464 vdd.n7463 35.2919
R9845 vdd.n7463 vdd.n7449 35.2919
R9846 vdd.n7786 vdd.n7777 35.2919
R9847 vdd.n7795 vdd.n7777 35.2919
R9848 vdd.n7796 vdd.n7795 35.2919
R9849 vdd.n7799 vdd.n7796 35.2919
R9850 vdd.n7799 vdd.n7798 35.2919
R9851 vdd.n7798 vdd.n7775 35.2919
R9852 vdd.n7831 vdd.n7822 35.2919
R9853 vdd.n7840 vdd.n7822 35.2919
R9854 vdd.n7841 vdd.n7840 35.2919
R9855 vdd.n7844 vdd.n7841 35.2919
R9856 vdd.n7844 vdd.n7843 35.2919
R9857 vdd.n7843 vdd.n7820 35.2919
R9858 vdd.n7877 vdd.n7868 35.2919
R9859 vdd.n7886 vdd.n7868 35.2919
R9860 vdd.n7887 vdd.n7886 35.2919
R9861 vdd.n7890 vdd.n7887 35.2919
R9862 vdd.n7890 vdd.n7889 35.2919
R9863 vdd.n7889 vdd.n7866 35.2919
R9864 vdd.n7928 vdd.n7919 35.2919
R9865 vdd.n7937 vdd.n7919 35.2919
R9866 vdd.n7938 vdd.n7937 35.2919
R9867 vdd.n7941 vdd.n7938 35.2919
R9868 vdd.n7941 vdd.n7940 35.2919
R9869 vdd.n7940 vdd.n7917 35.2919
R9870 vdd.n7974 vdd.n7965 35.2919
R9871 vdd.n7983 vdd.n7965 35.2919
R9872 vdd.n7984 vdd.n7983 35.2919
R9873 vdd.n7987 vdd.n7984 35.2919
R9874 vdd.n7987 vdd.n7986 35.2919
R9875 vdd.n7986 vdd.n7963 35.2919
R9876 vdd.n8022 vdd.n8013 35.2919
R9877 vdd.n8031 vdd.n8013 35.2919
R9878 vdd.n8032 vdd.n8031 35.2919
R9879 vdd.n8035 vdd.n8032 35.2919
R9880 vdd.n8035 vdd.n8034 35.2919
R9881 vdd.n8034 vdd.n8011 35.2919
R9882 vdd.n8068 vdd.n8059 35.2919
R9883 vdd.n8077 vdd.n8059 35.2919
R9884 vdd.n8078 vdd.n8077 35.2919
R9885 vdd.n8081 vdd.n8078 35.2919
R9886 vdd.n8081 vdd.n8080 35.2919
R9887 vdd.n8080 vdd.n8057 35.2919
R9888 vdd.n8113 vdd.n8104 35.2919
R9889 vdd.n8122 vdd.n8104 35.2919
R9890 vdd.n8123 vdd.n8122 35.2919
R9891 vdd.n8126 vdd.n8123 35.2919
R9892 vdd.n8126 vdd.n8125 35.2919
R9893 vdd.n8125 vdd.n8102 35.2919
R9894 vdd.n8163 vdd.n8154 35.2919
R9895 vdd.n8172 vdd.n8154 35.2919
R9896 vdd.n8173 vdd.n8172 35.2919
R9897 vdd.n8176 vdd.n8173 35.2919
R9898 vdd.n8176 vdd.n8175 35.2919
R9899 vdd.n8175 vdd.n8152 35.2919
R9900 vdd.n8209 vdd.n8200 35.2919
R9901 vdd.n8218 vdd.n8200 35.2919
R9902 vdd.n8219 vdd.n8218 35.2919
R9903 vdd.n8222 vdd.n8219 35.2919
R9904 vdd.n8222 vdd.n8221 35.2919
R9905 vdd.n8221 vdd.n8198 35.2919
R9906 vdd.n8257 vdd.n8248 35.2919
R9907 vdd.n8266 vdd.n8248 35.2919
R9908 vdd.n8267 vdd.n8266 35.2919
R9909 vdd.n8270 vdd.n8267 35.2919
R9910 vdd.n8270 vdd.n8269 35.2919
R9911 vdd.n8269 vdd.n8246 35.2919
R9912 vdd.n7221 vdd.n7219 35.2919
R9913 vdd.n7225 vdd.n7219 35.2919
R9914 vdd.n7226 vdd.n7225 35.2919
R9915 vdd.n7229 vdd.n7226 35.2919
R9916 vdd.n7229 vdd.n7228 35.2919
R9917 vdd.n7228 vdd.n7214 35.2919
R9918 vdd.n8304 vdd.n8295 35.2919
R9919 vdd.n8313 vdd.n8295 35.2919
R9920 vdd.n8314 vdd.n8313 35.2919
R9921 vdd.n8317 vdd.n8314 35.2919
R9922 vdd.n8317 vdd.n8316 35.2919
R9923 vdd.n8316 vdd.n8293 35.2919
R9924 vdd.n8349 vdd.n8340 35.2919
R9925 vdd.n8358 vdd.n8340 35.2919
R9926 vdd.n8359 vdd.n8358 35.2919
R9927 vdd.n8362 vdd.n8359 35.2919
R9928 vdd.n8362 vdd.n8361 35.2919
R9929 vdd.n8361 vdd.n8338 35.2919
R9930 vdd.n8399 vdd.n8390 35.2919
R9931 vdd.n8408 vdd.n8390 35.2919
R9932 vdd.n8409 vdd.n8408 35.2919
R9933 vdd.n8412 vdd.n8409 35.2919
R9934 vdd.n8412 vdd.n8411 35.2919
R9935 vdd.n8411 vdd.n8388 35.2919
R9936 vdd.n8445 vdd.n8436 35.2919
R9937 vdd.n8454 vdd.n8436 35.2919
R9938 vdd.n8455 vdd.n8454 35.2919
R9939 vdd.n8458 vdd.n8455 35.2919
R9940 vdd.n8458 vdd.n8457 35.2919
R9941 vdd.n8457 vdd.n8434 35.2919
R9942 vdd.n8493 vdd.n8484 35.2919
R9943 vdd.n8502 vdd.n8484 35.2919
R9944 vdd.n8503 vdd.n8502 35.2919
R9945 vdd.n8506 vdd.n8503 35.2919
R9946 vdd.n8506 vdd.n8505 35.2919
R9947 vdd.n8505 vdd.n8482 35.2919
R9948 vdd.n8630 vdd.n8623 35.2919
R9949 vdd.n8641 vdd.n8623 35.2919
R9950 vdd.n8642 vdd.n8641 35.2919
R9951 vdd.n8643 vdd.n8642 35.2919
R9952 vdd.n8644 vdd.n8643 35.2919
R9953 vdd.n8649 vdd.n8644 35.2919
R9954 vdd.n8584 vdd.n8577 35.2919
R9955 vdd.n8595 vdd.n8577 35.2919
R9956 vdd.n8596 vdd.n8595 35.2919
R9957 vdd.n8597 vdd.n8596 35.2919
R9958 vdd.n8598 vdd.n8597 35.2919
R9959 vdd.n8603 vdd.n8598 35.2919
R9960 vdd.n8677 vdd.n8670 35.2919
R9961 vdd.n8688 vdd.n8670 35.2919
R9962 vdd.n8689 vdd.n8688 35.2919
R9963 vdd.n8690 vdd.n8689 35.2919
R9964 vdd.n8691 vdd.n8690 35.2919
R9965 vdd.n8696 vdd.n8691 35.2919
R9966 vdd.n8725 vdd.n8718 35.2919
R9967 vdd.n8736 vdd.n8718 35.2919
R9968 vdd.n8737 vdd.n8736 35.2919
R9969 vdd.n8738 vdd.n8737 35.2919
R9970 vdd.n8739 vdd.n8738 35.2919
R9971 vdd.n8744 vdd.n8739 35.2919
R9972 vdd.n8771 vdd.n8764 35.2919
R9973 vdd.n8782 vdd.n8764 35.2919
R9974 vdd.n8783 vdd.n8782 35.2919
R9975 vdd.n8784 vdd.n8783 35.2919
R9976 vdd.n8785 vdd.n8784 35.2919
R9977 vdd.n8790 vdd.n8785 35.2919
R9978 vdd.n7037 vdd.n7036 35.2919
R9979 vdd.n7038 vdd.n7037 35.2919
R9980 vdd.n7039 vdd.n7038 35.2919
R9981 vdd.n7040 vdd.n7039 35.2919
R9982 vdd.n7040 vdd.n7015 35.2919
R9983 vdd.n7056 vdd.n7015 35.2919
R9984 vdd.n8913 vdd.n8906 35.2919
R9985 vdd.n8924 vdd.n8906 35.2919
R9986 vdd.n8925 vdd.n8924 35.2919
R9987 vdd.n8926 vdd.n8925 35.2919
R9988 vdd.n8927 vdd.n8926 35.2919
R9989 vdd.n8932 vdd.n8927 35.2919
R9990 vdd.n8866 vdd.n8859 35.2919
R9991 vdd.n8877 vdd.n8859 35.2919
R9992 vdd.n8878 vdd.n8877 35.2919
R9993 vdd.n8879 vdd.n8878 35.2919
R9994 vdd.n8880 vdd.n8879 35.2919
R9995 vdd.n8885 vdd.n8880 35.2919
R9996 vdd.n8820 vdd.n8813 35.2919
R9997 vdd.n8831 vdd.n8813 35.2919
R9998 vdd.n8832 vdd.n8831 35.2919
R9999 vdd.n8833 vdd.n8832 35.2919
R10000 vdd.n8834 vdd.n8833 35.2919
R10001 vdd.n8839 vdd.n8834 35.2919
R10002 vdd.n8960 vdd.n8953 35.2919
R10003 vdd.n8971 vdd.n8953 35.2919
R10004 vdd.n8972 vdd.n8971 35.2919
R10005 vdd.n8973 vdd.n8972 35.2919
R10006 vdd.n8974 vdd.n8973 35.2919
R10007 vdd.n8979 vdd.n8974 35.2919
R10008 vdd.n9008 vdd.n9001 35.2919
R10009 vdd.n9019 vdd.n9001 35.2919
R10010 vdd.n9020 vdd.n9019 35.2919
R10011 vdd.n9021 vdd.n9020 35.2919
R10012 vdd.n9022 vdd.n9021 35.2919
R10013 vdd.n9027 vdd.n9022 35.2919
R10014 vdd.n9054 vdd.n9047 35.2919
R10015 vdd.n9065 vdd.n9047 35.2919
R10016 vdd.n9066 vdd.n9065 35.2919
R10017 vdd.n9067 vdd.n9066 35.2919
R10018 vdd.n9068 vdd.n9067 35.2919
R10019 vdd.n9073 vdd.n9068 35.2919
R10020 vdd.n9148 vdd.n9141 35.2919
R10021 vdd.n9159 vdd.n9141 35.2919
R10022 vdd.n9160 vdd.n9159 35.2919
R10023 vdd.n9161 vdd.n9160 35.2919
R10024 vdd.n9162 vdd.n9161 35.2919
R10025 vdd.n9167 vdd.n9162 35.2919
R10026 vdd.n9102 vdd.n9095 35.2919
R10027 vdd.n9113 vdd.n9095 35.2919
R10028 vdd.n9114 vdd.n9113 35.2919
R10029 vdd.n9115 vdd.n9114 35.2919
R10030 vdd.n9116 vdd.n9115 35.2919
R10031 vdd.n9121 vdd.n9116 35.2919
R10032 vdd.n9195 vdd.n9188 35.2919
R10033 vdd.n9206 vdd.n9188 35.2919
R10034 vdd.n9207 vdd.n9206 35.2919
R10035 vdd.n9208 vdd.n9207 35.2919
R10036 vdd.n9209 vdd.n9208 35.2919
R10037 vdd.n9214 vdd.n9209 35.2919
R10038 vdd.n9243 vdd.n9236 35.2919
R10039 vdd.n9254 vdd.n9236 35.2919
R10040 vdd.n9255 vdd.n9254 35.2919
R10041 vdd.n9256 vdd.n9255 35.2919
R10042 vdd.n9257 vdd.n9256 35.2919
R10043 vdd.n9262 vdd.n9257 35.2919
R10044 vdd.n9289 vdd.n9282 35.2919
R10045 vdd.n9300 vdd.n9282 35.2919
R10046 vdd.n9301 vdd.n9300 35.2919
R10047 vdd.n9302 vdd.n9301 35.2919
R10048 vdd.n9303 vdd.n9302 35.2919
R10049 vdd.n9308 vdd.n9303 35.2919
R10050 vdd.n6801 vdd.n6800 35.2919
R10051 vdd.n6802 vdd.n6801 35.2919
R10052 vdd.n6803 vdd.n6802 35.2919
R10053 vdd.n6804 vdd.n6803 35.2919
R10054 vdd.n6804 vdd.n6779 35.2919
R10055 vdd.n6820 vdd.n6779 35.2919
R10056 vdd.n9384 vdd.n9377 35.2919
R10057 vdd.n9395 vdd.n9377 35.2919
R10058 vdd.n9396 vdd.n9395 35.2919
R10059 vdd.n9397 vdd.n9396 35.2919
R10060 vdd.n9398 vdd.n9397 35.2919
R10061 vdd.n9403 vdd.n9398 35.2919
R10062 vdd.n9338 vdd.n9331 35.2919
R10063 vdd.n9349 vdd.n9331 35.2919
R10064 vdd.n9350 vdd.n9349 35.2919
R10065 vdd.n9351 vdd.n9350 35.2919
R10066 vdd.n9352 vdd.n9351 35.2919
R10067 vdd.n9357 vdd.n9352 35.2919
R10068 vdd.n9431 vdd.n9424 35.2919
R10069 vdd.n9442 vdd.n9424 35.2919
R10070 vdd.n9443 vdd.n9442 35.2919
R10071 vdd.n9444 vdd.n9443 35.2919
R10072 vdd.n9445 vdd.n9444 35.2919
R10073 vdd.n9450 vdd.n9445 35.2919
R10074 vdd.n9479 vdd.n9472 35.2919
R10075 vdd.n9490 vdd.n9472 35.2919
R10076 vdd.n9491 vdd.n9490 35.2919
R10077 vdd.n9492 vdd.n9491 35.2919
R10078 vdd.n9493 vdd.n9492 35.2919
R10079 vdd.n9498 vdd.n9493 35.2919
R10080 vdd.n9525 vdd.n9518 35.2919
R10081 vdd.n9536 vdd.n9518 35.2919
R10082 vdd.n9537 vdd.n9536 35.2919
R10083 vdd.n9538 vdd.n9537 35.2919
R10084 vdd.n9539 vdd.n9538 35.2919
R10085 vdd.n9544 vdd.n9539 35.2919
R10086 vdd.n3685 vdd.n3678 35.2919
R10087 vdd.n3696 vdd.n3678 35.2919
R10088 vdd.n3697 vdd.n3696 35.2919
R10089 vdd.n3698 vdd.n3697 35.2919
R10090 vdd.n3699 vdd.n3698 35.2919
R10091 vdd.n3704 vdd.n3699 35.2919
R10092 vdd.n3731 vdd.n3724 35.2919
R10093 vdd.n3742 vdd.n3724 35.2919
R10094 vdd.n3743 vdd.n3742 35.2919
R10095 vdd.n3744 vdd.n3743 35.2919
R10096 vdd.n3745 vdd.n3744 35.2919
R10097 vdd.n3750 vdd.n3745 35.2919
R10098 vdd.n3829 vdd.n3822 35.2919
R10099 vdd.n3840 vdd.n3822 35.2919
R10100 vdd.n3841 vdd.n3840 35.2919
R10101 vdd.n3842 vdd.n3841 35.2919
R10102 vdd.n3843 vdd.n3842 35.2919
R10103 vdd.n3848 vdd.n3843 35.2919
R10104 vdd.n3875 vdd.n3868 35.2919
R10105 vdd.n3886 vdd.n3868 35.2919
R10106 vdd.n3887 vdd.n3886 35.2919
R10107 vdd.n3888 vdd.n3887 35.2919
R10108 vdd.n3889 vdd.n3888 35.2919
R10109 vdd.n3894 vdd.n3889 35.2919
R10110 vdd.n3921 vdd.n3914 35.2919
R10111 vdd.n3932 vdd.n3914 35.2919
R10112 vdd.n3933 vdd.n3932 35.2919
R10113 vdd.n3934 vdd.n3933 35.2919
R10114 vdd.n3935 vdd.n3934 35.2919
R10115 vdd.n3940 vdd.n3935 35.2919
R10116 vdd.n3967 vdd.n3960 35.2919
R10117 vdd.n3978 vdd.n3960 35.2919
R10118 vdd.n3979 vdd.n3978 35.2919
R10119 vdd.n3980 vdd.n3979 35.2919
R10120 vdd.n3981 vdd.n3980 35.2919
R10121 vdd.n3986 vdd.n3981 35.2919
R10122 vdd.n4065 vdd.n4058 35.2919
R10123 vdd.n4076 vdd.n4058 35.2919
R10124 vdd.n4077 vdd.n4076 35.2919
R10125 vdd.n4078 vdd.n4077 35.2919
R10126 vdd.n4079 vdd.n4078 35.2919
R10127 vdd.n4084 vdd.n4079 35.2919
R10128 vdd.n5523 vdd.n5516 35.2919
R10129 vdd.n5534 vdd.n5516 35.2919
R10130 vdd.n5535 vdd.n5534 35.2919
R10131 vdd.n5536 vdd.n5535 35.2919
R10132 vdd.n5537 vdd.n5536 35.2919
R10133 vdd.n5542 vdd.n5537 35.2919
R10134 vdd.n4114 vdd.n4105 35.2919
R10135 vdd.n4123 vdd.n4105 35.2919
R10136 vdd.n4124 vdd.n4123 35.2919
R10137 vdd.n4127 vdd.n4124 35.2919
R10138 vdd.n4127 vdd.n4126 35.2919
R10139 vdd.n4126 vdd.n4103 35.2919
R10140 vdd.n4160 vdd.n4151 35.2919
R10141 vdd.n4169 vdd.n4151 35.2919
R10142 vdd.n4170 vdd.n4169 35.2919
R10143 vdd.n4173 vdd.n4170 35.2919
R10144 vdd.n4173 vdd.n4172 35.2919
R10145 vdd.n4172 vdd.n4149 35.2919
R10146 vdd.n4257 vdd.n4248 35.2919
R10147 vdd.n4266 vdd.n4248 35.2919
R10148 vdd.n4267 vdd.n4266 35.2919
R10149 vdd.n4270 vdd.n4267 35.2919
R10150 vdd.n4270 vdd.n4269 35.2919
R10151 vdd.n4269 vdd.n4246 35.2919
R10152 vdd.n4303 vdd.n4294 35.2919
R10153 vdd.n4312 vdd.n4294 35.2919
R10154 vdd.n4313 vdd.n4312 35.2919
R10155 vdd.n4316 vdd.n4313 35.2919
R10156 vdd.n4316 vdd.n4315 35.2919
R10157 vdd.n4315 vdd.n4292 35.2919
R10158 vdd.n4349 vdd.n4340 35.2919
R10159 vdd.n4358 vdd.n4340 35.2919
R10160 vdd.n4359 vdd.n4358 35.2919
R10161 vdd.n4362 vdd.n4359 35.2919
R10162 vdd.n4362 vdd.n4361 35.2919
R10163 vdd.n4361 vdd.n4338 35.2919
R10164 vdd.n4395 vdd.n4386 35.2919
R10165 vdd.n4404 vdd.n4386 35.2919
R10166 vdd.n4405 vdd.n4404 35.2919
R10167 vdd.n4408 vdd.n4405 35.2919
R10168 vdd.n4408 vdd.n4407 35.2919
R10169 vdd.n4407 vdd.n4384 35.2919
R10170 vdd.n4492 vdd.n4483 35.2919
R10171 vdd.n4501 vdd.n4483 35.2919
R10172 vdd.n4502 vdd.n4501 35.2919
R10173 vdd.n4505 vdd.n4502 35.2919
R10174 vdd.n4505 vdd.n4504 35.2919
R10175 vdd.n4504 vdd.n4481 35.2919
R10176 vdd.n3641 vdd.n3632 35.2919
R10177 vdd.n3650 vdd.n3632 35.2919
R10178 vdd.n3651 vdd.n3650 35.2919
R10179 vdd.n3654 vdd.n3651 35.2919
R10180 vdd.n3654 vdd.n3653 35.2919
R10181 vdd.n3653 vdd.n3630 35.2919
R10182 vdd.n4536 vdd.n4527 35.2919
R10183 vdd.n4545 vdd.n4527 35.2919
R10184 vdd.n4546 vdd.n4545 35.2919
R10185 vdd.n4549 vdd.n4546 35.2919
R10186 vdd.n4549 vdd.n4548 35.2919
R10187 vdd.n4548 vdd.n4525 35.2919
R10188 vdd.n4581 vdd.n4572 35.2919
R10189 vdd.n4590 vdd.n4572 35.2919
R10190 vdd.n4591 vdd.n4590 35.2919
R10191 vdd.n4594 vdd.n4591 35.2919
R10192 vdd.n4594 vdd.n4593 35.2919
R10193 vdd.n4593 vdd.n4570 35.2919
R10194 vdd.n4631 vdd.n4622 35.2919
R10195 vdd.n4640 vdd.n4622 35.2919
R10196 vdd.n4641 vdd.n4640 35.2919
R10197 vdd.n4644 vdd.n4641 35.2919
R10198 vdd.n4644 vdd.n4643 35.2919
R10199 vdd.n4643 vdd.n4620 35.2919
R10200 vdd.n4677 vdd.n4668 35.2919
R10201 vdd.n4686 vdd.n4668 35.2919
R10202 vdd.n4687 vdd.n4686 35.2919
R10203 vdd.n4690 vdd.n4687 35.2919
R10204 vdd.n4690 vdd.n4689 35.2919
R10205 vdd.n4689 vdd.n4666 35.2919
R10206 vdd.n4725 vdd.n4716 35.2919
R10207 vdd.n4734 vdd.n4716 35.2919
R10208 vdd.n4735 vdd.n4734 35.2919
R10209 vdd.n4738 vdd.n4735 35.2919
R10210 vdd.n4738 vdd.n4737 35.2919
R10211 vdd.n4737 vdd.n4714 35.2919
R10212 vdd.n4442 vdd.n4440 35.2919
R10213 vdd.n4446 vdd.n4440 35.2919
R10214 vdd.n4447 vdd.n4446 35.2919
R10215 vdd.n4450 vdd.n4447 35.2919
R10216 vdd.n4450 vdd.n4449 35.2919
R10217 vdd.n4449 vdd.n4435 35.2919
R10218 vdd.n4772 vdd.n4763 35.2919
R10219 vdd.n4781 vdd.n4763 35.2919
R10220 vdd.n4782 vdd.n4781 35.2919
R10221 vdd.n4785 vdd.n4782 35.2919
R10222 vdd.n4785 vdd.n4784 35.2919
R10223 vdd.n4784 vdd.n4761 35.2919
R10224 vdd.n4817 vdd.n4808 35.2919
R10225 vdd.n4826 vdd.n4808 35.2919
R10226 vdd.n4827 vdd.n4826 35.2919
R10227 vdd.n4830 vdd.n4827 35.2919
R10228 vdd.n4830 vdd.n4829 35.2919
R10229 vdd.n4829 vdd.n4806 35.2919
R10230 vdd.n4863 vdd.n4854 35.2919
R10231 vdd.n4872 vdd.n4854 35.2919
R10232 vdd.n4873 vdd.n4872 35.2919
R10233 vdd.n4876 vdd.n4873 35.2919
R10234 vdd.n4876 vdd.n4875 35.2919
R10235 vdd.n4875 vdd.n4852 35.2919
R10236 vdd.n4914 vdd.n4905 35.2919
R10237 vdd.n4923 vdd.n4905 35.2919
R10238 vdd.n4924 vdd.n4923 35.2919
R10239 vdd.n4927 vdd.n4924 35.2919
R10240 vdd.n4927 vdd.n4926 35.2919
R10241 vdd.n4926 vdd.n4903 35.2919
R10242 vdd.n4960 vdd.n4951 35.2919
R10243 vdd.n4969 vdd.n4951 35.2919
R10244 vdd.n4970 vdd.n4969 35.2919
R10245 vdd.n4973 vdd.n4970 35.2919
R10246 vdd.n4973 vdd.n4972 35.2919
R10247 vdd.n4972 vdd.n4949 35.2919
R10248 vdd.n5008 vdd.n4999 35.2919
R10249 vdd.n5017 vdd.n4999 35.2919
R10250 vdd.n5018 vdd.n5017 35.2919
R10251 vdd.n5021 vdd.n5018 35.2919
R10252 vdd.n5021 vdd.n5020 35.2919
R10253 vdd.n5020 vdd.n4997 35.2919
R10254 vdd.n5054 vdd.n5045 35.2919
R10255 vdd.n5063 vdd.n5045 35.2919
R10256 vdd.n5064 vdd.n5063 35.2919
R10257 vdd.n5067 vdd.n5064 35.2919
R10258 vdd.n5067 vdd.n5066 35.2919
R10259 vdd.n5066 vdd.n5043 35.2919
R10260 vdd.n5099 vdd.n5090 35.2919
R10261 vdd.n5108 vdd.n5090 35.2919
R10262 vdd.n5109 vdd.n5108 35.2919
R10263 vdd.n5112 vdd.n5109 35.2919
R10264 vdd.n5112 vdd.n5111 35.2919
R10265 vdd.n5111 vdd.n5088 35.2919
R10266 vdd.n5149 vdd.n5140 35.2919
R10267 vdd.n5158 vdd.n5140 35.2919
R10268 vdd.n5159 vdd.n5158 35.2919
R10269 vdd.n5162 vdd.n5159 35.2919
R10270 vdd.n5162 vdd.n5161 35.2919
R10271 vdd.n5161 vdd.n5138 35.2919
R10272 vdd.n5195 vdd.n5186 35.2919
R10273 vdd.n5204 vdd.n5186 35.2919
R10274 vdd.n5205 vdd.n5204 35.2919
R10275 vdd.n5208 vdd.n5205 35.2919
R10276 vdd.n5208 vdd.n5207 35.2919
R10277 vdd.n5207 vdd.n5184 35.2919
R10278 vdd.n5243 vdd.n5234 35.2919
R10279 vdd.n5252 vdd.n5234 35.2919
R10280 vdd.n5253 vdd.n5252 35.2919
R10281 vdd.n5256 vdd.n5253 35.2919
R10282 vdd.n5256 vdd.n5255 35.2919
R10283 vdd.n5255 vdd.n5232 35.2919
R10284 vdd.n4207 vdd.n4205 35.2919
R10285 vdd.n4211 vdd.n4205 35.2919
R10286 vdd.n4212 vdd.n4211 35.2919
R10287 vdd.n4215 vdd.n4212 35.2919
R10288 vdd.n4215 vdd.n4214 35.2919
R10289 vdd.n4214 vdd.n4200 35.2919
R10290 vdd.n5290 vdd.n5281 35.2919
R10291 vdd.n5299 vdd.n5281 35.2919
R10292 vdd.n5300 vdd.n5299 35.2919
R10293 vdd.n5303 vdd.n5300 35.2919
R10294 vdd.n5303 vdd.n5302 35.2919
R10295 vdd.n5302 vdd.n5279 35.2919
R10296 vdd.n5335 vdd.n5326 35.2919
R10297 vdd.n5344 vdd.n5326 35.2919
R10298 vdd.n5345 vdd.n5344 35.2919
R10299 vdd.n5348 vdd.n5345 35.2919
R10300 vdd.n5348 vdd.n5347 35.2919
R10301 vdd.n5347 vdd.n5324 35.2919
R10302 vdd.n5385 vdd.n5376 35.2919
R10303 vdd.n5394 vdd.n5376 35.2919
R10304 vdd.n5395 vdd.n5394 35.2919
R10305 vdd.n5398 vdd.n5395 35.2919
R10306 vdd.n5398 vdd.n5397 35.2919
R10307 vdd.n5397 vdd.n5374 35.2919
R10308 vdd.n5431 vdd.n5422 35.2919
R10309 vdd.n5440 vdd.n5422 35.2919
R10310 vdd.n5441 vdd.n5440 35.2919
R10311 vdd.n5444 vdd.n5441 35.2919
R10312 vdd.n5444 vdd.n5443 35.2919
R10313 vdd.n5443 vdd.n5420 35.2919
R10314 vdd.n5479 vdd.n5470 35.2919
R10315 vdd.n5488 vdd.n5470 35.2919
R10316 vdd.n5489 vdd.n5488 35.2919
R10317 vdd.n5492 vdd.n5489 35.2919
R10318 vdd.n5492 vdd.n5491 35.2919
R10319 vdd.n5491 vdd.n5468 35.2919
R10320 vdd.n5616 vdd.n5609 35.2919
R10321 vdd.n5627 vdd.n5609 35.2919
R10322 vdd.n5628 vdd.n5627 35.2919
R10323 vdd.n5629 vdd.n5628 35.2919
R10324 vdd.n5630 vdd.n5629 35.2919
R10325 vdd.n5635 vdd.n5630 35.2919
R10326 vdd.n5570 vdd.n5563 35.2919
R10327 vdd.n5581 vdd.n5563 35.2919
R10328 vdd.n5582 vdd.n5581 35.2919
R10329 vdd.n5583 vdd.n5582 35.2919
R10330 vdd.n5584 vdd.n5583 35.2919
R10331 vdd.n5589 vdd.n5584 35.2919
R10332 vdd.n5663 vdd.n5656 35.2919
R10333 vdd.n5674 vdd.n5656 35.2919
R10334 vdd.n5675 vdd.n5674 35.2919
R10335 vdd.n5676 vdd.n5675 35.2919
R10336 vdd.n5677 vdd.n5676 35.2919
R10337 vdd.n5682 vdd.n5677 35.2919
R10338 vdd.n5711 vdd.n5704 35.2919
R10339 vdd.n5722 vdd.n5704 35.2919
R10340 vdd.n5723 vdd.n5722 35.2919
R10341 vdd.n5724 vdd.n5723 35.2919
R10342 vdd.n5725 vdd.n5724 35.2919
R10343 vdd.n5730 vdd.n5725 35.2919
R10344 vdd.n5757 vdd.n5750 35.2919
R10345 vdd.n5768 vdd.n5750 35.2919
R10346 vdd.n5769 vdd.n5768 35.2919
R10347 vdd.n5770 vdd.n5769 35.2919
R10348 vdd.n5771 vdd.n5770 35.2919
R10349 vdd.n5776 vdd.n5771 35.2919
R10350 vdd.n4023 vdd.n4022 35.2919
R10351 vdd.n4024 vdd.n4023 35.2919
R10352 vdd.n4025 vdd.n4024 35.2919
R10353 vdd.n4026 vdd.n4025 35.2919
R10354 vdd.n4026 vdd.n4001 35.2919
R10355 vdd.n4042 vdd.n4001 35.2919
R10356 vdd.n5899 vdd.n5892 35.2919
R10357 vdd.n5910 vdd.n5892 35.2919
R10358 vdd.n5911 vdd.n5910 35.2919
R10359 vdd.n5912 vdd.n5911 35.2919
R10360 vdd.n5913 vdd.n5912 35.2919
R10361 vdd.n5918 vdd.n5913 35.2919
R10362 vdd.n5852 vdd.n5845 35.2919
R10363 vdd.n5863 vdd.n5845 35.2919
R10364 vdd.n5864 vdd.n5863 35.2919
R10365 vdd.n5865 vdd.n5864 35.2919
R10366 vdd.n5866 vdd.n5865 35.2919
R10367 vdd.n5871 vdd.n5866 35.2919
R10368 vdd.n5806 vdd.n5799 35.2919
R10369 vdd.n5817 vdd.n5799 35.2919
R10370 vdd.n5818 vdd.n5817 35.2919
R10371 vdd.n5819 vdd.n5818 35.2919
R10372 vdd.n5820 vdd.n5819 35.2919
R10373 vdd.n5825 vdd.n5820 35.2919
R10374 vdd.n5946 vdd.n5939 35.2919
R10375 vdd.n5957 vdd.n5939 35.2919
R10376 vdd.n5958 vdd.n5957 35.2919
R10377 vdd.n5959 vdd.n5958 35.2919
R10378 vdd.n5960 vdd.n5959 35.2919
R10379 vdd.n5965 vdd.n5960 35.2919
R10380 vdd.n5994 vdd.n5987 35.2919
R10381 vdd.n6005 vdd.n5987 35.2919
R10382 vdd.n6006 vdd.n6005 35.2919
R10383 vdd.n6007 vdd.n6006 35.2919
R10384 vdd.n6008 vdd.n6007 35.2919
R10385 vdd.n6013 vdd.n6008 35.2919
R10386 vdd.n6040 vdd.n6033 35.2919
R10387 vdd.n6051 vdd.n6033 35.2919
R10388 vdd.n6052 vdd.n6051 35.2919
R10389 vdd.n6053 vdd.n6052 35.2919
R10390 vdd.n6054 vdd.n6053 35.2919
R10391 vdd.n6059 vdd.n6054 35.2919
R10392 vdd.n6134 vdd.n6127 35.2919
R10393 vdd.n6145 vdd.n6127 35.2919
R10394 vdd.n6146 vdd.n6145 35.2919
R10395 vdd.n6147 vdd.n6146 35.2919
R10396 vdd.n6148 vdd.n6147 35.2919
R10397 vdd.n6153 vdd.n6148 35.2919
R10398 vdd.n6088 vdd.n6081 35.2919
R10399 vdd.n6099 vdd.n6081 35.2919
R10400 vdd.n6100 vdd.n6099 35.2919
R10401 vdd.n6101 vdd.n6100 35.2919
R10402 vdd.n6102 vdd.n6101 35.2919
R10403 vdd.n6107 vdd.n6102 35.2919
R10404 vdd.n6181 vdd.n6174 35.2919
R10405 vdd.n6192 vdd.n6174 35.2919
R10406 vdd.n6193 vdd.n6192 35.2919
R10407 vdd.n6194 vdd.n6193 35.2919
R10408 vdd.n6195 vdd.n6194 35.2919
R10409 vdd.n6200 vdd.n6195 35.2919
R10410 vdd.n6229 vdd.n6222 35.2919
R10411 vdd.n6240 vdd.n6222 35.2919
R10412 vdd.n6241 vdd.n6240 35.2919
R10413 vdd.n6242 vdd.n6241 35.2919
R10414 vdd.n6243 vdd.n6242 35.2919
R10415 vdd.n6248 vdd.n6243 35.2919
R10416 vdd.n6275 vdd.n6268 35.2919
R10417 vdd.n6286 vdd.n6268 35.2919
R10418 vdd.n6287 vdd.n6286 35.2919
R10419 vdd.n6288 vdd.n6287 35.2919
R10420 vdd.n6289 vdd.n6288 35.2919
R10421 vdd.n6294 vdd.n6289 35.2919
R10422 vdd.n3787 vdd.n3786 35.2919
R10423 vdd.n3788 vdd.n3787 35.2919
R10424 vdd.n3789 vdd.n3788 35.2919
R10425 vdd.n3790 vdd.n3789 35.2919
R10426 vdd.n3790 vdd.n3765 35.2919
R10427 vdd.n3806 vdd.n3765 35.2919
R10428 vdd.n6370 vdd.n6363 35.2919
R10429 vdd.n6381 vdd.n6363 35.2919
R10430 vdd.n6382 vdd.n6381 35.2919
R10431 vdd.n6383 vdd.n6382 35.2919
R10432 vdd.n6384 vdd.n6383 35.2919
R10433 vdd.n6389 vdd.n6384 35.2919
R10434 vdd.n6324 vdd.n6317 35.2919
R10435 vdd.n6335 vdd.n6317 35.2919
R10436 vdd.n6336 vdd.n6335 35.2919
R10437 vdd.n6337 vdd.n6336 35.2919
R10438 vdd.n6338 vdd.n6337 35.2919
R10439 vdd.n6343 vdd.n6338 35.2919
R10440 vdd.n6417 vdd.n6410 35.2919
R10441 vdd.n6428 vdd.n6410 35.2919
R10442 vdd.n6429 vdd.n6428 35.2919
R10443 vdd.n6430 vdd.n6429 35.2919
R10444 vdd.n6431 vdd.n6430 35.2919
R10445 vdd.n6436 vdd.n6431 35.2919
R10446 vdd.n6465 vdd.n6458 35.2919
R10447 vdd.n6476 vdd.n6458 35.2919
R10448 vdd.n6477 vdd.n6476 35.2919
R10449 vdd.n6478 vdd.n6477 35.2919
R10450 vdd.n6479 vdd.n6478 35.2919
R10451 vdd.n6484 vdd.n6479 35.2919
R10452 vdd.n6511 vdd.n6504 35.2919
R10453 vdd.n6522 vdd.n6504 35.2919
R10454 vdd.n6523 vdd.n6522 35.2919
R10455 vdd.n6524 vdd.n6523 35.2919
R10456 vdd.n6525 vdd.n6524 35.2919
R10457 vdd.n6530 vdd.n6525 35.2919
R10458 vdd.n671 vdd.n664 35.2919
R10459 vdd.n682 vdd.n664 35.2919
R10460 vdd.n683 vdd.n682 35.2919
R10461 vdd.n684 vdd.n683 35.2919
R10462 vdd.n685 vdd.n684 35.2919
R10463 vdd.n690 vdd.n685 35.2919
R10464 vdd.n717 vdd.n710 35.2919
R10465 vdd.n728 vdd.n710 35.2919
R10466 vdd.n729 vdd.n728 35.2919
R10467 vdd.n730 vdd.n729 35.2919
R10468 vdd.n731 vdd.n730 35.2919
R10469 vdd.n736 vdd.n731 35.2919
R10470 vdd.n815 vdd.n808 35.2919
R10471 vdd.n826 vdd.n808 35.2919
R10472 vdd.n827 vdd.n826 35.2919
R10473 vdd.n828 vdd.n827 35.2919
R10474 vdd.n829 vdd.n828 35.2919
R10475 vdd.n834 vdd.n829 35.2919
R10476 vdd.n861 vdd.n854 35.2919
R10477 vdd.n872 vdd.n854 35.2919
R10478 vdd.n873 vdd.n872 35.2919
R10479 vdd.n874 vdd.n873 35.2919
R10480 vdd.n875 vdd.n874 35.2919
R10481 vdd.n880 vdd.n875 35.2919
R10482 vdd.n907 vdd.n900 35.2919
R10483 vdd.n918 vdd.n900 35.2919
R10484 vdd.n919 vdd.n918 35.2919
R10485 vdd.n920 vdd.n919 35.2919
R10486 vdd.n921 vdd.n920 35.2919
R10487 vdd.n926 vdd.n921 35.2919
R10488 vdd.n953 vdd.n946 35.2919
R10489 vdd.n964 vdd.n946 35.2919
R10490 vdd.n965 vdd.n964 35.2919
R10491 vdd.n966 vdd.n965 35.2919
R10492 vdd.n967 vdd.n966 35.2919
R10493 vdd.n972 vdd.n967 35.2919
R10494 vdd.n1051 vdd.n1044 35.2919
R10495 vdd.n1062 vdd.n1044 35.2919
R10496 vdd.n1063 vdd.n1062 35.2919
R10497 vdd.n1064 vdd.n1063 35.2919
R10498 vdd.n1065 vdd.n1064 35.2919
R10499 vdd.n1070 vdd.n1065 35.2919
R10500 vdd.n2509 vdd.n2502 35.2919
R10501 vdd.n2520 vdd.n2502 35.2919
R10502 vdd.n2521 vdd.n2520 35.2919
R10503 vdd.n2522 vdd.n2521 35.2919
R10504 vdd.n2523 vdd.n2522 35.2919
R10505 vdd.n2528 vdd.n2523 35.2919
R10506 vdd.n1100 vdd.n1091 35.2919
R10507 vdd.n1109 vdd.n1091 35.2919
R10508 vdd.n1110 vdd.n1109 35.2919
R10509 vdd.n1113 vdd.n1110 35.2919
R10510 vdd.n1113 vdd.n1112 35.2919
R10511 vdd.n1112 vdd.n1089 35.2919
R10512 vdd.n1146 vdd.n1137 35.2919
R10513 vdd.n1155 vdd.n1137 35.2919
R10514 vdd.n1156 vdd.n1155 35.2919
R10515 vdd.n1159 vdd.n1156 35.2919
R10516 vdd.n1159 vdd.n1158 35.2919
R10517 vdd.n1158 vdd.n1135 35.2919
R10518 vdd.n1243 vdd.n1234 35.2919
R10519 vdd.n1252 vdd.n1234 35.2919
R10520 vdd.n1253 vdd.n1252 35.2919
R10521 vdd.n1256 vdd.n1253 35.2919
R10522 vdd.n1256 vdd.n1255 35.2919
R10523 vdd.n1255 vdd.n1232 35.2919
R10524 vdd.n1289 vdd.n1280 35.2919
R10525 vdd.n1298 vdd.n1280 35.2919
R10526 vdd.n1299 vdd.n1298 35.2919
R10527 vdd.n1302 vdd.n1299 35.2919
R10528 vdd.n1302 vdd.n1301 35.2919
R10529 vdd.n1301 vdd.n1278 35.2919
R10530 vdd.n1335 vdd.n1326 35.2919
R10531 vdd.n1344 vdd.n1326 35.2919
R10532 vdd.n1345 vdd.n1344 35.2919
R10533 vdd.n1348 vdd.n1345 35.2919
R10534 vdd.n1348 vdd.n1347 35.2919
R10535 vdd.n1347 vdd.n1324 35.2919
R10536 vdd.n1381 vdd.n1372 35.2919
R10537 vdd.n1390 vdd.n1372 35.2919
R10538 vdd.n1391 vdd.n1390 35.2919
R10539 vdd.n1394 vdd.n1391 35.2919
R10540 vdd.n1394 vdd.n1393 35.2919
R10541 vdd.n1393 vdd.n1370 35.2919
R10542 vdd.n1478 vdd.n1469 35.2919
R10543 vdd.n1487 vdd.n1469 35.2919
R10544 vdd.n1488 vdd.n1487 35.2919
R10545 vdd.n1491 vdd.n1488 35.2919
R10546 vdd.n1491 vdd.n1490 35.2919
R10547 vdd.n1490 vdd.n1467 35.2919
R10548 vdd.n627 vdd.n618 35.2919
R10549 vdd.n636 vdd.n618 35.2919
R10550 vdd.n637 vdd.n636 35.2919
R10551 vdd.n640 vdd.n637 35.2919
R10552 vdd.n640 vdd.n639 35.2919
R10553 vdd.n639 vdd.n616 35.2919
R10554 vdd.n1522 vdd.n1513 35.2919
R10555 vdd.n1531 vdd.n1513 35.2919
R10556 vdd.n1532 vdd.n1531 35.2919
R10557 vdd.n1535 vdd.n1532 35.2919
R10558 vdd.n1535 vdd.n1534 35.2919
R10559 vdd.n1534 vdd.n1511 35.2919
R10560 vdd.n1567 vdd.n1558 35.2919
R10561 vdd.n1576 vdd.n1558 35.2919
R10562 vdd.n1577 vdd.n1576 35.2919
R10563 vdd.n1580 vdd.n1577 35.2919
R10564 vdd.n1580 vdd.n1579 35.2919
R10565 vdd.n1579 vdd.n1556 35.2919
R10566 vdd.n1617 vdd.n1608 35.2919
R10567 vdd.n1626 vdd.n1608 35.2919
R10568 vdd.n1627 vdd.n1626 35.2919
R10569 vdd.n1630 vdd.n1627 35.2919
R10570 vdd.n1630 vdd.n1629 35.2919
R10571 vdd.n1629 vdd.n1606 35.2919
R10572 vdd.n1663 vdd.n1654 35.2919
R10573 vdd.n1672 vdd.n1654 35.2919
R10574 vdd.n1673 vdd.n1672 35.2919
R10575 vdd.n1676 vdd.n1673 35.2919
R10576 vdd.n1676 vdd.n1675 35.2919
R10577 vdd.n1675 vdd.n1652 35.2919
R10578 vdd.n1711 vdd.n1702 35.2919
R10579 vdd.n1720 vdd.n1702 35.2919
R10580 vdd.n1721 vdd.n1720 35.2919
R10581 vdd.n1724 vdd.n1721 35.2919
R10582 vdd.n1724 vdd.n1723 35.2919
R10583 vdd.n1723 vdd.n1700 35.2919
R10584 vdd.n1428 vdd.n1426 35.2919
R10585 vdd.n1432 vdd.n1426 35.2919
R10586 vdd.n1433 vdd.n1432 35.2919
R10587 vdd.n1436 vdd.n1433 35.2919
R10588 vdd.n1436 vdd.n1435 35.2919
R10589 vdd.n1435 vdd.n1421 35.2919
R10590 vdd.n1758 vdd.n1749 35.2919
R10591 vdd.n1767 vdd.n1749 35.2919
R10592 vdd.n1768 vdd.n1767 35.2919
R10593 vdd.n1771 vdd.n1768 35.2919
R10594 vdd.n1771 vdd.n1770 35.2919
R10595 vdd.n1770 vdd.n1747 35.2919
R10596 vdd.n1803 vdd.n1794 35.2919
R10597 vdd.n1812 vdd.n1794 35.2919
R10598 vdd.n1813 vdd.n1812 35.2919
R10599 vdd.n1816 vdd.n1813 35.2919
R10600 vdd.n1816 vdd.n1815 35.2919
R10601 vdd.n1815 vdd.n1792 35.2919
R10602 vdd.n1849 vdd.n1840 35.2919
R10603 vdd.n1858 vdd.n1840 35.2919
R10604 vdd.n1859 vdd.n1858 35.2919
R10605 vdd.n1862 vdd.n1859 35.2919
R10606 vdd.n1862 vdd.n1861 35.2919
R10607 vdd.n1861 vdd.n1838 35.2919
R10608 vdd.n1900 vdd.n1891 35.2919
R10609 vdd.n1909 vdd.n1891 35.2919
R10610 vdd.n1910 vdd.n1909 35.2919
R10611 vdd.n1913 vdd.n1910 35.2919
R10612 vdd.n1913 vdd.n1912 35.2919
R10613 vdd.n1912 vdd.n1889 35.2919
R10614 vdd.n1946 vdd.n1937 35.2919
R10615 vdd.n1955 vdd.n1937 35.2919
R10616 vdd.n1956 vdd.n1955 35.2919
R10617 vdd.n1959 vdd.n1956 35.2919
R10618 vdd.n1959 vdd.n1958 35.2919
R10619 vdd.n1958 vdd.n1935 35.2919
R10620 vdd.n1994 vdd.n1985 35.2919
R10621 vdd.n2003 vdd.n1985 35.2919
R10622 vdd.n2004 vdd.n2003 35.2919
R10623 vdd.n2007 vdd.n2004 35.2919
R10624 vdd.n2007 vdd.n2006 35.2919
R10625 vdd.n2006 vdd.n1983 35.2919
R10626 vdd.n2040 vdd.n2031 35.2919
R10627 vdd.n2049 vdd.n2031 35.2919
R10628 vdd.n2050 vdd.n2049 35.2919
R10629 vdd.n2053 vdd.n2050 35.2919
R10630 vdd.n2053 vdd.n2052 35.2919
R10631 vdd.n2052 vdd.n2029 35.2919
R10632 vdd.n2085 vdd.n2076 35.2919
R10633 vdd.n2094 vdd.n2076 35.2919
R10634 vdd.n2095 vdd.n2094 35.2919
R10635 vdd.n2098 vdd.n2095 35.2919
R10636 vdd.n2098 vdd.n2097 35.2919
R10637 vdd.n2097 vdd.n2074 35.2919
R10638 vdd.n2135 vdd.n2126 35.2919
R10639 vdd.n2144 vdd.n2126 35.2919
R10640 vdd.n2145 vdd.n2144 35.2919
R10641 vdd.n2148 vdd.n2145 35.2919
R10642 vdd.n2148 vdd.n2147 35.2919
R10643 vdd.n2147 vdd.n2124 35.2919
R10644 vdd.n2181 vdd.n2172 35.2919
R10645 vdd.n2190 vdd.n2172 35.2919
R10646 vdd.n2191 vdd.n2190 35.2919
R10647 vdd.n2194 vdd.n2191 35.2919
R10648 vdd.n2194 vdd.n2193 35.2919
R10649 vdd.n2193 vdd.n2170 35.2919
R10650 vdd.n2229 vdd.n2220 35.2919
R10651 vdd.n2238 vdd.n2220 35.2919
R10652 vdd.n2239 vdd.n2238 35.2919
R10653 vdd.n2242 vdd.n2239 35.2919
R10654 vdd.n2242 vdd.n2241 35.2919
R10655 vdd.n2241 vdd.n2218 35.2919
R10656 vdd.n1193 vdd.n1191 35.2919
R10657 vdd.n1197 vdd.n1191 35.2919
R10658 vdd.n1198 vdd.n1197 35.2919
R10659 vdd.n1201 vdd.n1198 35.2919
R10660 vdd.n1201 vdd.n1200 35.2919
R10661 vdd.n1200 vdd.n1186 35.2919
R10662 vdd.n2276 vdd.n2267 35.2919
R10663 vdd.n2285 vdd.n2267 35.2919
R10664 vdd.n2286 vdd.n2285 35.2919
R10665 vdd.n2289 vdd.n2286 35.2919
R10666 vdd.n2289 vdd.n2288 35.2919
R10667 vdd.n2288 vdd.n2265 35.2919
R10668 vdd.n2321 vdd.n2312 35.2919
R10669 vdd.n2330 vdd.n2312 35.2919
R10670 vdd.n2331 vdd.n2330 35.2919
R10671 vdd.n2334 vdd.n2331 35.2919
R10672 vdd.n2334 vdd.n2333 35.2919
R10673 vdd.n2333 vdd.n2310 35.2919
R10674 vdd.n2371 vdd.n2362 35.2919
R10675 vdd.n2380 vdd.n2362 35.2919
R10676 vdd.n2381 vdd.n2380 35.2919
R10677 vdd.n2384 vdd.n2381 35.2919
R10678 vdd.n2384 vdd.n2383 35.2919
R10679 vdd.n2383 vdd.n2360 35.2919
R10680 vdd.n2417 vdd.n2408 35.2919
R10681 vdd.n2426 vdd.n2408 35.2919
R10682 vdd.n2427 vdd.n2426 35.2919
R10683 vdd.n2430 vdd.n2427 35.2919
R10684 vdd.n2430 vdd.n2429 35.2919
R10685 vdd.n2429 vdd.n2406 35.2919
R10686 vdd.n2465 vdd.n2456 35.2919
R10687 vdd.n2474 vdd.n2456 35.2919
R10688 vdd.n2475 vdd.n2474 35.2919
R10689 vdd.n2478 vdd.n2475 35.2919
R10690 vdd.n2478 vdd.n2477 35.2919
R10691 vdd.n2477 vdd.n2454 35.2919
R10692 vdd.n2602 vdd.n2595 35.2919
R10693 vdd.n2613 vdd.n2595 35.2919
R10694 vdd.n2614 vdd.n2613 35.2919
R10695 vdd.n2615 vdd.n2614 35.2919
R10696 vdd.n2616 vdd.n2615 35.2919
R10697 vdd.n2621 vdd.n2616 35.2919
R10698 vdd.n2556 vdd.n2549 35.2919
R10699 vdd.n2567 vdd.n2549 35.2919
R10700 vdd.n2568 vdd.n2567 35.2919
R10701 vdd.n2569 vdd.n2568 35.2919
R10702 vdd.n2570 vdd.n2569 35.2919
R10703 vdd.n2575 vdd.n2570 35.2919
R10704 vdd.n2649 vdd.n2642 35.2919
R10705 vdd.n2660 vdd.n2642 35.2919
R10706 vdd.n2661 vdd.n2660 35.2919
R10707 vdd.n2662 vdd.n2661 35.2919
R10708 vdd.n2663 vdd.n2662 35.2919
R10709 vdd.n2668 vdd.n2663 35.2919
R10710 vdd.n2697 vdd.n2690 35.2919
R10711 vdd.n2708 vdd.n2690 35.2919
R10712 vdd.n2709 vdd.n2708 35.2919
R10713 vdd.n2710 vdd.n2709 35.2919
R10714 vdd.n2711 vdd.n2710 35.2919
R10715 vdd.n2716 vdd.n2711 35.2919
R10716 vdd.n2743 vdd.n2736 35.2919
R10717 vdd.n2754 vdd.n2736 35.2919
R10718 vdd.n2755 vdd.n2754 35.2919
R10719 vdd.n2756 vdd.n2755 35.2919
R10720 vdd.n2757 vdd.n2756 35.2919
R10721 vdd.n2762 vdd.n2757 35.2919
R10722 vdd.n1009 vdd.n1008 35.2919
R10723 vdd.n1010 vdd.n1009 35.2919
R10724 vdd.n1011 vdd.n1010 35.2919
R10725 vdd.n1012 vdd.n1011 35.2919
R10726 vdd.n1012 vdd.n987 35.2919
R10727 vdd.n1028 vdd.n987 35.2919
R10728 vdd.n2885 vdd.n2878 35.2919
R10729 vdd.n2896 vdd.n2878 35.2919
R10730 vdd.n2897 vdd.n2896 35.2919
R10731 vdd.n2898 vdd.n2897 35.2919
R10732 vdd.n2899 vdd.n2898 35.2919
R10733 vdd.n2904 vdd.n2899 35.2919
R10734 vdd.n2838 vdd.n2831 35.2919
R10735 vdd.n2849 vdd.n2831 35.2919
R10736 vdd.n2850 vdd.n2849 35.2919
R10737 vdd.n2851 vdd.n2850 35.2919
R10738 vdd.n2852 vdd.n2851 35.2919
R10739 vdd.n2857 vdd.n2852 35.2919
R10740 vdd.n2792 vdd.n2785 35.2919
R10741 vdd.n2803 vdd.n2785 35.2919
R10742 vdd.n2804 vdd.n2803 35.2919
R10743 vdd.n2805 vdd.n2804 35.2919
R10744 vdd.n2806 vdd.n2805 35.2919
R10745 vdd.n2811 vdd.n2806 35.2919
R10746 vdd.n2932 vdd.n2925 35.2919
R10747 vdd.n2943 vdd.n2925 35.2919
R10748 vdd.n2944 vdd.n2943 35.2919
R10749 vdd.n2945 vdd.n2944 35.2919
R10750 vdd.n2946 vdd.n2945 35.2919
R10751 vdd.n2951 vdd.n2946 35.2919
R10752 vdd.n2980 vdd.n2973 35.2919
R10753 vdd.n2991 vdd.n2973 35.2919
R10754 vdd.n2992 vdd.n2991 35.2919
R10755 vdd.n2993 vdd.n2992 35.2919
R10756 vdd.n2994 vdd.n2993 35.2919
R10757 vdd.n2999 vdd.n2994 35.2919
R10758 vdd.n3026 vdd.n3019 35.2919
R10759 vdd.n3037 vdd.n3019 35.2919
R10760 vdd.n3038 vdd.n3037 35.2919
R10761 vdd.n3039 vdd.n3038 35.2919
R10762 vdd.n3040 vdd.n3039 35.2919
R10763 vdd.n3045 vdd.n3040 35.2919
R10764 vdd.n3120 vdd.n3113 35.2919
R10765 vdd.n3131 vdd.n3113 35.2919
R10766 vdd.n3132 vdd.n3131 35.2919
R10767 vdd.n3133 vdd.n3132 35.2919
R10768 vdd.n3134 vdd.n3133 35.2919
R10769 vdd.n3139 vdd.n3134 35.2919
R10770 vdd.n3074 vdd.n3067 35.2919
R10771 vdd.n3085 vdd.n3067 35.2919
R10772 vdd.n3086 vdd.n3085 35.2919
R10773 vdd.n3087 vdd.n3086 35.2919
R10774 vdd.n3088 vdd.n3087 35.2919
R10775 vdd.n3093 vdd.n3088 35.2919
R10776 vdd.n3167 vdd.n3160 35.2919
R10777 vdd.n3178 vdd.n3160 35.2919
R10778 vdd.n3179 vdd.n3178 35.2919
R10779 vdd.n3180 vdd.n3179 35.2919
R10780 vdd.n3181 vdd.n3180 35.2919
R10781 vdd.n3186 vdd.n3181 35.2919
R10782 vdd.n3215 vdd.n3208 35.2919
R10783 vdd.n3226 vdd.n3208 35.2919
R10784 vdd.n3227 vdd.n3226 35.2919
R10785 vdd.n3228 vdd.n3227 35.2919
R10786 vdd.n3229 vdd.n3228 35.2919
R10787 vdd.n3234 vdd.n3229 35.2919
R10788 vdd.n3261 vdd.n3254 35.2919
R10789 vdd.n3272 vdd.n3254 35.2919
R10790 vdd.n3273 vdd.n3272 35.2919
R10791 vdd.n3274 vdd.n3273 35.2919
R10792 vdd.n3275 vdd.n3274 35.2919
R10793 vdd.n3280 vdd.n3275 35.2919
R10794 vdd.n773 vdd.n772 35.2919
R10795 vdd.n774 vdd.n773 35.2919
R10796 vdd.n775 vdd.n774 35.2919
R10797 vdd.n776 vdd.n775 35.2919
R10798 vdd.n776 vdd.n751 35.2919
R10799 vdd.n792 vdd.n751 35.2919
R10800 vdd.n3356 vdd.n3349 35.2919
R10801 vdd.n3367 vdd.n3349 35.2919
R10802 vdd.n3368 vdd.n3367 35.2919
R10803 vdd.n3369 vdd.n3368 35.2919
R10804 vdd.n3370 vdd.n3369 35.2919
R10805 vdd.n3375 vdd.n3370 35.2919
R10806 vdd.n3310 vdd.n3303 35.2919
R10807 vdd.n3321 vdd.n3303 35.2919
R10808 vdd.n3322 vdd.n3321 35.2919
R10809 vdd.n3323 vdd.n3322 35.2919
R10810 vdd.n3324 vdd.n3323 35.2919
R10811 vdd.n3329 vdd.n3324 35.2919
R10812 vdd.n3403 vdd.n3396 35.2919
R10813 vdd.n3414 vdd.n3396 35.2919
R10814 vdd.n3415 vdd.n3414 35.2919
R10815 vdd.n3416 vdd.n3415 35.2919
R10816 vdd.n3417 vdd.n3416 35.2919
R10817 vdd.n3422 vdd.n3417 35.2919
R10818 vdd.n3451 vdd.n3444 35.2919
R10819 vdd.n3462 vdd.n3444 35.2919
R10820 vdd.n3463 vdd.n3462 35.2919
R10821 vdd.n3464 vdd.n3463 35.2919
R10822 vdd.n3465 vdd.n3464 35.2919
R10823 vdd.n3470 vdd.n3465 35.2919
R10824 vdd.n3497 vdd.n3490 35.2919
R10825 vdd.n3508 vdd.n3490 35.2919
R10826 vdd.n3509 vdd.n3508 35.2919
R10827 vdd.n3510 vdd.n3509 35.2919
R10828 vdd.n3511 vdd.n3510 35.2919
R10829 vdd.n3516 vdd.n3511 35.2919
R10830 vdd.n579 vdd.n572 35.2919
R10831 vdd.n590 vdd.n572 35.2919
R10832 vdd.n591 vdd.n590 35.2919
R10833 vdd.n592 vdd.n591 35.2919
R10834 vdd.n593 vdd.n592 35.2919
R10835 vdd.n598 vdd.n593 35.2919
R10836 vdd.n3592 vdd.n3585 35.2919
R10837 vdd.n3603 vdd.n3585 35.2919
R10838 vdd.n3604 vdd.n3603 35.2919
R10839 vdd.n3605 vdd.n3604 35.2919
R10840 vdd.n3606 vdd.n3605 35.2919
R10841 vdd.n3611 vdd.n3606 35.2919
R10842 vdd.n3546 vdd.n3539 35.2919
R10843 vdd.n3557 vdd.n3539 35.2919
R10844 vdd.n3558 vdd.n3557 35.2919
R10845 vdd.n3559 vdd.n3558 35.2919
R10846 vdd.n3560 vdd.n3559 35.2919
R10847 vdd.n3565 vdd.n3560 35.2919
R10848 vdd.n6606 vdd.n6599 35.2919
R10849 vdd.n6617 vdd.n6599 35.2919
R10850 vdd.n6618 vdd.n6617 35.2919
R10851 vdd.n6619 vdd.n6618 35.2919
R10852 vdd.n6620 vdd.n6619 35.2919
R10853 vdd.n6625 vdd.n6620 35.2919
R10854 vdd.n6560 vdd.n6553 35.2919
R10855 vdd.n6571 vdd.n6553 35.2919
R10856 vdd.n6572 vdd.n6571 35.2919
R10857 vdd.n6573 vdd.n6572 35.2919
R10858 vdd.n6574 vdd.n6573 35.2919
R10859 vdd.n6579 vdd.n6574 35.2919
R10860 vdd.n9620 vdd.n9613 35.2919
R10861 vdd.n9631 vdd.n9613 35.2919
R10862 vdd.n9632 vdd.n9631 35.2919
R10863 vdd.n9633 vdd.n9632 35.2919
R10864 vdd.n9634 vdd.n9633 35.2919
R10865 vdd.n9639 vdd.n9634 35.2919
R10866 vdd.n9574 vdd.n9567 35.2919
R10867 vdd.n9585 vdd.n9567 35.2919
R10868 vdd.n9586 vdd.n9585 35.2919
R10869 vdd.n9587 vdd.n9586 35.2919
R10870 vdd.n9588 vdd.n9587 35.2919
R10871 vdd.n9593 vdd.n9588 35.2919
R10872 vdd.n9666 vdd.n9659 35.2919
R10873 vdd.n9677 vdd.n9659 35.2919
R10874 vdd.n9678 vdd.n9677 35.2919
R10875 vdd.n9679 vdd.n9678 35.2919
R10876 vdd.n9680 vdd.n9679 35.2919
R10877 vdd.n9685 vdd.n9680 35.2919
R10878 vdd.n9712 vdd.n9705 35.2919
R10879 vdd.n9723 vdd.n9705 35.2919
R10880 vdd.n9724 vdd.n9723 35.2919
R10881 vdd.n9725 vdd.n9724 35.2919
R10882 vdd.n9726 vdd.n9725 35.2919
R10883 vdd.n9731 vdd.n9726 35.2919
R10884 vdd.n9810 vdd.n9803 35.2919
R10885 vdd.n9821 vdd.n9803 35.2919
R10886 vdd.n9822 vdd.n9821 35.2919
R10887 vdd.n9823 vdd.n9822 35.2919
R10888 vdd.n9824 vdd.n9823 35.2919
R10889 vdd.n9829 vdd.n9824 35.2919
R10890 vdd.n9856 vdd.n9849 35.2919
R10891 vdd.n9867 vdd.n9849 35.2919
R10892 vdd.n9868 vdd.n9867 35.2919
R10893 vdd.n9869 vdd.n9868 35.2919
R10894 vdd.n9870 vdd.n9869 35.2919
R10895 vdd.n9875 vdd.n9870 35.2919
R10896 vdd.n9902 vdd.n9895 35.2919
R10897 vdd.n9913 vdd.n9895 35.2919
R10898 vdd.n9914 vdd.n9913 35.2919
R10899 vdd.n9915 vdd.n9914 35.2919
R10900 vdd.n9916 vdd.n9915 35.2919
R10901 vdd.n9921 vdd.n9916 35.2919
R10902 vdd.n9948 vdd.n9941 35.2919
R10903 vdd.n9959 vdd.n9941 35.2919
R10904 vdd.n9960 vdd.n9959 35.2919
R10905 vdd.n9961 vdd.n9960 35.2919
R10906 vdd.n9962 vdd.n9961 35.2919
R10907 vdd.n9967 vdd.n9962 35.2919
R10908 vdd.n10046 vdd.n10039 35.2919
R10909 vdd.n10057 vdd.n10039 35.2919
R10910 vdd.n10058 vdd.n10057 35.2919
R10911 vdd.n10059 vdd.n10058 35.2919
R10912 vdd.n10060 vdd.n10059 35.2919
R10913 vdd.n10065 vdd.n10060 35.2919
R10914 vdd.n62 vdd.n55 35.2919
R10915 vdd.n73 vdd.n55 35.2919
R10916 vdd.n74 vdd.n73 35.2919
R10917 vdd.n75 vdd.n74 35.2919
R10918 vdd.n76 vdd.n75 35.2919
R10919 vdd.n81 vdd.n76 35.2919
R10920 vdd.n16 vdd.n9 35.2919
R10921 vdd.n27 vdd.n9 35.2919
R10922 vdd.n28 vdd.n27 35.2919
R10923 vdd.n29 vdd.n28 35.2919
R10924 vdd.n30 vdd.n29 35.2919
R10925 vdd.n35 vdd.n30 35.2919
R10926 vdd.n10092 vdd.n10085 35.2919
R10927 vdd.n10103 vdd.n10085 35.2919
R10928 vdd.n10104 vdd.n10103 35.2919
R10929 vdd.n10105 vdd.n10104 35.2919
R10930 vdd.n10106 vdd.n10105 35.2919
R10931 vdd.n10111 vdd.n10106 35.2919
R10932 vdd.n10140 vdd.n10133 35.2919
R10933 vdd.n10151 vdd.n10133 35.2919
R10934 vdd.n10152 vdd.n10151 35.2919
R10935 vdd.n10153 vdd.n10152 35.2919
R10936 vdd.n10154 vdd.n10153 35.2919
R10937 vdd.n10159 vdd.n10154 35.2919
R10938 vdd.n10186 vdd.n10179 35.2919
R10939 vdd.n10197 vdd.n10179 35.2919
R10940 vdd.n10198 vdd.n10197 35.2919
R10941 vdd.n10199 vdd.n10198 35.2919
R10942 vdd.n10200 vdd.n10199 35.2919
R10943 vdd.n10205 vdd.n10200 35.2919
R10944 vdd.n10004 vdd.n10003 35.2919
R10945 vdd.n10005 vdd.n10004 35.2919
R10946 vdd.n10006 vdd.n10005 35.2919
R10947 vdd.n10007 vdd.n10006 35.2919
R10948 vdd.n10007 vdd.n9982 35.2919
R10949 vdd.n10023 vdd.n9982 35.2919
R10950 vdd.n10328 vdd.n10321 35.2919
R10951 vdd.n10339 vdd.n10321 35.2919
R10952 vdd.n10340 vdd.n10339 35.2919
R10953 vdd.n10341 vdd.n10340 35.2919
R10954 vdd.n10342 vdd.n10341 35.2919
R10955 vdd.n10347 vdd.n10342 35.2919
R10956 vdd.n10281 vdd.n10274 35.2919
R10957 vdd.n10292 vdd.n10274 35.2919
R10958 vdd.n10293 vdd.n10292 35.2919
R10959 vdd.n10294 vdd.n10293 35.2919
R10960 vdd.n10295 vdd.n10294 35.2919
R10961 vdd.n10300 vdd.n10295 35.2919
R10962 vdd.n10235 vdd.n10228 35.2919
R10963 vdd.n10246 vdd.n10228 35.2919
R10964 vdd.n10247 vdd.n10246 35.2919
R10965 vdd.n10248 vdd.n10247 35.2919
R10966 vdd.n10249 vdd.n10248 35.2919
R10967 vdd.n10254 vdd.n10249 35.2919
R10968 vdd.n10375 vdd.n10368 35.2919
R10969 vdd.n10386 vdd.n10368 35.2919
R10970 vdd.n10387 vdd.n10386 35.2919
R10971 vdd.n10388 vdd.n10387 35.2919
R10972 vdd.n10389 vdd.n10388 35.2919
R10973 vdd.n10394 vdd.n10389 35.2919
R10974 vdd.n10423 vdd.n10416 35.2919
R10975 vdd.n10434 vdd.n10416 35.2919
R10976 vdd.n10435 vdd.n10434 35.2919
R10977 vdd.n10436 vdd.n10435 35.2919
R10978 vdd.n10437 vdd.n10436 35.2919
R10979 vdd.n10442 vdd.n10437 35.2919
R10980 vdd.n10469 vdd.n10462 35.2919
R10981 vdd.n10480 vdd.n10462 35.2919
R10982 vdd.n10481 vdd.n10480 35.2919
R10983 vdd.n10482 vdd.n10481 35.2919
R10984 vdd.n10483 vdd.n10482 35.2919
R10985 vdd.n10488 vdd.n10483 35.2919
R10986 vdd.n10563 vdd.n10556 35.2919
R10987 vdd.n10574 vdd.n10556 35.2919
R10988 vdd.n10575 vdd.n10574 35.2919
R10989 vdd.n10576 vdd.n10575 35.2919
R10990 vdd.n10577 vdd.n10576 35.2919
R10991 vdd.n10582 vdd.n10577 35.2919
R10992 vdd.n10517 vdd.n10510 35.2919
R10993 vdd.n10528 vdd.n10510 35.2919
R10994 vdd.n10529 vdd.n10528 35.2919
R10995 vdd.n10530 vdd.n10529 35.2919
R10996 vdd.n10531 vdd.n10530 35.2919
R10997 vdd.n10536 vdd.n10531 35.2919
R10998 vdd.n10610 vdd.n10603 35.2919
R10999 vdd.n10621 vdd.n10603 35.2919
R11000 vdd.n10622 vdd.n10621 35.2919
R11001 vdd.n10623 vdd.n10622 35.2919
R11002 vdd.n10624 vdd.n10623 35.2919
R11003 vdd.n10629 vdd.n10624 35.2919
R11004 vdd.n10658 vdd.n10651 35.2919
R11005 vdd.n10669 vdd.n10651 35.2919
R11006 vdd.n10670 vdd.n10669 35.2919
R11007 vdd.n10671 vdd.n10670 35.2919
R11008 vdd.n10672 vdd.n10671 35.2919
R11009 vdd.n10677 vdd.n10672 35.2919
R11010 vdd.n10704 vdd.n10697 35.2919
R11011 vdd.n10715 vdd.n10697 35.2919
R11012 vdd.n10716 vdd.n10715 35.2919
R11013 vdd.n10717 vdd.n10716 35.2919
R11014 vdd.n10718 vdd.n10717 35.2919
R11015 vdd.n10723 vdd.n10718 35.2919
R11016 vdd.n9768 vdd.n9767 35.2919
R11017 vdd.n9769 vdd.n9768 35.2919
R11018 vdd.n9770 vdd.n9769 35.2919
R11019 vdd.n9771 vdd.n9770 35.2919
R11020 vdd.n9771 vdd.n9746 35.2919
R11021 vdd.n9787 vdd.n9746 35.2919
R11022 vdd.n10799 vdd.n10792 35.2919
R11023 vdd.n10810 vdd.n10792 35.2919
R11024 vdd.n10811 vdd.n10810 35.2919
R11025 vdd.n10812 vdd.n10811 35.2919
R11026 vdd.n10813 vdd.n10812 35.2919
R11027 vdd.n10818 vdd.n10813 35.2919
R11028 vdd.n10753 vdd.n10746 35.2919
R11029 vdd.n10764 vdd.n10746 35.2919
R11030 vdd.n10765 vdd.n10764 35.2919
R11031 vdd.n10766 vdd.n10765 35.2919
R11032 vdd.n10767 vdd.n10766 35.2919
R11033 vdd.n10772 vdd.n10767 35.2919
R11034 vdd.n10846 vdd.n10839 35.2919
R11035 vdd.n10857 vdd.n10839 35.2919
R11036 vdd.n10858 vdd.n10857 35.2919
R11037 vdd.n10859 vdd.n10858 35.2919
R11038 vdd.n10860 vdd.n10859 35.2919
R11039 vdd.n10865 vdd.n10860 35.2919
R11040 vdd.n10894 vdd.n10887 35.2919
R11041 vdd.n10905 vdd.n10887 35.2919
R11042 vdd.n10906 vdd.n10905 35.2919
R11043 vdd.n10907 vdd.n10906 35.2919
R11044 vdd.n10908 vdd.n10907 35.2919
R11045 vdd.n10913 vdd.n10908 35.2919
R11046 vdd.n10940 vdd.n10933 35.2919
R11047 vdd.n10951 vdd.n10933 35.2919
R11048 vdd.n10952 vdd.n10951 35.2919
R11049 vdd.n10953 vdd.n10952 35.2919
R11050 vdd.n10954 vdd.n10953 35.2919
R11051 vdd.n10959 vdd.n10954 35.2919
R11052 vdd.n10990 vdd.n10981 35.2919
R11053 vdd.n10999 vdd.n10981 35.2919
R11054 vdd.n11000 vdd.n10999 35.2919
R11055 vdd.n11003 vdd.n11000 35.2919
R11056 vdd.n11003 vdd.n11002 35.2919
R11057 vdd.n11002 vdd.n10979 35.2919
R11058 vdd.n11035 vdd.n11026 35.2919
R11059 vdd.n11044 vdd.n11026 35.2919
R11060 vdd.n11045 vdd.n11044 35.2919
R11061 vdd.n11048 vdd.n11045 35.2919
R11062 vdd.n11048 vdd.n11047 35.2919
R11063 vdd.n11047 vdd.n11024 35.2919
R11064 vdd.n11085 vdd.n11076 35.2919
R11065 vdd.n11094 vdd.n11076 35.2919
R11066 vdd.n11095 vdd.n11094 35.2919
R11067 vdd.n11098 vdd.n11095 35.2919
R11068 vdd.n11098 vdd.n11097 35.2919
R11069 vdd.n11097 vdd.n11074 35.2919
R11070 vdd.n11131 vdd.n11122 35.2919
R11071 vdd.n11140 vdd.n11122 35.2919
R11072 vdd.n11141 vdd.n11140 35.2919
R11073 vdd.n11144 vdd.n11141 35.2919
R11074 vdd.n11144 vdd.n11143 35.2919
R11075 vdd.n11143 vdd.n11120 35.2919
R11076 vdd.n11179 vdd.n11170 35.2919
R11077 vdd.n11188 vdd.n11170 35.2919
R11078 vdd.n11189 vdd.n11188 35.2919
R11079 vdd.n11192 vdd.n11189 35.2919
R11080 vdd.n11192 vdd.n11191 35.2919
R11081 vdd.n11191 vdd.n11168 35.2919
R11082 vdd.n440 vdd.n438 35.2919
R11083 vdd.n444 vdd.n438 35.2919
R11084 vdd.n445 vdd.n444 35.2919
R11085 vdd.n448 vdd.n445 35.2919
R11086 vdd.n448 vdd.n447 35.2919
R11087 vdd.n447 vdd.n433 35.2919
R11088 vdd.n11226 vdd.n11217 35.2919
R11089 vdd.n11235 vdd.n11217 35.2919
R11090 vdd.n11236 vdd.n11235 35.2919
R11091 vdd.n11239 vdd.n11236 35.2919
R11092 vdd.n11239 vdd.n11238 35.2919
R11093 vdd.n11238 vdd.n11215 35.2919
R11094 vdd.n11271 vdd.n11262 35.2919
R11095 vdd.n11280 vdd.n11262 35.2919
R11096 vdd.n11281 vdd.n11280 35.2919
R11097 vdd.n11284 vdd.n11281 35.2919
R11098 vdd.n11284 vdd.n11283 35.2919
R11099 vdd.n11283 vdd.n11260 35.2919
R11100 vdd.n11317 vdd.n11308 35.2919
R11101 vdd.n11326 vdd.n11308 35.2919
R11102 vdd.n11327 vdd.n11326 35.2919
R11103 vdd.n11330 vdd.n11327 35.2919
R11104 vdd.n11330 vdd.n11329 35.2919
R11105 vdd.n11329 vdd.n11306 35.2919
R11106 vdd.n11368 vdd.n11359 35.2919
R11107 vdd.n11377 vdd.n11359 35.2919
R11108 vdd.n11378 vdd.n11377 35.2919
R11109 vdd.n11381 vdd.n11378 35.2919
R11110 vdd.n11381 vdd.n11380 35.2919
R11111 vdd.n11380 vdd.n11357 35.2919
R11112 vdd.n11414 vdd.n11405 35.2919
R11113 vdd.n11423 vdd.n11405 35.2919
R11114 vdd.n11424 vdd.n11423 35.2919
R11115 vdd.n11427 vdd.n11424 35.2919
R11116 vdd.n11427 vdd.n11426 35.2919
R11117 vdd.n11426 vdd.n11403 35.2919
R11118 vdd.n11462 vdd.n11453 35.2919
R11119 vdd.n11471 vdd.n11453 35.2919
R11120 vdd.n11472 vdd.n11471 35.2919
R11121 vdd.n11475 vdd.n11472 35.2919
R11122 vdd.n11475 vdd.n11474 35.2919
R11123 vdd.n11474 vdd.n11451 35.2919
R11124 vdd.n11508 vdd.n11499 35.2919
R11125 vdd.n11517 vdd.n11499 35.2919
R11126 vdd.n11518 vdd.n11517 35.2919
R11127 vdd.n11521 vdd.n11518 35.2919
R11128 vdd.n11521 vdd.n11520 35.2919
R11129 vdd.n11520 vdd.n11497 35.2919
R11130 vdd.n11553 vdd.n11544 35.2919
R11131 vdd.n11562 vdd.n11544 35.2919
R11132 vdd.n11563 vdd.n11562 35.2919
R11133 vdd.n11566 vdd.n11563 35.2919
R11134 vdd.n11566 vdd.n11565 35.2919
R11135 vdd.n11565 vdd.n11542 35.2919
R11136 vdd.n11603 vdd.n11594 35.2919
R11137 vdd.n11612 vdd.n11594 35.2919
R11138 vdd.n11613 vdd.n11612 35.2919
R11139 vdd.n11616 vdd.n11613 35.2919
R11140 vdd.n11616 vdd.n11615 35.2919
R11141 vdd.n11615 vdd.n11592 35.2919
R11142 vdd.n11649 vdd.n11640 35.2919
R11143 vdd.n11658 vdd.n11640 35.2919
R11144 vdd.n11659 vdd.n11658 35.2919
R11145 vdd.n11662 vdd.n11659 35.2919
R11146 vdd.n11662 vdd.n11661 35.2919
R11147 vdd.n11661 vdd.n11638 35.2919
R11148 vdd.n11697 vdd.n11688 35.2919
R11149 vdd.n11706 vdd.n11688 35.2919
R11150 vdd.n11707 vdd.n11706 35.2919
R11151 vdd.n11710 vdd.n11707 35.2919
R11152 vdd.n11710 vdd.n11709 35.2919
R11153 vdd.n11709 vdd.n11686 35.2919
R11154 vdd.n205 vdd.n203 35.2919
R11155 vdd.n209 vdd.n203 35.2919
R11156 vdd.n210 vdd.n209 35.2919
R11157 vdd.n213 vdd.n210 35.2919
R11158 vdd.n213 vdd.n212 35.2919
R11159 vdd.n212 vdd.n198 35.2919
R11160 vdd.n11744 vdd.n11735 35.2919
R11161 vdd.n11753 vdd.n11735 35.2919
R11162 vdd.n11754 vdd.n11753 35.2919
R11163 vdd.n11757 vdd.n11754 35.2919
R11164 vdd.n11757 vdd.n11756 35.2919
R11165 vdd.n11756 vdd.n11733 35.2919
R11166 vdd.n11789 vdd.n11780 35.2919
R11167 vdd.n11798 vdd.n11780 35.2919
R11168 vdd.n11799 vdd.n11798 35.2919
R11169 vdd.n11802 vdd.n11799 35.2919
R11170 vdd.n11802 vdd.n11801 35.2919
R11171 vdd.n11801 vdd.n11778 35.2919
R11172 vdd.n11839 vdd.n11830 35.2919
R11173 vdd.n11848 vdd.n11830 35.2919
R11174 vdd.n11849 vdd.n11848 35.2919
R11175 vdd.n11852 vdd.n11849 35.2919
R11176 vdd.n11852 vdd.n11851 35.2919
R11177 vdd.n11851 vdd.n11828 35.2919
R11178 vdd.n11885 vdd.n11876 35.2919
R11179 vdd.n11894 vdd.n11876 35.2919
R11180 vdd.n11895 vdd.n11894 35.2919
R11181 vdd.n11898 vdd.n11895 35.2919
R11182 vdd.n11898 vdd.n11897 35.2919
R11183 vdd.n11897 vdd.n11874 35.2919
R11184 vdd.n11933 vdd.n11924 35.2919
R11185 vdd.n11942 vdd.n11924 35.2919
R11186 vdd.n11943 vdd.n11942 35.2919
R11187 vdd.n11946 vdd.n11943 35.2919
R11188 vdd.n11946 vdd.n11945 35.2919
R11189 vdd.n11945 vdd.n11922 35.2919
R11190 vdd.n6637 vdd.t705 28.9836
R11191 vdd.n7623 vdd.t1274 28.9836
R11192 vdd.n7577 vdd.t887 28.9836
R11193 vdd.n7627 vdd.t224 28.9836
R11194 vdd.n7488 vdd.t932 28.9836
R11195 vdd.n7717 vdd.t252 28.9836
R11196 vdd.n7721 vdd.t1266 28.9836
R11197 vdd.n7445 vdd.t444 28.9836
R11198 vdd.n7391 vdd.t1254 28.9836
R11199 vdd.n7906 vdd.t519 28.9836
R11200 vdd.n7813 vdd.t240 28.9836
R11201 vdd.n7859 vdd.t542 28.9836
R11202 vdd.n7910 vdd.t69 28.9836
R11203 vdd.n7345 vdd.t1093 28.9836
R11204 vdd.n8000 vdd.t320 28.9836
R11205 vdd.n8004 vdd.t963 28.9836
R11206 vdd.n7299 vdd.t533 28.9836
R11207 vdd.n8141 vdd.t644 28.9836
R11208 vdd.n8095 vdd.t131 28.9836
R11209 vdd.n8145 vdd.t326 28.9836
R11210 vdd.n7253 vdd.t884 28.9836
R11211 vdd.n8235 vdd.t249 28.9836
R11212 vdd.n8239 vdd.t1449 28.9836
R11213 vdd.n7210 vdd.t1395 28.9836
R11214 vdd.n7156 vdd.t184 28.9836
R11215 vdd.n8377 vdd.t1177 28.9836
R11216 vdd.n8331 vdd.t451 28.9836
R11217 vdd.n8381 vdd.t880 28.9836
R11218 vdd.n7110 vdd.t522 28.9836
R11219 vdd.n8471 vdd.t1421 28.9836
R11220 vdd.n8475 vdd.t1065 28.9836
R11221 vdd.n8565 vdd.t1453 28.9836
R11222 vdd.n8658 vdd.t1081 28.9836
R11223 vdd.n8612 vdd.t763 28.9836
R11224 vdd.n8705 vdd.t256 28.9836
R11225 vdd.n7107 vdd.t304 28.9836
R11226 vdd.n8752 vdd.t935 28.9836
R11227 vdd.n8799 vdd.t189 28.9836
R11228 vdd.n7045 vdd.t81 28.9836
R11229 vdd.n7009 vdd.t808 28.9836
R11230 vdd.n8941 vdd.t138 28.9836
R11231 vdd.n8894 vdd.t586 28.9836
R11232 vdd.n8848 vdd.t1200 28.9836
R11233 vdd.n8988 vdd.t757 28.9836
R11234 vdd.n6963 vdd.t982 28.9836
R11235 vdd.n9035 vdd.t639 28.9836
R11236 vdd.n9082 vdd.t1525 28.9836
R11237 vdd.n6917 vdd.t219 28.9836
R11238 vdd.n9176 vdd.t79 28.9836
R11239 vdd.n9130 vdd.t784 28.9836
R11240 vdd.n9223 vdd.t1269 28.9836
R11241 vdd.n6871 vdd.t154 28.9836
R11242 vdd.n9270 vdd.t746 28.9836
R11243 vdd.n9317 vdd.t400 28.9836
R11244 vdd.n6809 vdd.t692 28.9836
R11245 vdd.n6773 vdd.t626 28.9836
R11246 vdd.n9412 vdd.t178 28.9836
R11247 vdd.n9366 vdd.t1030 28.9836
R11248 vdd.n9459 vdd.t545 28.9836
R11249 vdd.n6727 vdd.t364 28.9836
R11250 vdd.n9506 vdd.t663 28.9836
R11251 vdd.n9553 vdd.t1520 28.9836
R11252 vdd.n3623 vdd.t1035 28.9836
R11253 vdd.n4609 vdd.t697 28.9836
R11254 vdd.n4563 vdd.t448 28.9836
R11255 vdd.n4613 vdd.t150 28.9836
R11256 vdd.n4474 vdd.t1232 28.9836
R11257 vdd.n4703 vdd.t669 28.9836
R11258 vdd.n4707 vdd.t471 28.9836
R11259 vdd.n4431 vdd.t1240 28.9836
R11260 vdd.n4377 vdd.t1436 28.9836
R11261 vdd.n4892 vdd.t228 28.9836
R11262 vdd.n4799 vdd.t366 28.9836
R11263 vdd.n4845 vdd.t415 28.9836
R11264 vdd.n4896 vdd.t1228 28.9836
R11265 vdd.n4331 vdd.t1425 28.9836
R11266 vdd.n4986 vdd.t511 28.9836
R11267 vdd.n4990 vdd.t1100 28.9836
R11268 vdd.n4285 vdd.t420 28.9836
R11269 vdd.n5127 vdd.t1168 28.9836
R11270 vdd.n5081 vdd.t108 28.9836
R11271 vdd.n5131 vdd.t345 28.9836
R11272 vdd.n4239 vdd.t1184 28.9836
R11273 vdd.n5221 vdd.t323 28.9836
R11274 vdd.n5225 vdd.t701 28.9836
R11275 vdd.n4196 vdd.t711 28.9836
R11276 vdd.n4142 vdd.t622 28.9836
R11277 vdd.n5363 vdd.t1110 28.9836
R11278 vdd.n5317 vdd.t1504 28.9836
R11279 vdd.n5367 vdd.t720 28.9836
R11280 vdd.n4096 vdd.t395 28.9836
R11281 vdd.n5457 vdd.t501 28.9836
R11282 vdd.n5461 vdd.t505 28.9836
R11283 vdd.n5551 vdd.t761 28.9836
R11284 vdd.n5644 vdd.t715 28.9836
R11285 vdd.n5598 vdd.t187 28.9836
R11286 vdd.n5691 vdd.t398 28.9836
R11287 vdd.n4093 vdd.t1409 28.9836
R11288 vdd.n5738 vdd.t1216 28.9836
R11289 vdd.n5785 vdd.t582 28.9836
R11290 vdd.n4031 vdd.t1516 28.9836
R11291 vdd.n3995 vdd.t1209 28.9836
R11292 vdd.n5927 vdd.t329 28.9836
R11293 vdd.n5880 vdd.t1529 28.9836
R11294 vdd.n5834 vdd.t779 28.9836
R11295 vdd.n5974 vdd.t678 28.9836
R11296 vdd.n3949 vdd.t1134 28.9836
R11297 vdd.n6021 vdd.t1194 28.9836
R11298 vdd.n6068 vdd.t1 28.9836
R11299 vdd.n3903 vdd.t1281 28.9836
R11300 vdd.n6162 vdd.t633 28.9836
R11301 vdd.n6116 vdd.t1205 28.9836
R11302 vdd.n6209 vdd.t1159 28.9836
R11303 vdd.n3857 vdd.t194 28.9836
R11304 vdd.n6256 vdd.t1405 28.9836
R11305 vdd.n6303 vdd.t946 28.9836
R11306 vdd.n3795 vdd.t723 28.9836
R11307 vdd.n3759 vdd.t682 28.9836
R11308 vdd.n6398 vdd.t19 28.9836
R11309 vdd.n6352 vdd.t751 28.9836
R11310 vdd.n6445 vdd.t685 28.9836
R11311 vdd.n3713 vdd.t476 28.9836
R11312 vdd.n6492 vdd.t1171 28.9836
R11313 vdd.n6539 vdd.t120 28.9836
R11314 vdd.n609 vdd.t349 28.9836
R11315 vdd.n1595 vdd.t1223 28.9836
R11316 vdd.n1549 vdd.t1189 28.9836
R11317 vdd.n1599 vdd.t1069 28.9836
R11318 vdd.n1460 vdd.t410 28.9836
R11319 vdd.n1689 vdd.t954 28.9836
R11320 vdd.n1693 vdd.t84 28.9836
R11321 vdd.n1417 vdd.t1073 28.9836
R11322 vdd.n1363 vdd.t919 28.9836
R11323 vdd.n1878 vdd.t665 28.9836
R11324 vdd.n1785 vdd.t369 28.9836
R11325 vdd.n1831 vdd.t655 28.9836
R11326 vdd.n1882 vdd.t788 28.9836
R11327 vdd.n1317 vdd.t312 28.9836
R11328 vdd.n1972 vdd.t389 28.9836
R11329 vdd.n1976 vdd.t159 28.9836
R11330 vdd.n1271 vdd.t1104 28.9836
R11331 vdd.n2113 vdd.t1219 28.9836
R11332 vdd.n2067 vdd.t842 28.9836
R11333 vdd.n2117 vdd.t636 28.9836
R11334 vdd.n1225 vdd.t1369 28.9836
R11335 vdd.n2207 vdd.t233 28.9836
R11336 vdd.n2211 vdd.t1117 28.9836
R11337 vdd.n1182 vdd.t673 28.9836
R11338 vdd.n1128 vdd.t732 28.9836
R11339 vdd.n2349 vdd.t297 28.9836
R11340 vdd.n2303 vdd.t117 28.9836
R11341 vdd.n2353 vdd.t1039 28.9836
R11342 vdd.n1082 vdd.t112 28.9836
R11343 vdd.n2443 vdd.t876 28.9836
R11344 vdd.n2447 vdd.t1445 28.9836
R11345 vdd.n2537 vdd.t180 28.9836
R11346 vdd.n2630 vdd.t525 28.9836
R11347 vdd.n2584 vdd.t333 28.9836
R11348 vdd.n2677 vdd.t617 28.9836
R11349 vdd.n1079 vdd.t956 28.9836
R11350 vdd.n2724 vdd.t1097 28.9836
R11351 vdd.n2771 vdd.t1140 28.9836
R11352 vdd.n1017 vdd.t403 28.9836
R11353 vdd.n981 vdd.t922 28.9836
R11354 vdd.n2913 vdd.t74 28.9836
R11355 vdd.n2866 vdd.t135 28.9836
R11356 vdd.n2820 vdd.t613 28.9836
R11357 vdd.n2960 vdd.t221 28.9836
R11358 vdd.n935 vdd.t214 28.9836
R11359 vdd.n3007 vdd.t1385 28.9836
R11360 vdd.n3054 vdd.t453 28.9836
R11361 vdd.n889 vdd.t426 28.9836
R11362 vdd.n3148 vdd.t800 28.9836
R11363 vdd.n3102 vdd.t275 28.9836
R11364 vdd.n3195 vdd.t279 28.9836
R11365 vdd.n843 vdd.t290 28.9836
R11366 vdd.n3242 vdd.t1211 28.9836
R11367 vdd.n3289 vdd.t1276 28.9836
R11368 vdd.n781 vdd.t1432 28.9836
R11369 vdd.n745 vdd.t125 28.9836
R11370 vdd.n3384 vdd.t267 28.9836
R11371 vdd.n3338 vdd.t1510 28.9836
R11372 vdd.n3431 vdd.t1136 28.9836
R11373 vdd.n699 vdd.t48 28.9836
R11374 vdd.n3478 vdd.t650 28.9836
R11375 vdd.n3525 vdd.t832 28.9836
R11376 vdd.n9648 vdd.t911 28.9836
R11377 vdd.n9602 vdd.t1115 28.9836
R11378 vdd.n6634 vdd.t708 28.9836
R11379 vdd.n6588 vdd.t551 28.9836
R11380 vdd.n3620 vdd.t1430 28.9836
R11381 vdd.n3574 vdd.t1174 28.9836
R11382 vdd.n606 vdd.t1152 28.9836
R11383 vdd.n90 vdd.t244 28.9836
R11384 vdd.n44 vdd.t652 28.9836
R11385 vdd.n10120 vdd.t1086 28.9836
R11386 vdd.n10074 vdd.t339 28.9836
R11387 vdd.n10167 vdd.t782 28.9836
R11388 vdd.n10214 vdd.t1022 28.9836
R11389 vdd.n10012 vdd.t1399 28.9836
R11390 vdd.n9976 vdd.t61 28.9836
R11391 vdd.n10356 vdd.t689 28.9836
R11392 vdd.n10309 vdd.t301 28.9836
R11393 vdd.n10263 vdd.t1418 28.9836
R11394 vdd.n10403 vdd.t356 28.9836
R11395 vdd.n9930 vdd.t258 28.9836
R11396 vdd.n10450 vdd.t1402 28.9836
R11397 vdd.n10497 vdd.t805 28.9836
R11398 vdd.n9884 vdd.t1181 28.9836
R11399 vdd.n10591 vdd.t1262 28.9836
R11400 vdd.n10545 vdd.t263 28.9836
R11401 vdd.n10638 vdd.t1076 28.9836
R11402 vdd.n9838 vdd.t726 28.9836
R11403 vdd.n10685 vdd.t609 28.9836
R11404 vdd.n10732 vdd.t148 28.9836
R11405 vdd.n9776 vdd.t1365 28.9836
R11406 vdd.n9740 vdd.t1389 28.9836
R11407 vdd.n10827 vdd.t1236 28.9836
R11408 vdd.n10781 vdd.t1246 28.9836
R11409 vdd.n10874 vdd.t1161 28.9836
R11410 vdd.n9694 vdd.t1513 28.9836
R11411 vdd.n10921 vdd.t950 28.9836
R11412 vdd.n10968 vdd.t1198 28.9836
R11413 vdd.n518 vdd.t128 28.9836
R11414 vdd.n11063 vdd.t287 28.9836
R11415 vdd.n11017 vdd.t646 28.9836
R11416 vdd.n11067 vdd.t734 28.9836
R11417 vdd.n472 vdd.t926 28.9836
R11418 vdd.n11157 vdd.t295 28.9836
R11419 vdd.n11161 vdd.t351 28.9836
R11420 vdd.n429 vdd.t741 28.9836
R11421 vdd.n375 vdd.t1414 28.9836
R11422 vdd.n11346 vdd.t515 28.9836
R11423 vdd.n11253 vdd.t890 28.9836
R11424 vdd.n11299 vdd.t406 28.9836
R11425 vdd.n11350 vdd.t1146 28.9836
R11426 vdd.n329 vdd.t573 28.9836
R11427 vdd.n11440 vdd.t283 28.9836
R11428 vdd.n11444 vdd.t1522 28.9836
R11429 vdd.n283 vdd.t162 28.9836
R11430 vdd.n11581 vdd.t271 28.9836
R11431 vdd.n11535 vdd.t1440 28.9836
R11432 vdd.n11585 vdd.t1391 28.9836
R11433 vdd.n237 vdd.t737 28.9836
R11434 vdd.n11675 vdd.t1249 28.9836
R11435 vdd.n11679 vdd.t529 28.9836
R11436 vdd.n194 vdd.t142 28.9836
R11437 vdd.n140 vdd.t914 28.9836
R11438 vdd.n11817 vdd.t358 28.9836
R11439 vdd.n11771 vdd.t105 28.9836
R11440 vdd.n11821 vdd.t317 28.9836
R11441 vdd.n94 vdd.t508 28.9836
R11442 vdd.n11911 vdd.t753 28.9836
R11443 vdd.n11915 vdd.t341 28.9836
R11444 vdd.n12006 vdd.t1084 28.9836
R11445 vdd.n6636 vdd.t485 28.9065
R11446 vdd.n7624 vdd.t899 28.9065
R11447 vdd.n7576 vdd.t167 28.9065
R11448 vdd.n7626 vdd.t590 28.9065
R11449 vdd.n7487 vdd.t1327 28.9065
R11450 vdd.n7718 vdd.t863 28.9065
R11451 vdd.n7720 vdd.t1343 28.9065
R11452 vdd.n7437 vdd.t1155 28.9065
R11453 vdd.n7390 vdd.t380 28.9065
R11454 vdd.n7907 vdd.t897 28.9065
R11455 vdd.n7812 vdd.t838 28.9065
R11456 vdd.n7858 vdd.t1376 28.9065
R11457 vdd.n7909 vdd.t487 28.9065
R11458 vdd.n7344 vdd.t594 28.9065
R11459 vdd.n8001 vdd.t873 28.9065
R11460 vdd.n8003 vdd.t1331 28.9065
R11461 vdd.n7298 vdd.t1361 28.9065
R11462 vdd.n8142 vdd.t37 28.9065
R11463 vdd.n8094 vdd.t836 28.9065
R11464 vdd.n8144 vdd.t202 28.9065
R11465 vdd.n7252 vdd.t1050 28.9065
R11466 vdd.n8236 vdd.t974 28.9065
R11467 vdd.n8238 vdd.t1347 28.9065
R11468 vdd.n7202 vdd.t1460 28.9065
R11469 vdd.n7155 vdd.t1311 28.9065
R11470 vdd.n8378 vdd.t855 28.9065
R11471 vdd.n8330 vdd.t57 28.9065
R11472 vdd.n8380 vdd.t10 28.9065
R11473 vdd.n7109 vdd.t1464 28.9065
R11474 vdd.n8472 vdd.t41 28.9065
R11475 vdd.n8474 vdd.t212 28.9065
R11476 vdd.n8564 vdd.t483 28.9065
R11477 vdd.n8659 vdd.t849 28.9065
R11478 vdd.n8611 vdd.t774 28.9065
R11479 vdd.n8704 vdd.t1315 28.9065
R11480 vdd.n7106 vdd.t588 28.9065
R11481 vdd.n8753 vdd.t857 28.9065
R11482 vdd.n8798 vdd.t1468 28.9065
R11483 vdd.n7012 vdd.t98 28.9065
R11484 vdd.n7008 vdd.t378 28.9065
R11485 vdd.n8942 vdd.t826 28.9065
R11486 vdd.n8893 vdd.t766 28.9065
R11487 vdd.n8847 vdd.t1130 28.9065
R11488 vdd.n8987 vdd.t459 28.9065
R11489 vdd.n6962 vdd.t559 28.9065
R11490 vdd.n9036 vdd.t865 28.9065
R11491 vdd.n9081 vdd.t1478 28.9065
R11492 vdd.n6916 vdd.t206 28.9065
R11493 vdd.n9177 vdd.t1007 28.9065
R11494 vdd.n9129 vdd.t431 28.9065
R11495 vdd.n9222 vdd.t567 28.9065
R11496 vdd.n6870 vdd.t1319 28.9065
R11497 vdd.n9271 vdd.t43 28.9065
R11498 vdd.n9316 vdd.t1303 28.9065
R11499 vdd.n6776 vdd.t90 28.9065
R11500 vdd.n6772 vdd.t208 28.9065
R11501 vdd.n9413 vdd.t989 28.9065
R11502 vdd.n9365 vdd.t628 28.9065
R11503 vdd.n9458 vdd.t602 28.9065
R11504 vdd.n6726 vdd.t1289 28.9065
R11505 vdd.n9507 vdd.t861 28.9065
R11506 vdd.n9552 vdd.t1042 28.9065
R11507 vdd.n3622 vdd.t561 28.9065
R11508 vdd.n4610 vdd.t1001 28.9065
R11509 vdd.n4562 vdd.t175 28.9065
R11510 vdd.n4612 vdd.t198 28.9065
R11511 vdd.n4473 vdd.t1046 28.9065
R11512 vdd.n4704 vdd.t35 28.9065
R11513 vdd.n4706 vdd.t1474 28.9065
R11514 vdd.n4423 vdd.t1458 28.9065
R11515 vdd.n4376 vdd.t571 28.9065
R11516 vdd.n4893 vdd.t828 28.9065
R11517 vdd.n4798 vdd.t53 28.9065
R11518 vdd.n4844 vdd.t1372 28.9065
R11519 vdd.n4895 vdd.t1488 28.9065
R11520 vdd.n4330 vdd.t1056 28.9065
R11521 vdd.n4987 vdd.t859 28.9065
R11522 vdd.n4989 vdd.t1301 28.9065
R11523 vdd.n4284 vdd.t1317 28.9065
R11524 vdd.n5128 vdd.t1011 28.9065
R11525 vdd.n5080 vdd.t51 28.9065
R11526 vdd.n5130 vdd.t1044 28.9065
R11527 vdd.n4238 vdd.t1291 28.9065
R11528 vdd.n5222 vdd.t943 28.9065
R11529 vdd.n5224 vdd.t1305 28.9065
R11530 vdd.n4188 vdd.t1456 28.9065
R11531 vdd.n4141 vdd.t555 28.9065
R11532 vdd.n5364 vdd.t845 28.9065
R11533 vdd.n5316 vdd.t173 28.9065
R11534 vdd.n5366 vdd.t457 28.9065
R11535 vdd.n4095 vdd.t204 28.9065
R11536 vdd.n5458 vdd.t1013 28.9065
R11537 vdd.n5460 vdd.t1052 28.9065
R11538 vdd.n5550 vdd.t557 28.9065
R11539 vdd.n5645 vdd.t907 28.9065
R11540 vdd.n5597 vdd.t165 28.9065
R11541 vdd.n5690 vdd.t596 28.9065
R11542 vdd.n4092 vdd.t469 28.9065
R11543 vdd.n5739 vdd.t991 28.9065
R11544 vdd.n5784 vdd.t14 28.9065
R11545 vdd.n3998 vdd.t100 28.9065
R11546 vdd.n3994 vdd.t604 28.9065
R11547 vdd.n5928 vdd.t867 28.9065
R11548 vdd.n5879 vdd.t768 28.9065
R11549 vdd.n5833 vdd.t1374 28.9065
R11550 vdd.n5973 vdd.t1480 28.9065
R11551 vdd.n3948 vdd.t1058 28.9065
R11552 vdd.n6022 vdd.t1003 28.9065
R11553 vdd.n6067 vdd.t1490 28.9065
R11554 vdd.n3902 vdd.t461 28.9065
R11555 vdd.n6163 vdd.t970 28.9065
R11556 vdd.n6115 vdd.t435 28.9065
R11557 vdd.n6208 vdd.t1337 28.9065
R11558 vdd.n3856 vdd.t600 28.9065
R11559 vdd.n6257 vdd.t33 28.9065
R11560 vdd.n6302 vdd.t497 28.9065
R11561 vdd.n3762 vdd.t94 28.9065
R11562 vdd.n3758 vdd.t465 28.9065
R11563 vdd.n6399 vdd.t869 28.9065
R11564 vdd.n6351 vdd.t433 28.9065
R11565 vdd.n6444 vdd.t1054 28.9065
R11566 vdd.n3712 vdd.t1484 28.9065
R11567 vdd.n6493 vdd.t895 28.9065
R11568 vdd.n6538 vdd.t565 28.9065
R11569 vdd.n608 vdd.t553 28.9065
R11570 vdd.n1596 vdd.t824 28.9065
R11571 vdd.n1548 vdd.t834 28.9065
R11572 vdd.n1598 vdd.t467 28.9065
R11573 vdd.n1459 vdd.t386 28.9065
R11574 vdd.n1690 vdd.t999 28.9065
R11575 vdd.n1692 vdd.t1494 28.9065
R11576 vdd.n1409 vdd.t102 28.9065
R11577 vdd.n1362 vdd.t592 28.9065
R11578 vdd.n1879 vdd.t871 28.9065
R11579 vdd.n1784 vdd.t171 28.9065
R11580 vdd.n1830 vdd.t1128 28.9065
R11581 vdd.n1881 vdd.t1325 28.9065
R11582 vdd.n1316 vdd.t1357 28.9065
R11583 vdd.n1973 vdd.t993 28.9065
R11584 vdd.n1975 vdd.t372 28.9065
R11585 vdd.n1270 vdd.t1496 28.9065
R11586 vdd.n2114 vdd.t972 28.9065
R11587 vdd.n2066 vdd.t169 28.9065
R11588 vdd.n2116 vdd.t1345 28.9065
R11589 vdd.n1224 vdd.t1309 28.9065
R11590 vdd.n2208 vdd.t941 28.9065
R11591 vdd.n2210 vdd.t1482 28.9065
R11592 vdd.n1174 vdd.t96 28.9065
R11593 vdd.n1127 vdd.t196 28.9065
R11594 vdd.n2350 vdd.t901 28.9065
R11595 vdd.n2302 vdd.t772 28.9065
R11596 vdd.n2352 vdd.t493 28.9065
R11597 vdd.n1081 vdd.t4 28.9065
R11598 vdd.n2444 vdd.t976 28.9065
R11599 vdd.n2446 vdd.t1349 28.9065
R11600 vdd.n2536 vdd.t382 28.9065
R11601 vdd.n2631 vdd.t816 28.9065
R11602 vdd.n2583 vdd.t770 28.9065
R11603 vdd.n2676 vdd.t1351 28.9065
R11604 vdd.n1078 vdd.t1470 28.9065
R11605 vdd.n2725 vdd.t1017 28.9065
R11606 vdd.n2770 vdd.t495 28.9065
R11607 vdd.n984 vdd.t92 28.9065
R11608 vdd.n980 vdd.t463 28.9065
R11609 vdd.n2914 vdd.t45 28.9065
R11610 vdd.n2865 vdd.t439 28.9065
R11611 vdd.n2819 vdd.t1126 28.9065
R11612 vdd.n2959 vdd.t12 28.9065
R11613 vdd.n934 vdd.t1313 28.9065
R11614 vdd.n3008 vdd.t39 28.9065
R11615 vdd.n3053 vdd.t1297 28.9065
R11616 vdd.n888 vdd.t1498 28.9065
R11617 vdd.n3149 vdd.t853 28.9065
R11618 vdd.n3101 vdd.t791 28.9065
R11619 vdd.n3194 vdd.t374 28.9065
R11620 vdd.n842 vdd.t1359 28.9065
R11621 vdd.n3243 vdd.t968 28.9065
R11622 vdd.n3288 vdd.t1329 28.9065
R11623 vdd.n748 vdd.t88 28.9065
R11624 vdd.n744 vdd.t1502 28.9065
R11625 vdd.n3385 vdd.t820 28.9065
R11626 vdd.n3337 vdd.t437 28.9065
R11627 vdd.n3430 vdd.t1333 28.9065
R11628 vdd.n698 vdd.t1466 28.9065
R11629 vdd.n3479 vdd.t905 28.9065
R11630 vdd.n3524 vdd.t489 28.9065
R11631 vdd.n9649 vdd.t27 28.9065
R11632 vdd.n9603 vdd.t985 28.9065
R11633 vdd.n6635 vdd.t29 28.9065
R11634 vdd.n6589 vdd.t1187 28.9065
R11635 vdd.n3621 vdd.t25 28.9065
R11636 vdd.n3575 vdd.t987 28.9065
R11637 vdd.n607 vdd.t31 28.9065
R11638 vdd.n91 vdd.t1009 28.9065
R11639 vdd.n43 vdd.t840 28.9065
R11640 vdd.n10119 vdd.t569 28.9065
R11641 vdd.n10073 vdd.t1335 28.9065
R11642 vdd.n10168 vdd.t909 28.9065
R11643 vdd.n10213 vdd.t598 28.9065
R11644 vdd.n9979 vdd.t576 28.9065
R11645 vdd.n9975 vdd.t491 28.9065
R11646 vdd.n10357 vdd.t939 28.9065
R11647 vdd.n10308 vdd.t55 28.9065
R11648 vdd.n10262 vdd.t1380 28.9065
R11649 vdd.n10402 vdd.t384 28.9065
R11650 vdd.n9929 vdd.t16 28.9065
R11651 vdd.n10451 vdd.t847 28.9065
R11652 vdd.n10496 vdd.t1307 28.9065
R11653 vdd.n9883 vdd.t1060 28.9065
R11654 vdd.n10592 vdd.t1005 28.9065
R11655 vdd.n10544 vdd.t776 28.9065
R11656 vdd.n10637 vdd.t1492 28.9065
R11657 vdd.n9837 vdd.t479 28.9065
R11658 vdd.n10686 vdd.t818 28.9065
R11659 vdd.n10731 vdd.t1353 28.9065
R11660 vdd.n9743 vdd.t1462 28.9065
R11661 vdd.n9739 vdd.t1323 28.9065
R11662 vdd.n10828 vdd.t903 28.9065
R11663 vdd.n10780 vdd.t630 28.9065
R11664 vdd.n10873 vdd.t481 28.9065
R11665 vdd.n9693 vdd.t1355 28.9065
R11666 vdd.n10922 vdd.t937 28.9065
R11667 vdd.n10967 vdd.t6 28.9065
R11668 vdd.n517 vdd.t376 28.9065
R11669 vdd.n11064 vdd.t822 28.9065
R11670 vdd.n11016 vdd.t59 28.9065
R11671 vdd.n11066 vdd.t1500 28.9065
R11672 vdd.n471 vdd.t210 28.9065
R11673 vdd.n11158 vdd.t997 28.9065
R11674 vdd.n11160 vdd.t1295 28.9065
R11675 vdd.n421 vdd.t580 28.9065
R11676 vdd.n374 vdd.t1486 28.9065
R11677 vdd.n11347 vdd.t966 28.9065
R11678 vdd.n11252 vdd.t797 28.9065
R11679 vdd.n11298 vdd.t1378 28.9065
R11680 vdd.n11349 vdd.t200 28.9065
R11681 vdd.n328 vdd.t1299 28.9065
R11682 vdd.n11441 vdd.t851 28.9065
R11683 vdd.n11443 vdd.t1341 28.9065
R11684 vdd.n282 vdd.t563 28.9065
R11685 vdd.n11582 vdd.t812 28.9065
R11686 vdd.n11534 vdd.t795 28.9065
R11687 vdd.n11584 vdd.t1287 28.9065
R11688 vdd.n236 vdd.t1476 28.9065
R11689 vdd.n11676 vdd.t995 28.9065
R11690 vdd.n11678 vdd.t1339 28.9065
R11691 vdd.n186 vdd.t578 28.9065
R11692 vdd.n139 vdd.t8 28.9065
R11693 vdd.n11818 vdd.t1015 28.9065
R11694 vdd.n11770 vdd.t793 28.9065
R11695 vdd.n11820 vdd.t1321 28.9065
R11696 vdd.n93 vdd.t1048 28.9065
R11697 vdd.n11912 vdd.t814 28.9065
R11698 vdd.n11914 vdd.t1293 28.9065
R11699 vdd.n12005 vdd.t1472 28.9065
R11700 vdd.n11975 vdd.n11974 16.2531
R11701 vdd.n11983 vdd.n11975 16.2531
R11702 vdd.n12004 vdd.n11983 16.2531
R11703 vdd.n12004 vdd.n12003 16.2531
R11704 vdd.n12003 vdd.n11994 16.2531
R11705 vdd.n11994 vdd.n11993 16.2531
R11706 vdd.n116 vdd.n115 16.2531
R11707 vdd.n115 vdd.n96 16.2531
R11708 vdd.n137 vdd.n96 16.2531
R11709 vdd.n137 vdd.n136 16.2531
R11710 vdd.n136 vdd.n97 16.2531
R11711 vdd.n132 vdd.n97 16.2531
R11712 vdd.n162 vdd.n161 16.2531
R11713 vdd.n161 vdd.n142 16.2531
R11714 vdd.n183 vdd.n142 16.2531
R11715 vdd.n183 vdd.n182 16.2531
R11716 vdd.n182 vdd.n143 16.2531
R11717 vdd.n178 vdd.n143 16.2531
R11718 vdd.n259 vdd.n258 16.2531
R11719 vdd.n258 vdd.n239 16.2531
R11720 vdd.n280 vdd.n239 16.2531
R11721 vdd.n280 vdd.n279 16.2531
R11722 vdd.n279 vdd.n240 16.2531
R11723 vdd.n275 vdd.n240 16.2531
R11724 vdd.n305 vdd.n304 16.2531
R11725 vdd.n304 vdd.n285 16.2531
R11726 vdd.n326 vdd.n285 16.2531
R11727 vdd.n326 vdd.n325 16.2531
R11728 vdd.n325 vdd.n286 16.2531
R11729 vdd.n321 vdd.n286 16.2531
R11730 vdd.n351 vdd.n350 16.2531
R11731 vdd.n350 vdd.n331 16.2531
R11732 vdd.n372 vdd.n331 16.2531
R11733 vdd.n372 vdd.n371 16.2531
R11734 vdd.n371 vdd.n332 16.2531
R11735 vdd.n367 vdd.n332 16.2531
R11736 vdd.n397 vdd.n396 16.2531
R11737 vdd.n396 vdd.n377 16.2531
R11738 vdd.n418 vdd.n377 16.2531
R11739 vdd.n418 vdd.n417 16.2531
R11740 vdd.n417 vdd.n378 16.2531
R11741 vdd.n413 vdd.n378 16.2531
R11742 vdd.n494 vdd.n493 16.2531
R11743 vdd.n493 vdd.n474 16.2531
R11744 vdd.n515 vdd.n474 16.2531
R11745 vdd.n515 vdd.n514 16.2531
R11746 vdd.n514 vdd.n475 16.2531
R11747 vdd.n510 vdd.n475 16.2531
R11748 vdd.n540 vdd.n539 16.2531
R11749 vdd.n539 vdd.n520 16.2531
R11750 vdd.n561 vdd.n520 16.2531
R11751 vdd.n561 vdd.n560 16.2531
R11752 vdd.n560 vdd.n521 16.2531
R11753 vdd.n556 vdd.n521 16.2531
R11754 vdd.n6705 vdd.n6704 16.2531
R11755 vdd.n6704 vdd.n6684 16.2531
R11756 vdd.n6725 vdd.n6684 16.2531
R11757 vdd.n6725 vdd.n6724 16.2531
R11758 vdd.n6724 vdd.n6685 16.2531
R11759 vdd.n6714 vdd.n6685 16.2531
R11760 vdd.n6751 vdd.n6750 16.2531
R11761 vdd.n6750 vdd.n6730 16.2531
R11762 vdd.n6771 vdd.n6730 16.2531
R11763 vdd.n6771 vdd.n6770 16.2531
R11764 vdd.n6770 vdd.n6731 16.2531
R11765 vdd.n6760 vdd.n6731 16.2531
R11766 vdd.n6849 vdd.n6848 16.2531
R11767 vdd.n6848 vdd.n6828 16.2531
R11768 vdd.n6869 vdd.n6828 16.2531
R11769 vdd.n6869 vdd.n6868 16.2531
R11770 vdd.n6868 vdd.n6829 16.2531
R11771 vdd.n6858 vdd.n6829 16.2531
R11772 vdd.n6895 vdd.n6894 16.2531
R11773 vdd.n6894 vdd.n6874 16.2531
R11774 vdd.n6915 vdd.n6874 16.2531
R11775 vdd.n6915 vdd.n6914 16.2531
R11776 vdd.n6914 vdd.n6875 16.2531
R11777 vdd.n6904 vdd.n6875 16.2531
R11778 vdd.n6941 vdd.n6940 16.2531
R11779 vdd.n6940 vdd.n6920 16.2531
R11780 vdd.n6961 vdd.n6920 16.2531
R11781 vdd.n6961 vdd.n6960 16.2531
R11782 vdd.n6960 vdd.n6921 16.2531
R11783 vdd.n6950 vdd.n6921 16.2531
R11784 vdd.n6987 vdd.n6986 16.2531
R11785 vdd.n6986 vdd.n6966 16.2531
R11786 vdd.n7007 vdd.n6966 16.2531
R11787 vdd.n7007 vdd.n7006 16.2531
R11788 vdd.n7006 vdd.n6967 16.2531
R11789 vdd.n6996 vdd.n6967 16.2531
R11790 vdd.n7085 vdd.n7084 16.2531
R11791 vdd.n7084 vdd.n7064 16.2531
R11792 vdd.n7105 vdd.n7064 16.2531
R11793 vdd.n7105 vdd.n7104 16.2531
R11794 vdd.n7104 vdd.n7065 16.2531
R11795 vdd.n7094 vdd.n7065 16.2531
R11796 vdd.n8543 vdd.n8542 16.2531
R11797 vdd.n8542 vdd.n8522 16.2531
R11798 vdd.n8563 vdd.n8522 16.2531
R11799 vdd.n8563 vdd.n8562 16.2531
R11800 vdd.n8562 vdd.n8523 16.2531
R11801 vdd.n8552 vdd.n8523 16.2531
R11802 vdd.n7132 vdd.n7131 16.2531
R11803 vdd.n7131 vdd.n7112 16.2531
R11804 vdd.n7153 vdd.n7112 16.2531
R11805 vdd.n7153 vdd.n7152 16.2531
R11806 vdd.n7152 vdd.n7113 16.2531
R11807 vdd.n7148 vdd.n7113 16.2531
R11808 vdd.n7178 vdd.n7177 16.2531
R11809 vdd.n7177 vdd.n7158 16.2531
R11810 vdd.n7199 vdd.n7158 16.2531
R11811 vdd.n7199 vdd.n7198 16.2531
R11812 vdd.n7198 vdd.n7159 16.2531
R11813 vdd.n7194 vdd.n7159 16.2531
R11814 vdd.n7275 vdd.n7274 16.2531
R11815 vdd.n7274 vdd.n7255 16.2531
R11816 vdd.n7296 vdd.n7255 16.2531
R11817 vdd.n7296 vdd.n7295 16.2531
R11818 vdd.n7295 vdd.n7256 16.2531
R11819 vdd.n7291 vdd.n7256 16.2531
R11820 vdd.n7321 vdd.n7320 16.2531
R11821 vdd.n7320 vdd.n7301 16.2531
R11822 vdd.n7342 vdd.n7301 16.2531
R11823 vdd.n7342 vdd.n7341 16.2531
R11824 vdd.n7341 vdd.n7302 16.2531
R11825 vdd.n7337 vdd.n7302 16.2531
R11826 vdd.n7367 vdd.n7366 16.2531
R11827 vdd.n7366 vdd.n7347 16.2531
R11828 vdd.n7388 vdd.n7347 16.2531
R11829 vdd.n7388 vdd.n7387 16.2531
R11830 vdd.n7387 vdd.n7348 16.2531
R11831 vdd.n7383 vdd.n7348 16.2531
R11832 vdd.n7413 vdd.n7412 16.2531
R11833 vdd.n7412 vdd.n7393 16.2531
R11834 vdd.n7434 vdd.n7393 16.2531
R11835 vdd.n7434 vdd.n7433 16.2531
R11836 vdd.n7433 vdd.n7394 16.2531
R11837 vdd.n7429 vdd.n7394 16.2531
R11838 vdd.n7510 vdd.n7509 16.2531
R11839 vdd.n7509 vdd.n7490 16.2531
R11840 vdd.n7531 vdd.n7490 16.2531
R11841 vdd.n7531 vdd.n7530 16.2531
R11842 vdd.n7530 vdd.n7491 16.2531
R11843 vdd.n7526 vdd.n7491 16.2531
R11844 vdd.n6659 vdd.n6658 16.2531
R11845 vdd.n6658 vdd.n6639 16.2531
R11846 vdd.n6680 vdd.n6639 16.2531
R11847 vdd.n6680 vdd.n6679 16.2531
R11848 vdd.n6679 vdd.n6640 16.2531
R11849 vdd.n6675 vdd.n6640 16.2531
R11850 vdd.n7554 vdd.n7553 16.2531
R11851 vdd.n7553 vdd.n7534 16.2531
R11852 vdd.n7575 vdd.n7534 16.2531
R11853 vdd.n7575 vdd.n7574 16.2531
R11854 vdd.n7574 vdd.n7535 16.2531
R11855 vdd.n7570 vdd.n7535 16.2531
R11856 vdd.n7599 vdd.n7598 16.2531
R11857 vdd.n7598 vdd.n7579 16.2531
R11858 vdd.n7620 vdd.n7579 16.2531
R11859 vdd.n7620 vdd.n7619 16.2531
R11860 vdd.n7619 vdd.n7580 16.2531
R11861 vdd.n7615 vdd.n7580 16.2531
R11862 vdd.n7649 vdd.n7648 16.2531
R11863 vdd.n7648 vdd.n7629 16.2531
R11864 vdd.n7670 vdd.n7629 16.2531
R11865 vdd.n7670 vdd.n7669 16.2531
R11866 vdd.n7669 vdd.n7630 16.2531
R11867 vdd.n7665 vdd.n7630 16.2531
R11868 vdd.n7695 vdd.n7694 16.2531
R11869 vdd.n7694 vdd.n7675 16.2531
R11870 vdd.n7716 vdd.n7675 16.2531
R11871 vdd.n7716 vdd.n7715 16.2531
R11872 vdd.n7715 vdd.n7676 16.2531
R11873 vdd.n7711 vdd.n7676 16.2531
R11874 vdd.n7743 vdd.n7742 16.2531
R11875 vdd.n7742 vdd.n7723 16.2531
R11876 vdd.n7764 vdd.n7723 16.2531
R11877 vdd.n7764 vdd.n7763 16.2531
R11878 vdd.n7763 vdd.n7724 16.2531
R11879 vdd.n7759 vdd.n7724 16.2531
R11880 vdd.n7482 vdd.n7439 16.2531
R11881 vdd.n7478 vdd.n7439 16.2531
R11882 vdd.n7478 vdd.n7477 16.2531
R11883 vdd.n7475 vdd.n7446 16.2531
R11884 vdd.n7471 vdd.n7446 16.2531
R11885 vdd.n7790 vdd.n7789 16.2531
R11886 vdd.n7789 vdd.n7770 16.2531
R11887 vdd.n7811 vdd.n7770 16.2531
R11888 vdd.n7811 vdd.n7810 16.2531
R11889 vdd.n7810 vdd.n7771 16.2531
R11890 vdd.n7806 vdd.n7771 16.2531
R11891 vdd.n7835 vdd.n7834 16.2531
R11892 vdd.n7834 vdd.n7815 16.2531
R11893 vdd.n7856 vdd.n7815 16.2531
R11894 vdd.n7856 vdd.n7855 16.2531
R11895 vdd.n7855 vdd.n7816 16.2531
R11896 vdd.n7851 vdd.n7816 16.2531
R11897 vdd.n7881 vdd.n7880 16.2531
R11898 vdd.n7880 vdd.n7861 16.2531
R11899 vdd.n7902 vdd.n7861 16.2531
R11900 vdd.n7902 vdd.n7901 16.2531
R11901 vdd.n7901 vdd.n7862 16.2531
R11902 vdd.n7897 vdd.n7862 16.2531
R11903 vdd.n7932 vdd.n7931 16.2531
R11904 vdd.n7931 vdd.n7912 16.2531
R11905 vdd.n7953 vdd.n7912 16.2531
R11906 vdd.n7953 vdd.n7952 16.2531
R11907 vdd.n7952 vdd.n7913 16.2531
R11908 vdd.n7948 vdd.n7913 16.2531
R11909 vdd.n7978 vdd.n7977 16.2531
R11910 vdd.n7977 vdd.n7958 16.2531
R11911 vdd.n7999 vdd.n7958 16.2531
R11912 vdd.n7999 vdd.n7998 16.2531
R11913 vdd.n7998 vdd.n7959 16.2531
R11914 vdd.n7994 vdd.n7959 16.2531
R11915 vdd.n8026 vdd.n8025 16.2531
R11916 vdd.n8025 vdd.n8006 16.2531
R11917 vdd.n8047 vdd.n8006 16.2531
R11918 vdd.n8047 vdd.n8046 16.2531
R11919 vdd.n8046 vdd.n8007 16.2531
R11920 vdd.n8042 vdd.n8007 16.2531
R11921 vdd.n8072 vdd.n8071 16.2531
R11922 vdd.n8071 vdd.n8052 16.2531
R11923 vdd.n8093 vdd.n8052 16.2531
R11924 vdd.n8093 vdd.n8092 16.2531
R11925 vdd.n8092 vdd.n8053 16.2531
R11926 vdd.n8088 vdd.n8053 16.2531
R11927 vdd.n8117 vdd.n8116 16.2531
R11928 vdd.n8116 vdd.n8097 16.2531
R11929 vdd.n8138 vdd.n8097 16.2531
R11930 vdd.n8138 vdd.n8137 16.2531
R11931 vdd.n8137 vdd.n8098 16.2531
R11932 vdd.n8133 vdd.n8098 16.2531
R11933 vdd.n8167 vdd.n8166 16.2531
R11934 vdd.n8166 vdd.n8147 16.2531
R11935 vdd.n8188 vdd.n8147 16.2531
R11936 vdd.n8188 vdd.n8187 16.2531
R11937 vdd.n8187 vdd.n8148 16.2531
R11938 vdd.n8183 vdd.n8148 16.2531
R11939 vdd.n8213 vdd.n8212 16.2531
R11940 vdd.n8212 vdd.n8193 16.2531
R11941 vdd.n8234 vdd.n8193 16.2531
R11942 vdd.n8234 vdd.n8233 16.2531
R11943 vdd.n8233 vdd.n8194 16.2531
R11944 vdd.n8229 vdd.n8194 16.2531
R11945 vdd.n8261 vdd.n8260 16.2531
R11946 vdd.n8260 vdd.n8241 16.2531
R11947 vdd.n8282 vdd.n8241 16.2531
R11948 vdd.n8282 vdd.n8281 16.2531
R11949 vdd.n8281 vdd.n8242 16.2531
R11950 vdd.n8277 vdd.n8242 16.2531
R11951 vdd.n7247 vdd.n7204 16.2531
R11952 vdd.n7243 vdd.n7204 16.2531
R11953 vdd.n7243 vdd.n7242 16.2531
R11954 vdd.n7240 vdd.n7211 16.2531
R11955 vdd.n7236 vdd.n7211 16.2531
R11956 vdd.n8308 vdd.n8307 16.2531
R11957 vdd.n8307 vdd.n8288 16.2531
R11958 vdd.n8329 vdd.n8288 16.2531
R11959 vdd.n8329 vdd.n8328 16.2531
R11960 vdd.n8328 vdd.n8289 16.2531
R11961 vdd.n8324 vdd.n8289 16.2531
R11962 vdd.n8353 vdd.n8352 16.2531
R11963 vdd.n8352 vdd.n8333 16.2531
R11964 vdd.n8374 vdd.n8333 16.2531
R11965 vdd.n8374 vdd.n8373 16.2531
R11966 vdd.n8373 vdd.n8334 16.2531
R11967 vdd.n8369 vdd.n8334 16.2531
R11968 vdd.n8403 vdd.n8402 16.2531
R11969 vdd.n8402 vdd.n8383 16.2531
R11970 vdd.n8424 vdd.n8383 16.2531
R11971 vdd.n8424 vdd.n8423 16.2531
R11972 vdd.n8423 vdd.n8384 16.2531
R11973 vdd.n8419 vdd.n8384 16.2531
R11974 vdd.n8449 vdd.n8448 16.2531
R11975 vdd.n8448 vdd.n8429 16.2531
R11976 vdd.n8470 vdd.n8429 16.2531
R11977 vdd.n8470 vdd.n8469 16.2531
R11978 vdd.n8469 vdd.n8430 16.2531
R11979 vdd.n8465 vdd.n8430 16.2531
R11980 vdd.n8497 vdd.n8496 16.2531
R11981 vdd.n8496 vdd.n8477 16.2531
R11982 vdd.n8518 vdd.n8477 16.2531
R11983 vdd.n8518 vdd.n8517 16.2531
R11984 vdd.n8517 vdd.n8478 16.2531
R11985 vdd.n8513 vdd.n8478 16.2531
R11986 vdd.n8636 vdd.n8635 16.2531
R11987 vdd.n8635 vdd.n8615 16.2531
R11988 vdd.n8656 vdd.n8615 16.2531
R11989 vdd.n8656 vdd.n8655 16.2531
R11990 vdd.n8655 vdd.n8616 16.2531
R11991 vdd.n8645 vdd.n8616 16.2531
R11992 vdd.n8590 vdd.n8589 16.2531
R11993 vdd.n8589 vdd.n8569 16.2531
R11994 vdd.n8610 vdd.n8569 16.2531
R11995 vdd.n8610 vdd.n8609 16.2531
R11996 vdd.n8609 vdd.n8570 16.2531
R11997 vdd.n8599 vdd.n8570 16.2531
R11998 vdd.n8683 vdd.n8682 16.2531
R11999 vdd.n8682 vdd.n8662 16.2531
R12000 vdd.n8703 vdd.n8662 16.2531
R12001 vdd.n8703 vdd.n8702 16.2531
R12002 vdd.n8702 vdd.n8663 16.2531
R12003 vdd.n8692 vdd.n8663 16.2531
R12004 vdd.n8731 vdd.n8730 16.2531
R12005 vdd.n8730 vdd.n8710 16.2531
R12006 vdd.n8751 vdd.n8710 16.2531
R12007 vdd.n8751 vdd.n8750 16.2531
R12008 vdd.n8750 vdd.n8711 16.2531
R12009 vdd.n8740 vdd.n8711 16.2531
R12010 vdd.n8777 vdd.n8776 16.2531
R12011 vdd.n8776 vdd.n8756 16.2531
R12012 vdd.n8797 vdd.n8756 16.2531
R12013 vdd.n8797 vdd.n8796 16.2531
R12014 vdd.n8796 vdd.n8757 16.2531
R12015 vdd.n8786 vdd.n8757 16.2531
R12016 vdd.n7032 vdd.n7020 16.2531
R12017 vdd.n7044 vdd.n7020 16.2531
R12018 vdd.n7048 vdd.n7047 16.2531
R12019 vdd.n7049 vdd.n7048 16.2531
R12020 vdd.n7049 vdd.n7013 16.2531
R12021 vdd.n8919 vdd.n8918 16.2531
R12022 vdd.n8918 vdd.n8898 16.2531
R12023 vdd.n8939 vdd.n8898 16.2531
R12024 vdd.n8939 vdd.n8938 16.2531
R12025 vdd.n8938 vdd.n8899 16.2531
R12026 vdd.n8928 vdd.n8899 16.2531
R12027 vdd.n8872 vdd.n8871 16.2531
R12028 vdd.n8871 vdd.n8851 16.2531
R12029 vdd.n8892 vdd.n8851 16.2531
R12030 vdd.n8892 vdd.n8891 16.2531
R12031 vdd.n8891 vdd.n8852 16.2531
R12032 vdd.n8881 vdd.n8852 16.2531
R12033 vdd.n8826 vdd.n8825 16.2531
R12034 vdd.n8825 vdd.n8805 16.2531
R12035 vdd.n8846 vdd.n8805 16.2531
R12036 vdd.n8846 vdd.n8845 16.2531
R12037 vdd.n8845 vdd.n8806 16.2531
R12038 vdd.n8835 vdd.n8806 16.2531
R12039 vdd.n8966 vdd.n8965 16.2531
R12040 vdd.n8965 vdd.n8945 16.2531
R12041 vdd.n8986 vdd.n8945 16.2531
R12042 vdd.n8986 vdd.n8985 16.2531
R12043 vdd.n8985 vdd.n8946 16.2531
R12044 vdd.n8975 vdd.n8946 16.2531
R12045 vdd.n9014 vdd.n9013 16.2531
R12046 vdd.n9013 vdd.n8993 16.2531
R12047 vdd.n9034 vdd.n8993 16.2531
R12048 vdd.n9034 vdd.n9033 16.2531
R12049 vdd.n9033 vdd.n8994 16.2531
R12050 vdd.n9023 vdd.n8994 16.2531
R12051 vdd.n9060 vdd.n9059 16.2531
R12052 vdd.n9059 vdd.n9039 16.2531
R12053 vdd.n9080 vdd.n9039 16.2531
R12054 vdd.n9080 vdd.n9079 16.2531
R12055 vdd.n9079 vdd.n9040 16.2531
R12056 vdd.n9069 vdd.n9040 16.2531
R12057 vdd.n9154 vdd.n9153 16.2531
R12058 vdd.n9153 vdd.n9133 16.2531
R12059 vdd.n9174 vdd.n9133 16.2531
R12060 vdd.n9174 vdd.n9173 16.2531
R12061 vdd.n9173 vdd.n9134 16.2531
R12062 vdd.n9163 vdd.n9134 16.2531
R12063 vdd.n9108 vdd.n9107 16.2531
R12064 vdd.n9107 vdd.n9087 16.2531
R12065 vdd.n9128 vdd.n9087 16.2531
R12066 vdd.n9128 vdd.n9127 16.2531
R12067 vdd.n9127 vdd.n9088 16.2531
R12068 vdd.n9117 vdd.n9088 16.2531
R12069 vdd.n9201 vdd.n9200 16.2531
R12070 vdd.n9200 vdd.n9180 16.2531
R12071 vdd.n9221 vdd.n9180 16.2531
R12072 vdd.n9221 vdd.n9220 16.2531
R12073 vdd.n9220 vdd.n9181 16.2531
R12074 vdd.n9210 vdd.n9181 16.2531
R12075 vdd.n9249 vdd.n9248 16.2531
R12076 vdd.n9248 vdd.n9228 16.2531
R12077 vdd.n9269 vdd.n9228 16.2531
R12078 vdd.n9269 vdd.n9268 16.2531
R12079 vdd.n9268 vdd.n9229 16.2531
R12080 vdd.n9258 vdd.n9229 16.2531
R12081 vdd.n9295 vdd.n9294 16.2531
R12082 vdd.n9294 vdd.n9274 16.2531
R12083 vdd.n9315 vdd.n9274 16.2531
R12084 vdd.n9315 vdd.n9314 16.2531
R12085 vdd.n9314 vdd.n9275 16.2531
R12086 vdd.n9304 vdd.n9275 16.2531
R12087 vdd.n6796 vdd.n6784 16.2531
R12088 vdd.n6808 vdd.n6784 16.2531
R12089 vdd.n6812 vdd.n6811 16.2531
R12090 vdd.n6813 vdd.n6812 16.2531
R12091 vdd.n6813 vdd.n6777 16.2531
R12092 vdd.n9390 vdd.n9389 16.2531
R12093 vdd.n9389 vdd.n9369 16.2531
R12094 vdd.n9410 vdd.n9369 16.2531
R12095 vdd.n9410 vdd.n9409 16.2531
R12096 vdd.n9409 vdd.n9370 16.2531
R12097 vdd.n9399 vdd.n9370 16.2531
R12098 vdd.n9344 vdd.n9343 16.2531
R12099 vdd.n9343 vdd.n9323 16.2531
R12100 vdd.n9364 vdd.n9323 16.2531
R12101 vdd.n9364 vdd.n9363 16.2531
R12102 vdd.n9363 vdd.n9324 16.2531
R12103 vdd.n9353 vdd.n9324 16.2531
R12104 vdd.n9437 vdd.n9436 16.2531
R12105 vdd.n9436 vdd.n9416 16.2531
R12106 vdd.n9457 vdd.n9416 16.2531
R12107 vdd.n9457 vdd.n9456 16.2531
R12108 vdd.n9456 vdd.n9417 16.2531
R12109 vdd.n9446 vdd.n9417 16.2531
R12110 vdd.n9485 vdd.n9484 16.2531
R12111 vdd.n9484 vdd.n9464 16.2531
R12112 vdd.n9505 vdd.n9464 16.2531
R12113 vdd.n9505 vdd.n9504 16.2531
R12114 vdd.n9504 vdd.n9465 16.2531
R12115 vdd.n9494 vdd.n9465 16.2531
R12116 vdd.n9531 vdd.n9530 16.2531
R12117 vdd.n9530 vdd.n9510 16.2531
R12118 vdd.n9551 vdd.n9510 16.2531
R12119 vdd.n9551 vdd.n9550 16.2531
R12120 vdd.n9550 vdd.n9511 16.2531
R12121 vdd.n9540 vdd.n9511 16.2531
R12122 vdd.n3691 vdd.n3690 16.2531
R12123 vdd.n3690 vdd.n3670 16.2531
R12124 vdd.n3711 vdd.n3670 16.2531
R12125 vdd.n3711 vdd.n3710 16.2531
R12126 vdd.n3710 vdd.n3671 16.2531
R12127 vdd.n3700 vdd.n3671 16.2531
R12128 vdd.n3737 vdd.n3736 16.2531
R12129 vdd.n3736 vdd.n3716 16.2531
R12130 vdd.n3757 vdd.n3716 16.2531
R12131 vdd.n3757 vdd.n3756 16.2531
R12132 vdd.n3756 vdd.n3717 16.2531
R12133 vdd.n3746 vdd.n3717 16.2531
R12134 vdd.n3835 vdd.n3834 16.2531
R12135 vdd.n3834 vdd.n3814 16.2531
R12136 vdd.n3855 vdd.n3814 16.2531
R12137 vdd.n3855 vdd.n3854 16.2531
R12138 vdd.n3854 vdd.n3815 16.2531
R12139 vdd.n3844 vdd.n3815 16.2531
R12140 vdd.n3881 vdd.n3880 16.2531
R12141 vdd.n3880 vdd.n3860 16.2531
R12142 vdd.n3901 vdd.n3860 16.2531
R12143 vdd.n3901 vdd.n3900 16.2531
R12144 vdd.n3900 vdd.n3861 16.2531
R12145 vdd.n3890 vdd.n3861 16.2531
R12146 vdd.n3927 vdd.n3926 16.2531
R12147 vdd.n3926 vdd.n3906 16.2531
R12148 vdd.n3947 vdd.n3906 16.2531
R12149 vdd.n3947 vdd.n3946 16.2531
R12150 vdd.n3946 vdd.n3907 16.2531
R12151 vdd.n3936 vdd.n3907 16.2531
R12152 vdd.n3973 vdd.n3972 16.2531
R12153 vdd.n3972 vdd.n3952 16.2531
R12154 vdd.n3993 vdd.n3952 16.2531
R12155 vdd.n3993 vdd.n3992 16.2531
R12156 vdd.n3992 vdd.n3953 16.2531
R12157 vdd.n3982 vdd.n3953 16.2531
R12158 vdd.n4071 vdd.n4070 16.2531
R12159 vdd.n4070 vdd.n4050 16.2531
R12160 vdd.n4091 vdd.n4050 16.2531
R12161 vdd.n4091 vdd.n4090 16.2531
R12162 vdd.n4090 vdd.n4051 16.2531
R12163 vdd.n4080 vdd.n4051 16.2531
R12164 vdd.n5529 vdd.n5528 16.2531
R12165 vdd.n5528 vdd.n5508 16.2531
R12166 vdd.n5549 vdd.n5508 16.2531
R12167 vdd.n5549 vdd.n5548 16.2531
R12168 vdd.n5548 vdd.n5509 16.2531
R12169 vdd.n5538 vdd.n5509 16.2531
R12170 vdd.n4118 vdd.n4117 16.2531
R12171 vdd.n4117 vdd.n4098 16.2531
R12172 vdd.n4139 vdd.n4098 16.2531
R12173 vdd.n4139 vdd.n4138 16.2531
R12174 vdd.n4138 vdd.n4099 16.2531
R12175 vdd.n4134 vdd.n4099 16.2531
R12176 vdd.n4164 vdd.n4163 16.2531
R12177 vdd.n4163 vdd.n4144 16.2531
R12178 vdd.n4185 vdd.n4144 16.2531
R12179 vdd.n4185 vdd.n4184 16.2531
R12180 vdd.n4184 vdd.n4145 16.2531
R12181 vdd.n4180 vdd.n4145 16.2531
R12182 vdd.n4261 vdd.n4260 16.2531
R12183 vdd.n4260 vdd.n4241 16.2531
R12184 vdd.n4282 vdd.n4241 16.2531
R12185 vdd.n4282 vdd.n4281 16.2531
R12186 vdd.n4281 vdd.n4242 16.2531
R12187 vdd.n4277 vdd.n4242 16.2531
R12188 vdd.n4307 vdd.n4306 16.2531
R12189 vdd.n4306 vdd.n4287 16.2531
R12190 vdd.n4328 vdd.n4287 16.2531
R12191 vdd.n4328 vdd.n4327 16.2531
R12192 vdd.n4327 vdd.n4288 16.2531
R12193 vdd.n4323 vdd.n4288 16.2531
R12194 vdd.n4353 vdd.n4352 16.2531
R12195 vdd.n4352 vdd.n4333 16.2531
R12196 vdd.n4374 vdd.n4333 16.2531
R12197 vdd.n4374 vdd.n4373 16.2531
R12198 vdd.n4373 vdd.n4334 16.2531
R12199 vdd.n4369 vdd.n4334 16.2531
R12200 vdd.n4399 vdd.n4398 16.2531
R12201 vdd.n4398 vdd.n4379 16.2531
R12202 vdd.n4420 vdd.n4379 16.2531
R12203 vdd.n4420 vdd.n4419 16.2531
R12204 vdd.n4419 vdd.n4380 16.2531
R12205 vdd.n4415 vdd.n4380 16.2531
R12206 vdd.n4496 vdd.n4495 16.2531
R12207 vdd.n4495 vdd.n4476 16.2531
R12208 vdd.n4517 vdd.n4476 16.2531
R12209 vdd.n4517 vdd.n4516 16.2531
R12210 vdd.n4516 vdd.n4477 16.2531
R12211 vdd.n4512 vdd.n4477 16.2531
R12212 vdd.n3645 vdd.n3644 16.2531
R12213 vdd.n3644 vdd.n3625 16.2531
R12214 vdd.n3666 vdd.n3625 16.2531
R12215 vdd.n3666 vdd.n3665 16.2531
R12216 vdd.n3665 vdd.n3626 16.2531
R12217 vdd.n3661 vdd.n3626 16.2531
R12218 vdd.n4540 vdd.n4539 16.2531
R12219 vdd.n4539 vdd.n4520 16.2531
R12220 vdd.n4561 vdd.n4520 16.2531
R12221 vdd.n4561 vdd.n4560 16.2531
R12222 vdd.n4560 vdd.n4521 16.2531
R12223 vdd.n4556 vdd.n4521 16.2531
R12224 vdd.n4585 vdd.n4584 16.2531
R12225 vdd.n4584 vdd.n4565 16.2531
R12226 vdd.n4606 vdd.n4565 16.2531
R12227 vdd.n4606 vdd.n4605 16.2531
R12228 vdd.n4605 vdd.n4566 16.2531
R12229 vdd.n4601 vdd.n4566 16.2531
R12230 vdd.n4635 vdd.n4634 16.2531
R12231 vdd.n4634 vdd.n4615 16.2531
R12232 vdd.n4656 vdd.n4615 16.2531
R12233 vdd.n4656 vdd.n4655 16.2531
R12234 vdd.n4655 vdd.n4616 16.2531
R12235 vdd.n4651 vdd.n4616 16.2531
R12236 vdd.n4681 vdd.n4680 16.2531
R12237 vdd.n4680 vdd.n4661 16.2531
R12238 vdd.n4702 vdd.n4661 16.2531
R12239 vdd.n4702 vdd.n4701 16.2531
R12240 vdd.n4701 vdd.n4662 16.2531
R12241 vdd.n4697 vdd.n4662 16.2531
R12242 vdd.n4729 vdd.n4728 16.2531
R12243 vdd.n4728 vdd.n4709 16.2531
R12244 vdd.n4750 vdd.n4709 16.2531
R12245 vdd.n4750 vdd.n4749 16.2531
R12246 vdd.n4749 vdd.n4710 16.2531
R12247 vdd.n4745 vdd.n4710 16.2531
R12248 vdd.n4468 vdd.n4425 16.2531
R12249 vdd.n4464 vdd.n4425 16.2531
R12250 vdd.n4464 vdd.n4463 16.2531
R12251 vdd.n4461 vdd.n4432 16.2531
R12252 vdd.n4457 vdd.n4432 16.2531
R12253 vdd.n4776 vdd.n4775 16.2531
R12254 vdd.n4775 vdd.n4756 16.2531
R12255 vdd.n4797 vdd.n4756 16.2531
R12256 vdd.n4797 vdd.n4796 16.2531
R12257 vdd.n4796 vdd.n4757 16.2531
R12258 vdd.n4792 vdd.n4757 16.2531
R12259 vdd.n4821 vdd.n4820 16.2531
R12260 vdd.n4820 vdd.n4801 16.2531
R12261 vdd.n4842 vdd.n4801 16.2531
R12262 vdd.n4842 vdd.n4841 16.2531
R12263 vdd.n4841 vdd.n4802 16.2531
R12264 vdd.n4837 vdd.n4802 16.2531
R12265 vdd.n4867 vdd.n4866 16.2531
R12266 vdd.n4866 vdd.n4847 16.2531
R12267 vdd.n4888 vdd.n4847 16.2531
R12268 vdd.n4888 vdd.n4887 16.2531
R12269 vdd.n4887 vdd.n4848 16.2531
R12270 vdd.n4883 vdd.n4848 16.2531
R12271 vdd.n4918 vdd.n4917 16.2531
R12272 vdd.n4917 vdd.n4898 16.2531
R12273 vdd.n4939 vdd.n4898 16.2531
R12274 vdd.n4939 vdd.n4938 16.2531
R12275 vdd.n4938 vdd.n4899 16.2531
R12276 vdd.n4934 vdd.n4899 16.2531
R12277 vdd.n4964 vdd.n4963 16.2531
R12278 vdd.n4963 vdd.n4944 16.2531
R12279 vdd.n4985 vdd.n4944 16.2531
R12280 vdd.n4985 vdd.n4984 16.2531
R12281 vdd.n4984 vdd.n4945 16.2531
R12282 vdd.n4980 vdd.n4945 16.2531
R12283 vdd.n5012 vdd.n5011 16.2531
R12284 vdd.n5011 vdd.n4992 16.2531
R12285 vdd.n5033 vdd.n4992 16.2531
R12286 vdd.n5033 vdd.n5032 16.2531
R12287 vdd.n5032 vdd.n4993 16.2531
R12288 vdd.n5028 vdd.n4993 16.2531
R12289 vdd.n5058 vdd.n5057 16.2531
R12290 vdd.n5057 vdd.n5038 16.2531
R12291 vdd.n5079 vdd.n5038 16.2531
R12292 vdd.n5079 vdd.n5078 16.2531
R12293 vdd.n5078 vdd.n5039 16.2531
R12294 vdd.n5074 vdd.n5039 16.2531
R12295 vdd.n5103 vdd.n5102 16.2531
R12296 vdd.n5102 vdd.n5083 16.2531
R12297 vdd.n5124 vdd.n5083 16.2531
R12298 vdd.n5124 vdd.n5123 16.2531
R12299 vdd.n5123 vdd.n5084 16.2531
R12300 vdd.n5119 vdd.n5084 16.2531
R12301 vdd.n5153 vdd.n5152 16.2531
R12302 vdd.n5152 vdd.n5133 16.2531
R12303 vdd.n5174 vdd.n5133 16.2531
R12304 vdd.n5174 vdd.n5173 16.2531
R12305 vdd.n5173 vdd.n5134 16.2531
R12306 vdd.n5169 vdd.n5134 16.2531
R12307 vdd.n5199 vdd.n5198 16.2531
R12308 vdd.n5198 vdd.n5179 16.2531
R12309 vdd.n5220 vdd.n5179 16.2531
R12310 vdd.n5220 vdd.n5219 16.2531
R12311 vdd.n5219 vdd.n5180 16.2531
R12312 vdd.n5215 vdd.n5180 16.2531
R12313 vdd.n5247 vdd.n5246 16.2531
R12314 vdd.n5246 vdd.n5227 16.2531
R12315 vdd.n5268 vdd.n5227 16.2531
R12316 vdd.n5268 vdd.n5267 16.2531
R12317 vdd.n5267 vdd.n5228 16.2531
R12318 vdd.n5263 vdd.n5228 16.2531
R12319 vdd.n4233 vdd.n4190 16.2531
R12320 vdd.n4229 vdd.n4190 16.2531
R12321 vdd.n4229 vdd.n4228 16.2531
R12322 vdd.n4226 vdd.n4197 16.2531
R12323 vdd.n4222 vdd.n4197 16.2531
R12324 vdd.n5294 vdd.n5293 16.2531
R12325 vdd.n5293 vdd.n5274 16.2531
R12326 vdd.n5315 vdd.n5274 16.2531
R12327 vdd.n5315 vdd.n5314 16.2531
R12328 vdd.n5314 vdd.n5275 16.2531
R12329 vdd.n5310 vdd.n5275 16.2531
R12330 vdd.n5339 vdd.n5338 16.2531
R12331 vdd.n5338 vdd.n5319 16.2531
R12332 vdd.n5360 vdd.n5319 16.2531
R12333 vdd.n5360 vdd.n5359 16.2531
R12334 vdd.n5359 vdd.n5320 16.2531
R12335 vdd.n5355 vdd.n5320 16.2531
R12336 vdd.n5389 vdd.n5388 16.2531
R12337 vdd.n5388 vdd.n5369 16.2531
R12338 vdd.n5410 vdd.n5369 16.2531
R12339 vdd.n5410 vdd.n5409 16.2531
R12340 vdd.n5409 vdd.n5370 16.2531
R12341 vdd.n5405 vdd.n5370 16.2531
R12342 vdd.n5435 vdd.n5434 16.2531
R12343 vdd.n5434 vdd.n5415 16.2531
R12344 vdd.n5456 vdd.n5415 16.2531
R12345 vdd.n5456 vdd.n5455 16.2531
R12346 vdd.n5455 vdd.n5416 16.2531
R12347 vdd.n5451 vdd.n5416 16.2531
R12348 vdd.n5483 vdd.n5482 16.2531
R12349 vdd.n5482 vdd.n5463 16.2531
R12350 vdd.n5504 vdd.n5463 16.2531
R12351 vdd.n5504 vdd.n5503 16.2531
R12352 vdd.n5503 vdd.n5464 16.2531
R12353 vdd.n5499 vdd.n5464 16.2531
R12354 vdd.n5622 vdd.n5621 16.2531
R12355 vdd.n5621 vdd.n5601 16.2531
R12356 vdd.n5642 vdd.n5601 16.2531
R12357 vdd.n5642 vdd.n5641 16.2531
R12358 vdd.n5641 vdd.n5602 16.2531
R12359 vdd.n5631 vdd.n5602 16.2531
R12360 vdd.n5576 vdd.n5575 16.2531
R12361 vdd.n5575 vdd.n5555 16.2531
R12362 vdd.n5596 vdd.n5555 16.2531
R12363 vdd.n5596 vdd.n5595 16.2531
R12364 vdd.n5595 vdd.n5556 16.2531
R12365 vdd.n5585 vdd.n5556 16.2531
R12366 vdd.n5669 vdd.n5668 16.2531
R12367 vdd.n5668 vdd.n5648 16.2531
R12368 vdd.n5689 vdd.n5648 16.2531
R12369 vdd.n5689 vdd.n5688 16.2531
R12370 vdd.n5688 vdd.n5649 16.2531
R12371 vdd.n5678 vdd.n5649 16.2531
R12372 vdd.n5717 vdd.n5716 16.2531
R12373 vdd.n5716 vdd.n5696 16.2531
R12374 vdd.n5737 vdd.n5696 16.2531
R12375 vdd.n5737 vdd.n5736 16.2531
R12376 vdd.n5736 vdd.n5697 16.2531
R12377 vdd.n5726 vdd.n5697 16.2531
R12378 vdd.n5763 vdd.n5762 16.2531
R12379 vdd.n5762 vdd.n5742 16.2531
R12380 vdd.n5783 vdd.n5742 16.2531
R12381 vdd.n5783 vdd.n5782 16.2531
R12382 vdd.n5782 vdd.n5743 16.2531
R12383 vdd.n5772 vdd.n5743 16.2531
R12384 vdd.n4018 vdd.n4006 16.2531
R12385 vdd.n4030 vdd.n4006 16.2531
R12386 vdd.n4034 vdd.n4033 16.2531
R12387 vdd.n4035 vdd.n4034 16.2531
R12388 vdd.n4035 vdd.n3999 16.2531
R12389 vdd.n5905 vdd.n5904 16.2531
R12390 vdd.n5904 vdd.n5884 16.2531
R12391 vdd.n5925 vdd.n5884 16.2531
R12392 vdd.n5925 vdd.n5924 16.2531
R12393 vdd.n5924 vdd.n5885 16.2531
R12394 vdd.n5914 vdd.n5885 16.2531
R12395 vdd.n5858 vdd.n5857 16.2531
R12396 vdd.n5857 vdd.n5837 16.2531
R12397 vdd.n5878 vdd.n5837 16.2531
R12398 vdd.n5878 vdd.n5877 16.2531
R12399 vdd.n5877 vdd.n5838 16.2531
R12400 vdd.n5867 vdd.n5838 16.2531
R12401 vdd.n5812 vdd.n5811 16.2531
R12402 vdd.n5811 vdd.n5791 16.2531
R12403 vdd.n5832 vdd.n5791 16.2531
R12404 vdd.n5832 vdd.n5831 16.2531
R12405 vdd.n5831 vdd.n5792 16.2531
R12406 vdd.n5821 vdd.n5792 16.2531
R12407 vdd.n5952 vdd.n5951 16.2531
R12408 vdd.n5951 vdd.n5931 16.2531
R12409 vdd.n5972 vdd.n5931 16.2531
R12410 vdd.n5972 vdd.n5971 16.2531
R12411 vdd.n5971 vdd.n5932 16.2531
R12412 vdd.n5961 vdd.n5932 16.2531
R12413 vdd.n6000 vdd.n5999 16.2531
R12414 vdd.n5999 vdd.n5979 16.2531
R12415 vdd.n6020 vdd.n5979 16.2531
R12416 vdd.n6020 vdd.n6019 16.2531
R12417 vdd.n6019 vdd.n5980 16.2531
R12418 vdd.n6009 vdd.n5980 16.2531
R12419 vdd.n6046 vdd.n6045 16.2531
R12420 vdd.n6045 vdd.n6025 16.2531
R12421 vdd.n6066 vdd.n6025 16.2531
R12422 vdd.n6066 vdd.n6065 16.2531
R12423 vdd.n6065 vdd.n6026 16.2531
R12424 vdd.n6055 vdd.n6026 16.2531
R12425 vdd.n6140 vdd.n6139 16.2531
R12426 vdd.n6139 vdd.n6119 16.2531
R12427 vdd.n6160 vdd.n6119 16.2531
R12428 vdd.n6160 vdd.n6159 16.2531
R12429 vdd.n6159 vdd.n6120 16.2531
R12430 vdd.n6149 vdd.n6120 16.2531
R12431 vdd.n6094 vdd.n6093 16.2531
R12432 vdd.n6093 vdd.n6073 16.2531
R12433 vdd.n6114 vdd.n6073 16.2531
R12434 vdd.n6114 vdd.n6113 16.2531
R12435 vdd.n6113 vdd.n6074 16.2531
R12436 vdd.n6103 vdd.n6074 16.2531
R12437 vdd.n6187 vdd.n6186 16.2531
R12438 vdd.n6186 vdd.n6166 16.2531
R12439 vdd.n6207 vdd.n6166 16.2531
R12440 vdd.n6207 vdd.n6206 16.2531
R12441 vdd.n6206 vdd.n6167 16.2531
R12442 vdd.n6196 vdd.n6167 16.2531
R12443 vdd.n6235 vdd.n6234 16.2531
R12444 vdd.n6234 vdd.n6214 16.2531
R12445 vdd.n6255 vdd.n6214 16.2531
R12446 vdd.n6255 vdd.n6254 16.2531
R12447 vdd.n6254 vdd.n6215 16.2531
R12448 vdd.n6244 vdd.n6215 16.2531
R12449 vdd.n6281 vdd.n6280 16.2531
R12450 vdd.n6280 vdd.n6260 16.2531
R12451 vdd.n6301 vdd.n6260 16.2531
R12452 vdd.n6301 vdd.n6300 16.2531
R12453 vdd.n6300 vdd.n6261 16.2531
R12454 vdd.n6290 vdd.n6261 16.2531
R12455 vdd.n3782 vdd.n3770 16.2531
R12456 vdd.n3794 vdd.n3770 16.2531
R12457 vdd.n3798 vdd.n3797 16.2531
R12458 vdd.n3799 vdd.n3798 16.2531
R12459 vdd.n3799 vdd.n3763 16.2531
R12460 vdd.n6376 vdd.n6375 16.2531
R12461 vdd.n6375 vdd.n6355 16.2531
R12462 vdd.n6396 vdd.n6355 16.2531
R12463 vdd.n6396 vdd.n6395 16.2531
R12464 vdd.n6395 vdd.n6356 16.2531
R12465 vdd.n6385 vdd.n6356 16.2531
R12466 vdd.n6330 vdd.n6329 16.2531
R12467 vdd.n6329 vdd.n6309 16.2531
R12468 vdd.n6350 vdd.n6309 16.2531
R12469 vdd.n6350 vdd.n6349 16.2531
R12470 vdd.n6349 vdd.n6310 16.2531
R12471 vdd.n6339 vdd.n6310 16.2531
R12472 vdd.n6423 vdd.n6422 16.2531
R12473 vdd.n6422 vdd.n6402 16.2531
R12474 vdd.n6443 vdd.n6402 16.2531
R12475 vdd.n6443 vdd.n6442 16.2531
R12476 vdd.n6442 vdd.n6403 16.2531
R12477 vdd.n6432 vdd.n6403 16.2531
R12478 vdd.n6471 vdd.n6470 16.2531
R12479 vdd.n6470 vdd.n6450 16.2531
R12480 vdd.n6491 vdd.n6450 16.2531
R12481 vdd.n6491 vdd.n6490 16.2531
R12482 vdd.n6490 vdd.n6451 16.2531
R12483 vdd.n6480 vdd.n6451 16.2531
R12484 vdd.n6517 vdd.n6516 16.2531
R12485 vdd.n6516 vdd.n6496 16.2531
R12486 vdd.n6537 vdd.n6496 16.2531
R12487 vdd.n6537 vdd.n6536 16.2531
R12488 vdd.n6536 vdd.n6497 16.2531
R12489 vdd.n6526 vdd.n6497 16.2531
R12490 vdd.n677 vdd.n676 16.2531
R12491 vdd.n676 vdd.n656 16.2531
R12492 vdd.n697 vdd.n656 16.2531
R12493 vdd.n697 vdd.n696 16.2531
R12494 vdd.n696 vdd.n657 16.2531
R12495 vdd.n686 vdd.n657 16.2531
R12496 vdd.n723 vdd.n722 16.2531
R12497 vdd.n722 vdd.n702 16.2531
R12498 vdd.n743 vdd.n702 16.2531
R12499 vdd.n743 vdd.n742 16.2531
R12500 vdd.n742 vdd.n703 16.2531
R12501 vdd.n732 vdd.n703 16.2531
R12502 vdd.n821 vdd.n820 16.2531
R12503 vdd.n820 vdd.n800 16.2531
R12504 vdd.n841 vdd.n800 16.2531
R12505 vdd.n841 vdd.n840 16.2531
R12506 vdd.n840 vdd.n801 16.2531
R12507 vdd.n830 vdd.n801 16.2531
R12508 vdd.n867 vdd.n866 16.2531
R12509 vdd.n866 vdd.n846 16.2531
R12510 vdd.n887 vdd.n846 16.2531
R12511 vdd.n887 vdd.n886 16.2531
R12512 vdd.n886 vdd.n847 16.2531
R12513 vdd.n876 vdd.n847 16.2531
R12514 vdd.n913 vdd.n912 16.2531
R12515 vdd.n912 vdd.n892 16.2531
R12516 vdd.n933 vdd.n892 16.2531
R12517 vdd.n933 vdd.n932 16.2531
R12518 vdd.n932 vdd.n893 16.2531
R12519 vdd.n922 vdd.n893 16.2531
R12520 vdd.n959 vdd.n958 16.2531
R12521 vdd.n958 vdd.n938 16.2531
R12522 vdd.n979 vdd.n938 16.2531
R12523 vdd.n979 vdd.n978 16.2531
R12524 vdd.n978 vdd.n939 16.2531
R12525 vdd.n968 vdd.n939 16.2531
R12526 vdd.n1057 vdd.n1056 16.2531
R12527 vdd.n1056 vdd.n1036 16.2531
R12528 vdd.n1077 vdd.n1036 16.2531
R12529 vdd.n1077 vdd.n1076 16.2531
R12530 vdd.n1076 vdd.n1037 16.2531
R12531 vdd.n1066 vdd.n1037 16.2531
R12532 vdd.n2515 vdd.n2514 16.2531
R12533 vdd.n2514 vdd.n2494 16.2531
R12534 vdd.n2535 vdd.n2494 16.2531
R12535 vdd.n2535 vdd.n2534 16.2531
R12536 vdd.n2534 vdd.n2495 16.2531
R12537 vdd.n2524 vdd.n2495 16.2531
R12538 vdd.n1104 vdd.n1103 16.2531
R12539 vdd.n1103 vdd.n1084 16.2531
R12540 vdd.n1125 vdd.n1084 16.2531
R12541 vdd.n1125 vdd.n1124 16.2531
R12542 vdd.n1124 vdd.n1085 16.2531
R12543 vdd.n1120 vdd.n1085 16.2531
R12544 vdd.n1150 vdd.n1149 16.2531
R12545 vdd.n1149 vdd.n1130 16.2531
R12546 vdd.n1171 vdd.n1130 16.2531
R12547 vdd.n1171 vdd.n1170 16.2531
R12548 vdd.n1170 vdd.n1131 16.2531
R12549 vdd.n1166 vdd.n1131 16.2531
R12550 vdd.n1247 vdd.n1246 16.2531
R12551 vdd.n1246 vdd.n1227 16.2531
R12552 vdd.n1268 vdd.n1227 16.2531
R12553 vdd.n1268 vdd.n1267 16.2531
R12554 vdd.n1267 vdd.n1228 16.2531
R12555 vdd.n1263 vdd.n1228 16.2531
R12556 vdd.n1293 vdd.n1292 16.2531
R12557 vdd.n1292 vdd.n1273 16.2531
R12558 vdd.n1314 vdd.n1273 16.2531
R12559 vdd.n1314 vdd.n1313 16.2531
R12560 vdd.n1313 vdd.n1274 16.2531
R12561 vdd.n1309 vdd.n1274 16.2531
R12562 vdd.n1339 vdd.n1338 16.2531
R12563 vdd.n1338 vdd.n1319 16.2531
R12564 vdd.n1360 vdd.n1319 16.2531
R12565 vdd.n1360 vdd.n1359 16.2531
R12566 vdd.n1359 vdd.n1320 16.2531
R12567 vdd.n1355 vdd.n1320 16.2531
R12568 vdd.n1385 vdd.n1384 16.2531
R12569 vdd.n1384 vdd.n1365 16.2531
R12570 vdd.n1406 vdd.n1365 16.2531
R12571 vdd.n1406 vdd.n1405 16.2531
R12572 vdd.n1405 vdd.n1366 16.2531
R12573 vdd.n1401 vdd.n1366 16.2531
R12574 vdd.n1482 vdd.n1481 16.2531
R12575 vdd.n1481 vdd.n1462 16.2531
R12576 vdd.n1503 vdd.n1462 16.2531
R12577 vdd.n1503 vdd.n1502 16.2531
R12578 vdd.n1502 vdd.n1463 16.2531
R12579 vdd.n1498 vdd.n1463 16.2531
R12580 vdd.n631 vdd.n630 16.2531
R12581 vdd.n630 vdd.n611 16.2531
R12582 vdd.n652 vdd.n611 16.2531
R12583 vdd.n652 vdd.n651 16.2531
R12584 vdd.n651 vdd.n612 16.2531
R12585 vdd.n647 vdd.n612 16.2531
R12586 vdd.n1526 vdd.n1525 16.2531
R12587 vdd.n1525 vdd.n1506 16.2531
R12588 vdd.n1547 vdd.n1506 16.2531
R12589 vdd.n1547 vdd.n1546 16.2531
R12590 vdd.n1546 vdd.n1507 16.2531
R12591 vdd.n1542 vdd.n1507 16.2531
R12592 vdd.n1571 vdd.n1570 16.2531
R12593 vdd.n1570 vdd.n1551 16.2531
R12594 vdd.n1592 vdd.n1551 16.2531
R12595 vdd.n1592 vdd.n1591 16.2531
R12596 vdd.n1591 vdd.n1552 16.2531
R12597 vdd.n1587 vdd.n1552 16.2531
R12598 vdd.n1621 vdd.n1620 16.2531
R12599 vdd.n1620 vdd.n1601 16.2531
R12600 vdd.n1642 vdd.n1601 16.2531
R12601 vdd.n1642 vdd.n1641 16.2531
R12602 vdd.n1641 vdd.n1602 16.2531
R12603 vdd.n1637 vdd.n1602 16.2531
R12604 vdd.n1667 vdd.n1666 16.2531
R12605 vdd.n1666 vdd.n1647 16.2531
R12606 vdd.n1688 vdd.n1647 16.2531
R12607 vdd.n1688 vdd.n1687 16.2531
R12608 vdd.n1687 vdd.n1648 16.2531
R12609 vdd.n1683 vdd.n1648 16.2531
R12610 vdd.n1715 vdd.n1714 16.2531
R12611 vdd.n1714 vdd.n1695 16.2531
R12612 vdd.n1736 vdd.n1695 16.2531
R12613 vdd.n1736 vdd.n1735 16.2531
R12614 vdd.n1735 vdd.n1696 16.2531
R12615 vdd.n1731 vdd.n1696 16.2531
R12616 vdd.n1454 vdd.n1411 16.2531
R12617 vdd.n1450 vdd.n1411 16.2531
R12618 vdd.n1450 vdd.n1449 16.2531
R12619 vdd.n1447 vdd.n1418 16.2531
R12620 vdd.n1443 vdd.n1418 16.2531
R12621 vdd.n1762 vdd.n1761 16.2531
R12622 vdd.n1761 vdd.n1742 16.2531
R12623 vdd.n1783 vdd.n1742 16.2531
R12624 vdd.n1783 vdd.n1782 16.2531
R12625 vdd.n1782 vdd.n1743 16.2531
R12626 vdd.n1778 vdd.n1743 16.2531
R12627 vdd.n1807 vdd.n1806 16.2531
R12628 vdd.n1806 vdd.n1787 16.2531
R12629 vdd.n1828 vdd.n1787 16.2531
R12630 vdd.n1828 vdd.n1827 16.2531
R12631 vdd.n1827 vdd.n1788 16.2531
R12632 vdd.n1823 vdd.n1788 16.2531
R12633 vdd.n1853 vdd.n1852 16.2531
R12634 vdd.n1852 vdd.n1833 16.2531
R12635 vdd.n1874 vdd.n1833 16.2531
R12636 vdd.n1874 vdd.n1873 16.2531
R12637 vdd.n1873 vdd.n1834 16.2531
R12638 vdd.n1869 vdd.n1834 16.2531
R12639 vdd.n1904 vdd.n1903 16.2531
R12640 vdd.n1903 vdd.n1884 16.2531
R12641 vdd.n1925 vdd.n1884 16.2531
R12642 vdd.n1925 vdd.n1924 16.2531
R12643 vdd.n1924 vdd.n1885 16.2531
R12644 vdd.n1920 vdd.n1885 16.2531
R12645 vdd.n1950 vdd.n1949 16.2531
R12646 vdd.n1949 vdd.n1930 16.2531
R12647 vdd.n1971 vdd.n1930 16.2531
R12648 vdd.n1971 vdd.n1970 16.2531
R12649 vdd.n1970 vdd.n1931 16.2531
R12650 vdd.n1966 vdd.n1931 16.2531
R12651 vdd.n1998 vdd.n1997 16.2531
R12652 vdd.n1997 vdd.n1978 16.2531
R12653 vdd.n2019 vdd.n1978 16.2531
R12654 vdd.n2019 vdd.n2018 16.2531
R12655 vdd.n2018 vdd.n1979 16.2531
R12656 vdd.n2014 vdd.n1979 16.2531
R12657 vdd.n2044 vdd.n2043 16.2531
R12658 vdd.n2043 vdd.n2024 16.2531
R12659 vdd.n2065 vdd.n2024 16.2531
R12660 vdd.n2065 vdd.n2064 16.2531
R12661 vdd.n2064 vdd.n2025 16.2531
R12662 vdd.n2060 vdd.n2025 16.2531
R12663 vdd.n2089 vdd.n2088 16.2531
R12664 vdd.n2088 vdd.n2069 16.2531
R12665 vdd.n2110 vdd.n2069 16.2531
R12666 vdd.n2110 vdd.n2109 16.2531
R12667 vdd.n2109 vdd.n2070 16.2531
R12668 vdd.n2105 vdd.n2070 16.2531
R12669 vdd.n2139 vdd.n2138 16.2531
R12670 vdd.n2138 vdd.n2119 16.2531
R12671 vdd.n2160 vdd.n2119 16.2531
R12672 vdd.n2160 vdd.n2159 16.2531
R12673 vdd.n2159 vdd.n2120 16.2531
R12674 vdd.n2155 vdd.n2120 16.2531
R12675 vdd.n2185 vdd.n2184 16.2531
R12676 vdd.n2184 vdd.n2165 16.2531
R12677 vdd.n2206 vdd.n2165 16.2531
R12678 vdd.n2206 vdd.n2205 16.2531
R12679 vdd.n2205 vdd.n2166 16.2531
R12680 vdd.n2201 vdd.n2166 16.2531
R12681 vdd.n2233 vdd.n2232 16.2531
R12682 vdd.n2232 vdd.n2213 16.2531
R12683 vdd.n2254 vdd.n2213 16.2531
R12684 vdd.n2254 vdd.n2253 16.2531
R12685 vdd.n2253 vdd.n2214 16.2531
R12686 vdd.n2249 vdd.n2214 16.2531
R12687 vdd.n1219 vdd.n1176 16.2531
R12688 vdd.n1215 vdd.n1176 16.2531
R12689 vdd.n1215 vdd.n1214 16.2531
R12690 vdd.n1212 vdd.n1183 16.2531
R12691 vdd.n1208 vdd.n1183 16.2531
R12692 vdd.n2280 vdd.n2279 16.2531
R12693 vdd.n2279 vdd.n2260 16.2531
R12694 vdd.n2301 vdd.n2260 16.2531
R12695 vdd.n2301 vdd.n2300 16.2531
R12696 vdd.n2300 vdd.n2261 16.2531
R12697 vdd.n2296 vdd.n2261 16.2531
R12698 vdd.n2325 vdd.n2324 16.2531
R12699 vdd.n2324 vdd.n2305 16.2531
R12700 vdd.n2346 vdd.n2305 16.2531
R12701 vdd.n2346 vdd.n2345 16.2531
R12702 vdd.n2345 vdd.n2306 16.2531
R12703 vdd.n2341 vdd.n2306 16.2531
R12704 vdd.n2375 vdd.n2374 16.2531
R12705 vdd.n2374 vdd.n2355 16.2531
R12706 vdd.n2396 vdd.n2355 16.2531
R12707 vdd.n2396 vdd.n2395 16.2531
R12708 vdd.n2395 vdd.n2356 16.2531
R12709 vdd.n2391 vdd.n2356 16.2531
R12710 vdd.n2421 vdd.n2420 16.2531
R12711 vdd.n2420 vdd.n2401 16.2531
R12712 vdd.n2442 vdd.n2401 16.2531
R12713 vdd.n2442 vdd.n2441 16.2531
R12714 vdd.n2441 vdd.n2402 16.2531
R12715 vdd.n2437 vdd.n2402 16.2531
R12716 vdd.n2469 vdd.n2468 16.2531
R12717 vdd.n2468 vdd.n2449 16.2531
R12718 vdd.n2490 vdd.n2449 16.2531
R12719 vdd.n2490 vdd.n2489 16.2531
R12720 vdd.n2489 vdd.n2450 16.2531
R12721 vdd.n2485 vdd.n2450 16.2531
R12722 vdd.n2608 vdd.n2607 16.2531
R12723 vdd.n2607 vdd.n2587 16.2531
R12724 vdd.n2628 vdd.n2587 16.2531
R12725 vdd.n2628 vdd.n2627 16.2531
R12726 vdd.n2627 vdd.n2588 16.2531
R12727 vdd.n2617 vdd.n2588 16.2531
R12728 vdd.n2562 vdd.n2561 16.2531
R12729 vdd.n2561 vdd.n2541 16.2531
R12730 vdd.n2582 vdd.n2541 16.2531
R12731 vdd.n2582 vdd.n2581 16.2531
R12732 vdd.n2581 vdd.n2542 16.2531
R12733 vdd.n2571 vdd.n2542 16.2531
R12734 vdd.n2655 vdd.n2654 16.2531
R12735 vdd.n2654 vdd.n2634 16.2531
R12736 vdd.n2675 vdd.n2634 16.2531
R12737 vdd.n2675 vdd.n2674 16.2531
R12738 vdd.n2674 vdd.n2635 16.2531
R12739 vdd.n2664 vdd.n2635 16.2531
R12740 vdd.n2703 vdd.n2702 16.2531
R12741 vdd.n2702 vdd.n2682 16.2531
R12742 vdd.n2723 vdd.n2682 16.2531
R12743 vdd.n2723 vdd.n2722 16.2531
R12744 vdd.n2722 vdd.n2683 16.2531
R12745 vdd.n2712 vdd.n2683 16.2531
R12746 vdd.n2749 vdd.n2748 16.2531
R12747 vdd.n2748 vdd.n2728 16.2531
R12748 vdd.n2769 vdd.n2728 16.2531
R12749 vdd.n2769 vdd.n2768 16.2531
R12750 vdd.n2768 vdd.n2729 16.2531
R12751 vdd.n2758 vdd.n2729 16.2531
R12752 vdd.n1004 vdd.n992 16.2531
R12753 vdd.n1016 vdd.n992 16.2531
R12754 vdd.n1020 vdd.n1019 16.2531
R12755 vdd.n1021 vdd.n1020 16.2531
R12756 vdd.n1021 vdd.n985 16.2531
R12757 vdd.n2891 vdd.n2890 16.2531
R12758 vdd.n2890 vdd.n2870 16.2531
R12759 vdd.n2911 vdd.n2870 16.2531
R12760 vdd.n2911 vdd.n2910 16.2531
R12761 vdd.n2910 vdd.n2871 16.2531
R12762 vdd.n2900 vdd.n2871 16.2531
R12763 vdd.n2844 vdd.n2843 16.2531
R12764 vdd.n2843 vdd.n2823 16.2531
R12765 vdd.n2864 vdd.n2823 16.2531
R12766 vdd.n2864 vdd.n2863 16.2531
R12767 vdd.n2863 vdd.n2824 16.2531
R12768 vdd.n2853 vdd.n2824 16.2531
R12769 vdd.n2798 vdd.n2797 16.2531
R12770 vdd.n2797 vdd.n2777 16.2531
R12771 vdd.n2818 vdd.n2777 16.2531
R12772 vdd.n2818 vdd.n2817 16.2531
R12773 vdd.n2817 vdd.n2778 16.2531
R12774 vdd.n2807 vdd.n2778 16.2531
R12775 vdd.n2938 vdd.n2937 16.2531
R12776 vdd.n2937 vdd.n2917 16.2531
R12777 vdd.n2958 vdd.n2917 16.2531
R12778 vdd.n2958 vdd.n2957 16.2531
R12779 vdd.n2957 vdd.n2918 16.2531
R12780 vdd.n2947 vdd.n2918 16.2531
R12781 vdd.n2986 vdd.n2985 16.2531
R12782 vdd.n2985 vdd.n2965 16.2531
R12783 vdd.n3006 vdd.n2965 16.2531
R12784 vdd.n3006 vdd.n3005 16.2531
R12785 vdd.n3005 vdd.n2966 16.2531
R12786 vdd.n2995 vdd.n2966 16.2531
R12787 vdd.n3032 vdd.n3031 16.2531
R12788 vdd.n3031 vdd.n3011 16.2531
R12789 vdd.n3052 vdd.n3011 16.2531
R12790 vdd.n3052 vdd.n3051 16.2531
R12791 vdd.n3051 vdd.n3012 16.2531
R12792 vdd.n3041 vdd.n3012 16.2531
R12793 vdd.n3126 vdd.n3125 16.2531
R12794 vdd.n3125 vdd.n3105 16.2531
R12795 vdd.n3146 vdd.n3105 16.2531
R12796 vdd.n3146 vdd.n3145 16.2531
R12797 vdd.n3145 vdd.n3106 16.2531
R12798 vdd.n3135 vdd.n3106 16.2531
R12799 vdd.n3080 vdd.n3079 16.2531
R12800 vdd.n3079 vdd.n3059 16.2531
R12801 vdd.n3100 vdd.n3059 16.2531
R12802 vdd.n3100 vdd.n3099 16.2531
R12803 vdd.n3099 vdd.n3060 16.2531
R12804 vdd.n3089 vdd.n3060 16.2531
R12805 vdd.n3173 vdd.n3172 16.2531
R12806 vdd.n3172 vdd.n3152 16.2531
R12807 vdd.n3193 vdd.n3152 16.2531
R12808 vdd.n3193 vdd.n3192 16.2531
R12809 vdd.n3192 vdd.n3153 16.2531
R12810 vdd.n3182 vdd.n3153 16.2531
R12811 vdd.n3221 vdd.n3220 16.2531
R12812 vdd.n3220 vdd.n3200 16.2531
R12813 vdd.n3241 vdd.n3200 16.2531
R12814 vdd.n3241 vdd.n3240 16.2531
R12815 vdd.n3240 vdd.n3201 16.2531
R12816 vdd.n3230 vdd.n3201 16.2531
R12817 vdd.n3267 vdd.n3266 16.2531
R12818 vdd.n3266 vdd.n3246 16.2531
R12819 vdd.n3287 vdd.n3246 16.2531
R12820 vdd.n3287 vdd.n3286 16.2531
R12821 vdd.n3286 vdd.n3247 16.2531
R12822 vdd.n3276 vdd.n3247 16.2531
R12823 vdd.n768 vdd.n756 16.2531
R12824 vdd.n780 vdd.n756 16.2531
R12825 vdd.n784 vdd.n783 16.2531
R12826 vdd.n785 vdd.n784 16.2531
R12827 vdd.n785 vdd.n749 16.2531
R12828 vdd.n3362 vdd.n3361 16.2531
R12829 vdd.n3361 vdd.n3341 16.2531
R12830 vdd.n3382 vdd.n3341 16.2531
R12831 vdd.n3382 vdd.n3381 16.2531
R12832 vdd.n3381 vdd.n3342 16.2531
R12833 vdd.n3371 vdd.n3342 16.2531
R12834 vdd.n3316 vdd.n3315 16.2531
R12835 vdd.n3315 vdd.n3295 16.2531
R12836 vdd.n3336 vdd.n3295 16.2531
R12837 vdd.n3336 vdd.n3335 16.2531
R12838 vdd.n3335 vdd.n3296 16.2531
R12839 vdd.n3325 vdd.n3296 16.2531
R12840 vdd.n3409 vdd.n3408 16.2531
R12841 vdd.n3408 vdd.n3388 16.2531
R12842 vdd.n3429 vdd.n3388 16.2531
R12843 vdd.n3429 vdd.n3428 16.2531
R12844 vdd.n3428 vdd.n3389 16.2531
R12845 vdd.n3418 vdd.n3389 16.2531
R12846 vdd.n3457 vdd.n3456 16.2531
R12847 vdd.n3456 vdd.n3436 16.2531
R12848 vdd.n3477 vdd.n3436 16.2531
R12849 vdd.n3477 vdd.n3476 16.2531
R12850 vdd.n3476 vdd.n3437 16.2531
R12851 vdd.n3466 vdd.n3437 16.2531
R12852 vdd.n3503 vdd.n3502 16.2531
R12853 vdd.n3502 vdd.n3482 16.2531
R12854 vdd.n3523 vdd.n3482 16.2531
R12855 vdd.n3523 vdd.n3522 16.2531
R12856 vdd.n3522 vdd.n3483 16.2531
R12857 vdd.n3512 vdd.n3483 16.2531
R12858 vdd.n585 vdd.n584 16.2531
R12859 vdd.n584 vdd.n564 16.2531
R12860 vdd.n605 vdd.n564 16.2531
R12861 vdd.n605 vdd.n604 16.2531
R12862 vdd.n604 vdd.n565 16.2531
R12863 vdd.n594 vdd.n565 16.2531
R12864 vdd.n3598 vdd.n3597 16.2531
R12865 vdd.n3597 vdd.n3577 16.2531
R12866 vdd.n3618 vdd.n3577 16.2531
R12867 vdd.n3618 vdd.n3617 16.2531
R12868 vdd.n3617 vdd.n3578 16.2531
R12869 vdd.n3607 vdd.n3578 16.2531
R12870 vdd.n3552 vdd.n3551 16.2531
R12871 vdd.n3551 vdd.n3531 16.2531
R12872 vdd.n3572 vdd.n3531 16.2531
R12873 vdd.n3572 vdd.n3571 16.2531
R12874 vdd.n3571 vdd.n3532 16.2531
R12875 vdd.n3561 vdd.n3532 16.2531
R12876 vdd.n6612 vdd.n6611 16.2531
R12877 vdd.n6611 vdd.n6591 16.2531
R12878 vdd.n6632 vdd.n6591 16.2531
R12879 vdd.n6632 vdd.n6631 16.2531
R12880 vdd.n6631 vdd.n6592 16.2531
R12881 vdd.n6621 vdd.n6592 16.2531
R12882 vdd.n6566 vdd.n6565 16.2531
R12883 vdd.n6565 vdd.n6545 16.2531
R12884 vdd.n6586 vdd.n6545 16.2531
R12885 vdd.n6586 vdd.n6585 16.2531
R12886 vdd.n6585 vdd.n6546 16.2531
R12887 vdd.n6575 vdd.n6546 16.2531
R12888 vdd.n9626 vdd.n9625 16.2531
R12889 vdd.n9625 vdd.n9605 16.2531
R12890 vdd.n9646 vdd.n9605 16.2531
R12891 vdd.n9646 vdd.n9645 16.2531
R12892 vdd.n9645 vdd.n9606 16.2531
R12893 vdd.n9635 vdd.n9606 16.2531
R12894 vdd.n9580 vdd.n9579 16.2531
R12895 vdd.n9579 vdd.n9559 16.2531
R12896 vdd.n9600 vdd.n9559 16.2531
R12897 vdd.n9600 vdd.n9599 16.2531
R12898 vdd.n9599 vdd.n9560 16.2531
R12899 vdd.n9589 vdd.n9560 16.2531
R12900 vdd.n9672 vdd.n9671 16.2531
R12901 vdd.n9671 vdd.n9651 16.2531
R12902 vdd.n9692 vdd.n9651 16.2531
R12903 vdd.n9692 vdd.n9691 16.2531
R12904 vdd.n9691 vdd.n9652 16.2531
R12905 vdd.n9681 vdd.n9652 16.2531
R12906 vdd.n9718 vdd.n9717 16.2531
R12907 vdd.n9717 vdd.n9697 16.2531
R12908 vdd.n9738 vdd.n9697 16.2531
R12909 vdd.n9738 vdd.n9737 16.2531
R12910 vdd.n9737 vdd.n9698 16.2531
R12911 vdd.n9727 vdd.n9698 16.2531
R12912 vdd.n9816 vdd.n9815 16.2531
R12913 vdd.n9815 vdd.n9795 16.2531
R12914 vdd.n9836 vdd.n9795 16.2531
R12915 vdd.n9836 vdd.n9835 16.2531
R12916 vdd.n9835 vdd.n9796 16.2531
R12917 vdd.n9825 vdd.n9796 16.2531
R12918 vdd.n9862 vdd.n9861 16.2531
R12919 vdd.n9861 vdd.n9841 16.2531
R12920 vdd.n9882 vdd.n9841 16.2531
R12921 vdd.n9882 vdd.n9881 16.2531
R12922 vdd.n9881 vdd.n9842 16.2531
R12923 vdd.n9871 vdd.n9842 16.2531
R12924 vdd.n9908 vdd.n9907 16.2531
R12925 vdd.n9907 vdd.n9887 16.2531
R12926 vdd.n9928 vdd.n9887 16.2531
R12927 vdd.n9928 vdd.n9927 16.2531
R12928 vdd.n9927 vdd.n9888 16.2531
R12929 vdd.n9917 vdd.n9888 16.2531
R12930 vdd.n9954 vdd.n9953 16.2531
R12931 vdd.n9953 vdd.n9933 16.2531
R12932 vdd.n9974 vdd.n9933 16.2531
R12933 vdd.n9974 vdd.n9973 16.2531
R12934 vdd.n9973 vdd.n9934 16.2531
R12935 vdd.n9963 vdd.n9934 16.2531
R12936 vdd.n10052 vdd.n10051 16.2531
R12937 vdd.n10051 vdd.n10031 16.2531
R12938 vdd.n10072 vdd.n10031 16.2531
R12939 vdd.n10072 vdd.n10071 16.2531
R12940 vdd.n10071 vdd.n10032 16.2531
R12941 vdd.n10061 vdd.n10032 16.2531
R12942 vdd.n68 vdd.n67 16.2531
R12943 vdd.n67 vdd.n47 16.2531
R12944 vdd.n88 vdd.n47 16.2531
R12945 vdd.n88 vdd.n87 16.2531
R12946 vdd.n87 vdd.n48 16.2531
R12947 vdd.n77 vdd.n48 16.2531
R12948 vdd.n22 vdd.n21 16.2531
R12949 vdd.n21 vdd.n1 16.2531
R12950 vdd.n42 vdd.n1 16.2531
R12951 vdd.n42 vdd.n41 16.2531
R12952 vdd.n41 vdd.n2 16.2531
R12953 vdd.n31 vdd.n2 16.2531
R12954 vdd.n10098 vdd.n10097 16.2531
R12955 vdd.n10097 vdd.n10077 16.2531
R12956 vdd.n10118 vdd.n10077 16.2531
R12957 vdd.n10118 vdd.n10117 16.2531
R12958 vdd.n10117 vdd.n10078 16.2531
R12959 vdd.n10107 vdd.n10078 16.2531
R12960 vdd.n10146 vdd.n10145 16.2531
R12961 vdd.n10145 vdd.n10125 16.2531
R12962 vdd.n10166 vdd.n10125 16.2531
R12963 vdd.n10166 vdd.n10165 16.2531
R12964 vdd.n10165 vdd.n10126 16.2531
R12965 vdd.n10155 vdd.n10126 16.2531
R12966 vdd.n10192 vdd.n10191 16.2531
R12967 vdd.n10191 vdd.n10171 16.2531
R12968 vdd.n10212 vdd.n10171 16.2531
R12969 vdd.n10212 vdd.n10211 16.2531
R12970 vdd.n10211 vdd.n10172 16.2531
R12971 vdd.n10201 vdd.n10172 16.2531
R12972 vdd.n9999 vdd.n9987 16.2531
R12973 vdd.n10011 vdd.n9987 16.2531
R12974 vdd.n10015 vdd.n10014 16.2531
R12975 vdd.n10016 vdd.n10015 16.2531
R12976 vdd.n10016 vdd.n9980 16.2531
R12977 vdd.n10334 vdd.n10333 16.2531
R12978 vdd.n10333 vdd.n10313 16.2531
R12979 vdd.n10354 vdd.n10313 16.2531
R12980 vdd.n10354 vdd.n10353 16.2531
R12981 vdd.n10353 vdd.n10314 16.2531
R12982 vdd.n10343 vdd.n10314 16.2531
R12983 vdd.n10287 vdd.n10286 16.2531
R12984 vdd.n10286 vdd.n10266 16.2531
R12985 vdd.n10307 vdd.n10266 16.2531
R12986 vdd.n10307 vdd.n10306 16.2531
R12987 vdd.n10306 vdd.n10267 16.2531
R12988 vdd.n10296 vdd.n10267 16.2531
R12989 vdd.n10241 vdd.n10240 16.2531
R12990 vdd.n10240 vdd.n10220 16.2531
R12991 vdd.n10261 vdd.n10220 16.2531
R12992 vdd.n10261 vdd.n10260 16.2531
R12993 vdd.n10260 vdd.n10221 16.2531
R12994 vdd.n10250 vdd.n10221 16.2531
R12995 vdd.n10381 vdd.n10380 16.2531
R12996 vdd.n10380 vdd.n10360 16.2531
R12997 vdd.n10401 vdd.n10360 16.2531
R12998 vdd.n10401 vdd.n10400 16.2531
R12999 vdd.n10400 vdd.n10361 16.2531
R13000 vdd.n10390 vdd.n10361 16.2531
R13001 vdd.n10429 vdd.n10428 16.2531
R13002 vdd.n10428 vdd.n10408 16.2531
R13003 vdd.n10449 vdd.n10408 16.2531
R13004 vdd.n10449 vdd.n10448 16.2531
R13005 vdd.n10448 vdd.n10409 16.2531
R13006 vdd.n10438 vdd.n10409 16.2531
R13007 vdd.n10475 vdd.n10474 16.2531
R13008 vdd.n10474 vdd.n10454 16.2531
R13009 vdd.n10495 vdd.n10454 16.2531
R13010 vdd.n10495 vdd.n10494 16.2531
R13011 vdd.n10494 vdd.n10455 16.2531
R13012 vdd.n10484 vdd.n10455 16.2531
R13013 vdd.n10569 vdd.n10568 16.2531
R13014 vdd.n10568 vdd.n10548 16.2531
R13015 vdd.n10589 vdd.n10548 16.2531
R13016 vdd.n10589 vdd.n10588 16.2531
R13017 vdd.n10588 vdd.n10549 16.2531
R13018 vdd.n10578 vdd.n10549 16.2531
R13019 vdd.n10523 vdd.n10522 16.2531
R13020 vdd.n10522 vdd.n10502 16.2531
R13021 vdd.n10543 vdd.n10502 16.2531
R13022 vdd.n10543 vdd.n10542 16.2531
R13023 vdd.n10542 vdd.n10503 16.2531
R13024 vdd.n10532 vdd.n10503 16.2531
R13025 vdd.n10616 vdd.n10615 16.2531
R13026 vdd.n10615 vdd.n10595 16.2531
R13027 vdd.n10636 vdd.n10595 16.2531
R13028 vdd.n10636 vdd.n10635 16.2531
R13029 vdd.n10635 vdd.n10596 16.2531
R13030 vdd.n10625 vdd.n10596 16.2531
R13031 vdd.n10664 vdd.n10663 16.2531
R13032 vdd.n10663 vdd.n10643 16.2531
R13033 vdd.n10684 vdd.n10643 16.2531
R13034 vdd.n10684 vdd.n10683 16.2531
R13035 vdd.n10683 vdd.n10644 16.2531
R13036 vdd.n10673 vdd.n10644 16.2531
R13037 vdd.n10710 vdd.n10709 16.2531
R13038 vdd.n10709 vdd.n10689 16.2531
R13039 vdd.n10730 vdd.n10689 16.2531
R13040 vdd.n10730 vdd.n10729 16.2531
R13041 vdd.n10729 vdd.n10690 16.2531
R13042 vdd.n10719 vdd.n10690 16.2531
R13043 vdd.n9763 vdd.n9751 16.2531
R13044 vdd.n9775 vdd.n9751 16.2531
R13045 vdd.n9779 vdd.n9778 16.2531
R13046 vdd.n9780 vdd.n9779 16.2531
R13047 vdd.n9780 vdd.n9744 16.2531
R13048 vdd.n10805 vdd.n10804 16.2531
R13049 vdd.n10804 vdd.n10784 16.2531
R13050 vdd.n10825 vdd.n10784 16.2531
R13051 vdd.n10825 vdd.n10824 16.2531
R13052 vdd.n10824 vdd.n10785 16.2531
R13053 vdd.n10814 vdd.n10785 16.2531
R13054 vdd.n10759 vdd.n10758 16.2531
R13055 vdd.n10758 vdd.n10738 16.2531
R13056 vdd.n10779 vdd.n10738 16.2531
R13057 vdd.n10779 vdd.n10778 16.2531
R13058 vdd.n10778 vdd.n10739 16.2531
R13059 vdd.n10768 vdd.n10739 16.2531
R13060 vdd.n10852 vdd.n10851 16.2531
R13061 vdd.n10851 vdd.n10831 16.2531
R13062 vdd.n10872 vdd.n10831 16.2531
R13063 vdd.n10872 vdd.n10871 16.2531
R13064 vdd.n10871 vdd.n10832 16.2531
R13065 vdd.n10861 vdd.n10832 16.2531
R13066 vdd.n10900 vdd.n10899 16.2531
R13067 vdd.n10899 vdd.n10879 16.2531
R13068 vdd.n10920 vdd.n10879 16.2531
R13069 vdd.n10920 vdd.n10919 16.2531
R13070 vdd.n10919 vdd.n10880 16.2531
R13071 vdd.n10909 vdd.n10880 16.2531
R13072 vdd.n10946 vdd.n10945 16.2531
R13073 vdd.n10945 vdd.n10925 16.2531
R13074 vdd.n10966 vdd.n10925 16.2531
R13075 vdd.n10966 vdd.n10965 16.2531
R13076 vdd.n10965 vdd.n10926 16.2531
R13077 vdd.n10955 vdd.n10926 16.2531
R13078 vdd.n10994 vdd.n10993 16.2531
R13079 vdd.n10993 vdd.n10974 16.2531
R13080 vdd.n11015 vdd.n10974 16.2531
R13081 vdd.n11015 vdd.n11014 16.2531
R13082 vdd.n11014 vdd.n10975 16.2531
R13083 vdd.n11010 vdd.n10975 16.2531
R13084 vdd.n11039 vdd.n11038 16.2531
R13085 vdd.n11038 vdd.n11019 16.2531
R13086 vdd.n11060 vdd.n11019 16.2531
R13087 vdd.n11060 vdd.n11059 16.2531
R13088 vdd.n11059 vdd.n11020 16.2531
R13089 vdd.n11055 vdd.n11020 16.2531
R13090 vdd.n11089 vdd.n11088 16.2531
R13091 vdd.n11088 vdd.n11069 16.2531
R13092 vdd.n11110 vdd.n11069 16.2531
R13093 vdd.n11110 vdd.n11109 16.2531
R13094 vdd.n11109 vdd.n11070 16.2531
R13095 vdd.n11105 vdd.n11070 16.2531
R13096 vdd.n11135 vdd.n11134 16.2531
R13097 vdd.n11134 vdd.n11115 16.2531
R13098 vdd.n11156 vdd.n11115 16.2531
R13099 vdd.n11156 vdd.n11155 16.2531
R13100 vdd.n11155 vdd.n11116 16.2531
R13101 vdd.n11151 vdd.n11116 16.2531
R13102 vdd.n11183 vdd.n11182 16.2531
R13103 vdd.n11182 vdd.n11163 16.2531
R13104 vdd.n11204 vdd.n11163 16.2531
R13105 vdd.n11204 vdd.n11203 16.2531
R13106 vdd.n11203 vdd.n11164 16.2531
R13107 vdd.n11199 vdd.n11164 16.2531
R13108 vdd.n466 vdd.n423 16.2531
R13109 vdd.n462 vdd.n423 16.2531
R13110 vdd.n462 vdd.n461 16.2531
R13111 vdd.n459 vdd.n430 16.2531
R13112 vdd.n455 vdd.n430 16.2531
R13113 vdd.n11230 vdd.n11229 16.2531
R13114 vdd.n11229 vdd.n11210 16.2531
R13115 vdd.n11251 vdd.n11210 16.2531
R13116 vdd.n11251 vdd.n11250 16.2531
R13117 vdd.n11250 vdd.n11211 16.2531
R13118 vdd.n11246 vdd.n11211 16.2531
R13119 vdd.n11275 vdd.n11274 16.2531
R13120 vdd.n11274 vdd.n11255 16.2531
R13121 vdd.n11296 vdd.n11255 16.2531
R13122 vdd.n11296 vdd.n11295 16.2531
R13123 vdd.n11295 vdd.n11256 16.2531
R13124 vdd.n11291 vdd.n11256 16.2531
R13125 vdd.n11321 vdd.n11320 16.2531
R13126 vdd.n11320 vdd.n11301 16.2531
R13127 vdd.n11342 vdd.n11301 16.2531
R13128 vdd.n11342 vdd.n11341 16.2531
R13129 vdd.n11341 vdd.n11302 16.2531
R13130 vdd.n11337 vdd.n11302 16.2531
R13131 vdd.n11372 vdd.n11371 16.2531
R13132 vdd.n11371 vdd.n11352 16.2531
R13133 vdd.n11393 vdd.n11352 16.2531
R13134 vdd.n11393 vdd.n11392 16.2531
R13135 vdd.n11392 vdd.n11353 16.2531
R13136 vdd.n11388 vdd.n11353 16.2531
R13137 vdd.n11418 vdd.n11417 16.2531
R13138 vdd.n11417 vdd.n11398 16.2531
R13139 vdd.n11439 vdd.n11398 16.2531
R13140 vdd.n11439 vdd.n11438 16.2531
R13141 vdd.n11438 vdd.n11399 16.2531
R13142 vdd.n11434 vdd.n11399 16.2531
R13143 vdd.n11466 vdd.n11465 16.2531
R13144 vdd.n11465 vdd.n11446 16.2531
R13145 vdd.n11487 vdd.n11446 16.2531
R13146 vdd.n11487 vdd.n11486 16.2531
R13147 vdd.n11486 vdd.n11447 16.2531
R13148 vdd.n11482 vdd.n11447 16.2531
R13149 vdd.n11512 vdd.n11511 16.2531
R13150 vdd.n11511 vdd.n11492 16.2531
R13151 vdd.n11533 vdd.n11492 16.2531
R13152 vdd.n11533 vdd.n11532 16.2531
R13153 vdd.n11532 vdd.n11493 16.2531
R13154 vdd.n11528 vdd.n11493 16.2531
R13155 vdd.n11557 vdd.n11556 16.2531
R13156 vdd.n11556 vdd.n11537 16.2531
R13157 vdd.n11578 vdd.n11537 16.2531
R13158 vdd.n11578 vdd.n11577 16.2531
R13159 vdd.n11577 vdd.n11538 16.2531
R13160 vdd.n11573 vdd.n11538 16.2531
R13161 vdd.n11607 vdd.n11606 16.2531
R13162 vdd.n11606 vdd.n11587 16.2531
R13163 vdd.n11628 vdd.n11587 16.2531
R13164 vdd.n11628 vdd.n11627 16.2531
R13165 vdd.n11627 vdd.n11588 16.2531
R13166 vdd.n11623 vdd.n11588 16.2531
R13167 vdd.n11653 vdd.n11652 16.2531
R13168 vdd.n11652 vdd.n11633 16.2531
R13169 vdd.n11674 vdd.n11633 16.2531
R13170 vdd.n11674 vdd.n11673 16.2531
R13171 vdd.n11673 vdd.n11634 16.2531
R13172 vdd.n11669 vdd.n11634 16.2531
R13173 vdd.n11701 vdd.n11700 16.2531
R13174 vdd.n11700 vdd.n11681 16.2531
R13175 vdd.n11722 vdd.n11681 16.2531
R13176 vdd.n11722 vdd.n11721 16.2531
R13177 vdd.n11721 vdd.n11682 16.2531
R13178 vdd.n11717 vdd.n11682 16.2531
R13179 vdd.n231 vdd.n188 16.2531
R13180 vdd.n227 vdd.n188 16.2531
R13181 vdd.n227 vdd.n226 16.2531
R13182 vdd.n224 vdd.n195 16.2531
R13183 vdd.n220 vdd.n195 16.2531
R13184 vdd.n11748 vdd.n11747 16.2531
R13185 vdd.n11747 vdd.n11728 16.2531
R13186 vdd.n11769 vdd.n11728 16.2531
R13187 vdd.n11769 vdd.n11768 16.2531
R13188 vdd.n11768 vdd.n11729 16.2531
R13189 vdd.n11764 vdd.n11729 16.2531
R13190 vdd.n11793 vdd.n11792 16.2531
R13191 vdd.n11792 vdd.n11773 16.2531
R13192 vdd.n11814 vdd.n11773 16.2531
R13193 vdd.n11814 vdd.n11813 16.2531
R13194 vdd.n11813 vdd.n11774 16.2531
R13195 vdd.n11809 vdd.n11774 16.2531
R13196 vdd.n11843 vdd.n11842 16.2531
R13197 vdd.n11842 vdd.n11823 16.2531
R13198 vdd.n11864 vdd.n11823 16.2531
R13199 vdd.n11864 vdd.n11863 16.2531
R13200 vdd.n11863 vdd.n11824 16.2531
R13201 vdd.n11859 vdd.n11824 16.2531
R13202 vdd.n11889 vdd.n11888 16.2531
R13203 vdd.n11888 vdd.n11869 16.2531
R13204 vdd.n11910 vdd.n11869 16.2531
R13205 vdd.n11910 vdd.n11909 16.2531
R13206 vdd.n11909 vdd.n11870 16.2531
R13207 vdd.n11905 vdd.n11870 16.2531
R13208 vdd.n11937 vdd.n11936 16.2531
R13209 vdd.n11936 vdd.n11917 16.2531
R13210 vdd.n11958 vdd.n11917 16.2531
R13211 vdd.n11958 vdd.n11957 16.2531
R13212 vdd.n11957 vdd.n11918 16.2531
R13213 vdd.n11953 vdd.n11918 16.2531
R13214 vdd.n7476 vdd.n7475 13.9199
R13215 vdd.n7241 vdd.n7240 13.9199
R13216 vdd.n4462 vdd.n4461 13.9199
R13217 vdd.n4227 vdd.n4226 13.9199
R13218 vdd.n1448 vdd.n1447 13.9199
R13219 vdd.n1213 vdd.n1212 13.9199
R13220 vdd.n460 vdd.n459 13.9199
R13221 vdd.n225 vdd.n224 13.9199
R13222 vdd.n7046 vdd.n7044 13.9189
R13223 vdd.n6810 vdd.n6808 13.9189
R13224 vdd.n4032 vdd.n4030 13.9189
R13225 vdd.n3796 vdd.n3794 13.9189
R13226 vdd.n1018 vdd.n1016 13.9189
R13227 vdd.n782 vdd.n780 13.9189
R13228 vdd.n10013 vdd.n10011 13.9189
R13229 vdd.n9777 vdd.n9775 13.9189
R13230 vdd.n7483 vdd.n7482 12.4637
R13231 vdd.n7248 vdd.n7247 12.4637
R13232 vdd.n7058 vdd.n7013 12.4637
R13233 vdd.n6822 vdd.n6777 12.4637
R13234 vdd.n4469 vdd.n4468 12.4637
R13235 vdd.n4234 vdd.n4233 12.4637
R13236 vdd.n4044 vdd.n3999 12.4637
R13237 vdd.n3808 vdd.n3763 12.4637
R13238 vdd.n1455 vdd.n1454 12.4637
R13239 vdd.n1220 vdd.n1219 12.4637
R13240 vdd.n1030 vdd.n985 12.4637
R13241 vdd.n794 vdd.n749 12.4637
R13242 vdd.n10025 vdd.n9980 12.4637
R13243 vdd.n9789 vdd.n9744 12.4637
R13244 vdd.n467 vdd.n466 12.4637
R13245 vdd.n232 vdd.n231 12.4637
R13246 vdd vdd.n7436 9.01037
R13247 vdd vdd.n7201 9.01037
R13248 vdd vdd.n4422 9.01037
R13249 vdd vdd.n4187 9.01037
R13250 vdd vdd.n1408 9.01037
R13251 vdd vdd.n1173 9.01037
R13252 vdd vdd.n420 9.01037
R13253 vdd vdd.n185 9.01037
R13254 vdd.n7060 vdd.n7011 9.0005
R13255 vdd.n6824 vdd.n6775 9.0005
R13256 vdd.n4046 vdd.n3997 9.0005
R13257 vdd.n3810 vdd.n3761 9.0005
R13258 vdd.n1032 vdd.n983 9.0005
R13259 vdd.n796 vdd.n747 9.0005
R13260 vdd.n10027 vdd.n9978 9.0005
R13261 vdd.n9791 vdd.n9742 9.0005
R13262 vdd.n8567 vdd.n8520 6.24557
R13263 vdd.n5553 vdd.n5506 6.24557
R13264 vdd.n2539 vdd.n2492 6.24557
R13265 vdd.n11961 vdd.n11960 6.24557
R13266 vdd.n3619 vdd 5.95856
R13267 vdd.n9647 vdd 5.95856
R13268 vdd.n6633 vdd 5.76119
R13269 vdd.n9556 vdd.n6682 4.70938
R13270 vdd.n6542 vdd.n3668 4.70938
R13271 vdd.n3528 vdd.n654 4.70938
R13272 vdd.n10972 vdd.n10971 4.70938
R13273 vdd.n6587 vdd.n6543 4.23159
R13274 vdd.n7904 vdd.n7903 4.08685
R13275 vdd.n8896 vdd.n8849 4.08685
R13276 vdd.n4890 vdd.n4889 4.08685
R13277 vdd.n5882 vdd.n5835 4.08685
R13278 vdd.n1876 vdd.n1875 4.08685
R13279 vdd.n2868 vdd.n2821 4.08685
R13280 vdd.n10311 vdd.n10264 4.08685
R13281 vdd.n11344 vdd.n11343 4.08685
R13282 vdd.n3573 vdd.n3529 4.03422
R13283 vdd.n9601 vdd.n9557 4.03422
R13284 vdd.n7622 vdd.n7621 2.95445
R13285 vdd.n8140 vdd.n8139 2.95445
R13286 vdd.n8376 vdd.n8375 2.95445
R13287 vdd.n8657 vdd.n8613 2.95445
R13288 vdd.n9175 vdd.n9131 2.95445
R13289 vdd.n9411 vdd.n9367 2.95445
R13290 vdd.n4608 vdd.n4607 2.95445
R13291 vdd.n5126 vdd.n5125 2.95445
R13292 vdd.n5362 vdd.n5361 2.95445
R13293 vdd.n5643 vdd.n5599 2.95445
R13294 vdd.n6161 vdd.n6117 2.95445
R13295 vdd.n6397 vdd.n6353 2.95445
R13296 vdd.n1594 vdd.n1593 2.95445
R13297 vdd.n2112 vdd.n2111 2.95445
R13298 vdd.n2348 vdd.n2347 2.95445
R13299 vdd.n2629 vdd.n2585 2.95445
R13300 vdd.n3147 vdd.n3103 2.95445
R13301 vdd.n3383 vdd.n3339 2.95445
R13302 vdd.n89 vdd.n45 2.95445
R13303 vdd.n10590 vdd.n10546 2.95445
R13304 vdd.n10826 vdd.n10782 2.95445
R13305 vdd.n11062 vdd.n11061 2.95445
R13306 vdd.n11580 vdd.n11579 2.95445
R13307 vdd.n11816 vdd.n11815 2.95445
R13308 vdd.n7905 vdd.n7904 2.33849
R13309 vdd.n8940 vdd.n8896 2.33849
R13310 vdd.n4891 vdd.n4890 2.33849
R13311 vdd.n5926 vdd.n5882 2.33849
R13312 vdd.n1877 vdd.n1876 2.33849
R13313 vdd.n2912 vdd.n2868 2.33849
R13314 vdd.n10355 vdd.n10311 2.33849
R13315 vdd.n11345 vdd.n11344 2.33849
R13316 vdd.n10971 vdd 2.27025
R13317 vdd.n9557 vdd.n9556 1.54656
R13318 vdd.n6543 vdd.n6542 1.54656
R13319 vdd.n3529 vdd.n3528 1.54656
R13320 vdd.n9556 vdd.n9555 1.53669
R13321 vdd.n6542 vdd.n6541 1.53669
R13322 vdd.n3528 vdd.n3527 1.53669
R13323 vdd.n10971 vdd.n10970 1.53669
R13324 vdd.n7673 vdd.n7672 1.50544
R13325 vdd.n7956 vdd.n7955 1.50544
R13326 vdd.n8050 vdd.n8049 1.50544
R13327 vdd.n8191 vdd.n8190 1.50544
R13328 vdd.n8427 vdd.n8426 1.50544
R13329 vdd.n8708 vdd.n8707 1.50544
R13330 vdd.n8991 vdd.n8990 1.50544
R13331 vdd.n9085 vdd.n9084 1.50544
R13332 vdd.n9226 vdd.n9225 1.50544
R13333 vdd.n9462 vdd.n9461 1.50544
R13334 vdd.n4659 vdd.n4658 1.50544
R13335 vdd.n4942 vdd.n4941 1.50544
R13336 vdd.n5036 vdd.n5035 1.50544
R13337 vdd.n5177 vdd.n5176 1.50544
R13338 vdd.n5413 vdd.n5412 1.50544
R13339 vdd.n5694 vdd.n5693 1.50544
R13340 vdd.n5977 vdd.n5976 1.50544
R13341 vdd.n6071 vdd.n6070 1.50544
R13342 vdd.n6212 vdd.n6211 1.50544
R13343 vdd.n6448 vdd.n6447 1.50544
R13344 vdd.n1645 vdd.n1644 1.50544
R13345 vdd.n1928 vdd.n1927 1.50544
R13346 vdd.n2022 vdd.n2021 1.50544
R13347 vdd.n2163 vdd.n2162 1.50544
R13348 vdd.n2399 vdd.n2398 1.50544
R13349 vdd.n2680 vdd.n2679 1.50544
R13350 vdd.n2963 vdd.n2962 1.50544
R13351 vdd.n3057 vdd.n3056 1.50544
R13352 vdd.n3198 vdd.n3197 1.50544
R13353 vdd.n3434 vdd.n3433 1.50544
R13354 vdd.n10123 vdd.n10122 1.50544
R13355 vdd.n10406 vdd.n10405 1.50544
R13356 vdd.n10500 vdd.n10499 1.50544
R13357 vdd.n10641 vdd.n10640 1.50544
R13358 vdd.n10877 vdd.n10876 1.50544
R13359 vdd.n11113 vdd.n11112 1.50544
R13360 vdd.n11396 vdd.n11395 1.50544
R13361 vdd.n11490 vdd.n11489 1.50544
R13362 vdd.n11631 vdd.n11630 1.50544
R13363 vdd.n11867 vdd.n11866 1.50544
R13364 vdd.n7672 vdd.n7671 0.904283
R13365 vdd.n7673 vdd.n7532 0.904283
R13366 vdd.n7766 vdd.n7765 0.904283
R13367 vdd.n7955 vdd.n7954 0.904283
R13368 vdd.n7956 vdd.n7389 0.904283
R13369 vdd.n8049 vdd.n8048 0.904283
R13370 vdd.n8190 vdd.n8189 0.904283
R13371 vdd.n8191 vdd.n7297 0.904283
R13372 vdd.n8284 vdd.n8283 0.904283
R13373 vdd.n8426 vdd.n8425 0.904283
R13374 vdd.n8427 vdd.n7154 0.904283
R13375 vdd.n8520 vdd.n8519 0.904283
R13376 vdd.n8707 vdd.n8706 0.904283
R13377 vdd.n8708 vdd.n7108 0.904283
R13378 vdd.n8801 vdd.n8800 0.904283
R13379 vdd.n8990 vdd.n8989 0.904283
R13380 vdd.n8991 vdd.n6964 0.904283
R13381 vdd.n9084 vdd.n9083 0.904283
R13382 vdd.n9225 vdd.n9224 0.904283
R13383 vdd.n9226 vdd.n6872 0.904283
R13384 vdd.n9319 vdd.n9318 0.904283
R13385 vdd.n9461 vdd.n9460 0.904283
R13386 vdd.n9462 vdd.n6728 0.904283
R13387 vdd.n9555 vdd.n9554 0.904283
R13388 vdd.n4658 vdd.n4657 0.904283
R13389 vdd.n4659 vdd.n4518 0.904283
R13390 vdd.n4752 vdd.n4751 0.904283
R13391 vdd.n4941 vdd.n4940 0.904283
R13392 vdd.n4942 vdd.n4375 0.904283
R13393 vdd.n5035 vdd.n5034 0.904283
R13394 vdd.n5176 vdd.n5175 0.904283
R13395 vdd.n5177 vdd.n4283 0.904283
R13396 vdd.n5270 vdd.n5269 0.904283
R13397 vdd.n5412 vdd.n5411 0.904283
R13398 vdd.n5413 vdd.n4140 0.904283
R13399 vdd.n5506 vdd.n5505 0.904283
R13400 vdd.n5693 vdd.n5692 0.904283
R13401 vdd.n5694 vdd.n4094 0.904283
R13402 vdd.n5787 vdd.n5786 0.904283
R13403 vdd.n5976 vdd.n5975 0.904283
R13404 vdd.n5977 vdd.n3950 0.904283
R13405 vdd.n6070 vdd.n6069 0.904283
R13406 vdd.n6211 vdd.n6210 0.904283
R13407 vdd.n6212 vdd.n3858 0.904283
R13408 vdd.n6305 vdd.n6304 0.904283
R13409 vdd.n6447 vdd.n6446 0.904283
R13410 vdd.n6448 vdd.n3714 0.904283
R13411 vdd.n6541 vdd.n6540 0.904283
R13412 vdd.n1644 vdd.n1643 0.904283
R13413 vdd.n1645 vdd.n1504 0.904283
R13414 vdd.n1738 vdd.n1737 0.904283
R13415 vdd.n1927 vdd.n1926 0.904283
R13416 vdd.n1928 vdd.n1361 0.904283
R13417 vdd.n2021 vdd.n2020 0.904283
R13418 vdd.n2162 vdd.n2161 0.904283
R13419 vdd.n2163 vdd.n1269 0.904283
R13420 vdd.n2256 vdd.n2255 0.904283
R13421 vdd.n2398 vdd.n2397 0.904283
R13422 vdd.n2399 vdd.n1126 0.904283
R13423 vdd.n2492 vdd.n2491 0.904283
R13424 vdd.n2679 vdd.n2678 0.904283
R13425 vdd.n2680 vdd.n1080 0.904283
R13426 vdd.n2773 vdd.n2772 0.904283
R13427 vdd.n2962 vdd.n2961 0.904283
R13428 vdd.n2963 vdd.n936 0.904283
R13429 vdd.n3056 vdd.n3055 0.904283
R13430 vdd.n3197 vdd.n3196 0.904283
R13431 vdd.n3198 vdd.n844 0.904283
R13432 vdd.n3291 vdd.n3290 0.904283
R13433 vdd.n3433 vdd.n3432 0.904283
R13434 vdd.n3434 vdd.n700 0.904283
R13435 vdd.n3527 vdd.n3526 0.904283
R13436 vdd.n10122 vdd.n10121 0.904283
R13437 vdd.n10123 vdd.n10075 0.904283
R13438 vdd.n10216 vdd.n10215 0.904283
R13439 vdd.n10405 vdd.n10404 0.904283
R13440 vdd.n10406 vdd.n9931 0.904283
R13441 vdd.n10499 vdd.n10498 0.904283
R13442 vdd.n10640 vdd.n10639 0.904283
R13443 vdd.n10641 vdd.n9839 0.904283
R13444 vdd.n10734 vdd.n10733 0.904283
R13445 vdd.n10876 vdd.n10875 0.904283
R13446 vdd.n10877 vdd.n9695 0.904283
R13447 vdd.n10970 vdd.n10969 0.904283
R13448 vdd.n11112 vdd.n11111 0.904283
R13449 vdd.n11113 vdd.n516 0.904283
R13450 vdd.n11206 vdd.n11205 0.904283
R13451 vdd.n11395 vdd.n11394 0.904283
R13452 vdd.n11396 vdd.n373 0.904283
R13453 vdd.n11489 vdd.n11488 0.904283
R13454 vdd.n11630 vdd.n11629 0.904283
R13455 vdd.n11631 vdd.n281 0.904283
R13456 vdd.n11724 vdd.n11723 0.904283
R13457 vdd.n11866 vdd.n11865 0.904283
R13458 vdd.n11867 vdd.n138 0.904283
R13459 vdd.n11960 vdd.n11959 0.904283
R13460 vdd.n7767 vdd.n7766 0.854122
R13461 vdd.n8285 vdd.n8284 0.854122
R13462 vdd.n8802 vdd.n8801 0.854122
R13463 vdd.n9320 vdd.n9319 0.854122
R13464 vdd.n4753 vdd.n4752 0.854122
R13465 vdd.n5271 vdd.n5270 0.854122
R13466 vdd.n5788 vdd.n5787 0.854122
R13467 vdd.n6306 vdd.n6305 0.854122
R13468 vdd.n1739 vdd.n1738 0.854122
R13469 vdd.n2257 vdd.n2256 0.854122
R13470 vdd.n2774 vdd.n2773 0.854122
R13471 vdd.n3292 vdd.n3291 0.854122
R13472 vdd.n10217 vdd.n10216 0.854122
R13473 vdd.n10735 vdd.n10734 0.854122
R13474 vdd.n11207 vdd.n11206 0.854122
R13475 vdd.n11725 vdd.n11724 0.854122
R13476 vdd vdd.n7435 0.76448
R13477 vdd vdd.n7200 0.76448
R13478 vdd vdd.n4421 0.76448
R13479 vdd vdd.n4186 0.76448
R13480 vdd vdd.n1407 0.76448
R13481 vdd vdd.n1172 0.76448
R13482 vdd vdd.n419 0.76448
R13483 vdd vdd.n184 0.76448
R13484 vdd vdd.n6681 0.752967
R13485 vdd vdd.n7343 0.752967
R13486 vdd vdd.n3667 0.752967
R13487 vdd vdd.n4329 0.752967
R13488 vdd vdd.n653 0.752967
R13489 vdd vdd.n1315 0.752967
R13490 vdd vdd.n562 0.752967
R13491 vdd vdd.n327 0.752967
R13492 vdd.n3529 vdd 0.724184
R13493 vdd.n6543 vdd 0.724184
R13494 vdd.n9557 vdd 0.724184
R13495 vdd vdd.n12007 0.711849
R13496 vdd vdd.n8566 0.698691
R13497 vdd vdd.n7010 0.698691
R13498 vdd vdd.n6918 0.698691
R13499 vdd vdd.n6774 0.698691
R13500 vdd vdd.n5552 0.698691
R13501 vdd vdd.n3996 0.698691
R13502 vdd vdd.n3904 0.698691
R13503 vdd vdd.n3760 0.698691
R13504 vdd vdd.n2538 0.698691
R13505 vdd vdd.n982 0.698691
R13506 vdd vdd.n890 0.698691
R13507 vdd vdd.n746 0.698691
R13508 vdd vdd.n9977 0.698691
R13509 vdd vdd.n9885 0.698691
R13510 vdd vdd.n9741 0.698691
R13511 vdd.n7672 vdd.n7625 0.697868
R13512 vdd.n7766 vdd.n7719 0.697868
R13513 vdd.n7955 vdd.n7908 0.697868
R13514 vdd.n8049 vdd.n8002 0.697868
R13515 vdd.n8190 vdd.n8143 0.697868
R13516 vdd.n8284 vdd.n8237 0.697868
R13517 vdd.n8426 vdd.n8379 0.697868
R13518 vdd.n8520 vdd.n8473 0.697868
R13519 vdd.n8707 vdd.n8660 0.697868
R13520 vdd.n8801 vdd.n8754 0.697868
R13521 vdd.n8990 vdd.n8943 0.697868
R13522 vdd.n9084 vdd.n9037 0.697868
R13523 vdd.n9225 vdd.n9178 0.697868
R13524 vdd.n9319 vdd.n9272 0.697868
R13525 vdd.n9461 vdd.n9414 0.697868
R13526 vdd.n9555 vdd.n9508 0.697868
R13527 vdd.n4658 vdd.n4611 0.697868
R13528 vdd.n4752 vdd.n4705 0.697868
R13529 vdd.n4941 vdd.n4894 0.697868
R13530 vdd.n5035 vdd.n4988 0.697868
R13531 vdd.n5176 vdd.n5129 0.697868
R13532 vdd.n5270 vdd.n5223 0.697868
R13533 vdd.n5412 vdd.n5365 0.697868
R13534 vdd.n5506 vdd.n5459 0.697868
R13535 vdd.n5693 vdd.n5646 0.697868
R13536 vdd.n5787 vdd.n5740 0.697868
R13537 vdd.n5976 vdd.n5929 0.697868
R13538 vdd.n6070 vdd.n6023 0.697868
R13539 vdd.n6211 vdd.n6164 0.697868
R13540 vdd.n6305 vdd.n6258 0.697868
R13541 vdd.n6447 vdd.n6400 0.697868
R13542 vdd.n6541 vdd.n6494 0.697868
R13543 vdd.n1644 vdd.n1597 0.697868
R13544 vdd.n1738 vdd.n1691 0.697868
R13545 vdd.n1927 vdd.n1880 0.697868
R13546 vdd.n2021 vdd.n1974 0.697868
R13547 vdd.n2162 vdd.n2115 0.697868
R13548 vdd.n2256 vdd.n2209 0.697868
R13549 vdd.n2398 vdd.n2351 0.697868
R13550 vdd.n2492 vdd.n2445 0.697868
R13551 vdd.n2679 vdd.n2632 0.697868
R13552 vdd.n2773 vdd.n2726 0.697868
R13553 vdd.n2962 vdd.n2915 0.697868
R13554 vdd.n3056 vdd.n3009 0.697868
R13555 vdd.n3197 vdd.n3150 0.697868
R13556 vdd.n3291 vdd.n3244 0.697868
R13557 vdd.n3433 vdd.n3386 0.697868
R13558 vdd.n3527 vdd.n3480 0.697868
R13559 vdd.n10122 vdd.n92 0.697868
R13560 vdd.n10216 vdd.n10169 0.697868
R13561 vdd.n10405 vdd.n10358 0.697868
R13562 vdd.n10499 vdd.n10452 0.697868
R13563 vdd.n10640 vdd.n10593 0.697868
R13564 vdd.n10734 vdd.n10687 0.697868
R13565 vdd.n10876 vdd.n10829 0.697868
R13566 vdd.n10970 vdd.n10923 0.697868
R13567 vdd.n11112 vdd.n11065 0.697868
R13568 vdd.n11206 vdd.n11159 0.697868
R13569 vdd.n11395 vdd.n11348 0.697868
R13570 vdd.n11489 vdd.n11442 0.697868
R13571 vdd.n11630 vdd.n11583 0.697868
R13572 vdd.n11724 vdd.n11677 0.697868
R13573 vdd.n11866 vdd.n11819 0.697868
R13574 vdd.n11960 vdd.n11913 0.697868
R13575 vdd.n7767 vdd.n7486 0.628061
R13576 vdd.n8285 vdd.n7251 0.628061
R13577 vdd.n8802 vdd.n7062 0.628061
R13578 vdd.n9320 vdd.n6826 0.628061
R13579 vdd.n4753 vdd.n4472 0.628061
R13580 vdd.n5271 vdd.n4237 0.628061
R13581 vdd.n5788 vdd.n4048 0.628061
R13582 vdd.n6306 vdd.n3812 0.628061
R13583 vdd.n1739 vdd.n1458 0.628061
R13584 vdd.n2257 vdd.n1223 0.628061
R13585 vdd.n2774 vdd.n1034 0.628061
R13586 vdd.n3292 vdd.n798 0.628061
R13587 vdd.n10217 vdd.n10029 0.628061
R13588 vdd.n10735 vdd.n9793 0.628061
R13589 vdd.n11207 vdd.n470 0.628061
R13590 vdd.n11725 vdd.n235 0.628061
R13591 vdd.n7625 vdd.n6682 0.620566
R13592 vdd.n7719 vdd.n7673 0.620566
R13593 vdd.n7908 vdd.n7768 0.620566
R13594 vdd.n8002 vdd.n7956 0.620566
R13595 vdd.n8143 vdd.n8050 0.620566
R13596 vdd.n8237 vdd.n8191 0.620566
R13597 vdd.n8379 vdd.n8286 0.620566
R13598 vdd.n8473 vdd.n8427 0.620566
R13599 vdd.n8660 vdd.n8567 0.620566
R13600 vdd.n8754 vdd.n8708 0.620566
R13601 vdd.n8943 vdd.n8803 0.620566
R13602 vdd.n9037 vdd.n8991 0.620566
R13603 vdd.n9178 vdd.n9085 0.620566
R13604 vdd.n9272 vdd.n9226 0.620566
R13605 vdd.n9414 vdd.n9321 0.620566
R13606 vdd.n9508 vdd.n9462 0.620566
R13607 vdd.n4611 vdd.n3668 0.620566
R13608 vdd.n4705 vdd.n4659 0.620566
R13609 vdd.n4894 vdd.n4754 0.620566
R13610 vdd.n4988 vdd.n4942 0.620566
R13611 vdd.n5129 vdd.n5036 0.620566
R13612 vdd.n5223 vdd.n5177 0.620566
R13613 vdd.n5365 vdd.n5272 0.620566
R13614 vdd.n5459 vdd.n5413 0.620566
R13615 vdd.n5646 vdd.n5553 0.620566
R13616 vdd.n5740 vdd.n5694 0.620566
R13617 vdd.n5929 vdd.n5789 0.620566
R13618 vdd.n6023 vdd.n5977 0.620566
R13619 vdd.n6164 vdd.n6071 0.620566
R13620 vdd.n6258 vdd.n6212 0.620566
R13621 vdd.n6400 vdd.n6307 0.620566
R13622 vdd.n6494 vdd.n6448 0.620566
R13623 vdd.n1597 vdd.n654 0.620566
R13624 vdd.n1691 vdd.n1645 0.620566
R13625 vdd.n1880 vdd.n1740 0.620566
R13626 vdd.n1974 vdd.n1928 0.620566
R13627 vdd.n2115 vdd.n2022 0.620566
R13628 vdd.n2209 vdd.n2163 0.620566
R13629 vdd.n2351 vdd.n2258 0.620566
R13630 vdd.n2445 vdd.n2399 0.620566
R13631 vdd.n2632 vdd.n2539 0.620566
R13632 vdd.n2726 vdd.n2680 0.620566
R13633 vdd.n2915 vdd.n2775 0.620566
R13634 vdd.n3009 vdd.n2963 0.620566
R13635 vdd.n3150 vdd.n3057 0.620566
R13636 vdd.n3244 vdd.n3198 0.620566
R13637 vdd.n3386 vdd.n3293 0.620566
R13638 vdd.n3480 vdd.n3434 0.620566
R13639 vdd.n11961 vdd.n92 0.620566
R13640 vdd.n10169 vdd.n10123 0.620566
R13641 vdd.n10358 vdd.n10218 0.620566
R13642 vdd.n10452 vdd.n10406 0.620566
R13643 vdd.n10593 vdd.n10500 0.620566
R13644 vdd.n10687 vdd.n10641 0.620566
R13645 vdd.n10829 vdd.n10736 0.620566
R13646 vdd.n10923 vdd.n10877 0.620566
R13647 vdd.n11065 vdd.n10972 0.620566
R13648 vdd.n11159 vdd.n11113 0.620566
R13649 vdd.n11348 vdd.n11208 0.620566
R13650 vdd.n11442 vdd.n11396 0.620566
R13651 vdd.n11583 vdd.n11490 0.620566
R13652 vdd.n11677 vdd.n11631 0.620566
R13653 vdd.n11819 vdd.n11726 0.620566
R13654 vdd.n11913 vdd.n11867 0.620566
R13655 vdd.n7904 vdd.n7857 0.616454
R13656 vdd.n8896 vdd.n8895 0.616454
R13657 vdd.n4890 vdd.n4843 0.616454
R13658 vdd.n5882 vdd.n5881 0.616454
R13659 vdd.n1876 vdd.n1829 0.616454
R13660 vdd.n2868 vdd.n2867 0.616454
R13661 vdd.n10311 vdd.n10310 0.616454
R13662 vdd.n11344 vdd.n11297 0.616454
R13663 vdd.n7768 vdd.n7767 0.594253
R13664 vdd.n8286 vdd.n8285 0.594253
R13665 vdd.n8803 vdd.n8802 0.594253
R13666 vdd.n9321 vdd.n9320 0.594253
R13667 vdd.n4754 vdd.n4753 0.594253
R13668 vdd.n5272 vdd.n5271 0.594253
R13669 vdd.n5789 vdd.n5788 0.594253
R13670 vdd.n6307 vdd.n6306 0.594253
R13671 vdd.n1740 vdd.n1739 0.594253
R13672 vdd.n2258 vdd.n2257 0.594253
R13673 vdd.n2775 vdd.n2774 0.594253
R13674 vdd.n3293 vdd.n3292 0.594253
R13675 vdd.n10218 vdd.n10217 0.594253
R13676 vdd.n10736 vdd.n10735 0.594253
R13677 vdd.n11208 vdd.n11207 0.594253
R13678 vdd.n11726 vdd.n11725 0.594253
R13679 vdd.n6637 vdd.n6636 0.309711
R13680 vdd.n7577 vdd.n7576 0.309711
R13681 vdd.n7624 vdd.n7623 0.309711
R13682 vdd.n7627 vdd.n7626 0.309711
R13683 vdd.n7488 vdd.n7487 0.309711
R13684 vdd.n7718 vdd.n7717 0.309711
R13685 vdd.n7721 vdd.n7720 0.309711
R13686 vdd.n7445 vdd.n7437 0.309711
R13687 vdd.n7391 vdd.n7390 0.309711
R13688 vdd.n7859 vdd.n7858 0.309711
R13689 vdd.n7813 vdd.n7812 0.309711
R13690 vdd.n7907 vdd.n7906 0.309711
R13691 vdd.n7910 vdd.n7909 0.309711
R13692 vdd.n7345 vdd.n7344 0.309711
R13693 vdd.n8001 vdd.n8000 0.309711
R13694 vdd.n8004 vdd.n8003 0.309711
R13695 vdd.n7299 vdd.n7298 0.309711
R13696 vdd.n8095 vdd.n8094 0.309711
R13697 vdd.n8142 vdd.n8141 0.309711
R13698 vdd.n8145 vdd.n8144 0.309711
R13699 vdd.n7253 vdd.n7252 0.309711
R13700 vdd.n8236 vdd.n8235 0.309711
R13701 vdd.n8239 vdd.n8238 0.309711
R13702 vdd.n7210 vdd.n7202 0.309711
R13703 vdd.n7156 vdd.n7155 0.309711
R13704 vdd.n8331 vdd.n8330 0.309711
R13705 vdd.n8378 vdd.n8377 0.309711
R13706 vdd.n8381 vdd.n8380 0.309711
R13707 vdd.n7110 vdd.n7109 0.309711
R13708 vdd.n8472 vdd.n8471 0.309711
R13709 vdd.n8475 vdd.n8474 0.309711
R13710 vdd.n8565 vdd.n8564 0.309711
R13711 vdd.n8612 vdd.n8611 0.309711
R13712 vdd.n8659 vdd.n8658 0.309711
R13713 vdd.n8705 vdd.n8704 0.309711
R13714 vdd.n7107 vdd.n7106 0.309711
R13715 vdd.n8753 vdd.n8752 0.309711
R13716 vdd.n8799 vdd.n8798 0.309711
R13717 vdd.n7045 vdd.n7012 0.309711
R13718 vdd.n7009 vdd.n7008 0.309711
R13719 vdd.n8848 vdd.n8847 0.309711
R13720 vdd.n8894 vdd.n8893 0.309711
R13721 vdd.n8942 vdd.n8941 0.309711
R13722 vdd.n8988 vdd.n8987 0.309711
R13723 vdd.n6963 vdd.n6962 0.309711
R13724 vdd.n9036 vdd.n9035 0.309711
R13725 vdd.n9082 vdd.n9081 0.309711
R13726 vdd.n6917 vdd.n6916 0.309711
R13727 vdd.n9130 vdd.n9129 0.309711
R13728 vdd.n9177 vdd.n9176 0.309711
R13729 vdd.n9223 vdd.n9222 0.309711
R13730 vdd.n6871 vdd.n6870 0.309711
R13731 vdd.n9271 vdd.n9270 0.309711
R13732 vdd.n9317 vdd.n9316 0.309711
R13733 vdd.n6809 vdd.n6776 0.309711
R13734 vdd.n6773 vdd.n6772 0.309711
R13735 vdd.n9366 vdd.n9365 0.309711
R13736 vdd.n9413 vdd.n9412 0.309711
R13737 vdd.n9459 vdd.n9458 0.309711
R13738 vdd.n6727 vdd.n6726 0.309711
R13739 vdd.n9507 vdd.n9506 0.309711
R13740 vdd.n9553 vdd.n9552 0.309711
R13741 vdd.n3623 vdd.n3622 0.309711
R13742 vdd.n4563 vdd.n4562 0.309711
R13743 vdd.n4610 vdd.n4609 0.309711
R13744 vdd.n4613 vdd.n4612 0.309711
R13745 vdd.n4474 vdd.n4473 0.309711
R13746 vdd.n4704 vdd.n4703 0.309711
R13747 vdd.n4707 vdd.n4706 0.309711
R13748 vdd.n4431 vdd.n4423 0.309711
R13749 vdd.n4377 vdd.n4376 0.309711
R13750 vdd.n4845 vdd.n4844 0.309711
R13751 vdd.n4799 vdd.n4798 0.309711
R13752 vdd.n4893 vdd.n4892 0.309711
R13753 vdd.n4896 vdd.n4895 0.309711
R13754 vdd.n4331 vdd.n4330 0.309711
R13755 vdd.n4987 vdd.n4986 0.309711
R13756 vdd.n4990 vdd.n4989 0.309711
R13757 vdd.n4285 vdd.n4284 0.309711
R13758 vdd.n5081 vdd.n5080 0.309711
R13759 vdd.n5128 vdd.n5127 0.309711
R13760 vdd.n5131 vdd.n5130 0.309711
R13761 vdd.n4239 vdd.n4238 0.309711
R13762 vdd.n5222 vdd.n5221 0.309711
R13763 vdd.n5225 vdd.n5224 0.309711
R13764 vdd.n4196 vdd.n4188 0.309711
R13765 vdd.n4142 vdd.n4141 0.309711
R13766 vdd.n5317 vdd.n5316 0.309711
R13767 vdd.n5364 vdd.n5363 0.309711
R13768 vdd.n5367 vdd.n5366 0.309711
R13769 vdd.n4096 vdd.n4095 0.309711
R13770 vdd.n5458 vdd.n5457 0.309711
R13771 vdd.n5461 vdd.n5460 0.309711
R13772 vdd.n5551 vdd.n5550 0.309711
R13773 vdd.n5598 vdd.n5597 0.309711
R13774 vdd.n5645 vdd.n5644 0.309711
R13775 vdd.n5691 vdd.n5690 0.309711
R13776 vdd.n4093 vdd.n4092 0.309711
R13777 vdd.n5739 vdd.n5738 0.309711
R13778 vdd.n5785 vdd.n5784 0.309711
R13779 vdd.n4031 vdd.n3998 0.309711
R13780 vdd.n3995 vdd.n3994 0.309711
R13781 vdd.n5834 vdd.n5833 0.309711
R13782 vdd.n5880 vdd.n5879 0.309711
R13783 vdd.n5928 vdd.n5927 0.309711
R13784 vdd.n5974 vdd.n5973 0.309711
R13785 vdd.n3949 vdd.n3948 0.309711
R13786 vdd.n6022 vdd.n6021 0.309711
R13787 vdd.n6068 vdd.n6067 0.309711
R13788 vdd.n3903 vdd.n3902 0.309711
R13789 vdd.n6116 vdd.n6115 0.309711
R13790 vdd.n6163 vdd.n6162 0.309711
R13791 vdd.n6209 vdd.n6208 0.309711
R13792 vdd.n3857 vdd.n3856 0.309711
R13793 vdd.n6257 vdd.n6256 0.309711
R13794 vdd.n6303 vdd.n6302 0.309711
R13795 vdd.n3795 vdd.n3762 0.309711
R13796 vdd.n3759 vdd.n3758 0.309711
R13797 vdd.n6352 vdd.n6351 0.309711
R13798 vdd.n6399 vdd.n6398 0.309711
R13799 vdd.n6445 vdd.n6444 0.309711
R13800 vdd.n3713 vdd.n3712 0.309711
R13801 vdd.n6493 vdd.n6492 0.309711
R13802 vdd.n6539 vdd.n6538 0.309711
R13803 vdd.n609 vdd.n608 0.309711
R13804 vdd.n1549 vdd.n1548 0.309711
R13805 vdd.n1596 vdd.n1595 0.309711
R13806 vdd.n1599 vdd.n1598 0.309711
R13807 vdd.n1460 vdd.n1459 0.309711
R13808 vdd.n1690 vdd.n1689 0.309711
R13809 vdd.n1693 vdd.n1692 0.309711
R13810 vdd.n1417 vdd.n1409 0.309711
R13811 vdd.n1363 vdd.n1362 0.309711
R13812 vdd.n1831 vdd.n1830 0.309711
R13813 vdd.n1785 vdd.n1784 0.309711
R13814 vdd.n1879 vdd.n1878 0.309711
R13815 vdd.n1882 vdd.n1881 0.309711
R13816 vdd.n1317 vdd.n1316 0.309711
R13817 vdd.n1973 vdd.n1972 0.309711
R13818 vdd.n1976 vdd.n1975 0.309711
R13819 vdd.n1271 vdd.n1270 0.309711
R13820 vdd.n2067 vdd.n2066 0.309711
R13821 vdd.n2114 vdd.n2113 0.309711
R13822 vdd.n2117 vdd.n2116 0.309711
R13823 vdd.n1225 vdd.n1224 0.309711
R13824 vdd.n2208 vdd.n2207 0.309711
R13825 vdd.n2211 vdd.n2210 0.309711
R13826 vdd.n1182 vdd.n1174 0.309711
R13827 vdd.n1128 vdd.n1127 0.309711
R13828 vdd.n2303 vdd.n2302 0.309711
R13829 vdd.n2350 vdd.n2349 0.309711
R13830 vdd.n2353 vdd.n2352 0.309711
R13831 vdd.n1082 vdd.n1081 0.309711
R13832 vdd.n2444 vdd.n2443 0.309711
R13833 vdd.n2447 vdd.n2446 0.309711
R13834 vdd.n2537 vdd.n2536 0.309711
R13835 vdd.n2584 vdd.n2583 0.309711
R13836 vdd.n2631 vdd.n2630 0.309711
R13837 vdd.n2677 vdd.n2676 0.309711
R13838 vdd.n1079 vdd.n1078 0.309711
R13839 vdd.n2725 vdd.n2724 0.309711
R13840 vdd.n2771 vdd.n2770 0.309711
R13841 vdd.n1017 vdd.n984 0.309711
R13842 vdd.n981 vdd.n980 0.309711
R13843 vdd.n2820 vdd.n2819 0.309711
R13844 vdd.n2866 vdd.n2865 0.309711
R13845 vdd.n2914 vdd.n2913 0.309711
R13846 vdd.n2960 vdd.n2959 0.309711
R13847 vdd.n935 vdd.n934 0.309711
R13848 vdd.n3008 vdd.n3007 0.309711
R13849 vdd.n3054 vdd.n3053 0.309711
R13850 vdd.n889 vdd.n888 0.309711
R13851 vdd.n3102 vdd.n3101 0.309711
R13852 vdd.n3149 vdd.n3148 0.309711
R13853 vdd.n3195 vdd.n3194 0.309711
R13854 vdd.n843 vdd.n842 0.309711
R13855 vdd.n3243 vdd.n3242 0.309711
R13856 vdd.n3289 vdd.n3288 0.309711
R13857 vdd.n781 vdd.n748 0.309711
R13858 vdd.n745 vdd.n744 0.309711
R13859 vdd.n3338 vdd.n3337 0.309711
R13860 vdd.n3385 vdd.n3384 0.309711
R13861 vdd.n3431 vdd.n3430 0.309711
R13862 vdd.n699 vdd.n698 0.309711
R13863 vdd.n3479 vdd.n3478 0.309711
R13864 vdd.n3525 vdd.n3524 0.309711
R13865 vdd.n607 vdd.n606 0.309711
R13866 vdd.n3575 vdd.n3574 0.309711
R13867 vdd.n3621 vdd.n3620 0.309711
R13868 vdd.n6589 vdd.n6588 0.309711
R13869 vdd.n6635 vdd.n6634 0.309711
R13870 vdd.n9603 vdd.n9602 0.309711
R13871 vdd.n9649 vdd.n9648 0.309711
R13872 vdd.n44 vdd.n43 0.309711
R13873 vdd.n91 vdd.n90 0.309711
R13874 vdd.n10120 vdd.n10119 0.309711
R13875 vdd.n10074 vdd.n10073 0.309711
R13876 vdd.n10168 vdd.n10167 0.309711
R13877 vdd.n10214 vdd.n10213 0.309711
R13878 vdd.n10012 vdd.n9979 0.309711
R13879 vdd.n9976 vdd.n9975 0.309711
R13880 vdd.n10263 vdd.n10262 0.309711
R13881 vdd.n10309 vdd.n10308 0.309711
R13882 vdd.n10357 vdd.n10356 0.309711
R13883 vdd.n10403 vdd.n10402 0.309711
R13884 vdd.n9930 vdd.n9929 0.309711
R13885 vdd.n10451 vdd.n10450 0.309711
R13886 vdd.n10497 vdd.n10496 0.309711
R13887 vdd.n9884 vdd.n9883 0.309711
R13888 vdd.n10545 vdd.n10544 0.309711
R13889 vdd.n10592 vdd.n10591 0.309711
R13890 vdd.n10638 vdd.n10637 0.309711
R13891 vdd.n9838 vdd.n9837 0.309711
R13892 vdd.n10686 vdd.n10685 0.309711
R13893 vdd.n10732 vdd.n10731 0.309711
R13894 vdd.n9776 vdd.n9743 0.309711
R13895 vdd.n9740 vdd.n9739 0.309711
R13896 vdd.n10781 vdd.n10780 0.309711
R13897 vdd.n10828 vdd.n10827 0.309711
R13898 vdd.n10874 vdd.n10873 0.309711
R13899 vdd.n9694 vdd.n9693 0.309711
R13900 vdd.n10922 vdd.n10921 0.309711
R13901 vdd.n10968 vdd.n10967 0.309711
R13902 vdd.n518 vdd.n517 0.309711
R13903 vdd.n11017 vdd.n11016 0.309711
R13904 vdd.n11064 vdd.n11063 0.309711
R13905 vdd.n11067 vdd.n11066 0.309711
R13906 vdd.n472 vdd.n471 0.309711
R13907 vdd.n11158 vdd.n11157 0.309711
R13908 vdd.n11161 vdd.n11160 0.309711
R13909 vdd.n429 vdd.n421 0.309711
R13910 vdd.n375 vdd.n374 0.309711
R13911 vdd.n11299 vdd.n11298 0.309711
R13912 vdd.n11253 vdd.n11252 0.309711
R13913 vdd.n11347 vdd.n11346 0.309711
R13914 vdd.n11350 vdd.n11349 0.309711
R13915 vdd.n329 vdd.n328 0.309711
R13916 vdd.n11441 vdd.n11440 0.309711
R13917 vdd.n11444 vdd.n11443 0.309711
R13918 vdd.n283 vdd.n282 0.309711
R13919 vdd.n11535 vdd.n11534 0.309711
R13920 vdd.n11582 vdd.n11581 0.309711
R13921 vdd.n11585 vdd.n11584 0.309711
R13922 vdd.n237 vdd.n236 0.309711
R13923 vdd.n11676 vdd.n11675 0.309711
R13924 vdd.n11679 vdd.n11678 0.309711
R13925 vdd.n194 vdd.n186 0.309711
R13926 vdd.n140 vdd.n139 0.309711
R13927 vdd.n11771 vdd.n11770 0.309711
R13928 vdd.n11818 vdd.n11817 0.309711
R13929 vdd.n11821 vdd.n11820 0.309711
R13930 vdd.n94 vdd.n93 0.309711
R13931 vdd.n11912 vdd.n11911 0.309711
R13932 vdd.n11915 vdd.n11914 0.309711
R13933 vdd.n12006 vdd.n12005 0.309711
R13934 vdd.n7476 vdd.n7445 0.279783
R13935 vdd.n7241 vdd.n7210 0.279783
R13936 vdd.n7046 vdd.n7045 0.279783
R13937 vdd.n6810 vdd.n6809 0.279783
R13938 vdd.n4462 vdd.n4431 0.279783
R13939 vdd.n4227 vdd.n4196 0.279783
R13940 vdd.n4032 vdd.n4031 0.279783
R13941 vdd.n3796 vdd.n3795 0.279783
R13942 vdd.n1448 vdd.n1417 0.279783
R13943 vdd.n1213 vdd.n1182 0.279783
R13944 vdd.n1018 vdd.n1017 0.279783
R13945 vdd.n782 vdd.n781 0.279783
R13946 vdd.n10013 vdd.n10012 0.279783
R13947 vdd.n9777 vdd.n9776 0.279783
R13948 vdd.n460 vdd.n429 0.279783
R13949 vdd.n225 vdd.n194 0.279783
R13950 vdd.n7717 vdd.n7716 0.279284
R13951 vdd.n8000 vdd.n7999 0.279284
R13952 vdd.n8235 vdd.n8234 0.279284
R13953 vdd.n8471 vdd.n8470 0.279284
R13954 vdd.n8752 vdd.n8751 0.279284
R13955 vdd.n9035 vdd.n9034 0.279284
R13956 vdd.n9270 vdd.n9269 0.279284
R13957 vdd.n9506 vdd.n9505 0.279284
R13958 vdd.n4703 vdd.n4702 0.279284
R13959 vdd.n4986 vdd.n4985 0.279284
R13960 vdd.n5221 vdd.n5220 0.279284
R13961 vdd.n5457 vdd.n5456 0.279284
R13962 vdd.n5738 vdd.n5737 0.279284
R13963 vdd.n6021 vdd.n6020 0.279284
R13964 vdd.n6256 vdd.n6255 0.279284
R13965 vdd.n6492 vdd.n6491 0.279284
R13966 vdd.n1689 vdd.n1688 0.279284
R13967 vdd.n1972 vdd.n1971 0.279284
R13968 vdd.n2207 vdd.n2206 0.279284
R13969 vdd.n2443 vdd.n2442 0.279284
R13970 vdd.n2724 vdd.n2723 0.279284
R13971 vdd.n3007 vdd.n3006 0.279284
R13972 vdd.n3242 vdd.n3241 0.279284
R13973 vdd.n3478 vdd.n3477 0.279284
R13974 vdd.n606 vdd.n605 0.279284
R13975 vdd.n10167 vdd.n10166 0.279284
R13976 vdd.n10450 vdd.n10449 0.279284
R13977 vdd.n10685 vdd.n10684 0.279284
R13978 vdd.n10921 vdd.n10920 0.279284
R13979 vdd.n11157 vdd.n11156 0.279284
R13980 vdd.n11440 vdd.n11439 0.279284
R13981 vdd.n11675 vdd.n11674 0.279284
R13982 vdd.n11911 vdd.n11910 0.279284
R13983 vdd.n6681 vdd.n6637 0.279283
R13984 vdd.n7621 vdd.n7577 0.279283
R13985 vdd.n7623 vdd.n7622 0.279283
R13986 vdd.n7671 vdd.n7627 0.279283
R13987 vdd.n7532 vdd.n7488 0.279283
R13988 vdd.n7765 vdd.n7721 0.279283
R13989 vdd.n7435 vdd.n7391 0.279283
R13990 vdd.n7903 vdd.n7859 0.279283
R13991 vdd.n7857 vdd.n7813 0.279283
R13992 vdd.n7906 vdd.n7905 0.279283
R13993 vdd.n7954 vdd.n7910 0.279283
R13994 vdd.n7389 vdd.n7345 0.279283
R13995 vdd.n8048 vdd.n8004 0.279283
R13996 vdd.n7343 vdd.n7299 0.279283
R13997 vdd.n8139 vdd.n8095 0.279283
R13998 vdd.n8141 vdd.n8140 0.279283
R13999 vdd.n8189 vdd.n8145 0.279283
R14000 vdd.n7297 vdd.n7253 0.279283
R14001 vdd.n8283 vdd.n8239 0.279283
R14002 vdd.n7200 vdd.n7156 0.279283
R14003 vdd.n8375 vdd.n8331 0.279283
R14004 vdd.n8377 vdd.n8376 0.279283
R14005 vdd.n8425 vdd.n8381 0.279283
R14006 vdd.n7154 vdd.n7110 0.279283
R14007 vdd.n8519 vdd.n8475 0.279283
R14008 vdd.n8566 vdd.n8565 0.279283
R14009 vdd.n8613 vdd.n8612 0.279283
R14010 vdd.n8658 vdd.n8657 0.279283
R14011 vdd.n8706 vdd.n8705 0.279283
R14012 vdd.n7108 vdd.n7107 0.279283
R14013 vdd.n8800 vdd.n8799 0.279283
R14014 vdd.n7010 vdd.n7009 0.279283
R14015 vdd.n8849 vdd.n8848 0.279283
R14016 vdd.n8895 vdd.n8894 0.279283
R14017 vdd.n8941 vdd.n8940 0.279283
R14018 vdd.n8989 vdd.n8988 0.279283
R14019 vdd.n6964 vdd.n6963 0.279283
R14020 vdd.n9083 vdd.n9082 0.279283
R14021 vdd.n6918 vdd.n6917 0.279283
R14022 vdd.n9131 vdd.n9130 0.279283
R14023 vdd.n9176 vdd.n9175 0.279283
R14024 vdd.n9224 vdd.n9223 0.279283
R14025 vdd.n6872 vdd.n6871 0.279283
R14026 vdd.n9318 vdd.n9317 0.279283
R14027 vdd.n6774 vdd.n6773 0.279283
R14028 vdd.n9367 vdd.n9366 0.279283
R14029 vdd.n9412 vdd.n9411 0.279283
R14030 vdd.n9460 vdd.n9459 0.279283
R14031 vdd.n6728 vdd.n6727 0.279283
R14032 vdd.n9554 vdd.n9553 0.279283
R14033 vdd.n3667 vdd.n3623 0.279283
R14034 vdd.n4607 vdd.n4563 0.279283
R14035 vdd.n4609 vdd.n4608 0.279283
R14036 vdd.n4657 vdd.n4613 0.279283
R14037 vdd.n4518 vdd.n4474 0.279283
R14038 vdd.n4751 vdd.n4707 0.279283
R14039 vdd.n4421 vdd.n4377 0.279283
R14040 vdd.n4889 vdd.n4845 0.279283
R14041 vdd.n4843 vdd.n4799 0.279283
R14042 vdd.n4892 vdd.n4891 0.279283
R14043 vdd.n4940 vdd.n4896 0.279283
R14044 vdd.n4375 vdd.n4331 0.279283
R14045 vdd.n5034 vdd.n4990 0.279283
R14046 vdd.n4329 vdd.n4285 0.279283
R14047 vdd.n5125 vdd.n5081 0.279283
R14048 vdd.n5127 vdd.n5126 0.279283
R14049 vdd.n5175 vdd.n5131 0.279283
R14050 vdd.n4283 vdd.n4239 0.279283
R14051 vdd.n5269 vdd.n5225 0.279283
R14052 vdd.n4186 vdd.n4142 0.279283
R14053 vdd.n5361 vdd.n5317 0.279283
R14054 vdd.n5363 vdd.n5362 0.279283
R14055 vdd.n5411 vdd.n5367 0.279283
R14056 vdd.n4140 vdd.n4096 0.279283
R14057 vdd.n5505 vdd.n5461 0.279283
R14058 vdd.n5552 vdd.n5551 0.279283
R14059 vdd.n5599 vdd.n5598 0.279283
R14060 vdd.n5644 vdd.n5643 0.279283
R14061 vdd.n5692 vdd.n5691 0.279283
R14062 vdd.n4094 vdd.n4093 0.279283
R14063 vdd.n5786 vdd.n5785 0.279283
R14064 vdd.n3996 vdd.n3995 0.279283
R14065 vdd.n5835 vdd.n5834 0.279283
R14066 vdd.n5881 vdd.n5880 0.279283
R14067 vdd.n5927 vdd.n5926 0.279283
R14068 vdd.n5975 vdd.n5974 0.279283
R14069 vdd.n3950 vdd.n3949 0.279283
R14070 vdd.n6069 vdd.n6068 0.279283
R14071 vdd.n3904 vdd.n3903 0.279283
R14072 vdd.n6117 vdd.n6116 0.279283
R14073 vdd.n6162 vdd.n6161 0.279283
R14074 vdd.n6210 vdd.n6209 0.279283
R14075 vdd.n3858 vdd.n3857 0.279283
R14076 vdd.n6304 vdd.n6303 0.279283
R14077 vdd.n3760 vdd.n3759 0.279283
R14078 vdd.n6353 vdd.n6352 0.279283
R14079 vdd.n6398 vdd.n6397 0.279283
R14080 vdd.n6446 vdd.n6445 0.279283
R14081 vdd.n3714 vdd.n3713 0.279283
R14082 vdd.n6540 vdd.n6539 0.279283
R14083 vdd.n653 vdd.n609 0.279283
R14084 vdd.n1593 vdd.n1549 0.279283
R14085 vdd.n1595 vdd.n1594 0.279283
R14086 vdd.n1643 vdd.n1599 0.279283
R14087 vdd.n1504 vdd.n1460 0.279283
R14088 vdd.n1737 vdd.n1693 0.279283
R14089 vdd.n1407 vdd.n1363 0.279283
R14090 vdd.n1875 vdd.n1831 0.279283
R14091 vdd.n1829 vdd.n1785 0.279283
R14092 vdd.n1878 vdd.n1877 0.279283
R14093 vdd.n1926 vdd.n1882 0.279283
R14094 vdd.n1361 vdd.n1317 0.279283
R14095 vdd.n2020 vdd.n1976 0.279283
R14096 vdd.n1315 vdd.n1271 0.279283
R14097 vdd.n2111 vdd.n2067 0.279283
R14098 vdd.n2113 vdd.n2112 0.279283
R14099 vdd.n2161 vdd.n2117 0.279283
R14100 vdd.n1269 vdd.n1225 0.279283
R14101 vdd.n2255 vdd.n2211 0.279283
R14102 vdd.n1172 vdd.n1128 0.279283
R14103 vdd.n2347 vdd.n2303 0.279283
R14104 vdd.n2349 vdd.n2348 0.279283
R14105 vdd.n2397 vdd.n2353 0.279283
R14106 vdd.n1126 vdd.n1082 0.279283
R14107 vdd.n2491 vdd.n2447 0.279283
R14108 vdd.n2538 vdd.n2537 0.279283
R14109 vdd.n2585 vdd.n2584 0.279283
R14110 vdd.n2630 vdd.n2629 0.279283
R14111 vdd.n2678 vdd.n2677 0.279283
R14112 vdd.n1080 vdd.n1079 0.279283
R14113 vdd.n2772 vdd.n2771 0.279283
R14114 vdd.n982 vdd.n981 0.279283
R14115 vdd.n2821 vdd.n2820 0.279283
R14116 vdd.n2867 vdd.n2866 0.279283
R14117 vdd.n2913 vdd.n2912 0.279283
R14118 vdd.n2961 vdd.n2960 0.279283
R14119 vdd.n936 vdd.n935 0.279283
R14120 vdd.n3055 vdd.n3054 0.279283
R14121 vdd.n890 vdd.n889 0.279283
R14122 vdd.n3103 vdd.n3102 0.279283
R14123 vdd.n3148 vdd.n3147 0.279283
R14124 vdd.n3196 vdd.n3195 0.279283
R14125 vdd.n844 vdd.n843 0.279283
R14126 vdd.n3290 vdd.n3289 0.279283
R14127 vdd.n746 vdd.n745 0.279283
R14128 vdd.n3339 vdd.n3338 0.279283
R14129 vdd.n3384 vdd.n3383 0.279283
R14130 vdd.n3432 vdd.n3431 0.279283
R14131 vdd.n700 vdd.n699 0.279283
R14132 vdd.n3526 vdd.n3525 0.279283
R14133 vdd.n3574 vdd.n3573 0.279283
R14134 vdd.n3620 vdd.n3619 0.279283
R14135 vdd.n6588 vdd.n6587 0.279283
R14136 vdd.n6634 vdd.n6633 0.279283
R14137 vdd.n9602 vdd.n9601 0.279283
R14138 vdd.n9648 vdd.n9647 0.279283
R14139 vdd.n45 vdd.n44 0.279283
R14140 vdd.n90 vdd.n89 0.279283
R14141 vdd.n10121 vdd.n10120 0.279283
R14142 vdd.n10075 vdd.n10074 0.279283
R14143 vdd.n10215 vdd.n10214 0.279283
R14144 vdd.n9977 vdd.n9976 0.279283
R14145 vdd.n10264 vdd.n10263 0.279283
R14146 vdd.n10310 vdd.n10309 0.279283
R14147 vdd.n10356 vdd.n10355 0.279283
R14148 vdd.n10404 vdd.n10403 0.279283
R14149 vdd.n9931 vdd.n9930 0.279283
R14150 vdd.n10498 vdd.n10497 0.279283
R14151 vdd.n9885 vdd.n9884 0.279283
R14152 vdd.n10546 vdd.n10545 0.279283
R14153 vdd.n10591 vdd.n10590 0.279283
R14154 vdd.n10639 vdd.n10638 0.279283
R14155 vdd.n9839 vdd.n9838 0.279283
R14156 vdd.n10733 vdd.n10732 0.279283
R14157 vdd.n9741 vdd.n9740 0.279283
R14158 vdd.n10782 vdd.n10781 0.279283
R14159 vdd.n10827 vdd.n10826 0.279283
R14160 vdd.n10875 vdd.n10874 0.279283
R14161 vdd.n9695 vdd.n9694 0.279283
R14162 vdd.n10969 vdd.n10968 0.279283
R14163 vdd.n562 vdd.n518 0.279283
R14164 vdd.n11061 vdd.n11017 0.279283
R14165 vdd.n11063 vdd.n11062 0.279283
R14166 vdd.n11111 vdd.n11067 0.279283
R14167 vdd.n516 vdd.n472 0.279283
R14168 vdd.n11205 vdd.n11161 0.279283
R14169 vdd.n419 vdd.n375 0.279283
R14170 vdd.n11343 vdd.n11299 0.279283
R14171 vdd.n11297 vdd.n11253 0.279283
R14172 vdd.n11346 vdd.n11345 0.279283
R14173 vdd.n11394 vdd.n11350 0.279283
R14174 vdd.n373 vdd.n329 0.279283
R14175 vdd.n11488 vdd.n11444 0.279283
R14176 vdd.n327 vdd.n283 0.279283
R14177 vdd.n11579 vdd.n11535 0.279283
R14178 vdd.n11581 vdd.n11580 0.279283
R14179 vdd.n11629 vdd.n11585 0.279283
R14180 vdd.n281 vdd.n237 0.279283
R14181 vdd.n11723 vdd.n11679 0.279283
R14182 vdd.n184 vdd.n140 0.279283
R14183 vdd.n11815 vdd.n11771 0.279283
R14184 vdd.n11817 vdd.n11816 0.279283
R14185 vdd.n11865 vdd.n11821 0.279283
R14186 vdd.n138 vdd.n94 0.279283
R14187 vdd.n11959 vdd.n11915 0.279283
R14188 vdd.n12007 vdd.n12006 0.279283
R14189 vdd.n7625 vdd 0.276816
R14190 vdd.n7719 vdd 0.276816
R14191 vdd.n7908 vdd 0.276816
R14192 vdd.n8002 vdd 0.276816
R14193 vdd.n8143 vdd 0.276816
R14194 vdd.n8237 vdd 0.276816
R14195 vdd.n8379 vdd 0.276816
R14196 vdd.n8473 vdd 0.276816
R14197 vdd.n4611 vdd 0.276816
R14198 vdd.n4705 vdd 0.276816
R14199 vdd.n4894 vdd 0.276816
R14200 vdd.n4988 vdd 0.276816
R14201 vdd.n5129 vdd 0.276816
R14202 vdd.n5223 vdd 0.276816
R14203 vdd.n5365 vdd 0.276816
R14204 vdd.n5459 vdd 0.276816
R14205 vdd.n1597 vdd 0.276816
R14206 vdd.n1691 vdd 0.276816
R14207 vdd.n1880 vdd 0.276816
R14208 vdd.n1974 vdd 0.276816
R14209 vdd.n2115 vdd 0.276816
R14210 vdd.n2209 vdd 0.276816
R14211 vdd.n2351 vdd 0.276816
R14212 vdd.n2445 vdd 0.276816
R14213 vdd.n11065 vdd 0.276816
R14214 vdd.n11159 vdd 0.276816
R14215 vdd.n11348 vdd 0.276816
R14216 vdd.n11442 vdd 0.276816
R14217 vdd.n11583 vdd 0.276816
R14218 vdd.n11677 vdd 0.276816
R14219 vdd.n11819 vdd 0.276816
R14220 vdd.n11913 vdd 0.276816
R14221 vdd.n8660 vdd 0.243921
R14222 vdd.n8754 vdd 0.243921
R14223 vdd.n8943 vdd 0.243921
R14224 vdd.n9037 vdd 0.243921
R14225 vdd.n9178 vdd 0.243921
R14226 vdd.n9272 vdd 0.243921
R14227 vdd.n9414 vdd 0.243921
R14228 vdd.n9508 vdd 0.243921
R14229 vdd.n5646 vdd 0.243921
R14230 vdd.n5740 vdd 0.243921
R14231 vdd.n5929 vdd 0.243921
R14232 vdd.n6023 vdd 0.243921
R14233 vdd.n6164 vdd 0.243921
R14234 vdd.n6258 vdd 0.243921
R14235 vdd.n6400 vdd 0.243921
R14236 vdd.n6494 vdd 0.243921
R14237 vdd.n2632 vdd 0.243921
R14238 vdd.n2726 vdd 0.243921
R14239 vdd.n2915 vdd 0.243921
R14240 vdd.n3009 vdd 0.243921
R14241 vdd.n3150 vdd 0.243921
R14242 vdd.n3244 vdd 0.243921
R14243 vdd.n3386 vdd 0.243921
R14244 vdd.n3480 vdd 0.243921
R14245 vdd.n92 vdd 0.243921
R14246 vdd.n10169 vdd 0.243921
R14247 vdd.n10358 vdd 0.243921
R14248 vdd.n10452 vdd 0.243921
R14249 vdd.n10593 vdd 0.243921
R14250 vdd.n10687 vdd 0.243921
R14251 vdd.n10829 vdd 0.243921
R14252 vdd.n10923 vdd 0.243921
R14253 vdd.n8803 vdd 0.206092
R14254 vdd.n9321 vdd 0.206092
R14255 vdd.n5789 vdd 0.206092
R14256 vdd.n6307 vdd 0.206092
R14257 vdd.n2775 vdd 0.206092
R14258 vdd.n3293 vdd 0.206092
R14259 vdd.n10218 vdd 0.206092
R14260 vdd.n10736 vdd 0.206092
R14261 vdd.n8567 vdd 0.184711
R14262 vdd.n9085 vdd 0.184711
R14263 vdd.n5553 vdd 0.184711
R14264 vdd.n6071 vdd 0.184711
R14265 vdd.n2539 vdd 0.184711
R14266 vdd.n3057 vdd 0.184711
R14267 vdd.n10500 vdd 0.184711
R14268 vdd vdd.n11961 0.183066
R14269 vdd.n6682 vdd 0.140303
R14270 vdd.n7768 vdd 0.140303
R14271 vdd.n8050 vdd 0.140303
R14272 vdd.n8286 vdd 0.140303
R14273 vdd.n3668 vdd 0.140303
R14274 vdd.n4754 vdd 0.140303
R14275 vdd.n5036 vdd 0.140303
R14276 vdd.n5272 vdd 0.140303
R14277 vdd.n654 vdd 0.140303
R14278 vdd.n1740 vdd 0.140303
R14279 vdd.n2022 vdd 0.140303
R14280 vdd.n2258 vdd 0.140303
R14281 vdd.n10972 vdd 0.140303
R14282 vdd.n11208 vdd 0.140303
R14283 vdd.n11490 vdd 0.140303
R14284 vdd.n11726 vdd 0.140303
R14285 vdd.n8564 vdd 0.0745132
R14286 vdd.n8611 vdd 0.0745132
R14287 vdd vdd.n8659 0.0745132
R14288 vdd.n8704 vdd 0.0745132
R14289 vdd.n7106 vdd 0.0745132
R14290 vdd vdd.n8753 0.0745132
R14291 vdd.n8798 vdd 0.0745132
R14292 vdd.n7008 vdd 0.0745132
R14293 vdd.n8847 vdd 0.0745132
R14294 vdd.n8893 vdd 0.0745132
R14295 vdd vdd.n8942 0.0745132
R14296 vdd.n8987 vdd 0.0745132
R14297 vdd.n6962 vdd 0.0745132
R14298 vdd vdd.n9036 0.0745132
R14299 vdd.n9081 vdd 0.0745132
R14300 vdd.n6916 vdd 0.0745132
R14301 vdd.n9129 vdd 0.0745132
R14302 vdd vdd.n9177 0.0745132
R14303 vdd.n9222 vdd 0.0745132
R14304 vdd.n6870 vdd 0.0745132
R14305 vdd vdd.n9271 0.0745132
R14306 vdd.n9316 vdd 0.0745132
R14307 vdd.n6772 vdd 0.0745132
R14308 vdd.n9365 vdd 0.0745132
R14309 vdd vdd.n9413 0.0745132
R14310 vdd.n9458 vdd 0.0745132
R14311 vdd.n6726 vdd 0.0745132
R14312 vdd vdd.n9507 0.0745132
R14313 vdd.n9552 vdd 0.0745132
R14314 vdd.n5550 vdd 0.0745132
R14315 vdd.n5597 vdd 0.0745132
R14316 vdd vdd.n5645 0.0745132
R14317 vdd.n5690 vdd 0.0745132
R14318 vdd.n4092 vdd 0.0745132
R14319 vdd vdd.n5739 0.0745132
R14320 vdd.n5784 vdd 0.0745132
R14321 vdd.n3994 vdd 0.0745132
R14322 vdd.n5833 vdd 0.0745132
R14323 vdd.n5879 vdd 0.0745132
R14324 vdd vdd.n5928 0.0745132
R14325 vdd.n5973 vdd 0.0745132
R14326 vdd.n3948 vdd 0.0745132
R14327 vdd vdd.n6022 0.0745132
R14328 vdd.n6067 vdd 0.0745132
R14329 vdd.n3902 vdd 0.0745132
R14330 vdd.n6115 vdd 0.0745132
R14331 vdd vdd.n6163 0.0745132
R14332 vdd.n6208 vdd 0.0745132
R14333 vdd.n3856 vdd 0.0745132
R14334 vdd vdd.n6257 0.0745132
R14335 vdd.n6302 vdd 0.0745132
R14336 vdd.n3758 vdd 0.0745132
R14337 vdd.n6351 vdd 0.0745132
R14338 vdd vdd.n6399 0.0745132
R14339 vdd.n6444 vdd 0.0745132
R14340 vdd.n3712 vdd 0.0745132
R14341 vdd vdd.n6493 0.0745132
R14342 vdd.n6538 vdd 0.0745132
R14343 vdd.n2536 vdd 0.0745132
R14344 vdd.n2583 vdd 0.0745132
R14345 vdd vdd.n2631 0.0745132
R14346 vdd.n2676 vdd 0.0745132
R14347 vdd.n1078 vdd 0.0745132
R14348 vdd vdd.n2725 0.0745132
R14349 vdd.n2770 vdd 0.0745132
R14350 vdd.n980 vdd 0.0745132
R14351 vdd.n2819 vdd 0.0745132
R14352 vdd.n2865 vdd 0.0745132
R14353 vdd vdd.n2914 0.0745132
R14354 vdd.n2959 vdd 0.0745132
R14355 vdd.n934 vdd 0.0745132
R14356 vdd vdd.n3008 0.0745132
R14357 vdd.n3053 vdd 0.0745132
R14358 vdd.n888 vdd 0.0745132
R14359 vdd.n3101 vdd 0.0745132
R14360 vdd vdd.n3149 0.0745132
R14361 vdd.n3194 vdd 0.0745132
R14362 vdd.n842 vdd 0.0745132
R14363 vdd vdd.n3243 0.0745132
R14364 vdd.n3288 vdd 0.0745132
R14365 vdd.n744 vdd 0.0745132
R14366 vdd.n3337 vdd 0.0745132
R14367 vdd vdd.n3385 0.0745132
R14368 vdd.n3430 vdd 0.0745132
R14369 vdd.n698 vdd 0.0745132
R14370 vdd vdd.n3479 0.0745132
R14371 vdd.n3524 vdd 0.0745132
R14372 vdd vdd.n607 0.0745132
R14373 vdd vdd.n3575 0.0745132
R14374 vdd vdd.n3621 0.0745132
R14375 vdd vdd.n6589 0.0745132
R14376 vdd vdd.n6635 0.0745132
R14377 vdd vdd.n9603 0.0745132
R14378 vdd vdd.n9649 0.0745132
R14379 vdd.n43 vdd 0.0745132
R14380 vdd vdd.n91 0.0745132
R14381 vdd.n10119 vdd 0.0745132
R14382 vdd.n10073 vdd 0.0745132
R14383 vdd vdd.n10168 0.0745132
R14384 vdd.n10213 vdd 0.0745132
R14385 vdd.n9975 vdd 0.0745132
R14386 vdd.n10262 vdd 0.0745132
R14387 vdd.n10308 vdd 0.0745132
R14388 vdd vdd.n10357 0.0745132
R14389 vdd.n10402 vdd 0.0745132
R14390 vdd.n9929 vdd 0.0745132
R14391 vdd vdd.n10451 0.0745132
R14392 vdd.n10496 vdd 0.0745132
R14393 vdd.n9883 vdd 0.0745132
R14394 vdd.n10544 vdd 0.0745132
R14395 vdd vdd.n10592 0.0745132
R14396 vdd.n10637 vdd 0.0745132
R14397 vdd.n9837 vdd 0.0745132
R14398 vdd vdd.n10686 0.0745132
R14399 vdd.n10731 vdd 0.0745132
R14400 vdd.n9739 vdd 0.0745132
R14401 vdd.n10780 vdd 0.0745132
R14402 vdd vdd.n10828 0.0745132
R14403 vdd.n10873 vdd 0.0745132
R14404 vdd.n9693 vdd 0.0745132
R14405 vdd vdd.n10922 0.0745132
R14406 vdd.n10967 vdd 0.0745132
R14407 vdd.n12005 vdd 0.0745132
R14408 vdd.n7576 vdd 0.0416184
R14409 vdd vdd.n7624 0.0416184
R14410 vdd.n7626 vdd 0.0416184
R14411 vdd.n7487 vdd 0.0416184
R14412 vdd vdd.n7718 0.0416184
R14413 vdd.n7720 vdd 0.0416184
R14414 vdd.n7390 vdd 0.0416184
R14415 vdd.n7858 vdd 0.0416184
R14416 vdd.n7812 vdd 0.0416184
R14417 vdd vdd.n7907 0.0416184
R14418 vdd.n7909 vdd 0.0416184
R14419 vdd.n7344 vdd 0.0416184
R14420 vdd vdd.n8001 0.0416184
R14421 vdd.n8003 vdd 0.0416184
R14422 vdd.n7298 vdd 0.0416184
R14423 vdd.n8094 vdd 0.0416184
R14424 vdd vdd.n8142 0.0416184
R14425 vdd.n8144 vdd 0.0416184
R14426 vdd.n7252 vdd 0.0416184
R14427 vdd vdd.n8236 0.0416184
R14428 vdd.n8238 vdd 0.0416184
R14429 vdd.n7155 vdd 0.0416184
R14430 vdd.n8330 vdd 0.0416184
R14431 vdd vdd.n8378 0.0416184
R14432 vdd.n8380 vdd 0.0416184
R14433 vdd.n7109 vdd 0.0416184
R14434 vdd vdd.n8472 0.0416184
R14435 vdd.n8474 vdd 0.0416184
R14436 vdd.n4562 vdd 0.0416184
R14437 vdd vdd.n4610 0.0416184
R14438 vdd.n4612 vdd 0.0416184
R14439 vdd.n4473 vdd 0.0416184
R14440 vdd vdd.n4704 0.0416184
R14441 vdd.n4706 vdd 0.0416184
R14442 vdd.n4376 vdd 0.0416184
R14443 vdd.n4844 vdd 0.0416184
R14444 vdd.n4798 vdd 0.0416184
R14445 vdd vdd.n4893 0.0416184
R14446 vdd.n4895 vdd 0.0416184
R14447 vdd.n4330 vdd 0.0416184
R14448 vdd vdd.n4987 0.0416184
R14449 vdd.n4989 vdd 0.0416184
R14450 vdd.n4284 vdd 0.0416184
R14451 vdd.n5080 vdd 0.0416184
R14452 vdd vdd.n5128 0.0416184
R14453 vdd.n5130 vdd 0.0416184
R14454 vdd.n4238 vdd 0.0416184
R14455 vdd vdd.n5222 0.0416184
R14456 vdd.n5224 vdd 0.0416184
R14457 vdd.n4141 vdd 0.0416184
R14458 vdd.n5316 vdd 0.0416184
R14459 vdd vdd.n5364 0.0416184
R14460 vdd.n5366 vdd 0.0416184
R14461 vdd.n4095 vdd 0.0416184
R14462 vdd vdd.n5458 0.0416184
R14463 vdd.n5460 vdd 0.0416184
R14464 vdd.n1548 vdd 0.0416184
R14465 vdd vdd.n1596 0.0416184
R14466 vdd.n1598 vdd 0.0416184
R14467 vdd.n1459 vdd 0.0416184
R14468 vdd vdd.n1690 0.0416184
R14469 vdd.n1692 vdd 0.0416184
R14470 vdd.n1362 vdd 0.0416184
R14471 vdd.n1830 vdd 0.0416184
R14472 vdd.n1784 vdd 0.0416184
R14473 vdd vdd.n1879 0.0416184
R14474 vdd.n1881 vdd 0.0416184
R14475 vdd.n1316 vdd 0.0416184
R14476 vdd vdd.n1973 0.0416184
R14477 vdd.n1975 vdd 0.0416184
R14478 vdd.n1270 vdd 0.0416184
R14479 vdd.n2066 vdd 0.0416184
R14480 vdd vdd.n2114 0.0416184
R14481 vdd.n2116 vdd 0.0416184
R14482 vdd.n1224 vdd 0.0416184
R14483 vdd vdd.n2208 0.0416184
R14484 vdd.n2210 vdd 0.0416184
R14485 vdd.n1127 vdd 0.0416184
R14486 vdd.n2302 vdd 0.0416184
R14487 vdd vdd.n2350 0.0416184
R14488 vdd.n2352 vdd 0.0416184
R14489 vdd.n1081 vdd 0.0416184
R14490 vdd vdd.n2444 0.0416184
R14491 vdd.n2446 vdd 0.0416184
R14492 vdd.n11016 vdd 0.0416184
R14493 vdd vdd.n11064 0.0416184
R14494 vdd.n11066 vdd 0.0416184
R14495 vdd.n471 vdd 0.0416184
R14496 vdd vdd.n11158 0.0416184
R14497 vdd.n11160 vdd 0.0416184
R14498 vdd.n374 vdd 0.0416184
R14499 vdd.n11298 vdd 0.0416184
R14500 vdd.n11252 vdd 0.0416184
R14501 vdd vdd.n11347 0.0416184
R14502 vdd.n11349 vdd 0.0416184
R14503 vdd.n328 vdd 0.0416184
R14504 vdd vdd.n11441 0.0416184
R14505 vdd.n11443 vdd 0.0416184
R14506 vdd.n282 vdd 0.0416184
R14507 vdd.n11534 vdd 0.0416184
R14508 vdd vdd.n11582 0.0416184
R14509 vdd.n11584 vdd 0.0416184
R14510 vdd.n236 vdd 0.0416184
R14511 vdd vdd.n11676 0.0416184
R14512 vdd.n11678 vdd 0.0416184
R14513 vdd.n139 vdd 0.0416184
R14514 vdd.n11770 vdd 0.0416184
R14515 vdd vdd.n11818 0.0416184
R14516 vdd.n11820 vdd 0.0416184
R14517 vdd.n93 vdd 0.0416184
R14518 vdd vdd.n11912 0.0416184
R14519 vdd.n11914 vdd 0.0416184
R14520 vdd.n7486 vdd.n7436 0.02926
R14521 vdd.n7251 vdd.n7201 0.02926
R14522 vdd.n7062 vdd.n7011 0.02926
R14523 vdd.n6826 vdd.n6775 0.02926
R14524 vdd.n4472 vdd.n4422 0.02926
R14525 vdd.n4237 vdd.n4187 0.02926
R14526 vdd.n4048 vdd.n3997 0.02926
R14527 vdd.n3812 vdd.n3761 0.02926
R14528 vdd.n1458 vdd.n1408 0.02926
R14529 vdd.n1223 vdd.n1173 0.02926
R14530 vdd.n1034 vdd.n983 0.02926
R14531 vdd.n798 vdd.n747 0.02926
R14532 vdd.n10029 vdd.n9978 0.02926
R14533 vdd.n9793 vdd.n9742 0.02926
R14534 vdd.n470 vdd.n420 0.02926
R14535 vdd.n235 vdd.n185 0.02926
R14536 vdd.n6636 vdd 0.0251711
R14537 vdd.n3622 vdd 0.0251711
R14538 vdd.n608 vdd 0.0251711
R14539 vdd.n517 vdd 0.0251711
R14540 vdd.n7061 vdd.n7060 0.0235263
R14541 vdd.n7060 vdd 0.0235263
R14542 vdd.n6825 vdd.n6824 0.0235263
R14543 vdd.n6824 vdd 0.0235263
R14544 vdd.n4047 vdd.n4046 0.0235263
R14545 vdd.n4046 vdd 0.0235263
R14546 vdd.n3811 vdd.n3810 0.0235263
R14547 vdd.n3810 vdd 0.0235263
R14548 vdd.n1033 vdd.n1032 0.0235263
R14549 vdd.n1032 vdd 0.0235263
R14550 vdd.n797 vdd.n796 0.0235263
R14551 vdd.n796 vdd 0.0235263
R14552 vdd.n10028 vdd.n10027 0.0235263
R14553 vdd.n10027 vdd 0.0235263
R14554 vdd.n9792 vdd.n9791 0.0235263
R14555 vdd.n9791 vdd 0.0235263
R14556 vdd.n11971 vdd.n11970 0.0225448
R14557 vdd.t829 vdd.n11971 0.0225448
R14558 vdd.n11981 vdd.n11980 0.0225448
R14559 vdd.t1082 vdd.n11981 0.0225448
R14560 vdd.n12001 vdd.n12000 0.0225448
R14561 vdd.t1083 vdd.n12001 0.0225448
R14562 vdd.n11990 vdd.n11989 0.0225448
R14563 vdd.n11974 vdd.n11973 0.0225448
R14564 vdd.n11983 vdd.n11982 0.0225448
R14565 vdd.n11982 vdd.t1082 0.0225448
R14566 vdd.n12003 vdd.n12002 0.0225448
R14567 vdd.n12002 vdd.t1083 0.0225448
R14568 vdd.n11993 vdd.n11992 0.0225448
R14569 vdd.n11992 vdd.t1471 0.0225448
R14570 vdd.n112 vdd.n111 0.0225448
R14571 vdd.n121 vdd.n120 0.0225448
R14572 vdd.n120 vdd.t507 0.0225448
R14573 vdd.n126 vdd.n125 0.0225448
R14574 vdd.n126 vdd.t509 0.0225448
R14575 vdd.n129 vdd.n101 0.0225448
R14576 vdd.n129 vdd.t1182 0.0225448
R14577 vdd.n117 vdd.t1047 0.0225448
R14578 vdd.t507 vdd.n119 0.0225448
R14579 vdd.n135 vdd.t509 0.0225448
R14580 vdd.n133 vdd.n132 0.0225448
R14581 vdd.n136 vdd.n135 0.0225448
R14582 vdd.n119 vdd.n96 0.0225448
R14583 vdd.n117 vdd.n116 0.0225448
R14584 vdd.n158 vdd.n157 0.0225448
R14585 vdd.n167 vdd.n166 0.0225448
R14586 vdd.n166 vdd.t913 0.0225448
R14587 vdd.n172 vdd.n171 0.0225448
R14588 vdd.n172 vdd.t915 0.0225448
R14589 vdd.n175 vdd.n147 0.0225448
R14590 vdd.n175 vdd.t977 0.0225448
R14591 vdd.n163 vdd.t7 0.0225448
R14592 vdd.t913 vdd.n165 0.0225448
R14593 vdd.n181 vdd.t915 0.0225448
R14594 vdd.n179 vdd.n178 0.0225448
R14595 vdd.n182 vdd.n181 0.0225448
R14596 vdd.n165 vdd.n142 0.0225448
R14597 vdd.n163 vdd.n162 0.0225448
R14598 vdd.n255 vdd.n254 0.0225448
R14599 vdd.n264 vdd.n263 0.0225448
R14600 vdd.n263 vdd.t736 0.0225448
R14601 vdd.n269 vdd.n268 0.0225448
R14602 vdd.n269 vdd.t738 0.0225448
R14603 vdd.n272 vdd.n244 0.0225448
R14604 vdd.n272 vdd.t527 0.0225448
R14605 vdd.n260 vdd.t1475 0.0225448
R14606 vdd.t736 vdd.n262 0.0225448
R14607 vdd.n278 vdd.t738 0.0225448
R14608 vdd.n276 vdd.n275 0.0225448
R14609 vdd.n279 vdd.n278 0.0225448
R14610 vdd.n262 vdd.n239 0.0225448
R14611 vdd.n260 vdd.n259 0.0225448
R14612 vdd.n301 vdd.n300 0.0225448
R14613 vdd.n310 vdd.n309 0.0225448
R14614 vdd.n309 vdd.t161 0.0225448
R14615 vdd.n315 vdd.n314 0.0225448
R14616 vdd.n315 vdd.t163 0.0225448
R14617 vdd.n318 vdd.n290 0.0225448
R14618 vdd.n318 vdd.t1238 0.0225448
R14619 vdd.n306 vdd.t562 0.0225448
R14620 vdd.t161 vdd.n308 0.0225448
R14621 vdd.n324 vdd.t163 0.0225448
R14622 vdd.n322 vdd.n321 0.0225448
R14623 vdd.n325 vdd.n324 0.0225448
R14624 vdd.n308 vdd.n285 0.0225448
R14625 vdd.n306 vdd.n305 0.0225448
R14626 vdd.n347 vdd.n346 0.0225448
R14627 vdd.n356 vdd.n355 0.0225448
R14628 vdd.n355 vdd.t572 0.0225448
R14629 vdd.n361 vdd.n360 0.0225448
R14630 vdd.n361 vdd.t574 0.0225448
R14631 vdd.n364 vdd.n336 0.0225448
R14632 vdd.n364 vdd.t156 0.0225448
R14633 vdd.n352 vdd.t1298 0.0225448
R14634 vdd.t572 vdd.n354 0.0225448
R14635 vdd.n370 vdd.t574 0.0225448
R14636 vdd.n368 vdd.n367 0.0225448
R14637 vdd.n371 vdd.n370 0.0225448
R14638 vdd.n354 vdd.n331 0.0225448
R14639 vdd.n352 vdd.n351 0.0225448
R14640 vdd.n393 vdd.n392 0.0225448
R14641 vdd.n402 vdd.n401 0.0225448
R14642 vdd.n401 vdd.t1413 0.0225448
R14643 vdd.n407 vdd.n406 0.0225448
R14644 vdd.n407 vdd.t1415 0.0225448
R14645 vdd.n410 vdd.n382 0.0225448
R14646 vdd.n410 vdd.t959 0.0225448
R14647 vdd.n398 vdd.t1485 0.0225448
R14648 vdd.t1413 vdd.n400 0.0225448
R14649 vdd.n416 vdd.t1415 0.0225448
R14650 vdd.n414 vdd.n413 0.0225448
R14651 vdd.n417 vdd.n416 0.0225448
R14652 vdd.n400 vdd.n377 0.0225448
R14653 vdd.n398 vdd.n397 0.0225448
R14654 vdd.n490 vdd.n489 0.0225448
R14655 vdd.n499 vdd.n498 0.0225448
R14656 vdd.n498 vdd.t925 0.0225448
R14657 vdd.n504 vdd.n503 0.0225448
R14658 vdd.n504 vdd.t927 0.0225448
R14659 vdd.n507 vdd.n479 0.0225448
R14660 vdd.n507 vdd.t336 0.0225448
R14661 vdd.n495 vdd.t209 0.0225448
R14662 vdd.t925 vdd.n497 0.0225448
R14663 vdd.n513 vdd.t927 0.0225448
R14664 vdd.n511 vdd.n510 0.0225448
R14665 vdd.n514 vdd.n513 0.0225448
R14666 vdd.n497 vdd.n474 0.0225448
R14667 vdd.n495 vdd.n494 0.0225448
R14668 vdd.n536 vdd.n535 0.0225448
R14669 vdd.n545 vdd.n544 0.0225448
R14670 vdd.n544 vdd.t127 0.0225448
R14671 vdd.n550 vdd.n549 0.0225448
R14672 vdd.n550 vdd.t126 0.0225448
R14673 vdd.n553 vdd.n525 0.0225448
R14674 vdd.n553 vdd.t122 0.0225448
R14675 vdd.n541 vdd.t375 0.0225448
R14676 vdd.t127 vdd.n543 0.0225448
R14677 vdd.n559 vdd.t126 0.0225448
R14678 vdd.n557 vdd.n556 0.0225448
R14679 vdd.n560 vdd.n559 0.0225448
R14680 vdd.n543 vdd.n520 0.0225448
R14681 vdd.n541 vdd.n540 0.0225448
R14682 vdd.n6700 vdd.n6699 0.0225448
R14683 vdd.n6700 vdd.t728 0.0225448
R14684 vdd.n6710 vdd.n6709 0.0225448
R14685 vdd.n6709 vdd.t362 0.0225448
R14686 vdd.n6712 vdd.n6689 0.0225448
R14687 vdd.t363 vdd.n6689 0.0225448
R14688 vdd.n6719 vdd.n6718 0.0225448
R14689 vdd.n6715 vdd.n6714 0.0225448
R14690 vdd.n6715 vdd.t1288 0.0225448
R14691 vdd.n6724 vdd.n6723 0.0225448
R14692 vdd.n6723 vdd.t363 0.0225448
R14693 vdd.n6708 vdd.n6684 0.0225448
R14694 vdd.t362 vdd.n6708 0.0225448
R14695 vdd.n6706 vdd.n6705 0.0225448
R14696 vdd.n6746 vdd.n6745 0.0225448
R14697 vdd.n6746 vdd.t235 0.0225448
R14698 vdd.n6756 vdd.n6755 0.0225448
R14699 vdd.n6755 vdd.t624 0.0225448
R14700 vdd.n6758 vdd.n6735 0.0225448
R14701 vdd.t625 vdd.n6735 0.0225448
R14702 vdd.n6765 vdd.n6764 0.0225448
R14703 vdd.n6761 vdd.n6760 0.0225448
R14704 vdd.n6761 vdd.t207 0.0225448
R14705 vdd.n6770 vdd.n6769 0.0225448
R14706 vdd.n6769 vdd.t625 0.0225448
R14707 vdd.n6754 vdd.n6730 0.0225448
R14708 vdd.t624 vdd.n6754 0.0225448
R14709 vdd.n6752 vdd.n6751 0.0225448
R14710 vdd.n6844 vdd.n6843 0.0225448
R14711 vdd.n6844 vdd.t155 0.0225448
R14712 vdd.n6854 vdd.n6853 0.0225448
R14713 vdd.n6853 vdd.t152 0.0225448
R14714 vdd.n6856 vdd.n6833 0.0225448
R14715 vdd.t153 vdd.n6833 0.0225448
R14716 vdd.n6863 vdd.n6862 0.0225448
R14717 vdd.n6859 vdd.n6858 0.0225448
R14718 vdd.n6859 vdd.t1318 0.0225448
R14719 vdd.n6868 vdd.n6867 0.0225448
R14720 vdd.n6867 vdd.t153 0.0225448
R14721 vdd.n6852 vdd.n6828 0.0225448
R14722 vdd.t152 vdd.n6852 0.0225448
R14723 vdd.n6850 vdd.n6849 0.0225448
R14724 vdd.n6890 vdd.n6889 0.0225448
R14725 vdd.n6890 vdd.t413 0.0225448
R14726 vdd.n6900 vdd.n6899 0.0225448
R14727 vdd.n6899 vdd.t217 0.0225448
R14728 vdd.n6902 vdd.n6879 0.0225448
R14729 vdd.t218 vdd.n6879 0.0225448
R14730 vdd.n6909 vdd.n6908 0.0225448
R14731 vdd.n6905 vdd.n6904 0.0225448
R14732 vdd.n6905 vdd.t205 0.0225448
R14733 vdd.n6914 vdd.n6913 0.0225448
R14734 vdd.n6913 vdd.t218 0.0225448
R14735 vdd.n6898 vdd.n6874 0.0225448
R14736 vdd.t217 vdd.n6898 0.0225448
R14737 vdd.n6896 vdd.n6895 0.0225448
R14738 vdd.n6936 vdd.n6935 0.0225448
R14739 vdd.n6936 vdd.t983 0.0225448
R14740 vdd.n6946 vdd.n6945 0.0225448
R14741 vdd.n6945 vdd.t980 0.0225448
R14742 vdd.n6948 vdd.n6925 0.0225448
R14743 vdd.t981 vdd.n6925 0.0225448
R14744 vdd.n6955 vdd.n6954 0.0225448
R14745 vdd.n6951 vdd.n6950 0.0225448
R14746 vdd.n6951 vdd.t558 0.0225448
R14747 vdd.n6960 vdd.n6959 0.0225448
R14748 vdd.n6959 vdd.t981 0.0225448
R14749 vdd.n6944 vdd.n6920 0.0225448
R14750 vdd.t980 vdd.n6944 0.0225448
R14751 vdd.n6942 vdd.n6941 0.0225448
R14752 vdd.n6982 vdd.n6981 0.0225448
R14753 vdd.n6982 vdd.t1107 0.0225448
R14754 vdd.n6992 vdd.n6991 0.0225448
R14755 vdd.n6991 vdd.t806 0.0225448
R14756 vdd.n6994 vdd.n6971 0.0225448
R14757 vdd.t807 vdd.n6971 0.0225448
R14758 vdd.n7001 vdd.n7000 0.0225448
R14759 vdd.n6997 vdd.n6996 0.0225448
R14760 vdd.n6997 vdd.t377 0.0225448
R14761 vdd.n7006 vdd.n7005 0.0225448
R14762 vdd.n7005 vdd.t807 0.0225448
R14763 vdd.n6990 vdd.n6966 0.0225448
R14764 vdd.t806 vdd.n6990 0.0225448
R14765 vdd.n6988 vdd.n6987 0.0225448
R14766 vdd.n7080 vdd.n7079 0.0225448
R14767 vdd.n7080 vdd.t353 0.0225448
R14768 vdd.n7090 vdd.n7089 0.0225448
R14769 vdd.n7089 vdd.t302 0.0225448
R14770 vdd.n7092 vdd.n7069 0.0225448
R14771 vdd.t303 vdd.n7069 0.0225448
R14772 vdd.n7099 vdd.n7098 0.0225448
R14773 vdd.n7095 vdd.n7094 0.0225448
R14774 vdd.n7095 vdd.t587 0.0225448
R14775 vdd.n7104 vdd.n7103 0.0225448
R14776 vdd.n7103 vdd.t303 0.0225448
R14777 vdd.n7088 vdd.n7064 0.0225448
R14778 vdd.t302 vdd.n7088 0.0225448
R14779 vdd.n7086 vdd.n7085 0.0225448
R14780 vdd.n8538 vdd.n8537 0.0225448
R14781 vdd.n8538 vdd.t634 0.0225448
R14782 vdd.n8548 vdd.n8547 0.0225448
R14783 vdd.n8547 vdd.t1451 0.0225448
R14784 vdd.n8550 vdd.n8527 0.0225448
R14785 vdd.t1452 vdd.n8527 0.0225448
R14786 vdd.n8557 vdd.n8556 0.0225448
R14787 vdd.n8553 vdd.n8552 0.0225448
R14788 vdd.n8553 vdd.t482 0.0225448
R14789 vdd.n8562 vdd.n8561 0.0225448
R14790 vdd.n8561 vdd.t1452 0.0225448
R14791 vdd.n8546 vdd.n8522 0.0225448
R14792 vdd.t1451 vdd.n8546 0.0225448
R14793 vdd.n8544 vdd.n8543 0.0225448
R14794 vdd.n7128 vdd.n7127 0.0225448
R14795 vdd.n7137 vdd.n7136 0.0225448
R14796 vdd.n7136 vdd.t521 0.0225448
R14797 vdd.n7142 vdd.n7141 0.0225448
R14798 vdd.n7142 vdd.t520 0.0225448
R14799 vdd.n7145 vdd.n7117 0.0225448
R14800 vdd.n7145 vdd.t1025 0.0225448
R14801 vdd.n7133 vdd.t1463 0.0225448
R14802 vdd.t521 vdd.n7135 0.0225448
R14803 vdd.n7151 vdd.t520 0.0225448
R14804 vdd.n7149 vdd.n7148 0.0225448
R14805 vdd.n7152 vdd.n7151 0.0225448
R14806 vdd.n7135 vdd.n7112 0.0225448
R14807 vdd.n7133 vdd.n7132 0.0225448
R14808 vdd.n7174 vdd.n7173 0.0225448
R14809 vdd.n7183 vdd.n7182 0.0225448
R14810 vdd.n7182 vdd.t183 0.0225448
R14811 vdd.n7188 vdd.n7187 0.0225448
R14812 vdd.n7188 vdd.t182 0.0225448
R14813 vdd.n7191 vdd.n7163 0.0225448
R14814 vdd.n7191 vdd.t979 0.0225448
R14815 vdd.n7179 vdd.t1310 0.0225448
R14816 vdd.t183 vdd.n7181 0.0225448
R14817 vdd.n7197 vdd.t182 0.0225448
R14818 vdd.n7195 vdd.n7194 0.0225448
R14819 vdd.n7198 vdd.n7197 0.0225448
R14820 vdd.n7181 vdd.n7158 0.0225448
R14821 vdd.n7179 vdd.n7178 0.0225448
R14822 vdd.n7271 vdd.n7270 0.0225448
R14823 vdd.n7280 vdd.n7279 0.0225448
R14824 vdd.n7279 vdd.t883 0.0225448
R14825 vdd.n7285 vdd.n7284 0.0225448
R14826 vdd.n7285 vdd.t882 0.0225448
R14827 vdd.n7288 vdd.n7260 0.0225448
R14828 vdd.n7288 vdd.t1285 0.0225448
R14829 vdd.n7276 vdd.t1049 0.0225448
R14830 vdd.t883 vdd.n7278 0.0225448
R14831 vdd.n7294 vdd.t882 0.0225448
R14832 vdd.n7292 vdd.n7291 0.0225448
R14833 vdd.n7295 vdd.n7294 0.0225448
R14834 vdd.n7278 vdd.n7255 0.0225448
R14835 vdd.n7276 vdd.n7275 0.0225448
R14836 vdd.n7317 vdd.n7316 0.0225448
R14837 vdd.n7326 vdd.n7325 0.0225448
R14838 vdd.n7325 vdd.t532 0.0225448
R14839 vdd.n7331 vdd.n7330 0.0225448
R14840 vdd.n7331 vdd.t534 0.0225448
R14841 vdd.n7334 vdd.n7306 0.0225448
R14842 vdd.n7334 vdd.t536 0.0225448
R14843 vdd.n7322 vdd.t1360 0.0225448
R14844 vdd.t532 vdd.n7324 0.0225448
R14845 vdd.n7340 vdd.t534 0.0225448
R14846 vdd.n7338 vdd.n7337 0.0225448
R14847 vdd.n7341 vdd.n7340 0.0225448
R14848 vdd.n7324 vdd.n7301 0.0225448
R14849 vdd.n7322 vdd.n7321 0.0225448
R14850 vdd.n7363 vdd.n7362 0.0225448
R14851 vdd.n7372 vdd.n7371 0.0225448
R14852 vdd.n7371 vdd.t1092 0.0225448
R14853 vdd.n7377 vdd.n7376 0.0225448
R14854 vdd.n7377 vdd.t1091 0.0225448
R14855 vdd.n7380 vdd.n7352 0.0225448
R14856 vdd.n7380 vdd.t1094 0.0225448
R14857 vdd.n7368 vdd.t593 0.0225448
R14858 vdd.t1092 vdd.n7370 0.0225448
R14859 vdd.n7386 vdd.t1091 0.0225448
R14860 vdd.n7384 vdd.n7383 0.0225448
R14861 vdd.n7387 vdd.n7386 0.0225448
R14862 vdd.n7370 vdd.n7347 0.0225448
R14863 vdd.n7368 vdd.n7367 0.0225448
R14864 vdd.n7409 vdd.n7408 0.0225448
R14865 vdd.n7418 vdd.n7417 0.0225448
R14866 vdd.n7417 vdd.t1253 0.0225448
R14867 vdd.n7423 vdd.n7422 0.0225448
R14868 vdd.n7423 vdd.t1252 0.0225448
R14869 vdd.n7426 vdd.n7398 0.0225448
R14870 vdd.n7426 vdd.t1255 0.0225448
R14871 vdd.n7414 vdd.t379 0.0225448
R14872 vdd.t1253 vdd.n7416 0.0225448
R14873 vdd.n7432 vdd.t1252 0.0225448
R14874 vdd.n7430 vdd.n7429 0.0225448
R14875 vdd.n7433 vdd.n7432 0.0225448
R14876 vdd.n7416 vdd.n7393 0.0225448
R14877 vdd.n7414 vdd.n7413 0.0225448
R14878 vdd.n7506 vdd.n7505 0.0225448
R14879 vdd.n7515 vdd.n7514 0.0225448
R14880 vdd.n7514 vdd.t931 0.0225448
R14881 vdd.n7520 vdd.n7519 0.0225448
R14882 vdd.n7520 vdd.t930 0.0225448
R14883 vdd.n7523 vdd.n7495 0.0225448
R14884 vdd.n7523 vdd.t143 0.0225448
R14885 vdd.n7511 vdd.t1326 0.0225448
R14886 vdd.t931 vdd.n7513 0.0225448
R14887 vdd.n7529 vdd.t930 0.0225448
R14888 vdd.n7527 vdd.n7526 0.0225448
R14889 vdd.n7530 vdd.n7529 0.0225448
R14890 vdd.n7513 vdd.n7490 0.0225448
R14891 vdd.n7511 vdd.n7510 0.0225448
R14892 vdd.n6655 vdd.n6654 0.0225448
R14893 vdd.n6664 vdd.n6663 0.0225448
R14894 vdd.n6663 vdd.t704 0.0225448
R14895 vdd.n6669 vdd.n6668 0.0225448
R14896 vdd.n6669 vdd.t703 0.0225448
R14897 vdd.n6672 vdd.n6644 0.0225448
R14898 vdd.n6672 vdd.t1088 0.0225448
R14899 vdd.n6660 vdd.t484 0.0225448
R14900 vdd.t704 vdd.n6662 0.0225448
R14901 vdd.n6678 vdd.t703 0.0225448
R14902 vdd.n6676 vdd.n6675 0.0225448
R14903 vdd.n6679 vdd.n6678 0.0225448
R14904 vdd.n6662 vdd.n6639 0.0225448
R14905 vdd.n6660 vdd.n6659 0.0225448
R14906 vdd.n7550 vdd.n7549 0.0225448
R14907 vdd.n7559 vdd.n7558 0.0225448
R14908 vdd.n7558 vdd.t1273 0.0225448
R14909 vdd.n7564 vdd.n7563 0.0225448
R14910 vdd.n7564 vdd.t1272 0.0225448
R14911 vdd.n7567 vdd.n7539 0.0225448
R14912 vdd.n7567 vdd.t1263 0.0225448
R14913 vdd.n7555 vdd.t898 0.0225448
R14914 vdd.t1273 vdd.n7557 0.0225448
R14915 vdd.n7573 vdd.t1272 0.0225448
R14916 vdd.n7571 vdd.n7570 0.0225448
R14917 vdd.n7574 vdd.n7573 0.0225448
R14918 vdd.n7557 vdd.n7534 0.0225448
R14919 vdd.n7555 vdd.n7554 0.0225448
R14920 vdd.n7595 vdd.n7594 0.0225448
R14921 vdd.n7604 vdd.n7603 0.0225448
R14922 vdd.n7603 vdd.t886 0.0225448
R14923 vdd.n7609 vdd.n7608 0.0225448
R14924 vdd.n7609 vdd.t885 0.0225448
R14925 vdd.n7612 vdd.n7584 0.0225448
R14926 vdd.n7612 vdd.t809 0.0225448
R14927 vdd.n7600 vdd.t166 0.0225448
R14928 vdd.t886 vdd.n7602 0.0225448
R14929 vdd.n7618 vdd.t885 0.0225448
R14930 vdd.n7616 vdd.n7615 0.0225448
R14931 vdd.n7619 vdd.n7618 0.0225448
R14932 vdd.n7602 vdd.n7579 0.0225448
R14933 vdd.n7600 vdd.n7599 0.0225448
R14934 vdd.n7645 vdd.n7644 0.0225448
R14935 vdd.n7654 vdd.n7653 0.0225448
R14936 vdd.n7653 vdd.t223 0.0225448
R14937 vdd.n7659 vdd.n7658 0.0225448
R14938 vdd.n7659 vdd.t225 0.0225448
R14939 vdd.n7662 vdd.n7634 0.0225448
R14940 vdd.n7662 vdd.t1226 0.0225448
R14941 vdd.n7650 vdd.t589 0.0225448
R14942 vdd.t223 vdd.n7652 0.0225448
R14943 vdd.n7668 vdd.t225 0.0225448
R14944 vdd.n7666 vdd.n7665 0.0225448
R14945 vdd.n7669 vdd.n7668 0.0225448
R14946 vdd.n7652 vdd.n7629 0.0225448
R14947 vdd.n7650 vdd.n7649 0.0225448
R14948 vdd.n7691 vdd.n7690 0.0225448
R14949 vdd.n7700 vdd.n7699 0.0225448
R14950 vdd.n7699 vdd.t251 0.0225448
R14951 vdd.n7705 vdd.n7704 0.0225448
R14952 vdd.n7705 vdd.t250 0.0225448
R14953 vdd.n7708 vdd.n7680 0.0225448
R14954 vdd.n7708 vdd.t874 0.0225448
R14955 vdd.n7696 vdd.t862 0.0225448
R14956 vdd.t251 vdd.n7698 0.0225448
R14957 vdd.n7714 vdd.t250 0.0225448
R14958 vdd.n7712 vdd.n7711 0.0225448
R14959 vdd.n7715 vdd.n7714 0.0225448
R14960 vdd.n7698 vdd.n7675 0.0225448
R14961 vdd.n7696 vdd.n7695 0.0225448
R14962 vdd.n7739 vdd.n7738 0.0225448
R14963 vdd.n7748 vdd.n7747 0.0225448
R14964 vdd.n7747 vdd.t1265 0.0225448
R14965 vdd.n7753 vdd.n7752 0.0225448
R14966 vdd.n7753 vdd.t1264 0.0225448
R14967 vdd.n7756 vdd.n7728 0.0225448
R14968 vdd.n7756 vdd.t1078 0.0225448
R14969 vdd.n7744 vdd.t1342 0.0225448
R14970 vdd.t1265 vdd.n7746 0.0225448
R14971 vdd.n7762 vdd.t1264 0.0225448
R14972 vdd.n7760 vdd.n7759 0.0225448
R14973 vdd.n7763 vdd.n7762 0.0225448
R14974 vdd.n7746 vdd.n7723 0.0225448
R14975 vdd.n7744 vdd.n7743 0.0225448
R14976 vdd.n7457 vdd.n7456 0.0225448
R14977 vdd.n7460 vdd.n7459 0.0225448
R14978 vdd.n7459 vdd.t443 0.0225448
R14979 vdd.n7465 vdd.n7464 0.0225448
R14980 vdd.n7465 vdd.t442 0.0225448
R14981 vdd.n7468 vdd.n7449 0.0225448
R14982 vdd.n7468 vdd.t892 0.0225448
R14983 vdd.n7481 vdd.t1154 0.0225448
R14984 vdd.n7479 vdd.t443 0.0225448
R14985 vdd.n7474 vdd.t442 0.0225448
R14986 vdd.n7472 vdd.n7471 0.0225448
R14987 vdd.n7475 vdd.n7474 0.0225448
R14988 vdd.n7479 vdd.n7478 0.0225448
R14989 vdd.n7482 vdd.n7481 0.0225448
R14990 vdd.n7786 vdd.n7785 0.0225448
R14991 vdd.n7795 vdd.n7794 0.0225448
R14992 vdd.n7794 vdd.t518 0.0225448
R14993 vdd.n7800 vdd.n7799 0.0225448
R14994 vdd.n7800 vdd.t517 0.0225448
R14995 vdd.n7803 vdd.n7775 0.0225448
R14996 vdd.n7803 vdd.t1506 0.0225448
R14997 vdd.n7791 vdd.t896 0.0225448
R14998 vdd.t518 vdd.n7793 0.0225448
R14999 vdd.n7809 vdd.t517 0.0225448
R15000 vdd.n7807 vdd.n7806 0.0225448
R15001 vdd.n7810 vdd.n7809 0.0225448
R15002 vdd.n7793 vdd.n7770 0.0225448
R15003 vdd.n7791 vdd.n7790 0.0225448
R15004 vdd.n7831 vdd.n7830 0.0225448
R15005 vdd.n7840 vdd.n7839 0.0225448
R15006 vdd.n7839 vdd.t239 0.0225448
R15007 vdd.n7845 vdd.n7844 0.0225448
R15008 vdd.n7845 vdd.t238 0.0225448
R15009 vdd.n7848 vdd.n7820 0.0225448
R15010 vdd.n7848 vdd.t241 0.0225448
R15011 vdd.n7836 vdd.t837 0.0225448
R15012 vdd.t239 vdd.n7838 0.0225448
R15013 vdd.n7854 vdd.t238 0.0225448
R15014 vdd.n7852 vdd.n7851 0.0225448
R15015 vdd.n7855 vdd.n7854 0.0225448
R15016 vdd.n7838 vdd.n7815 0.0225448
R15017 vdd.n7836 vdd.n7835 0.0225448
R15018 vdd.n7877 vdd.n7876 0.0225448
R15019 vdd.n7886 vdd.n7885 0.0225448
R15020 vdd.n7885 vdd.t541 0.0225448
R15021 vdd.n7891 vdd.n7890 0.0225448
R15022 vdd.n7891 vdd.t540 0.0225448
R15023 vdd.n7894 vdd.n7866 0.0225448
R15024 vdd.n7894 vdd.t543 0.0225448
R15025 vdd.n7882 vdd.t1375 0.0225448
R15026 vdd.t541 vdd.n7884 0.0225448
R15027 vdd.n7900 vdd.t540 0.0225448
R15028 vdd.n7898 vdd.n7897 0.0225448
R15029 vdd.n7901 vdd.n7900 0.0225448
R15030 vdd.n7884 vdd.n7861 0.0225448
R15031 vdd.n7882 vdd.n7881 0.0225448
R15032 vdd.n7928 vdd.n7927 0.0225448
R15033 vdd.n7937 vdd.n7936 0.0225448
R15034 vdd.n7936 vdd.t68 0.0225448
R15035 vdd.n7942 vdd.n7941 0.0225448
R15036 vdd.n7942 vdd.t67 0.0225448
R15037 vdd.n7945 vdd.n7917 0.0225448
R15038 vdd.n7945 vdd.t306 0.0225448
R15039 vdd.n7933 vdd.t486 0.0225448
R15040 vdd.t68 vdd.n7935 0.0225448
R15041 vdd.n7951 vdd.t67 0.0225448
R15042 vdd.n7949 vdd.n7948 0.0225448
R15043 vdd.n7952 vdd.n7951 0.0225448
R15044 vdd.n7935 vdd.n7912 0.0225448
R15045 vdd.n7933 vdd.n7932 0.0225448
R15046 vdd.n7974 vdd.n7973 0.0225448
R15047 vdd.n7983 vdd.n7982 0.0225448
R15048 vdd.n7982 vdd.t319 0.0225448
R15049 vdd.n7988 vdd.n7987 0.0225448
R15050 vdd.n7988 vdd.t318 0.0225448
R15051 vdd.n7991 vdd.n7963 0.0225448
R15052 vdd.n7991 vdd.t620 0.0225448
R15053 vdd.n7979 vdd.t872 0.0225448
R15054 vdd.t319 vdd.n7981 0.0225448
R15055 vdd.n7997 vdd.t318 0.0225448
R15056 vdd.n7995 vdd.n7994 0.0225448
R15057 vdd.n7998 vdd.n7997 0.0225448
R15058 vdd.n7981 vdd.n7958 0.0225448
R15059 vdd.n7979 vdd.n7978 0.0225448
R15060 vdd.n8022 vdd.n8021 0.0225448
R15061 vdd.n8031 vdd.n8030 0.0225448
R15062 vdd.n8030 vdd.t962 0.0225448
R15063 vdd.n8036 vdd.n8035 0.0225448
R15064 vdd.n8036 vdd.t961 0.0225448
R15065 vdd.n8039 vdd.n8011 0.0225448
R15066 vdd.n8039 vdd.t978 0.0225448
R15067 vdd.n8027 vdd.t1330 0.0225448
R15068 vdd.t962 vdd.n8029 0.0225448
R15069 vdd.n8045 vdd.t961 0.0225448
R15070 vdd.n8043 vdd.n8042 0.0225448
R15071 vdd.n8046 vdd.n8045 0.0225448
R15072 vdd.n8029 vdd.n8006 0.0225448
R15073 vdd.n8027 vdd.n8026 0.0225448
R15074 vdd.n8068 vdd.n8067 0.0225448
R15075 vdd.n8077 vdd.n8076 0.0225448
R15076 vdd.n8076 vdd.t643 0.0225448
R15077 vdd.n8082 vdd.n8081 0.0225448
R15078 vdd.n8082 vdd.t642 0.0225448
R15079 vdd.n8085 vdd.n8057 0.0225448
R15080 vdd.n8085 vdd.t22 0.0225448
R15081 vdd.n8073 vdd.t36 0.0225448
R15082 vdd.t643 vdd.n8075 0.0225448
R15083 vdd.n8091 vdd.t642 0.0225448
R15084 vdd.n8089 vdd.n8088 0.0225448
R15085 vdd.n8092 vdd.n8091 0.0225448
R15086 vdd.n8075 vdd.n8052 0.0225448
R15087 vdd.n8073 vdd.n8072 0.0225448
R15088 vdd.n8113 vdd.n8112 0.0225448
R15089 vdd.n8122 vdd.n8121 0.0225448
R15090 vdd.n8121 vdd.t130 0.0225448
R15091 vdd.n8127 vdd.n8126 0.0225448
R15092 vdd.n8127 vdd.t129 0.0225448
R15093 vdd.n8130 vdd.n8102 0.0225448
R15094 vdd.n8130 vdd.t335 0.0225448
R15095 vdd.n8118 vdd.t835 0.0225448
R15096 vdd.t130 vdd.n8120 0.0225448
R15097 vdd.n8136 vdd.t129 0.0225448
R15098 vdd.n8134 vdd.n8133 0.0225448
R15099 vdd.n8137 vdd.n8136 0.0225448
R15100 vdd.n8120 vdd.n8097 0.0225448
R15101 vdd.n8118 vdd.n8117 0.0225448
R15102 vdd.n8163 vdd.n8162 0.0225448
R15103 vdd.n8172 vdd.n8171 0.0225448
R15104 vdd.n8171 vdd.t325 0.0225448
R15105 vdd.n8177 vdd.n8176 0.0225448
R15106 vdd.n8177 vdd.t324 0.0225448
R15107 vdd.n8180 vdd.n8152 0.0225448
R15108 vdd.n8180 vdd.t70 0.0225448
R15109 vdd.n8168 vdd.t201 0.0225448
R15110 vdd.t325 vdd.n8170 0.0225448
R15111 vdd.n8186 vdd.t324 0.0225448
R15112 vdd.n8184 vdd.n8183 0.0225448
R15113 vdd.n8187 vdd.n8186 0.0225448
R15114 vdd.n8170 vdd.n8147 0.0225448
R15115 vdd.n8168 vdd.n8167 0.0225448
R15116 vdd.n8209 vdd.n8208 0.0225448
R15117 vdd.n8218 vdd.n8217 0.0225448
R15118 vdd.n8217 vdd.t248 0.0225448
R15119 vdd.n8223 vdd.n8222 0.0225448
R15120 vdd.n8223 vdd.t247 0.0225448
R15121 vdd.n8226 vdd.n8198 0.0225448
R15122 vdd.n8226 vdd.t1442 0.0225448
R15123 vdd.n8214 vdd.t973 0.0225448
R15124 vdd.t248 vdd.n8216 0.0225448
R15125 vdd.n8232 vdd.t247 0.0225448
R15126 vdd.n8230 vdd.n8229 0.0225448
R15127 vdd.n8233 vdd.n8232 0.0225448
R15128 vdd.n8216 vdd.n8193 0.0225448
R15129 vdd.n8214 vdd.n8213 0.0225448
R15130 vdd.n8257 vdd.n8256 0.0225448
R15131 vdd.n8266 vdd.n8265 0.0225448
R15132 vdd.n8265 vdd.t1448 0.0225448
R15133 vdd.n8271 vdd.n8270 0.0225448
R15134 vdd.n8271 vdd.t1450 0.0225448
R15135 vdd.n8274 vdd.n8246 0.0225448
R15136 vdd.n8274 vdd.t743 0.0225448
R15137 vdd.n8262 vdd.t1346 0.0225448
R15138 vdd.t1448 vdd.n8264 0.0225448
R15139 vdd.n8280 vdd.t1450 0.0225448
R15140 vdd.n8278 vdd.n8277 0.0225448
R15141 vdd.n8281 vdd.n8280 0.0225448
R15142 vdd.n8264 vdd.n8241 0.0225448
R15143 vdd.n8262 vdd.n8261 0.0225448
R15144 vdd.n7222 vdd.n7221 0.0225448
R15145 vdd.n7225 vdd.n7224 0.0225448
R15146 vdd.n7224 vdd.t1394 0.0225448
R15147 vdd.n7230 vdd.n7229 0.0225448
R15148 vdd.n7230 vdd.t1393 0.0225448
R15149 vdd.n7233 vdd.n7214 0.0225448
R15150 vdd.n7233 vdd.t277 0.0225448
R15151 vdd.n7246 vdd.t1459 0.0225448
R15152 vdd.n7244 vdd.t1394 0.0225448
R15153 vdd.n7239 vdd.t1393 0.0225448
R15154 vdd.n7237 vdd.n7236 0.0225448
R15155 vdd.n7240 vdd.n7239 0.0225448
R15156 vdd.n7244 vdd.n7243 0.0225448
R15157 vdd.n7247 vdd.n7246 0.0225448
R15158 vdd.n8304 vdd.n8303 0.0225448
R15159 vdd.n8313 vdd.n8312 0.0225448
R15160 vdd.n8312 vdd.t1176 0.0225448
R15161 vdd.n8318 vdd.n8317 0.0225448
R15162 vdd.n8318 vdd.t1175 0.0225448
R15163 vdd.n8321 vdd.n8293 0.0225448
R15164 vdd.n8321 vdd.t1112 0.0225448
R15165 vdd.n8309 vdd.t854 0.0225448
R15166 vdd.t1176 vdd.n8311 0.0225448
R15167 vdd.n8327 vdd.t1175 0.0225448
R15168 vdd.n8325 vdd.n8324 0.0225448
R15169 vdd.n8328 vdd.n8327 0.0225448
R15170 vdd.n8311 vdd.n8288 0.0225448
R15171 vdd.n8309 vdd.n8308 0.0225448
R15172 vdd.n8349 vdd.n8348 0.0225448
R15173 vdd.n8358 vdd.n8357 0.0225448
R15174 vdd.n8357 vdd.t450 0.0225448
R15175 vdd.n8363 vdd.n8362 0.0225448
R15176 vdd.n8363 vdd.t449 0.0225448
R15177 vdd.n8366 vdd.n8338 0.0225448
R15178 vdd.n8366 vdd.t343 0.0225448
R15179 vdd.n8354 vdd.t56 0.0225448
R15180 vdd.t450 vdd.n8356 0.0225448
R15181 vdd.n8372 vdd.t449 0.0225448
R15182 vdd.n8370 vdd.n8369 0.0225448
R15183 vdd.n8373 vdd.n8372 0.0225448
R15184 vdd.n8356 vdd.n8333 0.0225448
R15185 vdd.n8354 vdd.n8353 0.0225448
R15186 vdd.n8399 vdd.n8398 0.0225448
R15187 vdd.n8408 vdd.n8407 0.0225448
R15188 vdd.n8407 vdd.t879 0.0225448
R15189 vdd.n8413 vdd.n8412 0.0225448
R15190 vdd.n8413 vdd.t878 0.0225448
R15191 vdd.n8416 vdd.n8388 0.0225448
R15192 vdd.n8416 vdd.t881 0.0225448
R15193 vdd.n8404 vdd.t9 0.0225448
R15194 vdd.t879 vdd.n8406 0.0225448
R15195 vdd.n8422 vdd.t878 0.0225448
R15196 vdd.n8420 vdd.n8419 0.0225448
R15197 vdd.n8423 vdd.n8422 0.0225448
R15198 vdd.n8406 vdd.n8383 0.0225448
R15199 vdd.n8404 vdd.n8403 0.0225448
R15200 vdd.n8445 vdd.n8444 0.0225448
R15201 vdd.n8454 vdd.n8453 0.0225448
R15202 vdd.n8453 vdd.t1420 0.0225448
R15203 vdd.n8459 vdd.n8458 0.0225448
R15204 vdd.n8459 vdd.t1419 0.0225448
R15205 vdd.n8462 vdd.n8434 0.0225448
R15206 vdd.n8462 vdd.t1149 0.0225448
R15207 vdd.n8450 vdd.t40 0.0225448
R15208 vdd.t1420 vdd.n8452 0.0225448
R15209 vdd.n8468 vdd.t1419 0.0225448
R15210 vdd.n8466 vdd.n8465 0.0225448
R15211 vdd.n8469 vdd.n8468 0.0225448
R15212 vdd.n8452 vdd.n8429 0.0225448
R15213 vdd.n8450 vdd.n8449 0.0225448
R15214 vdd.n8493 vdd.n8492 0.0225448
R15215 vdd.n8502 vdd.n8501 0.0225448
R15216 vdd.n8501 vdd.t1064 0.0225448
R15217 vdd.n8507 vdd.n8506 0.0225448
R15218 vdd.n8507 vdd.t1063 0.0225448
R15219 vdd.n8510 vdd.n8482 0.0225448
R15220 vdd.n8510 vdd.t1066 0.0225448
R15221 vdd.n8498 vdd.t211 0.0225448
R15222 vdd.t1064 vdd.n8500 0.0225448
R15223 vdd.n8516 vdd.t1063 0.0225448
R15224 vdd.n8514 vdd.n8513 0.0225448
R15225 vdd.n8517 vdd.n8516 0.0225448
R15226 vdd.n8500 vdd.n8477 0.0225448
R15227 vdd.n8498 vdd.n8497 0.0225448
R15228 vdd.n8631 vdd.n8630 0.0225448
R15229 vdd.n8631 vdd.t284 0.0225448
R15230 vdd.n8641 vdd.n8640 0.0225448
R15231 vdd.n8640 vdd.t1079 0.0225448
R15232 vdd.n8643 vdd.n8620 0.0225448
R15233 vdd.t1080 vdd.n8620 0.0225448
R15234 vdd.n8650 vdd.n8649 0.0225448
R15235 vdd.n8646 vdd.n8645 0.0225448
R15236 vdd.n8646 vdd.t848 0.0225448
R15237 vdd.n8655 vdd.n8654 0.0225448
R15238 vdd.n8654 vdd.t1080 0.0225448
R15239 vdd.n8639 vdd.n8615 0.0225448
R15240 vdd.t1079 vdd.n8639 0.0225448
R15241 vdd.n8637 vdd.n8636 0.0225448
R15242 vdd.n8585 vdd.n8584 0.0225448
R15243 vdd.n8585 vdd.t412 0.0225448
R15244 vdd.n8595 vdd.n8594 0.0225448
R15245 vdd.n8594 vdd.t764 0.0225448
R15246 vdd.n8597 vdd.n8574 0.0225448
R15247 vdd.t762 vdd.n8574 0.0225448
R15248 vdd.n8604 vdd.n8603 0.0225448
R15249 vdd.n8600 vdd.n8599 0.0225448
R15250 vdd.n8600 vdd.t773 0.0225448
R15251 vdd.n8609 vdd.n8608 0.0225448
R15252 vdd.n8608 vdd.t762 0.0225448
R15253 vdd.n8593 vdd.n8569 0.0225448
R15254 vdd.t764 vdd.n8593 0.0225448
R15255 vdd.n8591 vdd.n8590 0.0225448
R15256 vdd.n8678 vdd.n8677 0.0225448
R15257 vdd.n8678 vdd.t1143 0.0225448
R15258 vdd.n8688 vdd.n8687 0.0225448
R15259 vdd.n8687 vdd.t254 0.0225448
R15260 vdd.n8690 vdd.n8667 0.0225448
R15261 vdd.t255 vdd.n8667 0.0225448
R15262 vdd.n8697 vdd.n8696 0.0225448
R15263 vdd.n8693 vdd.n8692 0.0225448
R15264 vdd.n8693 vdd.t1314 0.0225448
R15265 vdd.n8702 vdd.n8701 0.0225448
R15266 vdd.n8701 vdd.t255 0.0225448
R15267 vdd.n8686 vdd.n8662 0.0225448
R15268 vdd.t254 vdd.n8686 0.0225448
R15269 vdd.n8684 vdd.n8683 0.0225448
R15270 vdd.n8726 vdd.n8725 0.0225448
R15271 vdd.n8726 vdd.t658 0.0225448
R15272 vdd.n8736 vdd.n8735 0.0225448
R15273 vdd.n8735 vdd.t933 0.0225448
R15274 vdd.n8738 vdd.n8715 0.0225448
R15275 vdd.t934 vdd.n8715 0.0225448
R15276 vdd.n8745 vdd.n8744 0.0225448
R15277 vdd.n8741 vdd.n8740 0.0225448
R15278 vdd.n8741 vdd.t856 0.0225448
R15279 vdd.n8750 vdd.n8749 0.0225448
R15280 vdd.n8749 vdd.t934 0.0225448
R15281 vdd.n8734 vdd.n8710 0.0225448
R15282 vdd.t933 vdd.n8734 0.0225448
R15283 vdd.n8732 vdd.n8731 0.0225448
R15284 vdd.n8772 vdd.n8771 0.0225448
R15285 vdd.n8772 vdd.t1507 0.0225448
R15286 vdd.n8782 vdd.n8781 0.0225448
R15287 vdd.n8781 vdd.t190 0.0225448
R15288 vdd.n8784 vdd.n8761 0.0225448
R15289 vdd.t188 vdd.n8761 0.0225448
R15290 vdd.n8791 vdd.n8790 0.0225448
R15291 vdd.n8787 vdd.n8786 0.0225448
R15292 vdd.n8787 vdd.t1467 0.0225448
R15293 vdd.n8796 vdd.n8795 0.0225448
R15294 vdd.n8795 vdd.t188 0.0225448
R15295 vdd.n8780 vdd.n8756 0.0225448
R15296 vdd.t190 vdd.n8780 0.0225448
R15297 vdd.n8778 vdd.n8777 0.0225448
R15298 vdd.n7036 vdd.n7035 0.0225448
R15299 vdd.n7035 vdd.t1089 0.0225448
R15300 vdd.n7038 vdd.n7024 0.0225448
R15301 vdd.t82 vdd.n7024 0.0225448
R15302 vdd.n7041 vdd.n7040 0.0225448
R15303 vdd.t80 vdd.n7041 0.0225448
R15304 vdd.n7056 vdd.n7055 0.0225448
R15305 vdd.n7053 vdd.n7013 0.0225448
R15306 vdd.t97 vdd.n7053 0.0225448
R15307 vdd.n7048 vdd.n7018 0.0225448
R15308 vdd.t80 vdd.n7018 0.0225448
R15309 vdd.n7044 vdd.n7043 0.0225448
R15310 vdd.n7043 vdd.t82 0.0225448
R15311 vdd.n7033 vdd.n7032 0.0225448
R15312 vdd.n8914 vdd.n8913 0.0225448
R15313 vdd.n8914 vdd.t66 0.0225448
R15314 vdd.n8924 vdd.n8923 0.0225448
R15315 vdd.n8923 vdd.t139 0.0225448
R15316 vdd.n8926 vdd.n8903 0.0225448
R15317 vdd.t137 vdd.n8903 0.0225448
R15318 vdd.n8933 vdd.n8932 0.0225448
R15319 vdd.n8929 vdd.n8928 0.0225448
R15320 vdd.n8929 vdd.t825 0.0225448
R15321 vdd.n8938 vdd.n8937 0.0225448
R15322 vdd.n8937 vdd.t137 0.0225448
R15323 vdd.n8922 vdd.n8898 0.0225448
R15324 vdd.t139 vdd.n8922 0.0225448
R15325 vdd.n8920 vdd.n8919 0.0225448
R15326 vdd.n8867 vdd.n8866 0.0225448
R15327 vdd.n8867 vdd.t1195 0.0225448
R15328 vdd.n8877 vdd.n8876 0.0225448
R15329 vdd.n8876 vdd.t584 0.0225448
R15330 vdd.n8879 vdd.n8856 0.0225448
R15331 vdd.t585 vdd.n8856 0.0225448
R15332 vdd.n8886 vdd.n8885 0.0225448
R15333 vdd.n8882 vdd.n8881 0.0225448
R15334 vdd.n8882 vdd.t765 0.0225448
R15335 vdd.n8891 vdd.n8890 0.0225448
R15336 vdd.n8890 vdd.t585 0.0225448
R15337 vdd.n8875 vdd.n8851 0.0225448
R15338 vdd.t584 vdd.n8875 0.0225448
R15339 vdd.n8873 vdd.n8872 0.0225448
R15340 vdd.n8821 vdd.n8820 0.0225448
R15341 vdd.n8821 vdd.t264 0.0225448
R15342 vdd.n8831 vdd.n8830 0.0225448
R15343 vdd.n8830 vdd.t1201 0.0225448
R15344 vdd.n8833 vdd.n8810 0.0225448
R15345 vdd.t1199 vdd.n8810 0.0225448
R15346 vdd.n8840 vdd.n8839 0.0225448
R15347 vdd.n8836 vdd.n8835 0.0225448
R15348 vdd.n8836 vdd.t1129 0.0225448
R15349 vdd.n8845 vdd.n8844 0.0225448
R15350 vdd.n8844 vdd.t1199 0.0225448
R15351 vdd.n8829 vdd.n8805 0.0225448
R15352 vdd.t1201 vdd.n8829 0.0225448
R15353 vdd.n8827 vdd.n8826 0.0225448
R15354 vdd.n8961 vdd.n8960 0.0225448
R15355 vdd.n8961 vdd.t758 0.0225448
R15356 vdd.n8971 vdd.n8970 0.0225448
R15357 vdd.n8970 vdd.t755 0.0225448
R15358 vdd.n8973 vdd.n8950 0.0225448
R15359 vdd.t756 vdd.n8950 0.0225448
R15360 vdd.n8980 vdd.n8979 0.0225448
R15361 vdd.n8976 vdd.n8975 0.0225448
R15362 vdd.n8976 vdd.t458 0.0225448
R15363 vdd.n8985 vdd.n8984 0.0225448
R15364 vdd.n8984 vdd.t756 0.0225448
R15365 vdd.n8969 vdd.n8945 0.0225448
R15366 vdd.t755 vdd.n8969 0.0225448
R15367 vdd.n8967 vdd.n8966 0.0225448
R15368 vdd.n9009 vdd.n9008 0.0225448
R15369 vdd.n9009 vdd.t1062 0.0225448
R15370 vdd.n9019 vdd.n9018 0.0225448
R15371 vdd.n9018 vdd.t640 0.0225448
R15372 vdd.n9021 vdd.n8998 0.0225448
R15373 vdd.t638 vdd.n8998 0.0225448
R15374 vdd.n9028 vdd.n9027 0.0225448
R15375 vdd.n9024 vdd.n9023 0.0225448
R15376 vdd.n9024 vdd.t864 0.0225448
R15377 vdd.n9033 vdd.n9032 0.0225448
R15378 vdd.n9032 vdd.t638 0.0225448
R15379 vdd.n9017 vdd.n8993 0.0225448
R15380 vdd.t640 vdd.n9017 0.0225448
R15381 vdd.n9015 vdd.n9014 0.0225448
R15382 vdd.n9055 vdd.n9054 0.0225448
R15383 vdd.n9055 vdd.t1108 0.0225448
R15384 vdd.n9065 vdd.n9064 0.0225448
R15385 vdd.n9064 vdd.t1526 0.0225448
R15386 vdd.n9067 vdd.n9044 0.0225448
R15387 vdd.t1524 vdd.n9044 0.0225448
R15388 vdd.n9074 vdd.n9073 0.0225448
R15389 vdd.n9070 vdd.n9069 0.0225448
R15390 vdd.n9070 vdd.t1477 0.0225448
R15391 vdd.n9079 vdd.n9078 0.0225448
R15392 vdd.n9078 vdd.t1524 0.0225448
R15393 vdd.n9063 vdd.n9039 0.0225448
R15394 vdd.t1526 vdd.n9063 0.0225448
R15395 vdd.n9061 vdd.n9060 0.0225448
R15396 vdd.n9149 vdd.n9148 0.0225448
R15397 vdd.n9149 vdd.t64 0.0225448
R15398 vdd.n9159 vdd.n9158 0.0225448
R15399 vdd.n9158 vdd.t77 0.0225448
R15400 vdd.n9161 vdd.n9138 0.0225448
R15401 vdd.t78 vdd.n9138 0.0225448
R15402 vdd.n9168 vdd.n9167 0.0225448
R15403 vdd.n9164 vdd.n9163 0.0225448
R15404 vdd.n9164 vdd.t1006 0.0225448
R15405 vdd.n9173 vdd.n9172 0.0225448
R15406 vdd.n9172 vdd.t78 0.0225448
R15407 vdd.n9157 vdd.n9133 0.0225448
R15408 vdd.t77 vdd.n9157 0.0225448
R15409 vdd.n9155 vdd.n9154 0.0225448
R15410 vdd.n9103 vdd.n9102 0.0225448
R15411 vdd.n9103 vdd.t1024 0.0225448
R15412 vdd.n9113 vdd.n9112 0.0225448
R15413 vdd.n9112 vdd.t785 0.0225448
R15414 vdd.n9115 vdd.n9092 0.0225448
R15415 vdd.t783 vdd.n9092 0.0225448
R15416 vdd.n9122 vdd.n9121 0.0225448
R15417 vdd.n9118 vdd.n9117 0.0225448
R15418 vdd.n9118 vdd.t430 0.0225448
R15419 vdd.n9127 vdd.n9126 0.0225448
R15420 vdd.n9126 vdd.t783 0.0225448
R15421 vdd.n9111 vdd.n9087 0.0225448
R15422 vdd.t785 vdd.n9111 0.0225448
R15423 vdd.n9109 vdd.n9108 0.0225448
R15424 vdd.n9196 vdd.n9195 0.0225448
R15425 vdd.n9196 vdd.t1270 0.0225448
R15426 vdd.n9206 vdd.n9205 0.0225448
R15427 vdd.n9205 vdd.t1267 0.0225448
R15428 vdd.n9208 vdd.n9185 0.0225448
R15429 vdd.t1268 vdd.n9185 0.0225448
R15430 vdd.n9215 vdd.n9214 0.0225448
R15431 vdd.n9211 vdd.n9210 0.0225448
R15432 vdd.n9211 vdd.t566 0.0225448
R15433 vdd.n9220 vdd.n9219 0.0225448
R15434 vdd.n9219 vdd.t1268 0.0225448
R15435 vdd.n9204 vdd.n9180 0.0225448
R15436 vdd.t1267 vdd.n9204 0.0225448
R15437 vdd.n9202 vdd.n9201 0.0225448
R15438 vdd.n9244 vdd.n9243 0.0225448
R15439 vdd.n9244 vdd.t675 0.0225448
R15440 vdd.n9254 vdd.n9253 0.0225448
R15441 vdd.n9253 vdd.t744 0.0225448
R15442 vdd.n9256 vdd.n9233 0.0225448
R15443 vdd.t745 vdd.n9233 0.0225448
R15444 vdd.n9263 vdd.n9262 0.0225448
R15445 vdd.n9259 vdd.n9258 0.0225448
R15446 vdd.n9259 vdd.t42 0.0225448
R15447 vdd.n9268 vdd.n9267 0.0225448
R15448 vdd.n9267 vdd.t745 0.0225448
R15449 vdd.n9252 vdd.n9228 0.0225448
R15450 vdd.t744 vdd.n9252 0.0225448
R15451 vdd.n9250 vdd.n9249 0.0225448
R15452 vdd.n9290 vdd.n9289 0.0225448
R15453 vdd.n9290 vdd.t547 0.0225448
R15454 vdd.n9300 vdd.n9299 0.0225448
R15455 vdd.n9299 vdd.t401 0.0225448
R15456 vdd.n9302 vdd.n9279 0.0225448
R15457 vdd.t399 vdd.n9279 0.0225448
R15458 vdd.n9309 vdd.n9308 0.0225448
R15459 vdd.n9305 vdd.n9304 0.0225448
R15460 vdd.n9305 vdd.t1302 0.0225448
R15461 vdd.n9314 vdd.n9313 0.0225448
R15462 vdd.n9313 vdd.t399 0.0225448
R15463 vdd.n9298 vdd.n9274 0.0225448
R15464 vdd.t401 vdd.n9298 0.0225448
R15465 vdd.n9296 vdd.n9295 0.0225448
R15466 vdd.n6800 vdd.n6799 0.0225448
R15467 vdd.n6799 vdd.t1362 0.0225448
R15468 vdd.n6802 vdd.n6788 0.0225448
R15469 vdd.t693 vdd.n6788 0.0225448
R15470 vdd.n6805 vdd.n6804 0.0225448
R15471 vdd.t691 vdd.n6805 0.0225448
R15472 vdd.n6820 vdd.n6819 0.0225448
R15473 vdd.n6817 vdd.n6777 0.0225448
R15474 vdd.t89 vdd.n6817 0.0225448
R15475 vdd.n6812 vdd.n6782 0.0225448
R15476 vdd.t691 vdd.n6782 0.0225448
R15477 vdd.n6808 vdd.n6807 0.0225448
R15478 vdd.n6807 vdd.t693 0.0225448
R15479 vdd.n6797 vdd.n6796 0.0225448
R15480 vdd.n9385 vdd.n9384 0.0225448
R15481 vdd.n9385 vdd.t523 0.0225448
R15482 vdd.n9395 vdd.n9394 0.0225448
R15483 vdd.n9394 vdd.t176 0.0225448
R15484 vdd.n9397 vdd.n9374 0.0225448
R15485 vdd.t177 vdd.n9374 0.0225448
R15486 vdd.n9404 vdd.n9403 0.0225448
R15487 vdd.n9400 vdd.n9399 0.0225448
R15488 vdd.n9400 vdd.t988 0.0225448
R15489 vdd.n9409 vdd.n9408 0.0225448
R15490 vdd.n9408 vdd.t177 0.0225448
R15491 vdd.n9393 vdd.n9369 0.0225448
R15492 vdd.t176 vdd.n9393 0.0225448
R15493 vdd.n9391 vdd.n9390 0.0225448
R15494 vdd.n9339 vdd.n9338 0.0225448
R15495 vdd.n9339 vdd.t1031 0.0225448
R15496 vdd.n9349 vdd.n9348 0.0225448
R15497 vdd.n9348 vdd.t1028 0.0225448
R15498 vdd.n9351 vdd.n9328 0.0225448
R15499 vdd.t1029 vdd.n9328 0.0225448
R15500 vdd.n9358 vdd.n9357 0.0225448
R15501 vdd.n9354 vdd.n9353 0.0225448
R15502 vdd.n9354 vdd.t627 0.0225448
R15503 vdd.n9363 vdd.n9362 0.0225448
R15504 vdd.n9362 vdd.t1029 0.0225448
R15505 vdd.n9347 vdd.n9323 0.0225448
R15506 vdd.t1028 vdd.n9347 0.0225448
R15507 vdd.n9345 vdd.n9344 0.0225448
R15508 vdd.n9432 vdd.n9431 0.0225448
R15509 vdd.n9432 vdd.t428 0.0225448
R15510 vdd.n9442 vdd.n9441 0.0225448
R15511 vdd.n9441 vdd.t546 0.0225448
R15512 vdd.n9444 vdd.n9421 0.0225448
R15513 vdd.t544 vdd.n9421 0.0225448
R15514 vdd.n9451 vdd.n9450 0.0225448
R15515 vdd.n9447 vdd.n9446 0.0225448
R15516 vdd.n9447 vdd.t601 0.0225448
R15517 vdd.n9456 vdd.n9455 0.0225448
R15518 vdd.n9455 vdd.t544 0.0225448
R15519 vdd.n9440 vdd.n9416 0.0225448
R15520 vdd.t546 vdd.n9440 0.0225448
R15521 vdd.n9438 vdd.n9437 0.0225448
R15522 vdd.n9480 vdd.n9479 0.0225448
R15523 vdd.n9480 vdd.t1191 0.0225448
R15524 vdd.n9490 vdd.n9489 0.0225448
R15525 vdd.n9489 vdd.t661 0.0225448
R15526 vdd.n9492 vdd.n9469 0.0225448
R15527 vdd.t662 vdd.n9469 0.0225448
R15528 vdd.n9499 vdd.n9498 0.0225448
R15529 vdd.n9495 vdd.n9494 0.0225448
R15530 vdd.n9495 vdd.t860 0.0225448
R15531 vdd.n9504 vdd.n9503 0.0225448
R15532 vdd.n9503 vdd.t662 0.0225448
R15533 vdd.n9488 vdd.n9464 0.0225448
R15534 vdd.t661 vdd.n9488 0.0225448
R15535 vdd.n9486 vdd.n9485 0.0225448
R15536 vdd.n9526 vdd.n9525 0.0225448
R15537 vdd.n9526 vdd.t76 0.0225448
R15538 vdd.n9536 vdd.n9535 0.0225448
R15539 vdd.n9535 vdd.t1518 0.0225448
R15540 vdd.n9538 vdd.n9515 0.0225448
R15541 vdd.t1519 vdd.n9515 0.0225448
R15542 vdd.n9545 vdd.n9544 0.0225448
R15543 vdd.n9541 vdd.n9540 0.0225448
R15544 vdd.n9541 vdd.t1041 0.0225448
R15545 vdd.n9550 vdd.n9549 0.0225448
R15546 vdd.n9549 vdd.t1519 0.0225448
R15547 vdd.n9534 vdd.n9510 0.0225448
R15548 vdd.t1518 vdd.n9534 0.0225448
R15549 vdd.n9532 vdd.n9531 0.0225448
R15550 vdd.n3686 vdd.n3685 0.0225448
R15551 vdd.n3686 vdd.t441 0.0225448
R15552 vdd.n3696 vdd.n3695 0.0225448
R15553 vdd.n3695 vdd.t474 0.0225448
R15554 vdd.n3698 vdd.n3675 0.0225448
R15555 vdd.t475 vdd.n3675 0.0225448
R15556 vdd.n3705 vdd.n3704 0.0225448
R15557 vdd.n3701 vdd.n3700 0.0225448
R15558 vdd.n3701 vdd.t1483 0.0225448
R15559 vdd.n3710 vdd.n3709 0.0225448
R15560 vdd.n3709 vdd.t475 0.0225448
R15561 vdd.n3694 vdd.n3670 0.0225448
R15562 vdd.t474 vdd.n3694 0.0225448
R15563 vdd.n3692 vdd.n3691 0.0225448
R15564 vdd.n3732 vdd.n3731 0.0225448
R15565 vdd.n3732 vdd.t234 0.0225448
R15566 vdd.n3742 vdd.n3741 0.0225448
R15567 vdd.n3741 vdd.t680 0.0225448
R15568 vdd.n3744 vdd.n3721 0.0225448
R15569 vdd.t681 vdd.n3721 0.0225448
R15570 vdd.n3751 vdd.n3750 0.0225448
R15571 vdd.n3747 vdd.n3746 0.0225448
R15572 vdd.n3747 vdd.t464 0.0225448
R15573 vdd.n3756 vdd.n3755 0.0225448
R15574 vdd.n3755 vdd.t681 0.0225448
R15575 vdd.n3740 vdd.n3716 0.0225448
R15576 vdd.t680 vdd.n3740 0.0225448
R15577 vdd.n3738 vdd.n3737 0.0225448
R15578 vdd.n3830 vdd.n3829 0.0225448
R15579 vdd.n3830 vdd.t503 0.0225448
R15580 vdd.n3840 vdd.n3839 0.0225448
R15581 vdd.n3839 vdd.t192 0.0225448
R15582 vdd.n3842 vdd.n3819 0.0225448
R15583 vdd.t193 vdd.n3819 0.0225448
R15584 vdd.n3849 vdd.n3848 0.0225448
R15585 vdd.n3845 vdd.n3844 0.0225448
R15586 vdd.n3845 vdd.t599 0.0225448
R15587 vdd.n3854 vdd.n3853 0.0225448
R15588 vdd.n3853 vdd.t193 0.0225448
R15589 vdd.n3838 vdd.n3814 0.0225448
R15590 vdd.t192 vdd.n3838 0.0225448
R15591 vdd.n3836 vdd.n3835 0.0225448
R15592 vdd.n3876 vdd.n3875 0.0225448
R15593 vdd.n3876 vdd.t136 0.0225448
R15594 vdd.n3886 vdd.n3885 0.0225448
R15595 vdd.n3885 vdd.t1279 0.0225448
R15596 vdd.n3888 vdd.n3865 0.0225448
R15597 vdd.t1280 vdd.n3865 0.0225448
R15598 vdd.n3895 vdd.n3894 0.0225448
R15599 vdd.n3891 vdd.n3890 0.0225448
R15600 vdd.n3891 vdd.t460 0.0225448
R15601 vdd.n3900 vdd.n3899 0.0225448
R15602 vdd.n3899 vdd.t1280 0.0225448
R15603 vdd.n3884 vdd.n3860 0.0225448
R15604 vdd.t1279 vdd.n3884 0.0225448
R15605 vdd.n3882 vdd.n3881 0.0225448
R15606 vdd.n3922 vdd.n3921 0.0225448
R15607 vdd.n3922 vdd.t611 0.0225448
R15608 vdd.n3932 vdd.n3931 0.0225448
R15609 vdd.n3931 vdd.t1132 0.0225448
R15610 vdd.n3934 vdd.n3911 0.0225448
R15611 vdd.t1133 vdd.n3911 0.0225448
R15612 vdd.n3941 vdd.n3940 0.0225448
R15613 vdd.n3937 vdd.n3936 0.0225448
R15614 vdd.n3937 vdd.t1057 0.0225448
R15615 vdd.n3946 vdd.n3945 0.0225448
R15616 vdd.n3945 vdd.t1133 0.0225448
R15617 vdd.n3930 vdd.n3906 0.0225448
R15618 vdd.t1132 vdd.n3930 0.0225448
R15619 vdd.n3928 vdd.n3927 0.0225448
R15620 vdd.n3968 vdd.n3967 0.0225448
R15621 vdd.n3968 vdd.t802 0.0225448
R15622 vdd.n3978 vdd.n3977 0.0225448
R15623 vdd.n3977 vdd.t1207 0.0225448
R15624 vdd.n3980 vdd.n3957 0.0225448
R15625 vdd.t1208 vdd.n3957 0.0225448
R15626 vdd.n3987 vdd.n3986 0.0225448
R15627 vdd.n3983 vdd.n3982 0.0225448
R15628 vdd.n3983 vdd.t603 0.0225448
R15629 vdd.n3992 vdd.n3991 0.0225448
R15630 vdd.n3991 vdd.t1208 0.0225448
R15631 vdd.n3976 vdd.n3952 0.0225448
R15632 vdd.t1207 vdd.n3976 0.0225448
R15633 vdd.n3974 vdd.n3973 0.0225448
R15634 vdd.n4066 vdd.n4065 0.0225448
R15635 vdd.n4066 vdd.t473 0.0225448
R15636 vdd.n4076 vdd.n4075 0.0225448
R15637 vdd.n4075 vdd.t1407 0.0225448
R15638 vdd.n4078 vdd.n4055 0.0225448
R15639 vdd.t1408 vdd.n4055 0.0225448
R15640 vdd.n4085 vdd.n4084 0.0225448
R15641 vdd.n4081 vdd.n4080 0.0225448
R15642 vdd.n4081 vdd.t468 0.0225448
R15643 vdd.n4090 vdd.n4089 0.0225448
R15644 vdd.n4089 vdd.t1408 0.0225448
R15645 vdd.n4074 vdd.n4050 0.0225448
R15646 vdd.t1407 vdd.n4074 0.0225448
R15647 vdd.n4072 vdd.n4071 0.0225448
R15648 vdd.n5524 vdd.n5523 0.0225448
R15649 vdd.n5524 vdd.t327 0.0225448
R15650 vdd.n5534 vdd.n5533 0.0225448
R15651 vdd.n5533 vdd.t759 0.0225448
R15652 vdd.n5536 vdd.n5513 0.0225448
R15653 vdd.t760 vdd.n5513 0.0225448
R15654 vdd.n5543 vdd.n5542 0.0225448
R15655 vdd.n5539 vdd.n5538 0.0225448
R15656 vdd.n5539 vdd.t556 0.0225448
R15657 vdd.n5548 vdd.n5547 0.0225448
R15658 vdd.n5547 vdd.t760 0.0225448
R15659 vdd.n5532 vdd.n5508 0.0225448
R15660 vdd.t759 vdd.n5532 0.0225448
R15661 vdd.n5530 vdd.n5529 0.0225448
R15662 vdd.n4114 vdd.n4113 0.0225448
R15663 vdd.n4123 vdd.n4122 0.0225448
R15664 vdd.n4122 vdd.t394 0.0225448
R15665 vdd.n4128 vdd.n4127 0.0225448
R15666 vdd.n4128 vdd.t393 0.0225448
R15667 vdd.n4131 vdd.n4103 0.0225448
R15668 vdd.n4131 vdd.t440 0.0225448
R15669 vdd.n4119 vdd.t203 0.0225448
R15670 vdd.t394 vdd.n4121 0.0225448
R15671 vdd.n4137 vdd.t393 0.0225448
R15672 vdd.n4135 vdd.n4134 0.0225448
R15673 vdd.n4138 vdd.n4137 0.0225448
R15674 vdd.n4121 vdd.n4098 0.0225448
R15675 vdd.n4119 vdd.n4118 0.0225448
R15676 vdd.n4160 vdd.n4159 0.0225448
R15677 vdd.n4169 vdd.n4168 0.0225448
R15678 vdd.n4168 vdd.t621 0.0225448
R15679 vdd.n4174 vdd.n4173 0.0225448
R15680 vdd.n4174 vdd.t623 0.0225448
R15681 vdd.n4177 vdd.n4149 0.0225448
R15682 vdd.n4177 vdd.t477 0.0225448
R15683 vdd.n4165 vdd.t554 0.0225448
R15684 vdd.t621 vdd.n4167 0.0225448
R15685 vdd.n4183 vdd.t623 0.0225448
R15686 vdd.n4181 vdd.n4180 0.0225448
R15687 vdd.n4184 vdd.n4183 0.0225448
R15688 vdd.n4167 vdd.n4144 0.0225448
R15689 vdd.n4165 vdd.n4164 0.0225448
R15690 vdd.n4257 vdd.n4256 0.0225448
R15691 vdd.n4266 vdd.n4265 0.0225448
R15692 vdd.n4265 vdd.t1183 0.0225448
R15693 vdd.n4271 vdd.n4270 0.0225448
R15694 vdd.n4271 vdd.t1185 0.0225448
R15695 vdd.n4274 vdd.n4246 0.0225448
R15696 vdd.n4274 vdd.t114 0.0225448
R15697 vdd.n4262 vdd.t1290 0.0225448
R15698 vdd.t1183 vdd.n4264 0.0225448
R15699 vdd.n4280 vdd.t1185 0.0225448
R15700 vdd.n4278 vdd.n4277 0.0225448
R15701 vdd.n4281 vdd.n4280 0.0225448
R15702 vdd.n4264 vdd.n4241 0.0225448
R15703 vdd.n4262 vdd.n4261 0.0225448
R15704 vdd.n4303 vdd.n4302 0.0225448
R15705 vdd.n4312 vdd.n4311 0.0225448
R15706 vdd.n4311 vdd.t419 0.0225448
R15707 vdd.n4317 vdd.n4316 0.0225448
R15708 vdd.n4317 vdd.t421 0.0225448
R15709 vdd.n4320 vdd.n4292 0.0225448
R15710 vdd.n4320 vdd.t810 0.0225448
R15711 vdd.n4308 vdd.t1316 0.0225448
R15712 vdd.t419 vdd.n4310 0.0225448
R15713 vdd.n4326 vdd.t421 0.0225448
R15714 vdd.n4324 vdd.n4323 0.0225448
R15715 vdd.n4327 vdd.n4326 0.0225448
R15716 vdd.n4310 vdd.n4287 0.0225448
R15717 vdd.n4308 vdd.n4307 0.0225448
R15718 vdd.n4349 vdd.n4348 0.0225448
R15719 vdd.n4358 vdd.n4357 0.0225448
R15720 vdd.n4357 vdd.t1424 0.0225448
R15721 vdd.n4363 vdd.n4362 0.0225448
R15722 vdd.n4363 vdd.t1426 0.0225448
R15723 vdd.n4366 vdd.n4338 0.0225448
R15724 vdd.n4366 vdd.t1427 0.0225448
R15725 vdd.n4354 vdd.t1055 0.0225448
R15726 vdd.t1424 vdd.n4356 0.0225448
R15727 vdd.n4372 vdd.t1426 0.0225448
R15728 vdd.n4370 vdd.n4369 0.0225448
R15729 vdd.n4373 vdd.n4372 0.0225448
R15730 vdd.n4356 vdd.n4333 0.0225448
R15731 vdd.n4354 vdd.n4353 0.0225448
R15732 vdd.n4395 vdd.n4394 0.0225448
R15733 vdd.n4404 vdd.n4403 0.0225448
R15734 vdd.n4403 vdd.t1435 0.0225448
R15735 vdd.n4409 vdd.n4408 0.0225448
R15736 vdd.n4409 vdd.t1437 0.0225448
R15737 vdd.n4412 vdd.n4384 0.0225448
R15738 vdd.n4412 vdd.t1225 0.0225448
R15739 vdd.n4400 vdd.t570 0.0225448
R15740 vdd.t1435 vdd.n4402 0.0225448
R15741 vdd.n4418 vdd.t1437 0.0225448
R15742 vdd.n4416 vdd.n4415 0.0225448
R15743 vdd.n4419 vdd.n4418 0.0225448
R15744 vdd.n4402 vdd.n4379 0.0225448
R15745 vdd.n4400 vdd.n4399 0.0225448
R15746 vdd.n4492 vdd.n4491 0.0225448
R15747 vdd.n4501 vdd.n4500 0.0225448
R15748 vdd.n4500 vdd.t1231 0.0225448
R15749 vdd.n4506 vdd.n4505 0.0225448
R15750 vdd.n4506 vdd.t1233 0.0225448
R15751 vdd.n4509 vdd.n4481 0.0225448
R15752 vdd.n4509 vdd.t951 0.0225448
R15753 vdd.n4497 vdd.t1045 0.0225448
R15754 vdd.t1231 vdd.n4499 0.0225448
R15755 vdd.n4515 vdd.t1233 0.0225448
R15756 vdd.n4513 vdd.n4512 0.0225448
R15757 vdd.n4516 vdd.n4515 0.0225448
R15758 vdd.n4499 vdd.n4476 0.0225448
R15759 vdd.n4497 vdd.n4496 0.0225448
R15760 vdd.n3641 vdd.n3640 0.0225448
R15761 vdd.n3650 vdd.n3649 0.0225448
R15762 vdd.n3649 vdd.t1034 0.0225448
R15763 vdd.n3655 vdd.n3654 0.0225448
R15764 vdd.n3655 vdd.t1036 0.0225448
R15765 vdd.n3658 vdd.n3630 0.0225448
R15766 vdd.n3658 vdd.t230 0.0225448
R15767 vdd.n3646 vdd.t560 0.0225448
R15768 vdd.t1034 vdd.n3648 0.0225448
R15769 vdd.n3664 vdd.t1036 0.0225448
R15770 vdd.n3662 vdd.n3661 0.0225448
R15771 vdd.n3665 vdd.n3664 0.0225448
R15772 vdd.n3648 vdd.n3625 0.0225448
R15773 vdd.n3646 vdd.n3645 0.0225448
R15774 vdd.n4536 vdd.n4535 0.0225448
R15775 vdd.n4545 vdd.n4544 0.0225448
R15776 vdd.n4544 vdd.t696 0.0225448
R15777 vdd.n4550 vdd.n4549 0.0225448
R15778 vdd.n4550 vdd.t698 0.0225448
R15779 vdd.n4553 vdd.n4525 0.0225448
R15780 vdd.n4553 vdd.t1148 0.0225448
R15781 vdd.n4541 vdd.t1000 0.0225448
R15782 vdd.t696 vdd.n4543 0.0225448
R15783 vdd.n4559 vdd.t698 0.0225448
R15784 vdd.n4557 vdd.n4556 0.0225448
R15785 vdd.n4560 vdd.n4559 0.0225448
R15786 vdd.n4543 vdd.n4520 0.0225448
R15787 vdd.n4541 vdd.n4540 0.0225448
R15788 vdd.n4581 vdd.n4580 0.0225448
R15789 vdd.n4590 vdd.n4589 0.0225448
R15790 vdd.n4589 vdd.t447 0.0225448
R15791 vdd.n4595 vdd.n4594 0.0225448
R15792 vdd.n4595 vdd.t446 0.0225448
R15793 vdd.n4598 vdd.n4570 0.0225448
R15794 vdd.n4598 vdd.t145 0.0225448
R15795 vdd.n4586 vdd.t174 0.0225448
R15796 vdd.t447 vdd.n4588 0.0225448
R15797 vdd.n4604 vdd.t446 0.0225448
R15798 vdd.n4602 vdd.n4601 0.0225448
R15799 vdd.n4605 vdd.n4604 0.0225448
R15800 vdd.n4588 vdd.n4565 0.0225448
R15801 vdd.n4586 vdd.n4585 0.0225448
R15802 vdd.n4631 vdd.n4630 0.0225448
R15803 vdd.n4640 vdd.n4639 0.0225448
R15804 vdd.n4639 vdd.t149 0.0225448
R15805 vdd.n4645 vdd.n4644 0.0225448
R15806 vdd.n4645 vdd.t151 0.0225448
R15807 vdd.n4648 vdd.n4620 0.0225448
R15808 vdd.n4648 vdd.t1178 0.0225448
R15809 vdd.n4636 vdd.t197 0.0225448
R15810 vdd.t149 vdd.n4638 0.0225448
R15811 vdd.n4654 vdd.t151 0.0225448
R15812 vdd.n4652 vdd.n4651 0.0225448
R15813 vdd.n4655 vdd.n4654 0.0225448
R15814 vdd.n4638 vdd.n4615 0.0225448
R15815 vdd.n4636 vdd.n4635 0.0225448
R15816 vdd.n4677 vdd.n4676 0.0225448
R15817 vdd.n4686 vdd.n4685 0.0225448
R15818 vdd.n4685 vdd.t668 0.0225448
R15819 vdd.n4691 vdd.n4690 0.0225448
R15820 vdd.n4691 vdd.t667 0.0225448
R15821 vdd.n4694 vdd.n4666 0.0225448
R15822 vdd.n4694 vdd.t670 0.0225448
R15823 vdd.n4682 vdd.t34 0.0225448
R15824 vdd.t668 vdd.n4684 0.0225448
R15825 vdd.n4700 vdd.t667 0.0225448
R15826 vdd.n4698 vdd.n4697 0.0225448
R15827 vdd.n4701 vdd.n4700 0.0225448
R15828 vdd.n4684 vdd.n4661 0.0225448
R15829 vdd.n4682 vdd.n4681 0.0225448
R15830 vdd.n4725 vdd.n4724 0.0225448
R15831 vdd.n4734 vdd.n4733 0.0225448
R15832 vdd.n4733 vdd.t470 0.0225448
R15833 vdd.n4739 vdd.n4738 0.0225448
R15834 vdd.n4739 vdd.t472 0.0225448
R15835 vdd.n4742 vdd.n4714 0.0225448
R15836 vdd.n4742 vdd.t1032 0.0225448
R15837 vdd.n4730 vdd.t1473 0.0225448
R15838 vdd.t470 vdd.n4732 0.0225448
R15839 vdd.n4748 vdd.t472 0.0225448
R15840 vdd.n4746 vdd.n4745 0.0225448
R15841 vdd.n4749 vdd.n4748 0.0225448
R15842 vdd.n4732 vdd.n4709 0.0225448
R15843 vdd.n4730 vdd.n4729 0.0225448
R15844 vdd.n4443 vdd.n4442 0.0225448
R15845 vdd.n4446 vdd.n4445 0.0225448
R15846 vdd.n4445 vdd.t1239 0.0225448
R15847 vdd.n4451 vdd.n4450 0.0225448
R15848 vdd.n4451 vdd.t1241 0.0225448
R15849 vdd.n4454 vdd.n4435 0.0225448
R15850 vdd.n4454 vdd.t455 0.0225448
R15851 vdd.n4467 vdd.t1457 0.0225448
R15852 vdd.n4465 vdd.t1239 0.0225448
R15853 vdd.n4460 vdd.t1241 0.0225448
R15854 vdd.n4458 vdd.n4457 0.0225448
R15855 vdd.n4461 vdd.n4460 0.0225448
R15856 vdd.n4465 vdd.n4464 0.0225448
R15857 vdd.n4468 vdd.n4467 0.0225448
R15858 vdd.n4772 vdd.n4771 0.0225448
R15859 vdd.n4781 vdd.n4780 0.0225448
R15860 vdd.n4780 vdd.t227 0.0225448
R15861 vdd.n4786 vdd.n4785 0.0225448
R15862 vdd.n4786 vdd.t229 0.0225448
R15863 vdd.n4789 vdd.n4761 0.0225448
R15864 vdd.n4789 vdd.t72 0.0225448
R15865 vdd.n4777 vdd.t827 0.0225448
R15866 vdd.t227 vdd.n4779 0.0225448
R15867 vdd.n4795 vdd.t229 0.0225448
R15868 vdd.n4793 vdd.n4792 0.0225448
R15869 vdd.n4796 vdd.n4795 0.0225448
R15870 vdd.n4779 vdd.n4756 0.0225448
R15871 vdd.n4777 vdd.n4776 0.0225448
R15872 vdd.n4817 vdd.n4816 0.0225448
R15873 vdd.n4826 vdd.n4825 0.0225448
R15874 vdd.n4825 vdd.t365 0.0225448
R15875 vdd.n4831 vdd.n4830 0.0225448
R15876 vdd.n4831 vdd.t367 0.0225448
R15877 vdd.n4834 vdd.n4806 0.0225448
R15878 vdd.n4834 vdd.t1256 0.0225448
R15879 vdd.n4822 vdd.t52 0.0225448
R15880 vdd.t365 vdd.n4824 0.0225448
R15881 vdd.n4840 vdd.t367 0.0225448
R15882 vdd.n4838 vdd.n4837 0.0225448
R15883 vdd.n4841 vdd.n4840 0.0225448
R15884 vdd.n4824 vdd.n4801 0.0225448
R15885 vdd.n4822 vdd.n4821 0.0225448
R15886 vdd.n4863 vdd.n4862 0.0225448
R15887 vdd.n4872 vdd.n4871 0.0225448
R15888 vdd.n4871 vdd.t414 0.0225448
R15889 vdd.n4877 vdd.n4876 0.0225448
R15890 vdd.n4877 vdd.t416 0.0225448
R15891 vdd.n4880 vdd.n4852 0.0225448
R15892 vdd.n4880 vdd.t411 0.0225448
R15893 vdd.n4868 vdd.t1371 0.0225448
R15894 vdd.t414 vdd.n4870 0.0225448
R15895 vdd.n4886 vdd.t416 0.0225448
R15896 vdd.n4884 vdd.n4883 0.0225448
R15897 vdd.n4887 vdd.n4886 0.0225448
R15898 vdd.n4870 vdd.n4847 0.0225448
R15899 vdd.n4868 vdd.n4867 0.0225448
R15900 vdd.n4914 vdd.n4913 0.0225448
R15901 vdd.n4923 vdd.n4922 0.0225448
R15902 vdd.n4922 vdd.t1227 0.0225448
R15903 vdd.n4928 vdd.n4927 0.0225448
R15904 vdd.n4928 vdd.t1229 0.0225448
R15905 vdd.n4931 vdd.n4903 0.0225448
R15906 vdd.n4931 vdd.t1090 0.0225448
R15907 vdd.n4919 vdd.t1487 0.0225448
R15908 vdd.t1227 vdd.n4921 0.0225448
R15909 vdd.n4937 vdd.t1229 0.0225448
R15910 vdd.n4935 vdd.n4934 0.0225448
R15911 vdd.n4938 vdd.n4937 0.0225448
R15912 vdd.n4921 vdd.n4898 0.0225448
R15913 vdd.n4919 vdd.n4918 0.0225448
R15914 vdd.n4960 vdd.n4959 0.0225448
R15915 vdd.n4969 vdd.n4968 0.0225448
R15916 vdd.n4968 vdd.t510 0.0225448
R15917 vdd.n4974 vdd.n4973 0.0225448
R15918 vdd.n4974 vdd.t512 0.0225448
R15919 vdd.n4977 vdd.n4949 0.0225448
R15920 vdd.n4977 vdd.t1165 0.0225448
R15921 vdd.n4965 vdd.t858 0.0225448
R15922 vdd.t510 vdd.n4967 0.0225448
R15923 vdd.n4983 vdd.t512 0.0225448
R15924 vdd.n4981 vdd.n4980 0.0225448
R15925 vdd.n4984 vdd.n4983 0.0225448
R15926 vdd.n4967 vdd.n4944 0.0225448
R15927 vdd.n4965 vdd.n4964 0.0225448
R15928 vdd.n5008 vdd.n5007 0.0225448
R15929 vdd.n5017 vdd.n5016 0.0225448
R15930 vdd.n5016 vdd.t1099 0.0225448
R15931 vdd.n5022 vdd.n5021 0.0225448
R15932 vdd.n5022 vdd.t1101 0.0225448
R15933 vdd.n5025 vdd.n4997 0.0225448
R15934 vdd.n5025 vdd.t308 0.0225448
R15935 vdd.n5013 vdd.t1300 0.0225448
R15936 vdd.t1099 vdd.n5015 0.0225448
R15937 vdd.n5031 vdd.t1101 0.0225448
R15938 vdd.n5029 vdd.n5028 0.0225448
R15939 vdd.n5032 vdd.n5031 0.0225448
R15940 vdd.n5015 vdd.n4992 0.0225448
R15941 vdd.n5013 vdd.n5012 0.0225448
R15942 vdd.n5054 vdd.n5053 0.0225448
R15943 vdd.n5063 vdd.n5062 0.0225448
R15944 vdd.n5062 vdd.t1167 0.0225448
R15945 vdd.n5068 vdd.n5067 0.0225448
R15946 vdd.n5068 vdd.t1166 0.0225448
R15947 vdd.n5071 vdd.n5043 0.0225448
R15948 vdd.n5071 vdd.t1412 0.0225448
R15949 vdd.n5059 vdd.t1010 0.0225448
R15950 vdd.t1167 vdd.n5061 0.0225448
R15951 vdd.n5077 vdd.t1166 0.0225448
R15952 vdd.n5075 vdd.n5074 0.0225448
R15953 vdd.n5078 vdd.n5077 0.0225448
R15954 vdd.n5061 vdd.n5038 0.0225448
R15955 vdd.n5059 vdd.n5058 0.0225448
R15956 vdd.n5099 vdd.n5098 0.0225448
R15957 vdd.n5108 vdd.n5107 0.0225448
R15958 vdd.n5107 vdd.t107 0.0225448
R15959 vdd.n5113 vdd.n5112 0.0225448
R15960 vdd.n5113 vdd.t109 0.0225448
R15961 vdd.n5116 vdd.n5088 0.0225448
R15962 vdd.n5116 vdd.t607 0.0225448
R15963 vdd.n5104 vdd.t50 0.0225448
R15964 vdd.t107 vdd.n5106 0.0225448
R15965 vdd.n5122 vdd.t109 0.0225448
R15966 vdd.n5120 vdd.n5119 0.0225448
R15967 vdd.n5123 vdd.n5122 0.0225448
R15968 vdd.n5106 vdd.n5083 0.0225448
R15969 vdd.n5104 vdd.n5103 0.0225448
R15970 vdd.n5149 vdd.n5148 0.0225448
R15971 vdd.n5158 vdd.n5157 0.0225448
R15972 vdd.n5157 vdd.t344 0.0225448
R15973 vdd.n5163 vdd.n5162 0.0225448
R15974 vdd.n5163 vdd.t346 0.0225448
R15975 vdd.n5166 vdd.n5138 0.0225448
R15976 vdd.n5166 vdd.t191 0.0225448
R15977 vdd.n5154 vdd.t1043 0.0225448
R15978 vdd.t344 vdd.n5156 0.0225448
R15979 vdd.n5172 vdd.t346 0.0225448
R15980 vdd.n5170 vdd.n5169 0.0225448
R15981 vdd.n5173 vdd.n5172 0.0225448
R15982 vdd.n5156 vdd.n5133 0.0225448
R15983 vdd.n5154 vdd.n5153 0.0225448
R15984 vdd.n5195 vdd.n5194 0.0225448
R15985 vdd.n5204 vdd.n5203 0.0225448
R15986 vdd.n5203 vdd.t322 0.0225448
R15987 vdd.n5209 vdd.n5208 0.0225448
R15988 vdd.n5209 vdd.t321 0.0225448
R15989 vdd.n5212 vdd.n5184 0.0225448
R15990 vdd.n5212 vdd.t1278 0.0225448
R15991 vdd.n5200 vdd.t942 0.0225448
R15992 vdd.t322 vdd.n5202 0.0225448
R15993 vdd.n5218 vdd.t321 0.0225448
R15994 vdd.n5216 vdd.n5215 0.0225448
R15995 vdd.n5219 vdd.n5218 0.0225448
R15996 vdd.n5202 vdd.n5179 0.0225448
R15997 vdd.n5200 vdd.n5199 0.0225448
R15998 vdd.n5243 vdd.n5242 0.0225448
R15999 vdd.n5252 vdd.n5251 0.0225448
R16000 vdd.n5251 vdd.t700 0.0225448
R16001 vdd.n5257 vdd.n5256 0.0225448
R16002 vdd.n5257 vdd.t699 0.0225448
R16003 vdd.n5260 vdd.n5232 0.0225448
R16004 vdd.n5260 vdd.t537 0.0225448
R16005 vdd.n5248 vdd.t1304 0.0225448
R16006 vdd.t700 vdd.n5250 0.0225448
R16007 vdd.n5266 vdd.t699 0.0225448
R16008 vdd.n5264 vdd.n5263 0.0225448
R16009 vdd.n5267 vdd.n5266 0.0225448
R16010 vdd.n5250 vdd.n5227 0.0225448
R16011 vdd.n5248 vdd.n5247 0.0225448
R16012 vdd.n4208 vdd.n4207 0.0225448
R16013 vdd.n4211 vdd.n4210 0.0225448
R16014 vdd.n4210 vdd.t710 0.0225448
R16015 vdd.n4216 vdd.n4215 0.0225448
R16016 vdd.n4216 vdd.t712 0.0225448
R16017 vdd.n4219 vdd.n4200 0.0225448
R16018 vdd.n4219 vdd.t1067 0.0225448
R16019 vdd.n4232 vdd.t1455 0.0225448
R16020 vdd.n4230 vdd.t710 0.0225448
R16021 vdd.n4225 vdd.t712 0.0225448
R16022 vdd.n4223 vdd.n4222 0.0225448
R16023 vdd.n4226 vdd.n4225 0.0225448
R16024 vdd.n4230 vdd.n4229 0.0225448
R16025 vdd.n4233 vdd.n4232 0.0225448
R16026 vdd.n5290 vdd.n5289 0.0225448
R16027 vdd.n5299 vdd.n5298 0.0225448
R16028 vdd.n5298 vdd.t1109 0.0225448
R16029 vdd.n5304 vdd.n5303 0.0225448
R16030 vdd.n5304 vdd.t1111 0.0225448
R16031 vdd.n5307 vdd.n5279 0.0225448
R16032 vdd.n5307 vdd.t888 0.0225448
R16033 vdd.n5295 vdd.t844 0.0225448
R16034 vdd.t1109 vdd.n5297 0.0225448
R16035 vdd.n5313 vdd.t1111 0.0225448
R16036 vdd.n5311 vdd.n5310 0.0225448
R16037 vdd.n5314 vdd.n5313 0.0225448
R16038 vdd.n5297 vdd.n5274 0.0225448
R16039 vdd.n5295 vdd.n5294 0.0225448
R16040 vdd.n5335 vdd.n5334 0.0225448
R16041 vdd.n5344 vdd.n5343 0.0225448
R16042 vdd.n5343 vdd.t1503 0.0225448
R16043 vdd.n5349 vdd.n5348 0.0225448
R16044 vdd.n5349 vdd.t1505 0.0225448
R16045 vdd.n5352 vdd.n5324 0.0225448
R16046 vdd.n5352 vdd.t660 0.0225448
R16047 vdd.n5340 vdd.t172 0.0225448
R16048 vdd.t1503 vdd.n5342 0.0225448
R16049 vdd.n5358 vdd.t1505 0.0225448
R16050 vdd.n5356 vdd.n5355 0.0225448
R16051 vdd.n5359 vdd.n5358 0.0225448
R16052 vdd.n5342 vdd.n5319 0.0225448
R16053 vdd.n5340 vdd.n5339 0.0225448
R16054 vdd.n5385 vdd.n5384 0.0225448
R16055 vdd.n5394 vdd.n5393 0.0225448
R16056 vdd.n5393 vdd.t719 0.0225448
R16057 vdd.n5399 vdd.n5398 0.0225448
R16058 vdd.n5399 vdd.t718 0.0225448
R16059 vdd.n5402 vdd.n5374 0.0225448
R16060 vdd.n5402 vdd.t63 0.0225448
R16061 vdd.n5390 vdd.t456 0.0225448
R16062 vdd.t719 vdd.n5392 0.0225448
R16063 vdd.n5408 vdd.t718 0.0225448
R16064 vdd.n5406 vdd.n5405 0.0225448
R16065 vdd.n5409 vdd.n5408 0.0225448
R16066 vdd.n5392 vdd.n5369 0.0225448
R16067 vdd.n5390 vdd.n5389 0.0225448
R16068 vdd.n5431 vdd.n5430 0.0225448
R16069 vdd.n5440 vdd.n5439 0.0225448
R16070 vdd.n5439 vdd.t500 0.0225448
R16071 vdd.n5445 vdd.n5444 0.0225448
R16072 vdd.n5445 vdd.t499 0.0225448
R16073 vdd.n5448 vdd.n5420 0.0225448
R16074 vdd.n5448 vdd.t1411 0.0225448
R16075 vdd.n5436 vdd.t1012 0.0225448
R16076 vdd.t500 vdd.n5438 0.0225448
R16077 vdd.n5454 vdd.t499 0.0225448
R16078 vdd.n5452 vdd.n5451 0.0225448
R16079 vdd.n5455 vdd.n5454 0.0225448
R16080 vdd.n5438 vdd.n5415 0.0225448
R16081 vdd.n5436 vdd.n5435 0.0225448
R16082 vdd.n5479 vdd.n5478 0.0225448
R16083 vdd.n5488 vdd.n5487 0.0225448
R16084 vdd.n5487 vdd.t504 0.0225448
R16085 vdd.n5493 vdd.n5492 0.0225448
R16086 vdd.n5493 vdd.t506 0.0225448
R16087 vdd.n5496 vdd.n5468 0.0225448
R16088 vdd.n5496 vdd.t269 0.0225448
R16089 vdd.n5484 vdd.t1051 0.0225448
R16090 vdd.t504 vdd.n5486 0.0225448
R16091 vdd.n5502 vdd.t506 0.0225448
R16092 vdd.n5500 vdd.n5499 0.0225448
R16093 vdd.n5503 vdd.n5502 0.0225448
R16094 vdd.n5486 vdd.n5463 0.0225448
R16095 vdd.n5484 vdd.n5483 0.0225448
R16096 vdd.n5617 vdd.n5616 0.0225448
R16097 vdd.n5617 vdd.t716 0.0225448
R16098 vdd.n5627 vdd.n5626 0.0225448
R16099 vdd.n5626 vdd.t713 0.0225448
R16100 vdd.n5629 vdd.n5606 0.0225448
R16101 vdd.t714 vdd.n5606 0.0225448
R16102 vdd.n5636 vdd.n5635 0.0225448
R16103 vdd.n5632 vdd.n5631 0.0225448
R16104 vdd.n5632 vdd.t906 0.0225448
R16105 vdd.n5641 vdd.n5640 0.0225448
R16106 vdd.n5640 vdd.t714 0.0225448
R16107 vdd.n5625 vdd.n5601 0.0225448
R16108 vdd.t713 vdd.n5625 0.0225448
R16109 vdd.n5623 vdd.n5622 0.0225448
R16110 vdd.n5571 vdd.n5570 0.0225448
R16111 vdd.n5571 vdd.t1237 0.0225448
R16112 vdd.n5581 vdd.n5580 0.0225448
R16113 vdd.n5580 vdd.t185 0.0225448
R16114 vdd.n5583 vdd.n5560 0.0225448
R16115 vdd.t186 vdd.n5560 0.0225448
R16116 vdd.n5590 vdd.n5589 0.0225448
R16117 vdd.n5586 vdd.n5585 0.0225448
R16118 vdd.n5586 vdd.t164 0.0225448
R16119 vdd.n5595 vdd.n5594 0.0225448
R16120 vdd.n5594 vdd.t186 0.0225448
R16121 vdd.n5579 vdd.n5555 0.0225448
R16122 vdd.t185 vdd.n5579 0.0225448
R16123 vdd.n5577 vdd.n5576 0.0225448
R16124 vdd.n5664 vdd.n5663 0.0225448
R16125 vdd.n5664 vdd.t144 0.0225448
R16126 vdd.n5674 vdd.n5673 0.0225448
R16127 vdd.n5673 vdd.t396 0.0225448
R16128 vdd.n5676 vdd.n5653 0.0225448
R16129 vdd.t397 vdd.n5653 0.0225448
R16130 vdd.n5683 vdd.n5682 0.0225448
R16131 vdd.n5679 vdd.n5678 0.0225448
R16132 vdd.n5679 vdd.t595 0.0225448
R16133 vdd.n5688 vdd.n5687 0.0225448
R16134 vdd.n5687 vdd.t397 0.0225448
R16135 vdd.n5672 vdd.n5648 0.0225448
R16136 vdd.t396 vdd.n5672 0.0225448
R16137 vdd.n5670 vdd.n5669 0.0225448
R16138 vdd.n5712 vdd.n5711 0.0225448
R16139 vdd.n5712 vdd.t924 0.0225448
R16140 vdd.n5722 vdd.n5721 0.0225448
R16141 vdd.n5721 vdd.t1214 0.0225448
R16142 vdd.n5724 vdd.n5701 0.0225448
R16143 vdd.t1215 vdd.n5701 0.0225448
R16144 vdd.n5731 vdd.n5730 0.0225448
R16145 vdd.n5727 vdd.n5726 0.0225448
R16146 vdd.n5727 vdd.t990 0.0225448
R16147 vdd.n5736 vdd.n5735 0.0225448
R16148 vdd.n5735 vdd.t1215 0.0225448
R16149 vdd.n5720 vdd.n5696 0.0225448
R16150 vdd.t1214 vdd.n5720 0.0225448
R16151 vdd.n5718 vdd.n5717 0.0225448
R16152 vdd.n5758 vdd.n5757 0.0225448
R16153 vdd.n5758 vdd.t424 0.0225448
R16154 vdd.n5768 vdd.n5767 0.0225448
R16155 vdd.n5767 vdd.t583 0.0225448
R16156 vdd.n5770 vdd.n5747 0.0225448
R16157 vdd.t581 vdd.n5747 0.0225448
R16158 vdd.n5777 vdd.n5776 0.0225448
R16159 vdd.n5773 vdd.n5772 0.0225448
R16160 vdd.n5773 vdd.t13 0.0225448
R16161 vdd.n5782 vdd.n5781 0.0225448
R16162 vdd.n5781 vdd.t581 0.0225448
R16163 vdd.n5766 vdd.n5742 0.0225448
R16164 vdd.t583 vdd.n5766 0.0225448
R16165 vdd.n5764 vdd.n5763 0.0225448
R16166 vdd.n4022 vdd.n4021 0.0225448
R16167 vdd.n4021 vdd.t1422 0.0225448
R16168 vdd.n4024 vdd.n4010 0.0225448
R16169 vdd.t1517 vdd.n4010 0.0225448
R16170 vdd.n4027 vdd.n4026 0.0225448
R16171 vdd.t1515 vdd.n4027 0.0225448
R16172 vdd.n4042 vdd.n4041 0.0225448
R16173 vdd.n4039 vdd.n3999 0.0225448
R16174 vdd.t99 vdd.n4039 0.0225448
R16175 vdd.n4034 vdd.n4004 0.0225448
R16176 vdd.t1515 vdd.n4004 0.0225448
R16177 vdd.n4030 vdd.n4029 0.0225448
R16178 vdd.n4029 vdd.t1517 0.0225448
R16179 vdd.n4019 vdd.n4018 0.0225448
R16180 vdd.n5900 vdd.n5899 0.0225448
R16181 vdd.n5900 vdd.t23 0.0225448
R16182 vdd.n5910 vdd.n5909 0.0225448
R16183 vdd.n5909 vdd.t330 0.0225448
R16184 vdd.n5912 vdd.n5889 0.0225448
R16185 vdd.t328 vdd.n5889 0.0225448
R16186 vdd.n5919 vdd.n5918 0.0225448
R16187 vdd.n5915 vdd.n5914 0.0225448
R16188 vdd.n5915 vdd.t866 0.0225448
R16189 vdd.n5924 vdd.n5923 0.0225448
R16190 vdd.n5923 vdd.t328 0.0225448
R16191 vdd.n5908 vdd.n5884 0.0225448
R16192 vdd.t330 vdd.n5908 0.0225448
R16193 vdd.n5906 vdd.n5905 0.0225448
R16194 vdd.n5853 vdd.n5852 0.0225448
R16195 vdd.n5853 vdd.t786 0.0225448
R16196 vdd.n5863 vdd.n5862 0.0225448
R16197 vdd.n5862 vdd.t1527 0.0225448
R16198 vdd.n5865 vdd.n5842 0.0225448
R16199 vdd.t1528 vdd.n5842 0.0225448
R16200 vdd.n5872 vdd.n5871 0.0225448
R16201 vdd.n5868 vdd.n5867 0.0225448
R16202 vdd.n5868 vdd.t767 0.0225448
R16203 vdd.n5877 vdd.n5876 0.0225448
R16204 vdd.n5876 vdd.t1528 0.0225448
R16205 vdd.n5861 vdd.n5837 0.0225448
R16206 vdd.t1527 vdd.n5861 0.0225448
R16207 vdd.n5859 vdd.n5858 0.0225448
R16208 vdd.n5807 vdd.n5806 0.0225448
R16209 vdd.n5807 vdd.t928 0.0225448
R16210 vdd.n5817 vdd.n5816 0.0225448
R16211 vdd.n5816 vdd.t777 0.0225448
R16212 vdd.n5819 vdd.n5796 0.0225448
R16213 vdd.t778 vdd.n5796 0.0225448
R16214 vdd.n5826 vdd.n5825 0.0225448
R16215 vdd.n5822 vdd.n5821 0.0225448
R16216 vdd.n5822 vdd.t1373 0.0225448
R16217 vdd.n5831 vdd.n5830 0.0225448
R16218 vdd.n5830 vdd.t778 0.0225448
R16219 vdd.n5815 vdd.n5791 0.0225448
R16220 vdd.t777 vdd.n5815 0.0225448
R16221 vdd.n5813 vdd.n5812 0.0225448
R16222 vdd.n5947 vdd.n5946 0.0225448
R16223 vdd.n5947 vdd.t679 0.0225448
R16224 vdd.n5957 vdd.n5956 0.0225448
R16225 vdd.n5956 vdd.t676 0.0225448
R16226 vdd.n5959 vdd.n5936 0.0225448
R16227 vdd.t677 vdd.n5936 0.0225448
R16228 vdd.n5966 vdd.n5965 0.0225448
R16229 vdd.n5962 vdd.n5961 0.0225448
R16230 vdd.n5962 vdd.t1479 0.0225448
R16231 vdd.n5971 vdd.n5970 0.0225448
R16232 vdd.n5970 vdd.t677 0.0225448
R16233 vdd.n5955 vdd.n5931 0.0225448
R16234 vdd.t676 vdd.n5955 0.0225448
R16235 vdd.n5953 vdd.n5952 0.0225448
R16236 vdd.n5995 vdd.n5994 0.0225448
R16237 vdd.n5995 vdd.t1258 0.0225448
R16238 vdd.n6005 vdd.n6004 0.0225448
R16239 vdd.n6004 vdd.t1192 0.0225448
R16240 vdd.n6007 vdd.n5984 0.0225448
R16241 vdd.t1193 vdd.n5984 0.0225448
R16242 vdd.n6014 vdd.n6013 0.0225448
R16243 vdd.n6010 vdd.n6009 0.0225448
R16244 vdd.n6010 vdd.t1002 0.0225448
R16245 vdd.n6019 vdd.n6018 0.0225448
R16246 vdd.n6018 vdd.t1193 0.0225448
R16247 vdd.n6003 vdd.n5979 0.0225448
R16248 vdd.t1192 vdd.n6003 0.0225448
R16249 vdd.n6001 vdd.n6000 0.0225448
R16250 vdd.n6041 vdd.n6040 0.0225448
R16251 vdd.n6041 vdd.t429 0.0225448
R16252 vdd.n6051 vdd.n6050 0.0225448
R16253 vdd.n6050 vdd.t2 0.0225448
R16254 vdd.n6053 vdd.n6030 0.0225448
R16255 vdd.t0 vdd.n6030 0.0225448
R16256 vdd.n6060 vdd.n6059 0.0225448
R16257 vdd.n6056 vdd.n6055 0.0225448
R16258 vdd.n6056 vdd.t1489 0.0225448
R16259 vdd.n6065 vdd.n6064 0.0225448
R16260 vdd.n6064 vdd.t0 0.0225448
R16261 vdd.n6049 vdd.n6025 0.0225448
R16262 vdd.t2 vdd.n6049 0.0225448
R16263 vdd.n6047 vdd.n6046 0.0225448
R16264 vdd.n6135 vdd.n6134 0.0225448
R16265 vdd.n6135 vdd.t305 0.0225448
R16266 vdd.n6145 vdd.n6144 0.0225448
R16267 vdd.n6144 vdd.t631 0.0225448
R16268 vdd.n6147 vdd.n6124 0.0225448
R16269 vdd.t632 vdd.n6124 0.0225448
R16270 vdd.n6154 vdd.n6153 0.0225448
R16271 vdd.n6150 vdd.n6149 0.0225448
R16272 vdd.n6150 vdd.t969 0.0225448
R16273 vdd.n6159 vdd.n6158 0.0225448
R16274 vdd.n6158 vdd.t632 0.0225448
R16275 vdd.n6143 vdd.n6119 0.0225448
R16276 vdd.t631 vdd.n6143 0.0225448
R16277 vdd.n6141 vdd.n6140 0.0225448
R16278 vdd.n6089 vdd.n6088 0.0225448
R16279 vdd.n6089 vdd.t671 0.0225448
R16280 vdd.n6099 vdd.n6098 0.0225448
R16281 vdd.n6098 vdd.t1206 0.0225448
R16282 vdd.n6101 vdd.n6078 0.0225448
R16283 vdd.t1204 vdd.n6078 0.0225448
R16284 vdd.n6108 vdd.n6107 0.0225448
R16285 vdd.n6104 vdd.n6103 0.0225448
R16286 vdd.n6104 vdd.t434 0.0225448
R16287 vdd.n6113 vdd.n6112 0.0225448
R16288 vdd.n6112 vdd.t1204 0.0225448
R16289 vdd.n6097 vdd.n6073 0.0225448
R16290 vdd.t1206 vdd.n6097 0.0225448
R16291 vdd.n6095 vdd.n6094 0.0225448
R16292 vdd.n6182 vdd.n6181 0.0225448
R16293 vdd.n6182 vdd.t387 0.0225448
R16294 vdd.n6192 vdd.n6191 0.0225448
R16295 vdd.n6191 vdd.t1157 0.0225448
R16296 vdd.n6194 vdd.n6171 0.0225448
R16297 vdd.t1158 vdd.n6171 0.0225448
R16298 vdd.n6201 vdd.n6200 0.0225448
R16299 vdd.n6197 vdd.n6196 0.0225448
R16300 vdd.n6197 vdd.t1336 0.0225448
R16301 vdd.n6206 vdd.n6205 0.0225448
R16302 vdd.n6205 vdd.t1158 0.0225448
R16303 vdd.n6190 vdd.n6166 0.0225448
R16304 vdd.t1157 vdd.n6190 0.0225448
R16305 vdd.n6188 vdd.n6187 0.0225448
R16306 vdd.n6230 vdd.n6229 0.0225448
R16307 vdd.n6230 vdd.t246 0.0225448
R16308 vdd.n6240 vdd.n6239 0.0225448
R16309 vdd.n6239 vdd.t1403 0.0225448
R16310 vdd.n6242 vdd.n6219 0.0225448
R16311 vdd.t1404 vdd.n6219 0.0225448
R16312 vdd.n6249 vdd.n6248 0.0225448
R16313 vdd.n6245 vdd.n6244 0.0225448
R16314 vdd.n6245 vdd.t32 0.0225448
R16315 vdd.n6254 vdd.n6253 0.0225448
R16316 vdd.n6253 vdd.t1404 0.0225448
R16317 vdd.n6238 vdd.n6214 0.0225448
R16318 vdd.t1403 vdd.n6238 0.0225448
R16319 vdd.n6236 vdd.n6235 0.0225448
R16320 vdd.n6276 vdd.n6275 0.0225448
R16321 vdd.n6276 vdd.t1026 0.0225448
R16322 vdd.n6286 vdd.n6285 0.0225448
R16323 vdd.n6285 vdd.t944 0.0225448
R16324 vdd.n6288 vdd.n6265 0.0225448
R16325 vdd.t945 vdd.n6265 0.0225448
R16326 vdd.n6295 vdd.n6294 0.0225448
R16327 vdd.n6291 vdd.n6290 0.0225448
R16328 vdd.n6291 vdd.t496 0.0225448
R16329 vdd.n6300 vdd.n6299 0.0225448
R16330 vdd.n6299 vdd.t945 0.0225448
R16331 vdd.n6284 vdd.n6260 0.0225448
R16332 vdd.t944 vdd.n6284 0.0225448
R16333 vdd.n6282 vdd.n6281 0.0225448
R16334 vdd.n3786 vdd.n3785 0.0225448
R16335 vdd.n3785 vdd.t724 0.0225448
R16336 vdd.n3788 vdd.n3774 0.0225448
R16337 vdd.t721 vdd.n3774 0.0225448
R16338 vdd.n3791 vdd.n3790 0.0225448
R16339 vdd.t722 vdd.n3791 0.0225448
R16340 vdd.n3806 vdd.n3805 0.0225448
R16341 vdd.n3803 vdd.n3763 0.0225448
R16342 vdd.t93 vdd.n3803 0.0225448
R16343 vdd.n3798 vdd.n3768 0.0225448
R16344 vdd.t722 vdd.n3768 0.0225448
R16345 vdd.n3794 vdd.n3793 0.0225448
R16346 vdd.n3793 vdd.t721 0.0225448
R16347 vdd.n3783 vdd.n3782 0.0225448
R16348 vdd.n6371 vdd.n6370 0.0225448
R16349 vdd.n6371 vdd.t20 0.0225448
R16350 vdd.n6381 vdd.n6380 0.0225448
R16351 vdd.n6380 vdd.t17 0.0225448
R16352 vdd.n6383 vdd.n6360 0.0225448
R16353 vdd.t18 vdd.n6360 0.0225448
R16354 vdd.n6390 vdd.n6389 0.0225448
R16355 vdd.n6386 vdd.n6385 0.0225448
R16356 vdd.n6386 vdd.t868 0.0225448
R16357 vdd.n6395 vdd.n6394 0.0225448
R16358 vdd.n6394 vdd.t18 0.0225448
R16359 vdd.n6379 vdd.n6355 0.0225448
R16360 vdd.t17 vdd.n6379 0.0225448
R16361 vdd.n6377 vdd.n6376 0.0225448
R16362 vdd.n6325 vdd.n6324 0.0225448
R16363 vdd.n6325 vdd.t331 0.0225448
R16364 vdd.n6335 vdd.n6334 0.0225448
R16365 vdd.n6334 vdd.t749 0.0225448
R16366 vdd.n6337 vdd.n6314 0.0225448
R16367 vdd.t750 vdd.n6314 0.0225448
R16368 vdd.n6344 vdd.n6343 0.0225448
R16369 vdd.n6340 vdd.n6339 0.0225448
R16370 vdd.n6340 vdd.t432 0.0225448
R16371 vdd.n6349 vdd.n6348 0.0225448
R16372 vdd.n6348 vdd.t750 0.0225448
R16373 vdd.n6333 vdd.n6309 0.0225448
R16374 vdd.t749 vdd.n6333 0.0225448
R16375 vdd.n6331 vdd.n6330 0.0225448
R16376 vdd.n6418 vdd.n6417 0.0225448
R16377 vdd.n6418 vdd.t615 0.0225448
R16378 vdd.n6428 vdd.n6427 0.0225448
R16379 vdd.n6427 vdd.t686 0.0225448
R16380 vdd.n6430 vdd.n6407 0.0225448
R16381 vdd.t684 vdd.n6407 0.0225448
R16382 vdd.n6437 vdd.n6436 0.0225448
R16383 vdd.n6433 vdd.n6432 0.0225448
R16384 vdd.n6433 vdd.t1053 0.0225448
R16385 vdd.n6442 vdd.n6441 0.0225448
R16386 vdd.n6441 vdd.t684 0.0225448
R16387 vdd.n6426 vdd.n6402 0.0225448
R16388 vdd.t686 vdd.n6426 0.0225448
R16389 vdd.n6424 vdd.n6423 0.0225448
R16390 vdd.n6466 vdd.n6465 0.0225448
R16391 vdd.n6466 vdd.t1367 0.0225448
R16392 vdd.n6476 vdd.n6475 0.0225448
R16393 vdd.n6475 vdd.t1169 0.0225448
R16394 vdd.n6478 vdd.n6455 0.0225448
R16395 vdd.t1170 vdd.n6455 0.0225448
R16396 vdd.n6485 vdd.n6484 0.0225448
R16397 vdd.n6481 vdd.n6480 0.0225448
R16398 vdd.n6481 vdd.t894 0.0225448
R16399 vdd.n6490 vdd.n6489 0.0225448
R16400 vdd.n6489 vdd.t1170 0.0225448
R16401 vdd.n6474 vdd.n6450 0.0225448
R16402 vdd.t1169 vdd.n6474 0.0225448
R16403 vdd.n6472 vdd.n6471 0.0225448
R16404 vdd.n6512 vdd.n6511 0.0225448
R16405 vdd.n6512 vdd.t314 0.0225448
R16406 vdd.n6522 vdd.n6521 0.0225448
R16407 vdd.n6521 vdd.t121 0.0225448
R16408 vdd.n6524 vdd.n6501 0.0225448
R16409 vdd.t119 vdd.n6501 0.0225448
R16410 vdd.n6531 vdd.n6530 0.0225448
R16411 vdd.n6527 vdd.n6526 0.0225448
R16412 vdd.n6527 vdd.t564 0.0225448
R16413 vdd.n6536 vdd.n6535 0.0225448
R16414 vdd.n6535 vdd.t119 0.0225448
R16415 vdd.n6520 vdd.n6496 0.0225448
R16416 vdd.t121 vdd.n6520 0.0225448
R16417 vdd.n6518 vdd.n6517 0.0225448
R16418 vdd.n672 vdd.n671 0.0225448
R16419 vdd.n672 vdd.t695 0.0225448
R16420 vdd.n682 vdd.n681 0.0225448
R16421 vdd.n681 vdd.t46 0.0225448
R16422 vdd.n684 vdd.n661 0.0225448
R16423 vdd.t47 vdd.n661 0.0225448
R16424 vdd.n691 vdd.n690 0.0225448
R16425 vdd.n687 vdd.n686 0.0225448
R16426 vdd.n687 vdd.t1465 0.0225448
R16427 vdd.n696 vdd.n695 0.0225448
R16428 vdd.n695 vdd.t47 0.0225448
R16429 vdd.n680 vdd.n656 0.0225448
R16430 vdd.t46 vdd.n680 0.0225448
R16431 vdd.n678 vdd.n677 0.0225448
R16432 vdd.n718 vdd.n717 0.0225448
R16433 vdd.n718 vdd.t1406 0.0225448
R16434 vdd.n728 vdd.n727 0.0225448
R16435 vdd.n727 vdd.t123 0.0225448
R16436 vdd.n730 vdd.n707 0.0225448
R16437 vdd.t124 vdd.n707 0.0225448
R16438 vdd.n737 vdd.n736 0.0225448
R16439 vdd.n733 vdd.n732 0.0225448
R16440 vdd.n733 vdd.t1501 0.0225448
R16441 vdd.n742 vdd.n741 0.0225448
R16442 vdd.n741 vdd.t124 0.0225448
R16443 vdd.n726 vdd.n702 0.0225448
R16444 vdd.t123 vdd.n726 0.0225448
R16445 vdd.n724 vdd.n723 0.0225448
R16446 vdd.n816 vdd.n815 0.0225448
R16447 vdd.n816 vdd.t1202 0.0225448
R16448 vdd.n826 vdd.n825 0.0225448
R16449 vdd.n825 vdd.t291 0.0225448
R16450 vdd.n828 vdd.n805 0.0225448
R16451 vdd.t289 vdd.n805 0.0225448
R16452 vdd.n835 vdd.n834 0.0225448
R16453 vdd.n831 vdd.n830 0.0225448
R16454 vdd.n831 vdd.t1358 0.0225448
R16455 vdd.n840 vdd.n839 0.0225448
R16456 vdd.n839 vdd.t289 0.0225448
R16457 vdd.n824 vdd.n800 0.0225448
R16458 vdd.t291 vdd.n824 0.0225448
R16459 vdd.n822 vdd.n821 0.0225448
R16460 vdd.n862 vdd.n861 0.0225448
R16461 vdd.n862 vdd.t1383 0.0225448
R16462 vdd.n872 vdd.n871 0.0225448
R16463 vdd.n871 vdd.t427 0.0225448
R16464 vdd.n874 vdd.n851 0.0225448
R16465 vdd.t425 vdd.n851 0.0225448
R16466 vdd.n881 vdd.n880 0.0225448
R16467 vdd.n877 vdd.n876 0.0225448
R16468 vdd.n877 vdd.t1497 0.0225448
R16469 vdd.n886 vdd.n885 0.0225448
R16470 vdd.n885 vdd.t425 0.0225448
R16471 vdd.n870 vdd.n846 0.0225448
R16472 vdd.t427 vdd.n870 0.0225448
R16473 vdd.n868 vdd.n867 0.0225448
R16474 vdd.n908 vdd.n907 0.0225448
R16475 vdd.n908 vdd.t361 0.0225448
R16476 vdd.n918 vdd.n917 0.0225448
R16477 vdd.n917 vdd.t215 0.0225448
R16478 vdd.n920 vdd.n897 0.0225448
R16479 vdd.t213 vdd.n897 0.0225448
R16480 vdd.n927 vdd.n926 0.0225448
R16481 vdd.n923 vdd.n922 0.0225448
R16482 vdd.n923 vdd.t1312 0.0225448
R16483 vdd.n932 vdd.n931 0.0225448
R16484 vdd.n931 vdd.t213 0.0225448
R16485 vdd.n916 vdd.n892 0.0225448
R16486 vdd.t215 vdd.n916 0.0225448
R16487 vdd.n914 vdd.n913 0.0225448
R16488 vdd.n954 vdd.n953 0.0225448
R16489 vdd.n954 vdd.t236 0.0225448
R16490 vdd.n964 vdd.n963 0.0225448
R16491 vdd.n963 vdd.t923 0.0225448
R16492 vdd.n966 vdd.n943 0.0225448
R16493 vdd.t921 vdd.n943 0.0225448
R16494 vdd.n973 vdd.n972 0.0225448
R16495 vdd.n969 vdd.n968 0.0225448
R16496 vdd.n969 vdd.t462 0.0225448
R16497 vdd.n978 vdd.n977 0.0225448
R16498 vdd.n977 vdd.t921 0.0225448
R16499 vdd.n962 vdd.n938 0.0225448
R16500 vdd.t923 vdd.n962 0.0225448
R16501 vdd.n960 vdd.n959 0.0225448
R16502 vdd.n1052 vdd.n1051 0.0225448
R16503 vdd.n1052 vdd.t1259 0.0225448
R16504 vdd.n1062 vdd.n1061 0.0225448
R16505 vdd.n1061 vdd.t957 0.0225448
R16506 vdd.n1064 vdd.n1041 0.0225448
R16507 vdd.t955 vdd.n1041 0.0225448
R16508 vdd.n1071 vdd.n1070 0.0225448
R16509 vdd.n1067 vdd.n1066 0.0225448
R16510 vdd.n1067 vdd.t1469 0.0225448
R16511 vdd.n1076 vdd.n1075 0.0225448
R16512 vdd.n1075 vdd.t955 0.0225448
R16513 vdd.n1060 vdd.n1036 0.0225448
R16514 vdd.t957 vdd.n1060 0.0225448
R16515 vdd.n1058 vdd.n1057 0.0225448
R16516 vdd.n2510 vdd.n2509 0.0225448
R16517 vdd.n2510 vdd.t1213 0.0225448
R16518 vdd.n2520 vdd.n2519 0.0225448
R16519 vdd.n2519 vdd.t181 0.0225448
R16520 vdd.n2522 vdd.n2499 0.0225448
R16521 vdd.t179 vdd.n2499 0.0225448
R16522 vdd.n2529 vdd.n2528 0.0225448
R16523 vdd.n2525 vdd.n2524 0.0225448
R16524 vdd.n2525 vdd.t381 0.0225448
R16525 vdd.n2534 vdd.n2533 0.0225448
R16526 vdd.n2533 vdd.t179 0.0225448
R16527 vdd.n2518 vdd.n2494 0.0225448
R16528 vdd.t181 vdd.n2518 0.0225448
R16529 vdd.n2516 vdd.n2515 0.0225448
R16530 vdd.n1100 vdd.n1099 0.0225448
R16531 vdd.n1109 vdd.n1108 0.0225448
R16532 vdd.n1108 vdd.t111 0.0225448
R16533 vdd.n1114 vdd.n1113 0.0225448
R16534 vdd.n1114 vdd.t113 0.0225448
R16535 vdd.n1117 vdd.n1089 0.0225448
R16536 vdd.n1117 vdd.t947 0.0225448
R16537 vdd.n1105 vdd.t3 0.0225448
R16538 vdd.t111 vdd.n1107 0.0225448
R16539 vdd.n1123 vdd.t113 0.0225448
R16540 vdd.n1121 vdd.n1120 0.0225448
R16541 vdd.n1124 vdd.n1123 0.0225448
R16542 vdd.n1107 vdd.n1084 0.0225448
R16543 vdd.n1105 vdd.n1104 0.0225448
R16544 vdd.n1146 vdd.n1145 0.0225448
R16545 vdd.n1155 vdd.n1154 0.0225448
R16546 vdd.n1154 vdd.t731 0.0225448
R16547 vdd.n1160 vdd.n1159 0.0225448
R16548 vdd.n1160 vdd.t730 0.0225448
R16549 vdd.n1163 vdd.n1135 0.0225448
R16550 vdd.n1163 vdd.t747 0.0225448
R16551 vdd.n1151 vdd.t195 0.0225448
R16552 vdd.t731 vdd.n1153 0.0225448
R16553 vdd.n1169 vdd.t730 0.0225448
R16554 vdd.n1167 vdd.n1166 0.0225448
R16555 vdd.n1170 vdd.n1169 0.0225448
R16556 vdd.n1153 vdd.n1130 0.0225448
R16557 vdd.n1151 vdd.n1150 0.0225448
R16558 vdd.n1243 vdd.n1242 0.0225448
R16559 vdd.n1252 vdd.n1251 0.0225448
R16560 vdd.n1251 vdd.t1368 0.0225448
R16561 vdd.n1257 vdd.n1256 0.0225448
R16562 vdd.n1257 vdd.t1370 0.0225448
R16563 vdd.n1260 vdd.n1232 0.0225448
R16564 vdd.n1260 vdd.t86 0.0225448
R16565 vdd.n1248 vdd.t1308 0.0225448
R16566 vdd.t1368 vdd.n1250 0.0225448
R16567 vdd.n1266 vdd.t1370 0.0225448
R16568 vdd.n1264 vdd.n1263 0.0225448
R16569 vdd.n1267 vdd.n1266 0.0225448
R16570 vdd.n1250 vdd.n1227 0.0225448
R16571 vdd.n1248 vdd.n1247 0.0225448
R16572 vdd.n1289 vdd.n1288 0.0225448
R16573 vdd.n1298 vdd.n1297 0.0225448
R16574 vdd.n1297 vdd.t1103 0.0225448
R16575 vdd.n1303 vdd.n1302 0.0225448
R16576 vdd.n1303 vdd.t1105 0.0225448
R16577 vdd.n1306 vdd.n1278 0.0225448
R16578 vdd.n1306 vdd.t157 0.0225448
R16579 vdd.n1294 vdd.t1495 0.0225448
R16580 vdd.t1103 vdd.n1296 0.0225448
R16581 vdd.n1312 vdd.t1105 0.0225448
R16582 vdd.n1310 vdd.n1309 0.0225448
R16583 vdd.n1313 vdd.n1312 0.0225448
R16584 vdd.n1296 vdd.n1273 0.0225448
R16585 vdd.n1294 vdd.n1293 0.0225448
R16586 vdd.n1335 vdd.n1334 0.0225448
R16587 vdd.n1344 vdd.n1343 0.0225448
R16588 vdd.n1343 vdd.t311 0.0225448
R16589 vdd.n1349 vdd.n1348 0.0225448
R16590 vdd.n1349 vdd.t313 0.0225448
R16591 vdd.n1352 vdd.n1324 0.0225448
R16592 vdd.n1352 vdd.t65 0.0225448
R16593 vdd.n1340 vdd.t1356 0.0225448
R16594 vdd.t311 vdd.n1342 0.0225448
R16595 vdd.n1358 vdd.t313 0.0225448
R16596 vdd.n1356 vdd.n1355 0.0225448
R16597 vdd.n1359 vdd.n1358 0.0225448
R16598 vdd.n1342 vdd.n1319 0.0225448
R16599 vdd.n1340 vdd.n1339 0.0225448
R16600 vdd.n1381 vdd.n1380 0.0225448
R16601 vdd.n1390 vdd.n1389 0.0225448
R16602 vdd.n1389 vdd.t918 0.0225448
R16603 vdd.n1395 vdd.n1394 0.0225448
R16604 vdd.n1395 vdd.t917 0.0225448
R16605 vdd.n1398 vdd.n1370 0.0225448
R16606 vdd.n1398 vdd.t920 0.0225448
R16607 vdd.n1386 vdd.t591 0.0225448
R16608 vdd.t918 vdd.n1388 0.0225448
R16609 vdd.n1404 vdd.t917 0.0225448
R16610 vdd.n1402 vdd.n1401 0.0225448
R16611 vdd.n1405 vdd.n1404 0.0225448
R16612 vdd.n1388 vdd.n1365 0.0225448
R16613 vdd.n1386 vdd.n1385 0.0225448
R16614 vdd.n1478 vdd.n1477 0.0225448
R16615 vdd.n1487 vdd.n1486 0.0225448
R16616 vdd.n1486 vdd.t409 0.0225448
R16617 vdd.n1492 vdd.n1491 0.0225448
R16618 vdd.n1492 vdd.t408 0.0225448
R16619 vdd.n1495 vdd.n1467 0.0225448
R16620 vdd.n1495 vdd.t1447 0.0225448
R16621 vdd.n1483 vdd.t385 0.0225448
R16622 vdd.t409 vdd.n1485 0.0225448
R16623 vdd.n1501 vdd.t408 0.0225448
R16624 vdd.n1499 vdd.n1498 0.0225448
R16625 vdd.n1502 vdd.n1501 0.0225448
R16626 vdd.n1485 vdd.n1462 0.0225448
R16627 vdd.n1483 vdd.n1482 0.0225448
R16628 vdd.n627 vdd.n626 0.0225448
R16629 vdd.n636 vdd.n635 0.0225448
R16630 vdd.n635 vdd.t348 0.0225448
R16631 vdd.n641 vdd.n640 0.0225448
R16632 vdd.n641 vdd.t347 0.0225448
R16633 vdd.n644 vdd.n616 0.0225448
R16634 vdd.n644 vdd.t893 0.0225448
R16635 vdd.n632 vdd.t552 0.0225448
R16636 vdd.t348 vdd.n634 0.0225448
R16637 vdd.n650 vdd.t347 0.0225448
R16638 vdd.n648 vdd.n647 0.0225448
R16639 vdd.n651 vdd.n650 0.0225448
R16640 vdd.n634 vdd.n611 0.0225448
R16641 vdd.n632 vdd.n631 0.0225448
R16642 vdd.n1522 vdd.n1521 0.0225448
R16643 vdd.n1531 vdd.n1530 0.0225448
R16644 vdd.n1530 vdd.t1222 0.0225448
R16645 vdd.n1536 vdd.n1535 0.0225448
R16646 vdd.n1536 vdd.t1224 0.0225448
R16647 vdd.n1539 vdd.n1511 0.0225448
R16648 vdd.n1539 vdd.t1142 0.0225448
R16649 vdd.n1527 vdd.t823 0.0225448
R16650 vdd.t1222 vdd.n1529 0.0225448
R16651 vdd.n1545 vdd.t1224 0.0225448
R16652 vdd.n1543 vdd.n1542 0.0225448
R16653 vdd.n1546 vdd.n1545 0.0225448
R16654 vdd.n1529 vdd.n1506 0.0225448
R16655 vdd.n1527 vdd.n1526 0.0225448
R16656 vdd.n1567 vdd.n1566 0.0225448
R16657 vdd.n1576 vdd.n1575 0.0225448
R16658 vdd.n1575 vdd.t1188 0.0225448
R16659 vdd.n1581 vdd.n1580 0.0225448
R16660 vdd.n1581 vdd.t1190 0.0225448
R16661 vdd.n1584 vdd.n1556 0.0225448
R16662 vdd.n1584 vdd.t1121 0.0225448
R16663 vdd.n1572 vdd.t833 0.0225448
R16664 vdd.t1188 vdd.n1574 0.0225448
R16665 vdd.n1590 vdd.t1190 0.0225448
R16666 vdd.n1588 vdd.n1587 0.0225448
R16667 vdd.n1591 vdd.n1590 0.0225448
R16668 vdd.n1574 vdd.n1551 0.0225448
R16669 vdd.n1572 vdd.n1571 0.0225448
R16670 vdd.n1617 vdd.n1616 0.0225448
R16671 vdd.n1626 vdd.n1625 0.0225448
R16672 vdd.n1625 vdd.t1068 0.0225448
R16673 vdd.n1631 vdd.n1630 0.0225448
R16674 vdd.n1631 vdd.t1070 0.0225448
R16675 vdd.n1634 vdd.n1606 0.0225448
R16676 vdd.n1634 vdd.t1033 0.0225448
R16677 vdd.n1622 vdd.t466 0.0225448
R16678 vdd.t1068 vdd.n1624 0.0225448
R16679 vdd.n1640 vdd.t1070 0.0225448
R16680 vdd.n1638 vdd.n1637 0.0225448
R16681 vdd.n1641 vdd.n1640 0.0225448
R16682 vdd.n1624 vdd.n1601 0.0225448
R16683 vdd.n1622 vdd.n1621 0.0225448
R16684 vdd.n1663 vdd.n1662 0.0225448
R16685 vdd.n1672 vdd.n1671 0.0225448
R16686 vdd.n1671 vdd.t953 0.0225448
R16687 vdd.n1677 vdd.n1676 0.0225448
R16688 vdd.n1677 vdd.t952 0.0225448
R16689 vdd.n1680 vdd.n1652 0.0225448
R16690 vdd.n1680 vdd.t309 0.0225448
R16691 vdd.n1668 vdd.t998 0.0225448
R16692 vdd.t953 vdd.n1670 0.0225448
R16693 vdd.n1686 vdd.t952 0.0225448
R16694 vdd.n1684 vdd.n1683 0.0225448
R16695 vdd.n1687 vdd.n1686 0.0225448
R16696 vdd.n1670 vdd.n1647 0.0225448
R16697 vdd.n1668 vdd.n1667 0.0225448
R16698 vdd.n1711 vdd.n1710 0.0225448
R16699 vdd.n1720 vdd.n1719 0.0225448
R16700 vdd.n1719 vdd.t83 0.0225448
R16701 vdd.n1725 vdd.n1724 0.0225448
R16702 vdd.n1725 vdd.t85 0.0225448
R16703 vdd.n1728 vdd.n1700 0.0225448
R16704 vdd.n1728 vdd.t1018 0.0225448
R16705 vdd.n1716 vdd.t1493 0.0225448
R16706 vdd.t83 vdd.n1718 0.0225448
R16707 vdd.n1734 vdd.t85 0.0225448
R16708 vdd.n1732 vdd.n1731 0.0225448
R16709 vdd.n1735 vdd.n1734 0.0225448
R16710 vdd.n1718 vdd.n1695 0.0225448
R16711 vdd.n1716 vdd.n1715 0.0225448
R16712 vdd.n1429 vdd.n1428 0.0225448
R16713 vdd.n1432 vdd.n1431 0.0225448
R16714 vdd.n1431 vdd.t1072 0.0225448
R16715 vdd.n1437 vdd.n1436 0.0225448
R16716 vdd.n1437 vdd.t1074 0.0225448
R16717 vdd.n1440 vdd.n1421 0.0225448
R16718 vdd.n1440 vdd.t1443 0.0225448
R16719 vdd.n1453 vdd.t101 0.0225448
R16720 vdd.n1451 vdd.t1072 0.0225448
R16721 vdd.n1446 vdd.t1074 0.0225448
R16722 vdd.n1444 vdd.n1443 0.0225448
R16723 vdd.n1447 vdd.n1446 0.0225448
R16724 vdd.n1451 vdd.n1450 0.0225448
R16725 vdd.n1454 vdd.n1453 0.0225448
R16726 vdd.n1758 vdd.n1757 0.0225448
R16727 vdd.n1767 vdd.n1766 0.0225448
R16728 vdd.n1766 vdd.t664 0.0225448
R16729 vdd.n1772 vdd.n1771 0.0225448
R16730 vdd.n1772 vdd.t666 0.0225448
R16731 vdd.n1775 vdd.n1747 0.0225448
R16732 vdd.n1775 vdd.t683 0.0225448
R16733 vdd.n1763 vdd.t870 0.0225448
R16734 vdd.t664 vdd.n1765 0.0225448
R16735 vdd.n1781 vdd.t666 0.0225448
R16736 vdd.n1779 vdd.n1778 0.0225448
R16737 vdd.n1782 vdd.n1781 0.0225448
R16738 vdd.n1765 vdd.n1742 0.0225448
R16739 vdd.n1763 vdd.n1762 0.0225448
R16740 vdd.n1803 vdd.n1802 0.0225448
R16741 vdd.n1812 vdd.n1811 0.0225448
R16742 vdd.n1811 vdd.t368 0.0225448
R16743 vdd.n1817 vdd.n1816 0.0225448
R16744 vdd.n1817 vdd.t370 0.0225448
R16745 vdd.n1820 vdd.n1792 0.0225448
R16746 vdd.n1820 vdd.t132 0.0225448
R16747 vdd.n1808 vdd.t170 0.0225448
R16748 vdd.t368 vdd.n1810 0.0225448
R16749 vdd.n1826 vdd.t370 0.0225448
R16750 vdd.n1824 vdd.n1823 0.0225448
R16751 vdd.n1827 vdd.n1826 0.0225448
R16752 vdd.n1810 vdd.n1787 0.0225448
R16753 vdd.n1808 vdd.n1807 0.0225448
R16754 vdd.n1849 vdd.n1848 0.0225448
R16755 vdd.n1858 vdd.n1857 0.0225448
R16756 vdd.n1857 vdd.t654 0.0225448
R16757 vdd.n1863 vdd.n1862 0.0225448
R16758 vdd.n1863 vdd.t656 0.0225448
R16759 vdd.n1866 vdd.n1838 0.0225448
R16760 vdd.n1866 vdd.t657 0.0225448
R16761 vdd.n1854 vdd.t1127 0.0225448
R16762 vdd.t654 vdd.n1856 0.0225448
R16763 vdd.n1872 vdd.t656 0.0225448
R16764 vdd.n1870 vdd.n1869 0.0225448
R16765 vdd.n1873 vdd.n1872 0.0225448
R16766 vdd.n1856 vdd.n1833 0.0225448
R16767 vdd.n1854 vdd.n1853 0.0225448
R16768 vdd.n1900 vdd.n1899 0.0225448
R16769 vdd.n1909 vdd.n1908 0.0225448
R16770 vdd.n1908 vdd.t787 0.0225448
R16771 vdd.n1914 vdd.n1913 0.0225448
R16772 vdd.n1914 vdd.t789 0.0225448
R16773 vdd.n1917 vdd.n1889 0.0225448
R16774 vdd.n1917 vdd.t1283 0.0225448
R16775 vdd.n1905 vdd.t1324 0.0225448
R16776 vdd.t787 vdd.n1907 0.0225448
R16777 vdd.n1923 vdd.t789 0.0225448
R16778 vdd.n1921 vdd.n1920 0.0225448
R16779 vdd.n1924 vdd.n1923 0.0225448
R16780 vdd.n1907 vdd.n1884 0.0225448
R16781 vdd.n1905 vdd.n1904 0.0225448
R16782 vdd.n1946 vdd.n1945 0.0225448
R16783 vdd.n1955 vdd.n1954 0.0225448
R16784 vdd.n1954 vdd.t388 0.0225448
R16785 vdd.n1960 vdd.n1959 0.0225448
R16786 vdd.n1960 vdd.t390 0.0225448
R16787 vdd.n1963 vdd.n1935 0.0225448
R16788 vdd.n1963 vdd.t391 0.0225448
R16789 vdd.n1951 vdd.t992 0.0225448
R16790 vdd.t388 vdd.n1953 0.0225448
R16791 vdd.n1969 vdd.t390 0.0225448
R16792 vdd.n1967 vdd.n1966 0.0225448
R16793 vdd.n1970 vdd.n1969 0.0225448
R16794 vdd.n1953 vdd.n1930 0.0225448
R16795 vdd.n1951 vdd.n1950 0.0225448
R16796 vdd.n1994 vdd.n1993 0.0225448
R16797 vdd.n2003 vdd.n2002 0.0225448
R16798 vdd.n2002 vdd.t158 0.0225448
R16799 vdd.n2008 vdd.n2007 0.0225448
R16800 vdd.n2008 vdd.t160 0.0225448
R16801 vdd.n2011 vdd.n1983 0.0225448
R16802 vdd.n2011 vdd.t268 0.0225448
R16803 vdd.n1999 vdd.t371 0.0225448
R16804 vdd.t158 vdd.n2001 0.0225448
R16805 vdd.n2017 vdd.t160 0.0225448
R16806 vdd.n2015 vdd.n2014 0.0225448
R16807 vdd.n2018 vdd.n2017 0.0225448
R16808 vdd.n2001 vdd.n1978 0.0225448
R16809 vdd.n1999 vdd.n1998 0.0225448
R16810 vdd.n2040 vdd.n2039 0.0225448
R16811 vdd.n2049 vdd.n2048 0.0225448
R16812 vdd.n2048 vdd.t1218 0.0225448
R16813 vdd.n2054 vdd.n2053 0.0225448
R16814 vdd.n2054 vdd.t1217 0.0225448
R16815 vdd.n2057 vdd.n2029 0.0225448
R16816 vdd.n2057 vdd.t1220 0.0225448
R16817 vdd.n2045 vdd.t971 0.0225448
R16818 vdd.t1218 vdd.n2047 0.0225448
R16819 vdd.n2063 vdd.t1217 0.0225448
R16820 vdd.n2061 vdd.n2060 0.0225448
R16821 vdd.n2064 vdd.n2063 0.0225448
R16822 vdd.n2047 vdd.n2024 0.0225448
R16823 vdd.n2045 vdd.n2044 0.0225448
R16824 vdd.n2085 vdd.n2084 0.0225448
R16825 vdd.n2094 vdd.n2093 0.0225448
R16826 vdd.n2093 vdd.t841 0.0225448
R16827 vdd.n2099 vdd.n2098 0.0225448
R16828 vdd.n2099 vdd.t843 0.0225448
R16829 vdd.n2102 vdd.n2074 0.0225448
R16830 vdd.n2102 vdd.t226 0.0225448
R16831 vdd.n2090 vdd.t168 0.0225448
R16832 vdd.t841 vdd.n2092 0.0225448
R16833 vdd.n2108 vdd.t843 0.0225448
R16834 vdd.n2106 vdd.n2105 0.0225448
R16835 vdd.n2109 vdd.n2108 0.0225448
R16836 vdd.n2092 vdd.n2069 0.0225448
R16837 vdd.n2090 vdd.n2089 0.0225448
R16838 vdd.n2135 vdd.n2134 0.0225448
R16839 vdd.n2144 vdd.n2143 0.0225448
R16840 vdd.n2143 vdd.t635 0.0225448
R16841 vdd.n2149 vdd.n2148 0.0225448
R16842 vdd.n2149 vdd.t637 0.0225448
R16843 vdd.n2152 vdd.n2124 0.0225448
R16844 vdd.n2152 vdd.t110 0.0225448
R16845 vdd.n2140 vdd.t1344 0.0225448
R16846 vdd.t635 vdd.n2142 0.0225448
R16847 vdd.n2158 vdd.t637 0.0225448
R16848 vdd.n2156 vdd.n2155 0.0225448
R16849 vdd.n2159 vdd.n2158 0.0225448
R16850 vdd.n2142 vdd.n2119 0.0225448
R16851 vdd.n2140 vdd.n2139 0.0225448
R16852 vdd.n2181 vdd.n2180 0.0225448
R16853 vdd.n2190 vdd.n2189 0.0225448
R16854 vdd.n2189 vdd.t232 0.0225448
R16855 vdd.n2195 vdd.n2194 0.0225448
R16856 vdd.n2195 vdd.t231 0.0225448
R16857 vdd.n2198 vdd.n2170 0.0225448
R16858 vdd.n2198 vdd.t1131 0.0225448
R16859 vdd.n2186 vdd.t940 0.0225448
R16860 vdd.t232 vdd.n2188 0.0225448
R16861 vdd.n2204 vdd.t231 0.0225448
R16862 vdd.n2202 vdd.n2201 0.0225448
R16863 vdd.n2205 vdd.n2204 0.0225448
R16864 vdd.n2188 vdd.n2165 0.0225448
R16865 vdd.n2186 vdd.n2185 0.0225448
R16866 vdd.n2229 vdd.n2228 0.0225448
R16867 vdd.n2238 vdd.n2237 0.0225448
R16868 vdd.n2237 vdd.t1116 0.0225448
R16869 vdd.n2243 vdd.n2242 0.0225448
R16870 vdd.n2243 vdd.t1118 0.0225448
R16871 vdd.n2246 vdd.n2218 0.0225448
R16872 vdd.n2246 vdd.t1119 0.0225448
R16873 vdd.n2234 vdd.t1481 0.0225448
R16874 vdd.t1116 vdd.n2236 0.0225448
R16875 vdd.n2252 vdd.t1118 0.0225448
R16876 vdd.n2250 vdd.n2249 0.0225448
R16877 vdd.n2253 vdd.n2252 0.0225448
R16878 vdd.n2236 vdd.n2213 0.0225448
R16879 vdd.n2234 vdd.n2233 0.0225448
R16880 vdd.n1194 vdd.n1193 0.0225448
R16881 vdd.n1197 vdd.n1196 0.0225448
R16882 vdd.n1196 vdd.t672 0.0225448
R16883 vdd.n1202 vdd.n1201 0.0225448
R16884 vdd.n1202 vdd.t674 0.0225448
R16885 vdd.n1205 vdd.n1186 0.0225448
R16886 vdd.n1205 vdd.t1163 0.0225448
R16887 vdd.n1218 vdd.t95 0.0225448
R16888 vdd.n1216 vdd.t672 0.0225448
R16889 vdd.n1211 vdd.t674 0.0225448
R16890 vdd.n1209 vdd.n1208 0.0225448
R16891 vdd.n1212 vdd.n1211 0.0225448
R16892 vdd.n1216 vdd.n1215 0.0225448
R16893 vdd.n1219 vdd.n1218 0.0225448
R16894 vdd.n2276 vdd.n2275 0.0225448
R16895 vdd.n2285 vdd.n2284 0.0225448
R16896 vdd.n2284 vdd.t296 0.0225448
R16897 vdd.n2290 vdd.n2289 0.0225448
R16898 vdd.n2290 vdd.t298 0.0225448
R16899 vdd.n2293 vdd.n2265 0.0225448
R16900 vdd.n2293 vdd.t929 0.0225448
R16901 vdd.n2281 vdd.t900 0.0225448
R16902 vdd.t296 vdd.n2283 0.0225448
R16903 vdd.n2299 vdd.t298 0.0225448
R16904 vdd.n2297 vdd.n2296 0.0225448
R16905 vdd.n2300 vdd.n2299 0.0225448
R16906 vdd.n2283 vdd.n2260 0.0225448
R16907 vdd.n2281 vdd.n2280 0.0225448
R16908 vdd.n2321 vdd.n2320 0.0225448
R16909 vdd.n2330 vdd.n2329 0.0225448
R16910 vdd.n2329 vdd.t116 0.0225448
R16911 vdd.n2335 vdd.n2334 0.0225448
R16912 vdd.n2335 vdd.t118 0.0225448
R16913 vdd.n2338 vdd.n2310 0.0225448
R16914 vdd.n2338 vdd.t516 0.0225448
R16915 vdd.n2326 vdd.t771 0.0225448
R16916 vdd.t116 vdd.n2328 0.0225448
R16917 vdd.n2344 vdd.t118 0.0225448
R16918 vdd.n2342 vdd.n2341 0.0225448
R16919 vdd.n2345 vdd.n2344 0.0225448
R16920 vdd.n2328 vdd.n2305 0.0225448
R16921 vdd.n2326 vdd.n2325 0.0225448
R16922 vdd.n2371 vdd.n2370 0.0225448
R16923 vdd.n2380 vdd.n2379 0.0225448
R16924 vdd.n2379 vdd.t1038 0.0225448
R16925 vdd.n2385 vdd.n2384 0.0225448
R16926 vdd.n2385 vdd.t1040 0.0225448
R16927 vdd.n2388 vdd.n2360 0.0225448
R16928 vdd.n2388 vdd.t103 0.0225448
R16929 vdd.n2376 vdd.t492 0.0225448
R16930 vdd.t1038 vdd.n2378 0.0225448
R16931 vdd.n2394 vdd.t1040 0.0225448
R16932 vdd.n2392 vdd.n2391 0.0225448
R16933 vdd.n2395 vdd.n2394 0.0225448
R16934 vdd.n2378 vdd.n2355 0.0225448
R16935 vdd.n2376 vdd.n2375 0.0225448
R16936 vdd.n2417 vdd.n2416 0.0225448
R16937 vdd.n2426 vdd.n2425 0.0225448
R16938 vdd.n2425 vdd.t875 0.0225448
R16939 vdd.n2431 vdd.n2430 0.0225448
R16940 vdd.n2431 vdd.t877 0.0225448
R16941 vdd.n2434 vdd.n2406 0.0225448
R16942 vdd.n2434 vdd.t606 0.0225448
R16943 vdd.n2422 vdd.t975 0.0225448
R16944 vdd.t875 vdd.n2424 0.0225448
R16945 vdd.n2440 vdd.t877 0.0225448
R16946 vdd.n2438 vdd.n2437 0.0225448
R16947 vdd.n2441 vdd.n2440 0.0225448
R16948 vdd.n2424 vdd.n2401 0.0225448
R16949 vdd.n2422 vdd.n2421 0.0225448
R16950 vdd.n2465 vdd.n2464 0.0225448
R16951 vdd.n2474 vdd.n2473 0.0225448
R16952 vdd.n2473 vdd.t1444 0.0225448
R16953 vdd.n2479 vdd.n2478 0.0225448
R16954 vdd.n2479 vdd.t1446 0.0225448
R16955 vdd.n2482 vdd.n2454 0.0225448
R16956 vdd.n2482 vdd.t1423 0.0225448
R16957 vdd.n2470 vdd.t1348 0.0225448
R16958 vdd.t1444 vdd.n2472 0.0225448
R16959 vdd.n2488 vdd.t1446 0.0225448
R16960 vdd.n2486 vdd.n2485 0.0225448
R16961 vdd.n2489 vdd.n2488 0.0225448
R16962 vdd.n2472 vdd.n2449 0.0225448
R16963 vdd.n2470 vdd.n2469 0.0225448
R16964 vdd.n2603 vdd.n2602 0.0225448
R16965 vdd.n2603 vdd.t423 0.0225448
R16966 vdd.n2613 vdd.n2612 0.0225448
R16967 vdd.n2612 vdd.t526 0.0225448
R16968 vdd.n2615 vdd.n2592 0.0225448
R16969 vdd.t524 vdd.n2592 0.0225448
R16970 vdd.n2622 vdd.n2621 0.0225448
R16971 vdd.n2618 vdd.n2617 0.0225448
R16972 vdd.n2618 vdd.t815 0.0225448
R16973 vdd.n2627 vdd.n2626 0.0225448
R16974 vdd.n2626 vdd.t524 0.0225448
R16975 vdd.n2611 vdd.n2587 0.0225448
R16976 vdd.t526 vdd.n2611 0.0225448
R16977 vdd.n2609 vdd.n2608 0.0225448
R16978 vdd.n2557 vdd.n2556 0.0225448
R16979 vdd.n2557 vdd.t1027 0.0225448
R16980 vdd.n2567 vdd.n2566 0.0225448
R16981 vdd.n2566 vdd.t334 0.0225448
R16982 vdd.n2569 vdd.n2546 0.0225448
R16983 vdd.t332 vdd.n2546 0.0225448
R16984 vdd.n2576 vdd.n2575 0.0225448
R16985 vdd.n2572 vdd.n2571 0.0225448
R16986 vdd.n2572 vdd.t769 0.0225448
R16987 vdd.n2581 vdd.n2580 0.0225448
R16988 vdd.n2580 vdd.t332 0.0225448
R16989 vdd.n2565 vdd.n2541 0.0225448
R16990 vdd.t334 vdd.n2565 0.0225448
R16991 vdd.n2563 vdd.n2562 0.0225448
R16992 vdd.n2650 vdd.n2649 0.0225448
R16993 vdd.n2650 vdd.t916 0.0225448
R16994 vdd.n2660 vdd.n2659 0.0225448
R16995 vdd.n2659 vdd.t618 0.0225448
R16996 vdd.n2662 vdd.n2639 0.0225448
R16997 vdd.t616 vdd.n2639 0.0225448
R16998 vdd.n2669 vdd.n2668 0.0225448
R16999 vdd.n2665 vdd.n2664 0.0225448
R17000 vdd.n2665 vdd.t1350 0.0225448
R17001 vdd.n2674 vdd.n2673 0.0225448
R17002 vdd.n2673 vdd.t616 0.0225448
R17003 vdd.n2658 vdd.n2634 0.0225448
R17004 vdd.t618 vdd.n2658 0.0225448
R17005 vdd.n2656 vdd.n2655 0.0225448
R17006 vdd.n2698 vdd.n2697 0.0225448
R17007 vdd.n2698 vdd.t717 0.0225448
R17008 vdd.n2708 vdd.n2707 0.0225448
R17009 vdd.n2707 vdd.t1098 0.0225448
R17010 vdd.n2710 vdd.n2687 0.0225448
R17011 vdd.t1096 vdd.n2687 0.0225448
R17012 vdd.n2717 vdd.n2716 0.0225448
R17013 vdd.n2713 vdd.n2712 0.0225448
R17014 vdd.n2713 vdd.t1016 0.0225448
R17015 vdd.n2722 vdd.n2721 0.0225448
R17016 vdd.n2721 vdd.t1096 0.0225448
R17017 vdd.n2706 vdd.n2682 0.0225448
R17018 vdd.t1098 vdd.n2706 0.0225448
R17019 vdd.n2704 vdd.n2703 0.0225448
R17020 vdd.n2744 vdd.n2743 0.0225448
R17021 vdd.n2744 vdd.t392 0.0225448
R17022 vdd.n2754 vdd.n2753 0.0225448
R17023 vdd.n2753 vdd.t1141 0.0225448
R17024 vdd.n2756 vdd.n2733 0.0225448
R17025 vdd.t1139 vdd.n2733 0.0225448
R17026 vdd.n2763 vdd.n2762 0.0225448
R17027 vdd.n2759 vdd.n2758 0.0225448
R17028 vdd.n2759 vdd.t494 0.0225448
R17029 vdd.n2768 vdd.n2767 0.0225448
R17030 vdd.n2767 vdd.t1139 0.0225448
R17031 vdd.n2752 vdd.n2728 0.0225448
R17032 vdd.t1141 vdd.n2752 0.0225448
R17033 vdd.n2750 vdd.n2749 0.0225448
R17034 vdd.n1008 vdd.n1007 0.0225448
R17035 vdd.n1007 vdd.t1230 0.0225448
R17036 vdd.n1010 vdd.n996 0.0225448
R17037 vdd.t404 vdd.n996 0.0225448
R17038 vdd.n1013 vdd.n1012 0.0225448
R17039 vdd.t402 vdd.n1013 0.0225448
R17040 vdd.n1028 vdd.n1027 0.0225448
R17041 vdd.n1025 vdd.n985 0.0225448
R17042 vdd.t91 vdd.n1025 0.0225448
R17043 vdd.n1020 vdd.n990 0.0225448
R17044 vdd.t402 vdd.n990 0.0225448
R17045 vdd.n1016 vdd.n1015 0.0225448
R17046 vdd.n1015 vdd.t404 0.0225448
R17047 vdd.n1005 vdd.n1004 0.0225448
R17048 vdd.n2886 vdd.n2885 0.0225448
R17049 vdd.n2886 vdd.t445 0.0225448
R17050 vdd.n2896 vdd.n2895 0.0225448
R17051 vdd.n2895 vdd.t75 0.0225448
R17052 vdd.n2898 vdd.n2875 0.0225448
R17053 vdd.t73 vdd.n2875 0.0225448
R17054 vdd.n2905 vdd.n2904 0.0225448
R17055 vdd.n2901 vdd.n2900 0.0225448
R17056 vdd.n2901 vdd.t44 0.0225448
R17057 vdd.n2910 vdd.n2909 0.0225448
R17058 vdd.n2909 vdd.t73 0.0225448
R17059 vdd.n2894 vdd.n2870 0.0225448
R17060 vdd.t75 vdd.n2894 0.0225448
R17061 vdd.n2892 vdd.n2891 0.0225448
R17062 vdd.n2839 vdd.n2838 0.0225448
R17063 vdd.n2839 vdd.t1106 0.0225448
R17064 vdd.n2849 vdd.n2848 0.0225448
R17065 vdd.n2848 vdd.t133 0.0225448
R17066 vdd.n2851 vdd.n2828 0.0225448
R17067 vdd.t134 vdd.n2828 0.0225448
R17068 vdd.n2858 vdd.n2857 0.0225448
R17069 vdd.n2854 vdd.n2853 0.0225448
R17070 vdd.n2854 vdd.t438 0.0225448
R17071 vdd.n2863 vdd.n2862 0.0225448
R17072 vdd.n2862 vdd.t134 0.0225448
R17073 vdd.n2847 vdd.n2823 0.0225448
R17074 vdd.t133 vdd.n2847 0.0225448
R17075 vdd.n2845 vdd.n2844 0.0225448
R17076 vdd.n2793 vdd.n2792 0.0225448
R17077 vdd.n2793 vdd.t729 0.0225448
R17078 vdd.n2803 vdd.n2802 0.0225448
R17079 vdd.n2802 vdd.t614 0.0225448
R17080 vdd.n2805 vdd.n2782 0.0225448
R17081 vdd.t612 vdd.n2782 0.0225448
R17082 vdd.n2812 vdd.n2811 0.0225448
R17083 vdd.n2808 vdd.n2807 0.0225448
R17084 vdd.n2808 vdd.t1125 0.0225448
R17085 vdd.n2817 vdd.n2816 0.0225448
R17086 vdd.n2816 vdd.t612 0.0225448
R17087 vdd.n2801 vdd.n2777 0.0225448
R17088 vdd.t614 vdd.n2801 0.0225448
R17089 vdd.n2799 vdd.n2798 0.0225448
R17090 vdd.n2933 vdd.n2932 0.0225448
R17091 vdd.n2933 vdd.t605 0.0225448
R17092 vdd.n2943 vdd.n2942 0.0225448
R17093 vdd.n2942 vdd.t222 0.0225448
R17094 vdd.n2945 vdd.n2922 0.0225448
R17095 vdd.t220 vdd.n2922 0.0225448
R17096 vdd.n2952 vdd.n2951 0.0225448
R17097 vdd.n2948 vdd.n2947 0.0225448
R17098 vdd.n2948 vdd.t11 0.0225448
R17099 vdd.n2957 vdd.n2956 0.0225448
R17100 vdd.n2956 vdd.t220 0.0225448
R17101 vdd.n2941 vdd.n2917 0.0225448
R17102 vdd.t222 vdd.n2941 0.0225448
R17103 vdd.n2939 vdd.n2938 0.0225448
R17104 vdd.n2981 vdd.n2980 0.0225448
R17105 vdd.n2981 vdd.t1221 0.0225448
R17106 vdd.n2991 vdd.n2990 0.0225448
R17107 vdd.n2990 vdd.t1386 0.0225448
R17108 vdd.n2993 vdd.n2970 0.0225448
R17109 vdd.t1384 vdd.n2970 0.0225448
R17110 vdd.n3000 vdd.n2999 0.0225448
R17111 vdd.n2996 vdd.n2995 0.0225448
R17112 vdd.n2996 vdd.t38 0.0225448
R17113 vdd.n3005 vdd.n3004 0.0225448
R17114 vdd.n3004 vdd.t1384 0.0225448
R17115 vdd.n2989 vdd.n2965 0.0225448
R17116 vdd.t1386 vdd.n2989 0.0225448
R17117 vdd.n2987 vdd.n2986 0.0225448
R17118 vdd.n3027 vdd.n3026 0.0225448
R17119 vdd.n3027 vdd.t1434 0.0225448
R17120 vdd.n3037 vdd.n3036 0.0225448
R17121 vdd.n3036 vdd.t454 0.0225448
R17122 vdd.n3039 vdd.n3016 0.0225448
R17123 vdd.t452 vdd.n3016 0.0225448
R17124 vdd.n3046 vdd.n3045 0.0225448
R17125 vdd.n3042 vdd.n3041 0.0225448
R17126 vdd.n3042 vdd.t1296 0.0225448
R17127 vdd.n3051 vdd.n3050 0.0225448
R17128 vdd.n3050 vdd.t452 0.0225448
R17129 vdd.n3035 vdd.n3011 0.0225448
R17130 vdd.t454 vdd.n3035 0.0225448
R17131 vdd.n3033 vdd.n3032 0.0225448
R17132 vdd.n3121 vdd.n3120 0.0225448
R17133 vdd.n3121 vdd.t1156 0.0225448
R17134 vdd.n3131 vdd.n3130 0.0225448
R17135 vdd.n3130 vdd.t801 0.0225448
R17136 vdd.n3133 vdd.n3110 0.0225448
R17137 vdd.t799 vdd.n3110 0.0225448
R17138 vdd.n3140 vdd.n3139 0.0225448
R17139 vdd.n3136 vdd.n3135 0.0225448
R17140 vdd.n3136 vdd.t852 0.0225448
R17141 vdd.n3145 vdd.n3144 0.0225448
R17142 vdd.n3144 vdd.t799 0.0225448
R17143 vdd.n3129 vdd.n3105 0.0225448
R17144 vdd.t801 vdd.n3129 0.0225448
R17145 vdd.n3127 vdd.n3126 0.0225448
R17146 vdd.n3075 vdd.n3074 0.0225448
R17147 vdd.n3075 vdd.t21 0.0225448
R17148 vdd.n3085 vdd.n3084 0.0225448
R17149 vdd.n3084 vdd.t276 0.0225448
R17150 vdd.n3087 vdd.n3064 0.0225448
R17151 vdd.t274 vdd.n3064 0.0225448
R17152 vdd.n3094 vdd.n3093 0.0225448
R17153 vdd.n3090 vdd.n3089 0.0225448
R17154 vdd.n3090 vdd.t790 0.0225448
R17155 vdd.n3099 vdd.n3098 0.0225448
R17156 vdd.n3098 vdd.t274 0.0225448
R17157 vdd.n3083 vdd.n3059 0.0225448
R17158 vdd.t276 vdd.n3083 0.0225448
R17159 vdd.n3081 vdd.n3080 0.0225448
R17160 vdd.n3168 vdd.n3167 0.0225448
R17161 vdd.n3168 vdd.t245 0.0225448
R17162 vdd.n3178 vdd.n3177 0.0225448
R17163 vdd.n3177 vdd.t280 0.0225448
R17164 vdd.n3180 vdd.n3157 0.0225448
R17165 vdd.t278 vdd.n3157 0.0225448
R17166 vdd.n3187 vdd.n3186 0.0225448
R17167 vdd.n3183 vdd.n3182 0.0225448
R17168 vdd.n3183 vdd.t373 0.0225448
R17169 vdd.n3192 vdd.n3191 0.0225448
R17170 vdd.n3191 vdd.t278 0.0225448
R17171 vdd.n3176 vdd.n3152 0.0225448
R17172 vdd.t280 vdd.n3176 0.0225448
R17173 vdd.n3174 vdd.n3173 0.0225448
R17174 vdd.n3216 vdd.n3215 0.0225448
R17175 vdd.n3216 vdd.t1282 0.0225448
R17176 vdd.n3226 vdd.n3225 0.0225448
R17177 vdd.n3225 vdd.t1212 0.0225448
R17178 vdd.n3228 vdd.n3205 0.0225448
R17179 vdd.t1210 vdd.n3205 0.0225448
R17180 vdd.n3235 vdd.n3234 0.0225448
R17181 vdd.n3231 vdd.n3230 0.0225448
R17182 vdd.n3231 vdd.t967 0.0225448
R17183 vdd.n3240 vdd.n3239 0.0225448
R17184 vdd.n3239 vdd.t1210 0.0225448
R17185 vdd.n3224 vdd.n3200 0.0225448
R17186 vdd.t1212 vdd.n3224 0.0225448
R17187 vdd.n3222 vdd.n3221 0.0225448
R17188 vdd.n3262 vdd.n3261 0.0225448
R17189 vdd.n3262 vdd.t798 0.0225448
R17190 vdd.n3272 vdd.n3271 0.0225448
R17191 vdd.n3271 vdd.t1277 0.0225448
R17192 vdd.n3274 vdd.n3251 0.0225448
R17193 vdd.t1275 vdd.n3251 0.0225448
R17194 vdd.n3281 vdd.n3280 0.0225448
R17195 vdd.n3277 vdd.n3276 0.0225448
R17196 vdd.n3277 vdd.t1328 0.0225448
R17197 vdd.n3286 vdd.n3285 0.0225448
R17198 vdd.n3285 vdd.t1275 0.0225448
R17199 vdd.n3270 vdd.n3246 0.0225448
R17200 vdd.t1277 vdd.n3270 0.0225448
R17201 vdd.n3268 vdd.n3267 0.0225448
R17202 vdd.n772 vdd.n771 0.0225448
R17203 vdd.n771 vdd.t1410 0.0225448
R17204 vdd.n774 vdd.n760 0.0225448
R17205 vdd.t1433 vdd.n760 0.0225448
R17206 vdd.n777 vdd.n776 0.0225448
R17207 vdd.t1431 vdd.n777 0.0225448
R17208 vdd.n792 vdd.n791 0.0225448
R17209 vdd.n789 vdd.n749 0.0225448
R17210 vdd.t87 vdd.n789 0.0225448
R17211 vdd.n784 vdd.n754 0.0225448
R17212 vdd.t1431 vdd.n754 0.0225448
R17213 vdd.n780 vdd.n779 0.0225448
R17214 vdd.n779 vdd.t1433 0.0225448
R17215 vdd.n769 vdd.n768 0.0225448
R17216 vdd.n3357 vdd.n3356 0.0225448
R17217 vdd.n3357 vdd.t1203 0.0225448
R17218 vdd.n3367 vdd.n3366 0.0225448
R17219 vdd.n3366 vdd.t265 0.0225448
R17220 vdd.n3369 vdd.n3346 0.0225448
R17221 vdd.t266 vdd.n3346 0.0225448
R17222 vdd.n3376 vdd.n3375 0.0225448
R17223 vdd.n3372 vdd.n3371 0.0225448
R17224 vdd.n3372 vdd.t819 0.0225448
R17225 vdd.n3381 vdd.n3380 0.0225448
R17226 vdd.n3380 vdd.t266 0.0225448
R17227 vdd.n3365 vdd.n3341 0.0225448
R17228 vdd.t265 vdd.n3365 0.0225448
R17229 vdd.n3363 vdd.n3362 0.0225448
R17230 vdd.n3311 vdd.n3310 0.0225448
R17231 vdd.n3311 vdd.t310 0.0225448
R17232 vdd.n3321 vdd.n3320 0.0225448
R17233 vdd.n3320 vdd.t1508 0.0225448
R17234 vdd.n3323 vdd.n3300 0.0225448
R17235 vdd.t1509 vdd.n3300 0.0225448
R17236 vdd.n3330 vdd.n3329 0.0225448
R17237 vdd.n3326 vdd.n3325 0.0225448
R17238 vdd.n3326 vdd.t436 0.0225448
R17239 vdd.n3335 vdd.n3334 0.0225448
R17240 vdd.n3334 vdd.t1509 0.0225448
R17241 vdd.n3319 vdd.n3295 0.0225448
R17242 vdd.t1508 vdd.n3319 0.0225448
R17243 vdd.n3317 vdd.n3316 0.0225448
R17244 vdd.n3404 vdd.n3403 0.0225448
R17245 vdd.n3404 vdd.t1124 0.0225448
R17246 vdd.n3414 vdd.n3413 0.0225448
R17247 vdd.n3413 vdd.t1137 0.0225448
R17248 vdd.n3416 vdd.n3393 0.0225448
R17249 vdd.t1135 vdd.n3393 0.0225448
R17250 vdd.n3423 vdd.n3422 0.0225448
R17251 vdd.n3419 vdd.n3418 0.0225448
R17252 vdd.n3419 vdd.t1332 0.0225448
R17253 vdd.n3428 vdd.n3427 0.0225448
R17254 vdd.n3427 vdd.t1135 0.0225448
R17255 vdd.n3412 vdd.n3388 0.0225448
R17256 vdd.t1137 vdd.n3412 0.0225448
R17257 vdd.n3410 vdd.n3409 0.0225448
R17258 vdd.n3452 vdd.n3451 0.0225448
R17259 vdd.n3452 vdd.t1061 0.0225448
R17260 vdd.n3462 vdd.n3461 0.0225448
R17261 vdd.n3461 vdd.t648 0.0225448
R17262 vdd.n3464 vdd.n3441 0.0225448
R17263 vdd.t649 vdd.n3441 0.0225448
R17264 vdd.n3471 vdd.n3470 0.0225448
R17265 vdd.n3467 vdd.n3466 0.0225448
R17266 vdd.n3467 vdd.t904 0.0225448
R17267 vdd.n3476 vdd.n3475 0.0225448
R17268 vdd.n3475 vdd.t649 0.0225448
R17269 vdd.n3460 vdd.n3436 0.0225448
R17270 vdd.t648 vdd.n3460 0.0225448
R17271 vdd.n3458 vdd.n3457 0.0225448
R17272 vdd.n3498 vdd.n3497 0.0225448
R17273 vdd.n3498 vdd.t1123 0.0225448
R17274 vdd.n3508 vdd.n3507 0.0225448
R17275 vdd.n3507 vdd.t830 0.0225448
R17276 vdd.n3510 vdd.n3487 0.0225448
R17277 vdd.t831 vdd.n3487 0.0225448
R17278 vdd.n3517 vdd.n3516 0.0225448
R17279 vdd.n3513 vdd.n3512 0.0225448
R17280 vdd.n3513 vdd.t488 0.0225448
R17281 vdd.n3522 vdd.n3521 0.0225448
R17282 vdd.n3521 vdd.t831 0.0225448
R17283 vdd.n3506 vdd.n3482 0.0225448
R17284 vdd.t830 vdd.n3506 0.0225448
R17285 vdd.n3504 vdd.n3503 0.0225448
R17286 vdd.n580 vdd.n579 0.0225448
R17287 vdd.n580 vdd.t748 0.0225448
R17288 vdd.n590 vdd.n589 0.0225448
R17289 vdd.n589 vdd.t1153 0.0225448
R17290 vdd.n592 vdd.n569 0.0225448
R17291 vdd.t1151 vdd.n569 0.0225448
R17292 vdd.n599 vdd.n598 0.0225448
R17293 vdd.n595 vdd.n594 0.0225448
R17294 vdd.n595 vdd.t30 0.0225448
R17295 vdd.n604 vdd.n603 0.0225448
R17296 vdd.n603 vdd.t1151 0.0225448
R17297 vdd.n588 vdd.n564 0.0225448
R17298 vdd.t1153 vdd.n588 0.0225448
R17299 vdd.n586 vdd.n585 0.0225448
R17300 vdd.n3593 vdd.n3592 0.0225448
R17301 vdd.n3593 vdd.t1382 0.0225448
R17302 vdd.n3603 vdd.n3602 0.0225448
R17303 vdd.n3602 vdd.t1428 0.0225448
R17304 vdd.n3605 vdd.n3582 0.0225448
R17305 vdd.t1429 vdd.n3582 0.0225448
R17306 vdd.n3612 vdd.n3611 0.0225448
R17307 vdd.n3608 vdd.n3607 0.0225448
R17308 vdd.n3608 vdd.t24 0.0225448
R17309 vdd.n3617 vdd.n3616 0.0225448
R17310 vdd.n3616 vdd.t1429 0.0225448
R17311 vdd.n3601 vdd.n3577 0.0225448
R17312 vdd.t1428 vdd.n3601 0.0225448
R17313 vdd.n3599 vdd.n3598 0.0225448
R17314 vdd.n3547 vdd.n3546 0.0225448
R17315 vdd.n3547 vdd.t1150 0.0225448
R17316 vdd.n3557 vdd.n3556 0.0225448
R17317 vdd.n3556 vdd.t1172 0.0225448
R17318 vdd.n3559 vdd.n3536 0.0225448
R17319 vdd.t1173 vdd.n3536 0.0225448
R17320 vdd.n3566 vdd.n3565 0.0225448
R17321 vdd.n3562 vdd.n3561 0.0225448
R17322 vdd.n3562 vdd.t986 0.0225448
R17323 vdd.n3571 vdd.n3570 0.0225448
R17324 vdd.n3570 vdd.t1173 0.0225448
R17325 vdd.n3555 vdd.n3531 0.0225448
R17326 vdd.t1172 vdd.n3555 0.0225448
R17327 vdd.n3553 vdd.n3552 0.0225448
R17328 vdd.n6607 vdd.n6606 0.0225448
R17329 vdd.n6607 vdd.t1095 0.0225448
R17330 vdd.n6617 vdd.n6616 0.0225448
R17331 vdd.n6616 vdd.t709 0.0225448
R17332 vdd.n6619 vdd.n6596 0.0225448
R17333 vdd.t707 vdd.n6596 0.0225448
R17334 vdd.n6626 vdd.n6625 0.0225448
R17335 vdd.n6622 vdd.n6621 0.0225448
R17336 vdd.n6622 vdd.t28 0.0225448
R17337 vdd.n6631 vdd.n6630 0.0225448
R17338 vdd.n6630 vdd.t707 0.0225448
R17339 vdd.n6615 vdd.n6591 0.0225448
R17340 vdd.t709 vdd.n6615 0.0225448
R17341 vdd.n6613 vdd.n6612 0.0225448
R17342 vdd.n6561 vdd.n6560 0.0225448
R17343 vdd.n6561 vdd.t1243 0.0225448
R17344 vdd.n6571 vdd.n6570 0.0225448
R17345 vdd.n6570 vdd.t549 0.0225448
R17346 vdd.n6573 vdd.n6550 0.0225448
R17347 vdd.t550 vdd.n6550 0.0225448
R17348 vdd.n6580 vdd.n6579 0.0225448
R17349 vdd.n6576 vdd.n6575 0.0225448
R17350 vdd.n6576 vdd.t1186 0.0225448
R17351 vdd.n6585 vdd.n6584 0.0225448
R17352 vdd.n6584 vdd.t550 0.0225448
R17353 vdd.n6569 vdd.n6545 0.0225448
R17354 vdd.t549 vdd.n6569 0.0225448
R17355 vdd.n6567 vdd.n6566 0.0225448
R17356 vdd.n9621 vdd.n9620 0.0225448
R17357 vdd.n9621 vdd.t706 0.0225448
R17358 vdd.n9631 vdd.n9630 0.0225448
R17359 vdd.n9630 vdd.t912 0.0225448
R17360 vdd.n9633 vdd.n9610 0.0225448
R17361 vdd.t910 vdd.n9610 0.0225448
R17362 vdd.n9640 vdd.n9639 0.0225448
R17363 vdd.n9636 vdd.n9635 0.0225448
R17364 vdd.n9636 vdd.t26 0.0225448
R17365 vdd.n9645 vdd.n9644 0.0225448
R17366 vdd.n9644 vdd.t910 0.0225448
R17367 vdd.n9629 vdd.n9605 0.0225448
R17368 vdd.t912 vdd.n9629 0.0225448
R17369 vdd.n9627 vdd.n9626 0.0225448
R17370 vdd.n9575 vdd.n9574 0.0225448
R17371 vdd.n9575 vdd.t237 0.0225448
R17372 vdd.n9585 vdd.n9584 0.0225448
R17373 vdd.n9584 vdd.t1113 0.0225448
R17374 vdd.n9587 vdd.n9564 0.0225448
R17375 vdd.t1114 vdd.n9564 0.0225448
R17376 vdd.n9594 vdd.n9593 0.0225448
R17377 vdd.n9590 vdd.n9589 0.0225448
R17378 vdd.n9590 vdd.t984 0.0225448
R17379 vdd.n9599 vdd.n9598 0.0225448
R17380 vdd.n9598 vdd.t1114 0.0225448
R17381 vdd.n9583 vdd.n9559 0.0225448
R17382 vdd.t1113 vdd.n9583 0.0225448
R17383 vdd.n9581 vdd.n9580 0.0225448
R17384 vdd.n9667 vdd.n9666 0.0225448
R17385 vdd.n9667 vdd.t1514 0.0225448
R17386 vdd.n9677 vdd.n9676 0.0225448
R17387 vdd.n9676 vdd.t1511 0.0225448
R17388 vdd.n9679 vdd.n9656 0.0225448
R17389 vdd.t1512 vdd.n9656 0.0225448
R17390 vdd.n9686 vdd.n9685 0.0225448
R17391 vdd.n9682 vdd.n9681 0.0225448
R17392 vdd.n9682 vdd.t1354 0.0225448
R17393 vdd.n9691 vdd.n9690 0.0225448
R17394 vdd.n9690 vdd.t1512 0.0225448
R17395 vdd.n9675 vdd.n9651 0.0225448
R17396 vdd.t1511 vdd.n9675 0.0225448
R17397 vdd.n9673 vdd.n9672 0.0225448
R17398 vdd.n9713 vdd.n9712 0.0225448
R17399 vdd.n9713 vdd.t71 0.0225448
R17400 vdd.n9723 vdd.n9722 0.0225448
R17401 vdd.n9722 vdd.t1387 0.0225448
R17402 vdd.n9725 vdd.n9702 0.0225448
R17403 vdd.t1388 vdd.n9702 0.0225448
R17404 vdd.n9732 vdd.n9731 0.0225448
R17405 vdd.n9728 vdd.n9727 0.0225448
R17406 vdd.n9728 vdd.t1322 0.0225448
R17407 vdd.n9737 vdd.n9736 0.0225448
R17408 vdd.n9736 vdd.t1388 0.0225448
R17409 vdd.n9721 vdd.n9697 0.0225448
R17410 vdd.t1387 vdd.n9721 0.0225448
R17411 vdd.n9719 vdd.n9718 0.0225448
R17412 vdd.n9811 vdd.n9810 0.0225448
R17413 vdd.n9811 vdd.t360 0.0225448
R17414 vdd.n9821 vdd.n9820 0.0225448
R17415 vdd.n9820 vdd.t727 0.0225448
R17416 vdd.n9823 vdd.n9800 0.0225448
R17417 vdd.t725 vdd.n9800 0.0225448
R17418 vdd.n9830 vdd.n9829 0.0225448
R17419 vdd.n9826 vdd.n9825 0.0225448
R17420 vdd.n9826 vdd.t478 0.0225448
R17421 vdd.n9835 vdd.n9834 0.0225448
R17422 vdd.n9834 vdd.t725 0.0225448
R17423 vdd.n9819 vdd.n9795 0.0225448
R17424 vdd.t727 vdd.n9819 0.0225448
R17425 vdd.n9817 vdd.n9816 0.0225448
R17426 vdd.n9857 vdd.n9856 0.0225448
R17427 vdd.n9857 vdd.t1284 0.0225448
R17428 vdd.n9867 vdd.n9866 0.0225448
R17429 vdd.n9866 vdd.t1179 0.0225448
R17430 vdd.n9869 vdd.n9846 0.0225448
R17431 vdd.t1180 vdd.n9846 0.0225448
R17432 vdd.n9876 vdd.n9875 0.0225448
R17433 vdd.n9872 vdd.n9871 0.0225448
R17434 vdd.n9872 vdd.t1059 0.0225448
R17435 vdd.n9881 vdd.n9880 0.0225448
R17436 vdd.n9880 vdd.t1180 0.0225448
R17437 vdd.n9865 vdd.n9841 0.0225448
R17438 vdd.t1179 vdd.n9865 0.0225448
R17439 vdd.n9863 vdd.n9862 0.0225448
R17440 vdd.n9903 vdd.n9902 0.0225448
R17441 vdd.n9903 vdd.t1023 0.0225448
R17442 vdd.n9913 vdd.n9912 0.0225448
R17443 vdd.n9912 vdd.t259 0.0225448
R17444 vdd.n9915 vdd.n9892 0.0225448
R17445 vdd.t257 vdd.n9892 0.0225448
R17446 vdd.n9922 vdd.n9921 0.0225448
R17447 vdd.n9918 vdd.n9917 0.0225448
R17448 vdd.n9918 vdd.t15 0.0225448
R17449 vdd.n9927 vdd.n9926 0.0225448
R17450 vdd.n9926 vdd.t257 0.0225448
R17451 vdd.n9911 vdd.n9887 0.0225448
R17452 vdd.t259 vdd.n9911 0.0225448
R17453 vdd.n9909 vdd.n9908 0.0225448
R17454 vdd.n9949 vdd.n9948 0.0225448
R17455 vdd.n9949 vdd.t960 0.0225448
R17456 vdd.n9959 vdd.n9958 0.0225448
R17457 vdd.n9958 vdd.t62 0.0225448
R17458 vdd.n9961 vdd.n9938 0.0225448
R17459 vdd.t60 vdd.n9938 0.0225448
R17460 vdd.n9968 vdd.n9967 0.0225448
R17461 vdd.n9964 vdd.n9963 0.0225448
R17462 vdd.n9964 vdd.t490 0.0225448
R17463 vdd.n9973 vdd.n9972 0.0225448
R17464 vdd.n9972 vdd.t60 0.0225448
R17465 vdd.n9957 vdd.n9933 0.0225448
R17466 vdd.t62 vdd.n9957 0.0225448
R17467 vdd.n9955 vdd.n9954 0.0225448
R17468 vdd.n10047 vdd.n10046 0.0225448
R17469 vdd.n10047 vdd.t548 0.0225448
R17470 vdd.n10057 vdd.n10056 0.0225448
R17471 vdd.n10056 vdd.t337 0.0225448
R17472 vdd.n10059 vdd.n10036 0.0225448
R17473 vdd.t338 vdd.n10036 0.0225448
R17474 vdd.n10066 vdd.n10065 0.0225448
R17475 vdd.n10062 vdd.n10061 0.0225448
R17476 vdd.n10062 vdd.t1334 0.0225448
R17477 vdd.n10071 vdd.n10070 0.0225448
R17478 vdd.n10070 vdd.t338 0.0225448
R17479 vdd.n10055 vdd.n10031 0.0225448
R17480 vdd.t337 vdd.n10055 0.0225448
R17481 vdd.n10053 vdd.n10052 0.0225448
R17482 vdd.n63 vdd.n62 0.0225448
R17483 vdd.n63 vdd.t422 0.0225448
R17484 vdd.n73 vdd.n72 0.0225448
R17485 vdd.n72 vdd.t242 0.0225448
R17486 vdd.n75 vdd.n52 0.0225448
R17487 vdd.t243 vdd.n52 0.0225448
R17488 vdd.n82 vdd.n81 0.0225448
R17489 vdd.n78 vdd.n77 0.0225448
R17490 vdd.n78 vdd.t1008 0.0225448
R17491 vdd.n87 vdd.n86 0.0225448
R17492 vdd.n86 vdd.t243 0.0225448
R17493 vdd.n71 vdd.n47 0.0225448
R17494 vdd.t242 vdd.n71 0.0225448
R17495 vdd.n69 vdd.n68 0.0225448
R17496 vdd.n17 vdd.n16 0.0225448
R17497 vdd.n17 vdd.t260 0.0225448
R17498 vdd.n27 vdd.n26 0.0225448
R17499 vdd.n26 vdd.t653 0.0225448
R17500 vdd.n29 vdd.n6 0.0225448
R17501 vdd.t651 vdd.n6 0.0225448
R17502 vdd.n36 vdd.n35 0.0225448
R17503 vdd.n32 vdd.n31 0.0225448
R17504 vdd.n32 vdd.t839 0.0225448
R17505 vdd.n41 vdd.n40 0.0225448
R17506 vdd.n40 vdd.t651 0.0225448
R17507 vdd.n25 vdd.n1 0.0225448
R17508 vdd.t653 vdd.n25 0.0225448
R17509 vdd.n23 vdd.n22 0.0225448
R17510 vdd.n10093 vdd.n10092 0.0225448
R17511 vdd.n10093 vdd.t1164 0.0225448
R17512 vdd.n10103 vdd.n10102 0.0225448
R17513 vdd.n10102 vdd.t1087 0.0225448
R17514 vdd.n10105 vdd.n10082 0.0225448
R17515 vdd.t1085 vdd.n10082 0.0225448
R17516 vdd.n10112 vdd.n10111 0.0225448
R17517 vdd.n10108 vdd.n10107 0.0225448
R17518 vdd.n10108 vdd.t568 0.0225448
R17519 vdd.n10117 vdd.n10116 0.0225448
R17520 vdd.n10116 vdd.t1085 0.0225448
R17521 vdd.n10101 vdd.n10077 0.0225448
R17522 vdd.t1087 vdd.n10101 0.0225448
R17523 vdd.n10099 vdd.n10098 0.0225448
R17524 vdd.n10141 vdd.n10140 0.0225448
R17525 vdd.n10141 vdd.t1438 0.0225448
R17526 vdd.n10151 vdd.n10150 0.0225448
R17527 vdd.n10150 vdd.t780 0.0225448
R17528 vdd.n10153 vdd.n10130 0.0225448
R17529 vdd.t781 vdd.n10130 0.0225448
R17530 vdd.n10160 vdd.n10159 0.0225448
R17531 vdd.n10156 vdd.n10155 0.0225448
R17532 vdd.n10156 vdd.t908 0.0225448
R17533 vdd.n10165 vdd.n10164 0.0225448
R17534 vdd.n10164 vdd.t781 0.0225448
R17535 vdd.n10149 vdd.n10125 0.0225448
R17536 vdd.t780 vdd.n10149 0.0225448
R17537 vdd.n10147 vdd.n10146 0.0225448
R17538 vdd.n10187 vdd.n10186 0.0225448
R17539 vdd.n10187 vdd.t418 0.0225448
R17540 vdd.n10197 vdd.n10196 0.0225448
R17541 vdd.n10196 vdd.t1020 0.0225448
R17542 vdd.n10199 vdd.n10176 0.0225448
R17543 vdd.t1021 vdd.n10176 0.0225448
R17544 vdd.n10206 vdd.n10205 0.0225448
R17545 vdd.n10202 vdd.n10201 0.0225448
R17546 vdd.n10202 vdd.t597 0.0225448
R17547 vdd.n10211 vdd.n10210 0.0225448
R17548 vdd.n10210 vdd.t1021 0.0225448
R17549 vdd.n10195 vdd.n10171 0.0225448
R17550 vdd.t1020 vdd.n10195 0.0225448
R17551 vdd.n10193 vdd.n10192 0.0225448
R17552 vdd.n10003 vdd.n10002 0.0225448
R17553 vdd.n10002 vdd.t694 0.0225448
R17554 vdd.n10005 vdd.n9991 0.0225448
R17555 vdd.t1397 vdd.n9991 0.0225448
R17556 vdd.n10008 vdd.n10007 0.0225448
R17557 vdd.t1398 vdd.n10008 0.0225448
R17558 vdd.n10023 vdd.n10022 0.0225448
R17559 vdd.n10020 vdd.n9980 0.0225448
R17560 vdd.t575 vdd.n10020 0.0225448
R17561 vdd.n10015 vdd.n9985 0.0225448
R17562 vdd.t1398 vdd.n9985 0.0225448
R17563 vdd.n10011 vdd.n10010 0.0225448
R17564 vdd.n10010 vdd.t1397 0.0225448
R17565 vdd.n10000 vdd.n9999 0.0225448
R17566 vdd.n10329 vdd.n10328 0.0225448
R17567 vdd.n10329 vdd.t702 0.0225448
R17568 vdd.n10339 vdd.n10338 0.0225448
R17569 vdd.n10338 vdd.t687 0.0225448
R17570 vdd.n10341 vdd.n10318 0.0225448
R17571 vdd.t688 vdd.n10318 0.0225448
R17572 vdd.n10348 vdd.n10347 0.0225448
R17573 vdd.n10344 vdd.n10343 0.0225448
R17574 vdd.n10344 vdd.t938 0.0225448
R17575 vdd.n10353 vdd.n10352 0.0225448
R17576 vdd.n10352 vdd.t688 0.0225448
R17577 vdd.n10337 vdd.n10313 0.0225448
R17578 vdd.t687 vdd.n10337 0.0225448
R17579 vdd.n10335 vdd.n10334 0.0225448
R17580 vdd.n10282 vdd.n10281 0.0225448
R17581 vdd.n10282 vdd.t502 0.0225448
R17582 vdd.n10292 vdd.n10291 0.0225448
R17583 vdd.n10291 vdd.t299 0.0225448
R17584 vdd.n10294 vdd.n10271 0.0225448
R17585 vdd.t300 vdd.n10271 0.0225448
R17586 vdd.n10301 vdd.n10300 0.0225448
R17587 vdd.n10297 vdd.n10296 0.0225448
R17588 vdd.n10297 vdd.t54 0.0225448
R17589 vdd.n10306 vdd.n10305 0.0225448
R17590 vdd.n10305 vdd.t300 0.0225448
R17591 vdd.n10290 vdd.n10266 0.0225448
R17592 vdd.t299 vdd.n10290 0.0225448
R17593 vdd.n10288 vdd.n10287 0.0225448
R17594 vdd.n10236 vdd.n10235 0.0225448
R17595 vdd.n10236 vdd.t659 0.0225448
R17596 vdd.n10246 vdd.n10245 0.0225448
R17597 vdd.n10245 vdd.t1416 0.0225448
R17598 vdd.n10248 vdd.n10225 0.0225448
R17599 vdd.t1417 vdd.n10225 0.0225448
R17600 vdd.n10255 vdd.n10254 0.0225448
R17601 vdd.n10251 vdd.n10250 0.0225448
R17602 vdd.n10251 vdd.t1379 0.0225448
R17603 vdd.n10260 vdd.n10259 0.0225448
R17604 vdd.n10259 vdd.t1417 0.0225448
R17605 vdd.n10244 vdd.n10220 0.0225448
R17606 vdd.t1416 vdd.n10244 0.0225448
R17607 vdd.n10242 vdd.n10241 0.0225448
R17608 vdd.n10376 vdd.n10375 0.0225448
R17609 vdd.n10376 vdd.t1138 0.0225448
R17610 vdd.n10386 vdd.n10385 0.0225448
R17611 vdd.n10385 vdd.t354 0.0225448
R17612 vdd.n10388 vdd.n10365 0.0225448
R17613 vdd.t355 vdd.n10365 0.0225448
R17614 vdd.n10395 vdd.n10394 0.0225448
R17615 vdd.n10391 vdd.n10390 0.0225448
R17616 vdd.n10391 vdd.t383 0.0225448
R17617 vdd.n10400 vdd.n10399 0.0225448
R17618 vdd.n10399 vdd.t355 0.0225448
R17619 vdd.n10384 vdd.n10360 0.0225448
R17620 vdd.t354 vdd.n10384 0.0225448
R17621 vdd.n10382 vdd.n10381 0.0225448
R17622 vdd.n10424 vdd.n10423 0.0225448
R17623 vdd.n10424 vdd.t1454 0.0225448
R17624 vdd.n10434 vdd.n10433 0.0225448
R17625 vdd.n10433 vdd.t1400 0.0225448
R17626 vdd.n10436 vdd.n10413 0.0225448
R17627 vdd.t1401 vdd.n10413 0.0225448
R17628 vdd.n10443 vdd.n10442 0.0225448
R17629 vdd.n10439 vdd.n10438 0.0225448
R17630 vdd.n10439 vdd.t846 0.0225448
R17631 vdd.n10448 vdd.n10447 0.0225448
R17632 vdd.n10447 vdd.t1401 0.0225448
R17633 vdd.n10432 vdd.n10408 0.0225448
R17634 vdd.t1400 vdd.n10432 0.0225448
R17635 vdd.n10430 vdd.n10429 0.0225448
R17636 vdd.n10470 vdd.n10469 0.0225448
R17637 vdd.n10470 vdd.t1257 0.0225448
R17638 vdd.n10480 vdd.n10479 0.0225448
R17639 vdd.n10479 vdd.t803 0.0225448
R17640 vdd.n10482 vdd.n10459 0.0225448
R17641 vdd.t804 vdd.n10459 0.0225448
R17642 vdd.n10489 vdd.n10488 0.0225448
R17643 vdd.n10485 vdd.n10484 0.0225448
R17644 vdd.n10485 vdd.t1306 0.0225448
R17645 vdd.n10494 vdd.n10493 0.0225448
R17646 vdd.n10493 vdd.t804 0.0225448
R17647 vdd.n10478 vdd.n10454 0.0225448
R17648 vdd.t803 vdd.n10478 0.0225448
R17649 vdd.n10476 vdd.n10475 0.0225448
R17650 vdd.n10564 vdd.n10563 0.0225448
R17651 vdd.n10564 vdd.t1366 0.0225448
R17652 vdd.n10574 vdd.n10573 0.0225448
R17653 vdd.n10573 vdd.t1260 0.0225448
R17654 vdd.n10576 vdd.n10553 0.0225448
R17655 vdd.t1261 vdd.n10553 0.0225448
R17656 vdd.n10583 vdd.n10582 0.0225448
R17657 vdd.n10579 vdd.n10578 0.0225448
R17658 vdd.n10579 vdd.t1004 0.0225448
R17659 vdd.n10588 vdd.n10587 0.0225448
R17660 vdd.n10587 vdd.t1261 0.0225448
R17661 vdd.n10572 vdd.n10548 0.0225448
R17662 vdd.t1260 vdd.n10572 0.0225448
R17663 vdd.n10570 vdd.n10569 0.0225448
R17664 vdd.n10518 vdd.n10517 0.0225448
R17665 vdd.n10518 vdd.t1102 0.0225448
R17666 vdd.n10528 vdd.n10527 0.0225448
R17667 vdd.n10527 vdd.t261 0.0225448
R17668 vdd.n10530 vdd.n10507 0.0225448
R17669 vdd.t262 vdd.n10507 0.0225448
R17670 vdd.n10537 vdd.n10536 0.0225448
R17671 vdd.n10533 vdd.n10532 0.0225448
R17672 vdd.n10533 vdd.t775 0.0225448
R17673 vdd.n10542 vdd.n10541 0.0225448
R17674 vdd.n10541 vdd.t262 0.0225448
R17675 vdd.n10526 vdd.n10502 0.0225448
R17676 vdd.t261 vdd.n10526 0.0225448
R17677 vdd.n10524 vdd.n10523 0.0225448
R17678 vdd.n10611 vdd.n10610 0.0225448
R17679 vdd.n10611 vdd.t1019 0.0225448
R17680 vdd.n10621 vdd.n10620 0.0225448
R17681 vdd.n10620 vdd.t1077 0.0225448
R17682 vdd.n10623 vdd.n10600 0.0225448
R17683 vdd.t1075 vdd.n10600 0.0225448
R17684 vdd.n10630 vdd.n10629 0.0225448
R17685 vdd.n10626 vdd.n10625 0.0225448
R17686 vdd.n10626 vdd.t1491 0.0225448
R17687 vdd.n10635 vdd.n10634 0.0225448
R17688 vdd.n10634 vdd.t1075 0.0225448
R17689 vdd.n10619 vdd.n10595 0.0225448
R17690 vdd.t1077 vdd.n10619 0.0225448
R17691 vdd.n10617 vdd.n10616 0.0225448
R17692 vdd.n10659 vdd.n10658 0.0225448
R17693 vdd.n10659 vdd.t253 0.0225448
R17694 vdd.n10669 vdd.n10668 0.0225448
R17695 vdd.n10668 vdd.t610 0.0225448
R17696 vdd.n10671 vdd.n10648 0.0225448
R17697 vdd.t608 vdd.n10648 0.0225448
R17698 vdd.n10678 vdd.n10677 0.0225448
R17699 vdd.n10674 vdd.n10673 0.0225448
R17700 vdd.n10674 vdd.t817 0.0225448
R17701 vdd.n10683 vdd.n10682 0.0225448
R17702 vdd.n10682 vdd.t608 0.0225448
R17703 vdd.n10667 vdd.n10643 0.0225448
R17704 vdd.t610 vdd.n10667 0.0225448
R17705 vdd.n10665 vdd.n10664 0.0225448
R17706 vdd.n10705 vdd.n10704 0.0225448
R17707 vdd.n10705 vdd.t292 0.0225448
R17708 vdd.n10715 vdd.n10714 0.0225448
R17709 vdd.n10714 vdd.t146 0.0225448
R17710 vdd.n10717 vdd.n10694 0.0225448
R17711 vdd.t147 vdd.n10694 0.0225448
R17712 vdd.n10724 vdd.n10723 0.0225448
R17713 vdd.n10720 vdd.n10719 0.0225448
R17714 vdd.n10720 vdd.t1352 0.0225448
R17715 vdd.n10729 vdd.n10728 0.0225448
R17716 vdd.n10728 vdd.t147 0.0225448
R17717 vdd.n10713 vdd.n10689 0.0225448
R17718 vdd.t146 vdd.n10713 0.0225448
R17719 vdd.n10711 vdd.n10710 0.0225448
R17720 vdd.n9767 vdd.n9766 0.0225448
R17721 vdd.n9766 vdd.t964 0.0225448
R17722 vdd.n9769 vdd.n9755 0.0225448
R17723 vdd.t1363 vdd.n9755 0.0225448
R17724 vdd.n9772 vdd.n9771 0.0225448
R17725 vdd.t1364 vdd.n9772 0.0225448
R17726 vdd.n9787 vdd.n9786 0.0225448
R17727 vdd.n9784 vdd.n9744 0.0225448
R17728 vdd.t1461 vdd.n9784 0.0225448
R17729 vdd.n9779 vdd.n9749 0.0225448
R17730 vdd.t1364 vdd.n9749 0.0225448
R17731 vdd.n9775 vdd.n9774 0.0225448
R17732 vdd.n9774 vdd.t1363 0.0225448
R17733 vdd.n9764 vdd.n9763 0.0225448
R17734 vdd.n10800 vdd.n10799 0.0225448
R17735 vdd.n10800 vdd.t742 0.0225448
R17736 vdd.n10810 vdd.n10809 0.0225448
R17737 vdd.n10809 vdd.t1234 0.0225448
R17738 vdd.n10812 vdd.n10789 0.0225448
R17739 vdd.t1235 vdd.n10789 0.0225448
R17740 vdd.n10819 vdd.n10818 0.0225448
R17741 vdd.n10815 vdd.n10814 0.0225448
R17742 vdd.n10815 vdd.t902 0.0225448
R17743 vdd.n10824 vdd.n10823 0.0225448
R17744 vdd.n10823 vdd.t1235 0.0225448
R17745 vdd.n10808 vdd.n10784 0.0225448
R17746 vdd.t1234 vdd.n10808 0.0225448
R17747 vdd.n10806 vdd.n10805 0.0225448
R17748 vdd.n10754 vdd.n10753 0.0225448
R17749 vdd.n10754 vdd.t1247 0.0225448
R17750 vdd.n10764 vdd.n10763 0.0225448
R17751 vdd.n10763 vdd.t1244 0.0225448
R17752 vdd.n10766 vdd.n10743 0.0225448
R17753 vdd.t1245 vdd.n10743 0.0225448
R17754 vdd.n10773 vdd.n10772 0.0225448
R17755 vdd.n10769 vdd.n10768 0.0225448
R17756 vdd.n10769 vdd.t629 0.0225448
R17757 vdd.n10778 vdd.n10777 0.0225448
R17758 vdd.n10777 vdd.t1245 0.0225448
R17759 vdd.n10762 vdd.n10738 0.0225448
R17760 vdd.t1244 vdd.n10762 0.0225448
R17761 vdd.n10760 vdd.n10759 0.0225448
R17762 vdd.n10847 vdd.n10846 0.0225448
R17763 vdd.n10847 vdd.t417 0.0225448
R17764 vdd.n10857 vdd.n10856 0.0225448
R17765 vdd.n10856 vdd.t1162 0.0225448
R17766 vdd.n10859 vdd.n10836 0.0225448
R17767 vdd.t1160 vdd.n10836 0.0225448
R17768 vdd.n10866 vdd.n10865 0.0225448
R17769 vdd.n10862 vdd.n10861 0.0225448
R17770 vdd.n10862 vdd.t480 0.0225448
R17771 vdd.n10871 vdd.n10870 0.0225448
R17772 vdd.n10870 vdd.t1160 0.0225448
R17773 vdd.n10855 vdd.n10831 0.0225448
R17774 vdd.t1162 vdd.n10855 0.0225448
R17775 vdd.n10853 vdd.n10852 0.0225448
R17776 vdd.n10895 vdd.n10894 0.0225448
R17777 vdd.n10895 vdd.t285 0.0225448
R17778 vdd.n10905 vdd.n10904 0.0225448
R17779 vdd.n10904 vdd.t948 0.0225448
R17780 vdd.n10907 vdd.n10884 0.0225448
R17781 vdd.t949 vdd.n10884 0.0225448
R17782 vdd.n10914 vdd.n10913 0.0225448
R17783 vdd.n10910 vdd.n10909 0.0225448
R17784 vdd.n10910 vdd.t936 0.0225448
R17785 vdd.n10919 vdd.n10918 0.0225448
R17786 vdd.n10918 vdd.t949 0.0225448
R17787 vdd.n10903 vdd.n10879 0.0225448
R17788 vdd.t948 vdd.n10903 0.0225448
R17789 vdd.n10901 vdd.n10900 0.0225448
R17790 vdd.n10941 vdd.n10940 0.0225448
R17791 vdd.n10941 vdd.t690 0.0225448
R17792 vdd.n10951 vdd.n10950 0.0225448
R17793 vdd.n10950 vdd.t1196 0.0225448
R17794 vdd.n10953 vdd.n10930 0.0225448
R17795 vdd.t1197 vdd.n10930 0.0225448
R17796 vdd.n10960 vdd.n10959 0.0225448
R17797 vdd.n10956 vdd.n10955 0.0225448
R17798 vdd.n10956 vdd.t5 0.0225448
R17799 vdd.n10965 vdd.n10964 0.0225448
R17800 vdd.n10964 vdd.t1197 0.0225448
R17801 vdd.n10949 vdd.n10925 0.0225448
R17802 vdd.t1196 vdd.n10949 0.0225448
R17803 vdd.n10947 vdd.n10946 0.0225448
R17804 vdd.n10990 vdd.n10989 0.0225448
R17805 vdd.n10999 vdd.n10998 0.0225448
R17806 vdd.n10998 vdd.t286 0.0225448
R17807 vdd.n11004 vdd.n11003 0.0225448
R17808 vdd.n11004 vdd.t288 0.0225448
R17809 vdd.n11007 vdd.n10979 0.0225448
R17810 vdd.n11007 vdd.t498 0.0225448
R17811 vdd.n10995 vdd.t821 0.0225448
R17812 vdd.t286 vdd.n10997 0.0225448
R17813 vdd.n11013 vdd.t288 0.0225448
R17814 vdd.n11011 vdd.n11010 0.0225448
R17815 vdd.n11014 vdd.n11013 0.0225448
R17816 vdd.n10997 vdd.n10974 0.0225448
R17817 vdd.n10995 vdd.n10994 0.0225448
R17818 vdd.n11035 vdd.n11034 0.0225448
R17819 vdd.n11044 vdd.n11043 0.0225448
R17820 vdd.n11043 vdd.t645 0.0225448
R17821 vdd.n11049 vdd.n11048 0.0225448
R17822 vdd.n11049 vdd.t647 0.0225448
R17823 vdd.n11052 vdd.n11024 0.0225448
R17824 vdd.n11052 vdd.t1251 0.0225448
R17825 vdd.n11040 vdd.t58 0.0225448
R17826 vdd.t645 vdd.n11042 0.0225448
R17827 vdd.n11058 vdd.t647 0.0225448
R17828 vdd.n11056 vdd.n11055 0.0225448
R17829 vdd.n11059 vdd.n11058 0.0225448
R17830 vdd.n11042 vdd.n11019 0.0225448
R17831 vdd.n11040 vdd.n11039 0.0225448
R17832 vdd.n11085 vdd.n11084 0.0225448
R17833 vdd.n11094 vdd.n11093 0.0225448
R17834 vdd.n11093 vdd.t733 0.0225448
R17835 vdd.n11099 vdd.n11098 0.0225448
R17836 vdd.n11099 vdd.t735 0.0225448
R17837 vdd.n11102 vdd.n11074 0.0225448
R17838 vdd.n11102 vdd.t538 0.0225448
R17839 vdd.n11090 vdd.t1499 0.0225448
R17840 vdd.t733 vdd.n11092 0.0225448
R17841 vdd.n11108 vdd.t735 0.0225448
R17842 vdd.n11106 vdd.n11105 0.0225448
R17843 vdd.n11109 vdd.n11108 0.0225448
R17844 vdd.n11092 vdd.n11069 0.0225448
R17845 vdd.n11090 vdd.n11089 0.0225448
R17846 vdd.n11131 vdd.n11130 0.0225448
R17847 vdd.n11140 vdd.n11139 0.0225448
R17848 vdd.n11139 vdd.t294 0.0225448
R17849 vdd.n11145 vdd.n11144 0.0225448
R17850 vdd.n11145 vdd.t293 0.0225448
R17851 vdd.n11148 vdd.n11120 0.0225448
R17852 vdd.n11148 vdd.t539 0.0225448
R17853 vdd.n11136 vdd.t996 0.0225448
R17854 vdd.t294 vdd.n11138 0.0225448
R17855 vdd.n11154 vdd.t293 0.0225448
R17856 vdd.n11152 vdd.n11151 0.0225448
R17857 vdd.n11155 vdd.n11154 0.0225448
R17858 vdd.n11138 vdd.n11115 0.0225448
R17859 vdd.n11136 vdd.n11135 0.0225448
R17860 vdd.n11179 vdd.n11178 0.0225448
R17861 vdd.n11188 vdd.n11187 0.0225448
R17862 vdd.n11187 vdd.t350 0.0225448
R17863 vdd.n11193 vdd.n11192 0.0225448
R17864 vdd.n11193 vdd.t352 0.0225448
R17865 vdd.n11196 vdd.n11168 0.0225448
R17866 vdd.n11196 vdd.t216 0.0225448
R17867 vdd.n11184 vdd.t1294 0.0225448
R17868 vdd.t350 vdd.n11186 0.0225448
R17869 vdd.n11202 vdd.t352 0.0225448
R17870 vdd.n11200 vdd.n11199 0.0225448
R17871 vdd.n11203 vdd.n11202 0.0225448
R17872 vdd.n11186 vdd.n11163 0.0225448
R17873 vdd.n11184 vdd.n11183 0.0225448
R17874 vdd.n441 vdd.n440 0.0225448
R17875 vdd.n444 vdd.n443 0.0225448
R17876 vdd.n443 vdd.t740 0.0225448
R17877 vdd.n449 vdd.n448 0.0225448
R17878 vdd.n449 vdd.t739 0.0225448
R17879 vdd.n452 vdd.n433 0.0225448
R17880 vdd.n452 vdd.t1122 0.0225448
R17881 vdd.n465 vdd.t579 0.0225448
R17882 vdd.n463 vdd.t740 0.0225448
R17883 vdd.n458 vdd.t739 0.0225448
R17884 vdd.n456 vdd.n455 0.0225448
R17885 vdd.n459 vdd.n458 0.0225448
R17886 vdd.n463 vdd.n462 0.0225448
R17887 vdd.n466 vdd.n465 0.0225448
R17888 vdd.n11226 vdd.n11225 0.0225448
R17889 vdd.n11235 vdd.n11234 0.0225448
R17890 vdd.n11234 vdd.t514 0.0225448
R17891 vdd.n11240 vdd.n11239 0.0225448
R17892 vdd.n11240 vdd.t513 0.0225448
R17893 vdd.n11243 vdd.n11215 0.0225448
R17894 vdd.n11243 vdd.t115 0.0225448
R17895 vdd.n11231 vdd.t965 0.0225448
R17896 vdd.t514 vdd.n11233 0.0225448
R17897 vdd.n11249 vdd.t513 0.0225448
R17898 vdd.n11247 vdd.n11246 0.0225448
R17899 vdd.n11250 vdd.n11249 0.0225448
R17900 vdd.n11233 vdd.n11210 0.0225448
R17901 vdd.n11231 vdd.n11230 0.0225448
R17902 vdd.n11271 vdd.n11270 0.0225448
R17903 vdd.n11280 vdd.n11279 0.0225448
R17904 vdd.n11279 vdd.t889 0.0225448
R17905 vdd.n11285 vdd.n11284 0.0225448
R17906 vdd.n11285 vdd.t891 0.0225448
R17907 vdd.n11288 vdd.n11260 0.0225448
R17908 vdd.n11288 vdd.t531 0.0225448
R17909 vdd.n11276 vdd.t796 0.0225448
R17910 vdd.t889 vdd.n11278 0.0225448
R17911 vdd.n11294 vdd.t891 0.0225448
R17912 vdd.n11292 vdd.n11291 0.0225448
R17913 vdd.n11295 vdd.n11294 0.0225448
R17914 vdd.n11278 vdd.n11255 0.0225448
R17915 vdd.n11276 vdd.n11275 0.0225448
R17916 vdd.n11317 vdd.n11316 0.0225448
R17917 vdd.n11326 vdd.n11325 0.0225448
R17918 vdd.n11325 vdd.t405 0.0225448
R17919 vdd.n11331 vdd.n11330 0.0225448
R17920 vdd.n11331 vdd.t407 0.0225448
R17921 vdd.n11334 vdd.n11306 0.0225448
R17922 vdd.n11334 vdd.t1037 0.0225448
R17923 vdd.n11322 vdd.t1377 0.0225448
R17924 vdd.t405 vdd.n11324 0.0225448
R17925 vdd.n11340 vdd.t407 0.0225448
R17926 vdd.n11338 vdd.n11337 0.0225448
R17927 vdd.n11341 vdd.n11340 0.0225448
R17928 vdd.n11324 vdd.n11301 0.0225448
R17929 vdd.n11322 vdd.n11321 0.0225448
R17930 vdd.n11368 vdd.n11367 0.0225448
R17931 vdd.n11377 vdd.n11376 0.0225448
R17932 vdd.n11376 vdd.t1145 0.0225448
R17933 vdd.n11382 vdd.n11381 0.0225448
R17934 vdd.n11382 vdd.t1144 0.0225448
R17935 vdd.n11385 vdd.n11357 0.0225448
R17936 vdd.n11385 vdd.t1147 0.0225448
R17937 vdd.n11373 vdd.t199 0.0225448
R17938 vdd.t1145 vdd.n11375 0.0225448
R17939 vdd.n11391 vdd.t1144 0.0225448
R17940 vdd.n11389 vdd.n11388 0.0225448
R17941 vdd.n11392 vdd.n11391 0.0225448
R17942 vdd.n11375 vdd.n11352 0.0225448
R17943 vdd.n11373 vdd.n11372 0.0225448
R17944 vdd.n11414 vdd.n11413 0.0225448
R17945 vdd.n11423 vdd.n11422 0.0225448
R17946 vdd.n11422 vdd.t282 0.0225448
R17947 vdd.n11428 vdd.n11427 0.0225448
R17948 vdd.n11428 vdd.t281 0.0225448
R17949 vdd.n11431 vdd.n11403 0.0225448
R17950 vdd.n11431 vdd.t958 0.0225448
R17951 vdd.n11419 vdd.t850 0.0225448
R17952 vdd.t282 vdd.n11421 0.0225448
R17953 vdd.n11437 vdd.t281 0.0225448
R17954 vdd.n11435 vdd.n11434 0.0225448
R17955 vdd.n11438 vdd.n11437 0.0225448
R17956 vdd.n11421 vdd.n11398 0.0225448
R17957 vdd.n11419 vdd.n11418 0.0225448
R17958 vdd.n11462 vdd.n11461 0.0225448
R17959 vdd.n11471 vdd.n11470 0.0225448
R17960 vdd.n11470 vdd.t1521 0.0225448
R17961 vdd.n11476 vdd.n11475 0.0225448
R17962 vdd.n11476 vdd.t1523 0.0225448
R17963 vdd.n11479 vdd.n11451 0.0225448
R17964 vdd.n11479 vdd.t1242 0.0225448
R17965 vdd.n11467 vdd.t1340 0.0225448
R17966 vdd.t1521 vdd.n11469 0.0225448
R17967 vdd.n11485 vdd.t1523 0.0225448
R17968 vdd.n11483 vdd.n11482 0.0225448
R17969 vdd.n11486 vdd.n11485 0.0225448
R17970 vdd.n11469 vdd.n11446 0.0225448
R17971 vdd.n11467 vdd.n11466 0.0225448
R17972 vdd.n11508 vdd.n11507 0.0225448
R17973 vdd.n11517 vdd.n11516 0.0225448
R17974 vdd.n11516 vdd.t270 0.0225448
R17975 vdd.n11522 vdd.n11521 0.0225448
R17976 vdd.n11522 vdd.t272 0.0225448
R17977 vdd.n11525 vdd.n11497 0.0225448
R17978 vdd.n11525 vdd.t273 0.0225448
R17979 vdd.n11513 vdd.t811 0.0225448
R17980 vdd.t270 vdd.n11515 0.0225448
R17981 vdd.n11531 vdd.t272 0.0225448
R17982 vdd.n11529 vdd.n11528 0.0225448
R17983 vdd.n11532 vdd.n11531 0.0225448
R17984 vdd.n11515 vdd.n11492 0.0225448
R17985 vdd.n11513 vdd.n11512 0.0225448
R17986 vdd.n11553 vdd.n11552 0.0225448
R17987 vdd.n11562 vdd.n11561 0.0225448
R17988 vdd.n11561 vdd.t1439 0.0225448
R17989 vdd.n11567 vdd.n11566 0.0225448
R17990 vdd.n11567 vdd.t1441 0.0225448
R17991 vdd.n11570 vdd.n11542 0.0225448
R17992 vdd.n11570 vdd.t307 0.0225448
R17993 vdd.n11558 vdd.t794 0.0225448
R17994 vdd.t1439 vdd.n11560 0.0225448
R17995 vdd.n11576 vdd.t1441 0.0225448
R17996 vdd.n11574 vdd.n11573 0.0225448
R17997 vdd.n11577 vdd.n11576 0.0225448
R17998 vdd.n11560 vdd.n11537 0.0225448
R17999 vdd.n11558 vdd.n11557 0.0225448
R18000 vdd.n11603 vdd.n11602 0.0225448
R18001 vdd.n11612 vdd.n11611 0.0225448
R18002 vdd.n11611 vdd.t1390 0.0225448
R18003 vdd.n11617 vdd.n11616 0.0225448
R18004 vdd.n11617 vdd.t1392 0.0225448
R18005 vdd.n11620 vdd.n11592 0.0225448
R18006 vdd.n11620 vdd.t535 0.0225448
R18007 vdd.n11608 vdd.t1286 0.0225448
R18008 vdd.t1390 vdd.n11610 0.0225448
R18009 vdd.n11626 vdd.t1392 0.0225448
R18010 vdd.n11624 vdd.n11623 0.0225448
R18011 vdd.n11627 vdd.n11626 0.0225448
R18012 vdd.n11610 vdd.n11587 0.0225448
R18013 vdd.n11608 vdd.n11607 0.0225448
R18014 vdd.n11649 vdd.n11648 0.0225448
R18015 vdd.n11658 vdd.n11657 0.0225448
R18016 vdd.n11657 vdd.t1248 0.0225448
R18017 vdd.n11663 vdd.n11662 0.0225448
R18018 vdd.n11663 vdd.t1250 0.0225448
R18019 vdd.n11666 vdd.n11638 0.0225448
R18020 vdd.n11666 vdd.t641 0.0225448
R18021 vdd.n11654 vdd.t994 0.0225448
R18022 vdd.t1248 vdd.n11656 0.0225448
R18023 vdd.n11672 vdd.t1250 0.0225448
R18024 vdd.n11670 vdd.n11669 0.0225448
R18025 vdd.n11673 vdd.n11672 0.0225448
R18026 vdd.n11656 vdd.n11633 0.0225448
R18027 vdd.n11654 vdd.n11653 0.0225448
R18028 vdd.n11697 vdd.n11696 0.0225448
R18029 vdd.n11706 vdd.n11705 0.0225448
R18030 vdd.n11705 vdd.t528 0.0225448
R18031 vdd.n11711 vdd.n11710 0.0225448
R18032 vdd.n11711 vdd.t530 0.0225448
R18033 vdd.n11714 vdd.n11686 0.0225448
R18034 vdd.n11714 vdd.t1120 0.0225448
R18035 vdd.n11702 vdd.t1338 0.0225448
R18036 vdd.t528 vdd.n11704 0.0225448
R18037 vdd.n11720 vdd.t530 0.0225448
R18038 vdd.n11718 vdd.n11717 0.0225448
R18039 vdd.n11721 vdd.n11720 0.0225448
R18040 vdd.n11704 vdd.n11681 0.0225448
R18041 vdd.n11702 vdd.n11701 0.0225448
R18042 vdd.n206 vdd.n205 0.0225448
R18043 vdd.n209 vdd.n208 0.0225448
R18044 vdd.n208 vdd.t141 0.0225448
R18045 vdd.n214 vdd.n213 0.0225448
R18046 vdd.n214 vdd.t140 0.0225448
R18047 vdd.n217 vdd.n198 0.0225448
R18048 vdd.n217 vdd.t1381 0.0225448
R18049 vdd.n230 vdd.t577 0.0225448
R18050 vdd.n228 vdd.t141 0.0225448
R18051 vdd.n223 vdd.t140 0.0225448
R18052 vdd.n221 vdd.n220 0.0225448
R18053 vdd.n224 vdd.n223 0.0225448
R18054 vdd.n228 vdd.n227 0.0225448
R18055 vdd.n231 vdd.n230 0.0225448
R18056 vdd.n11744 vdd.n11743 0.0225448
R18057 vdd.n11753 vdd.n11752 0.0225448
R18058 vdd.n11752 vdd.t357 0.0225448
R18059 vdd.n11758 vdd.n11757 0.0225448
R18060 vdd.n11758 vdd.t359 0.0225448
R18061 vdd.n11761 vdd.n11733 0.0225448
R18062 vdd.n11761 vdd.t49 0.0225448
R18063 vdd.n11749 vdd.t1014 0.0225448
R18064 vdd.t357 vdd.n11751 0.0225448
R18065 vdd.n11767 vdd.t359 0.0225448
R18066 vdd.n11765 vdd.n11764 0.0225448
R18067 vdd.n11768 vdd.n11767 0.0225448
R18068 vdd.n11751 vdd.n11728 0.0225448
R18069 vdd.n11749 vdd.n11748 0.0225448
R18070 vdd.n11789 vdd.n11788 0.0225448
R18071 vdd.n11798 vdd.n11797 0.0225448
R18072 vdd.n11797 vdd.t104 0.0225448
R18073 vdd.n11803 vdd.n11802 0.0225448
R18074 vdd.n11803 vdd.t106 0.0225448
R18075 vdd.n11806 vdd.n11778 0.0225448
R18076 vdd.n11806 vdd.t1396 0.0225448
R18077 vdd.n11794 vdd.t792 0.0225448
R18078 vdd.t104 vdd.n11796 0.0225448
R18079 vdd.n11812 vdd.t106 0.0225448
R18080 vdd.n11810 vdd.n11809 0.0225448
R18081 vdd.n11813 vdd.n11812 0.0225448
R18082 vdd.n11796 vdd.n11773 0.0225448
R18083 vdd.n11794 vdd.n11793 0.0225448
R18084 vdd.n11839 vdd.n11838 0.0225448
R18085 vdd.n11848 vdd.n11847 0.0225448
R18086 vdd.n11847 vdd.t316 0.0225448
R18087 vdd.n11853 vdd.n11852 0.0225448
R18088 vdd.n11853 vdd.t315 0.0225448
R18089 vdd.n11856 vdd.n11828 0.0225448
R18090 vdd.n11856 vdd.t1271 0.0225448
R18091 vdd.n11844 vdd.t1320 0.0225448
R18092 vdd.t316 vdd.n11846 0.0225448
R18093 vdd.n11862 vdd.t315 0.0225448
R18094 vdd.n11860 vdd.n11859 0.0225448
R18095 vdd.n11863 vdd.n11862 0.0225448
R18096 vdd.n11846 vdd.n11823 0.0225448
R18097 vdd.n11844 vdd.n11843 0.0225448
R18098 vdd.n11885 vdd.n11884 0.0225448
R18099 vdd.n11894 vdd.n11893 0.0225448
R18100 vdd.n11893 vdd.t752 0.0225448
R18101 vdd.n11899 vdd.n11898 0.0225448
R18102 vdd.n11899 vdd.t754 0.0225448
R18103 vdd.n11902 vdd.n11874 0.0225448
R18104 vdd.n11902 vdd.t619 0.0225448
R18105 vdd.n11890 vdd.t813 0.0225448
R18106 vdd.t752 vdd.n11892 0.0225448
R18107 vdd.n11908 vdd.t754 0.0225448
R18108 vdd.n11906 vdd.n11905 0.0225448
R18109 vdd.n11909 vdd.n11908 0.0225448
R18110 vdd.n11892 vdd.n11869 0.0225448
R18111 vdd.n11890 vdd.n11889 0.0225448
R18112 vdd.n11933 vdd.n11932 0.0225448
R18113 vdd.n11942 vdd.n11941 0.0225448
R18114 vdd.n11941 vdd.t340 0.0225448
R18115 vdd.n11947 vdd.n11946 0.0225448
R18116 vdd.n11947 vdd.t342 0.0225448
R18117 vdd.n11950 vdd.n11922 0.0225448
R18118 vdd.n11950 vdd.t1071 0.0225448
R18119 vdd.n11938 vdd.t1292 0.0225448
R18120 vdd.t340 vdd.n11940 0.0225448
R18121 vdd.n11956 vdd.t342 0.0225448
R18122 vdd.n11954 vdd.n11953 0.0225448
R18123 vdd.n11957 vdd.n11956 0.0225448
R18124 vdd.n11940 vdd.n11917 0.0225448
R18125 vdd.n11938 vdd.n11937 0.0225448
R18126 vdd.n7484 vdd.n7436 0.0216765
R18127 vdd.n7484 vdd.n7483 0.0216765
R18128 vdd.n7249 vdd.n7201 0.0216765
R18129 vdd.n7249 vdd.n7248 0.0216765
R18130 vdd.n7059 vdd.n7011 0.0216765
R18131 vdd.n7059 vdd.n7058 0.0216765
R18132 vdd.n6823 vdd.n6775 0.0216765
R18133 vdd.n6823 vdd.n6822 0.0216765
R18134 vdd.n4470 vdd.n4422 0.0216765
R18135 vdd.n4470 vdd.n4469 0.0216765
R18136 vdd.n4235 vdd.n4187 0.0216765
R18137 vdd.n4235 vdd.n4234 0.0216765
R18138 vdd.n4045 vdd.n3997 0.0216765
R18139 vdd.n4045 vdd.n4044 0.0216765
R18140 vdd.n3809 vdd.n3761 0.0216765
R18141 vdd.n3809 vdd.n3808 0.0216765
R18142 vdd.n1456 vdd.n1408 0.0216765
R18143 vdd.n1456 vdd.n1455 0.0216765
R18144 vdd.n1221 vdd.n1173 0.0216765
R18145 vdd.n1221 vdd.n1220 0.0216765
R18146 vdd.n1031 vdd.n983 0.0216765
R18147 vdd.n1031 vdd.n1030 0.0216765
R18148 vdd.n795 vdd.n747 0.0216765
R18149 vdd.n795 vdd.n794 0.0216765
R18150 vdd.n10026 vdd.n9978 0.0216765
R18151 vdd.n10026 vdd.n10025 0.0216765
R18152 vdd.n9790 vdd.n9742 0.0216765
R18153 vdd.n9790 vdd.n9789 0.0216765
R18154 vdd.n468 vdd.n420 0.0216765
R18155 vdd.n468 vdd.n467 0.0216765
R18156 vdd.n233 vdd.n185 0.0216765
R18157 vdd.n233 vdd.n232 0.0216765
R18158 vdd.n111 vdd.n110 0.0196536
R18159 vdd.n157 vdd.n156 0.0196536
R18160 vdd.n254 vdd.n253 0.0196536
R18161 vdd.n300 vdd.n299 0.0196536
R18162 vdd.n346 vdd.n345 0.0196536
R18163 vdd.n392 vdd.n391 0.0196536
R18164 vdd.n489 vdd.n488 0.0196536
R18165 vdd.n535 vdd.n534 0.0196536
R18166 vdd.n7127 vdd.n7126 0.0196536
R18167 vdd.n7173 vdd.n7172 0.0196536
R18168 vdd.n7270 vdd.n7269 0.0196536
R18169 vdd.n7316 vdd.n7315 0.0196536
R18170 vdd.n7362 vdd.n7361 0.0196536
R18171 vdd.n7408 vdd.n7407 0.0196536
R18172 vdd.n7505 vdd.n7504 0.0196536
R18173 vdd.n6654 vdd.n6653 0.0196536
R18174 vdd.n7549 vdd.n7548 0.0196536
R18175 vdd.n7594 vdd.n7593 0.0196536
R18176 vdd.n7644 vdd.n7643 0.0196536
R18177 vdd.n7690 vdd.n7689 0.0196536
R18178 vdd.n7738 vdd.n7737 0.0196536
R18179 vdd.n7457 vdd.n7455 0.0196536
R18180 vdd.n7785 vdd.n7784 0.0196536
R18181 vdd.n7830 vdd.n7829 0.0196536
R18182 vdd.n7876 vdd.n7875 0.0196536
R18183 vdd.n7927 vdd.n7926 0.0196536
R18184 vdd.n7973 vdd.n7972 0.0196536
R18185 vdd.n8021 vdd.n8020 0.0196536
R18186 vdd.n8067 vdd.n8066 0.0196536
R18187 vdd.n8112 vdd.n8111 0.0196536
R18188 vdd.n8162 vdd.n8161 0.0196536
R18189 vdd.n8208 vdd.n8207 0.0196536
R18190 vdd.n8256 vdd.n8255 0.0196536
R18191 vdd.n7222 vdd.n7220 0.0196536
R18192 vdd.n8303 vdd.n8302 0.0196536
R18193 vdd.n8348 vdd.n8347 0.0196536
R18194 vdd.n8398 vdd.n8397 0.0196536
R18195 vdd.n8444 vdd.n8443 0.0196536
R18196 vdd.n8492 vdd.n8491 0.0196536
R18197 vdd.n4113 vdd.n4112 0.0196536
R18198 vdd.n4159 vdd.n4158 0.0196536
R18199 vdd.n4256 vdd.n4255 0.0196536
R18200 vdd.n4302 vdd.n4301 0.0196536
R18201 vdd.n4348 vdd.n4347 0.0196536
R18202 vdd.n4394 vdd.n4393 0.0196536
R18203 vdd.n4491 vdd.n4490 0.0196536
R18204 vdd.n3640 vdd.n3639 0.0196536
R18205 vdd.n4535 vdd.n4534 0.0196536
R18206 vdd.n4580 vdd.n4579 0.0196536
R18207 vdd.n4630 vdd.n4629 0.0196536
R18208 vdd.n4676 vdd.n4675 0.0196536
R18209 vdd.n4724 vdd.n4723 0.0196536
R18210 vdd.n4443 vdd.n4441 0.0196536
R18211 vdd.n4771 vdd.n4770 0.0196536
R18212 vdd.n4816 vdd.n4815 0.0196536
R18213 vdd.n4862 vdd.n4861 0.0196536
R18214 vdd.n4913 vdd.n4912 0.0196536
R18215 vdd.n4959 vdd.n4958 0.0196536
R18216 vdd.n5007 vdd.n5006 0.0196536
R18217 vdd.n5053 vdd.n5052 0.0196536
R18218 vdd.n5098 vdd.n5097 0.0196536
R18219 vdd.n5148 vdd.n5147 0.0196536
R18220 vdd.n5194 vdd.n5193 0.0196536
R18221 vdd.n5242 vdd.n5241 0.0196536
R18222 vdd.n4208 vdd.n4206 0.0196536
R18223 vdd.n5289 vdd.n5288 0.0196536
R18224 vdd.n5334 vdd.n5333 0.0196536
R18225 vdd.n5384 vdd.n5383 0.0196536
R18226 vdd.n5430 vdd.n5429 0.0196536
R18227 vdd.n5478 vdd.n5477 0.0196536
R18228 vdd.n1099 vdd.n1098 0.0196536
R18229 vdd.n1145 vdd.n1144 0.0196536
R18230 vdd.n1242 vdd.n1241 0.0196536
R18231 vdd.n1288 vdd.n1287 0.0196536
R18232 vdd.n1334 vdd.n1333 0.0196536
R18233 vdd.n1380 vdd.n1379 0.0196536
R18234 vdd.n1477 vdd.n1476 0.0196536
R18235 vdd.n626 vdd.n625 0.0196536
R18236 vdd.n1521 vdd.n1520 0.0196536
R18237 vdd.n1566 vdd.n1565 0.0196536
R18238 vdd.n1616 vdd.n1615 0.0196536
R18239 vdd.n1662 vdd.n1661 0.0196536
R18240 vdd.n1710 vdd.n1709 0.0196536
R18241 vdd.n1429 vdd.n1427 0.0196536
R18242 vdd.n1757 vdd.n1756 0.0196536
R18243 vdd.n1802 vdd.n1801 0.0196536
R18244 vdd.n1848 vdd.n1847 0.0196536
R18245 vdd.n1899 vdd.n1898 0.0196536
R18246 vdd.n1945 vdd.n1944 0.0196536
R18247 vdd.n1993 vdd.n1992 0.0196536
R18248 vdd.n2039 vdd.n2038 0.0196536
R18249 vdd.n2084 vdd.n2083 0.0196536
R18250 vdd.n2134 vdd.n2133 0.0196536
R18251 vdd.n2180 vdd.n2179 0.0196536
R18252 vdd.n2228 vdd.n2227 0.0196536
R18253 vdd.n1194 vdd.n1192 0.0196536
R18254 vdd.n2275 vdd.n2274 0.0196536
R18255 vdd.n2320 vdd.n2319 0.0196536
R18256 vdd.n2370 vdd.n2369 0.0196536
R18257 vdd.n2416 vdd.n2415 0.0196536
R18258 vdd.n2464 vdd.n2463 0.0196536
R18259 vdd.n10989 vdd.n10988 0.0196536
R18260 vdd.n11034 vdd.n11033 0.0196536
R18261 vdd.n11084 vdd.n11083 0.0196536
R18262 vdd.n11130 vdd.n11129 0.0196536
R18263 vdd.n11178 vdd.n11177 0.0196536
R18264 vdd.n441 vdd.n439 0.0196536
R18265 vdd.n11225 vdd.n11224 0.0196536
R18266 vdd.n11270 vdd.n11269 0.0196536
R18267 vdd.n11316 vdd.n11315 0.0196536
R18268 vdd.n11367 vdd.n11366 0.0196536
R18269 vdd.n11413 vdd.n11412 0.0196536
R18270 vdd.n11461 vdd.n11460 0.0196536
R18271 vdd.n11507 vdd.n11506 0.0196536
R18272 vdd.n11552 vdd.n11551 0.0196536
R18273 vdd.n11602 vdd.n11601 0.0196536
R18274 vdd.n11648 vdd.n11647 0.0196536
R18275 vdd.n11696 vdd.n11695 0.0196536
R18276 vdd.n206 vdd.n204 0.0196536
R18277 vdd.n11743 vdd.n11742 0.0196536
R18278 vdd.n11788 vdd.n11787 0.0196536
R18279 vdd.n11838 vdd.n11837 0.0196536
R18280 vdd.n11884 vdd.n11883 0.0196536
R18281 vdd.n11932 vdd.n11931 0.0196536
R18282 vdd.n11973 vdd.n11972 0.0196151
R18283 vdd.n11991 vdd.n11990 0.0196151
R18284 vdd.n133 vdd.n100 0.0196151
R18285 vdd.n179 vdd.n146 0.0196151
R18286 vdd.n276 vdd.n243 0.0196151
R18287 vdd.n322 vdd.n289 0.0196151
R18288 vdd.n368 vdd.n335 0.0196151
R18289 vdd.n414 vdd.n381 0.0196151
R18290 vdd.n511 vdd.n478 0.0196151
R18291 vdd.n557 vdd.n524 0.0196151
R18292 vdd.n6706 vdd.n6698 0.0196151
R18293 vdd.n6719 vdd.n6691 0.0196151
R18294 vdd.n6752 vdd.n6744 0.0196151
R18295 vdd.n6765 vdd.n6737 0.0196151
R18296 vdd.n6850 vdd.n6842 0.0196151
R18297 vdd.n6863 vdd.n6835 0.0196151
R18298 vdd.n6896 vdd.n6888 0.0196151
R18299 vdd.n6909 vdd.n6881 0.0196151
R18300 vdd.n6942 vdd.n6934 0.0196151
R18301 vdd.n6955 vdd.n6927 0.0196151
R18302 vdd.n6988 vdd.n6980 0.0196151
R18303 vdd.n7001 vdd.n6973 0.0196151
R18304 vdd.n7086 vdd.n7078 0.0196151
R18305 vdd.n7099 vdd.n7071 0.0196151
R18306 vdd.n8544 vdd.n8536 0.0196151
R18307 vdd.n8557 vdd.n8529 0.0196151
R18308 vdd.n7149 vdd.n7116 0.0196151
R18309 vdd.n7195 vdd.n7162 0.0196151
R18310 vdd.n7292 vdd.n7259 0.0196151
R18311 vdd.n7338 vdd.n7305 0.0196151
R18312 vdd.n7384 vdd.n7351 0.0196151
R18313 vdd.n7430 vdd.n7397 0.0196151
R18314 vdd.n7527 vdd.n7494 0.0196151
R18315 vdd.n6676 vdd.n6643 0.0196151
R18316 vdd.n7571 vdd.n7538 0.0196151
R18317 vdd.n7616 vdd.n7583 0.0196151
R18318 vdd.n7666 vdd.n7633 0.0196151
R18319 vdd.n7712 vdd.n7679 0.0196151
R18320 vdd.n7760 vdd.n7727 0.0196151
R18321 vdd.n7472 vdd.n7448 0.0196151
R18322 vdd.n7807 vdd.n7774 0.0196151
R18323 vdd.n7852 vdd.n7819 0.0196151
R18324 vdd.n7898 vdd.n7865 0.0196151
R18325 vdd.n7949 vdd.n7916 0.0196151
R18326 vdd.n7995 vdd.n7962 0.0196151
R18327 vdd.n8043 vdd.n8010 0.0196151
R18328 vdd.n8089 vdd.n8056 0.0196151
R18329 vdd.n8134 vdd.n8101 0.0196151
R18330 vdd.n8184 vdd.n8151 0.0196151
R18331 vdd.n8230 vdd.n8197 0.0196151
R18332 vdd.n8278 vdd.n8245 0.0196151
R18333 vdd.n7237 vdd.n7213 0.0196151
R18334 vdd.n8325 vdd.n8292 0.0196151
R18335 vdd.n8370 vdd.n8337 0.0196151
R18336 vdd.n8420 vdd.n8387 0.0196151
R18337 vdd.n8466 vdd.n8433 0.0196151
R18338 vdd.n8514 vdd.n8481 0.0196151
R18339 vdd.n8637 vdd.n8629 0.0196151
R18340 vdd.n8650 vdd.n8622 0.0196151
R18341 vdd.n8591 vdd.n8583 0.0196151
R18342 vdd.n8604 vdd.n8576 0.0196151
R18343 vdd.n8684 vdd.n8676 0.0196151
R18344 vdd.n8697 vdd.n8669 0.0196151
R18345 vdd.n8732 vdd.n8724 0.0196151
R18346 vdd.n8745 vdd.n8717 0.0196151
R18347 vdd.n8778 vdd.n8770 0.0196151
R18348 vdd.n8791 vdd.n8763 0.0196151
R18349 vdd.n7034 vdd.n7033 0.0196151
R18350 vdd.n7055 vdd.n7054 0.0196151
R18351 vdd.n8920 vdd.n8912 0.0196151
R18352 vdd.n8933 vdd.n8905 0.0196151
R18353 vdd.n8873 vdd.n8865 0.0196151
R18354 vdd.n8886 vdd.n8858 0.0196151
R18355 vdd.n8827 vdd.n8819 0.0196151
R18356 vdd.n8840 vdd.n8812 0.0196151
R18357 vdd.n8967 vdd.n8959 0.0196151
R18358 vdd.n8980 vdd.n8952 0.0196151
R18359 vdd.n9015 vdd.n9007 0.0196151
R18360 vdd.n9028 vdd.n9000 0.0196151
R18361 vdd.n9061 vdd.n9053 0.0196151
R18362 vdd.n9074 vdd.n9046 0.0196151
R18363 vdd.n9155 vdd.n9147 0.0196151
R18364 vdd.n9168 vdd.n9140 0.0196151
R18365 vdd.n9109 vdd.n9101 0.0196151
R18366 vdd.n9122 vdd.n9094 0.0196151
R18367 vdd.n9202 vdd.n9194 0.0196151
R18368 vdd.n9215 vdd.n9187 0.0196151
R18369 vdd.n9250 vdd.n9242 0.0196151
R18370 vdd.n9263 vdd.n9235 0.0196151
R18371 vdd.n9296 vdd.n9288 0.0196151
R18372 vdd.n9309 vdd.n9281 0.0196151
R18373 vdd.n6798 vdd.n6797 0.0196151
R18374 vdd.n6819 vdd.n6818 0.0196151
R18375 vdd.n9391 vdd.n9383 0.0196151
R18376 vdd.n9404 vdd.n9376 0.0196151
R18377 vdd.n9345 vdd.n9337 0.0196151
R18378 vdd.n9358 vdd.n9330 0.0196151
R18379 vdd.n9438 vdd.n9430 0.0196151
R18380 vdd.n9451 vdd.n9423 0.0196151
R18381 vdd.n9486 vdd.n9478 0.0196151
R18382 vdd.n9499 vdd.n9471 0.0196151
R18383 vdd.n9532 vdd.n9524 0.0196151
R18384 vdd.n9545 vdd.n9517 0.0196151
R18385 vdd.n3692 vdd.n3684 0.0196151
R18386 vdd.n3705 vdd.n3677 0.0196151
R18387 vdd.n3738 vdd.n3730 0.0196151
R18388 vdd.n3751 vdd.n3723 0.0196151
R18389 vdd.n3836 vdd.n3828 0.0196151
R18390 vdd.n3849 vdd.n3821 0.0196151
R18391 vdd.n3882 vdd.n3874 0.0196151
R18392 vdd.n3895 vdd.n3867 0.0196151
R18393 vdd.n3928 vdd.n3920 0.0196151
R18394 vdd.n3941 vdd.n3913 0.0196151
R18395 vdd.n3974 vdd.n3966 0.0196151
R18396 vdd.n3987 vdd.n3959 0.0196151
R18397 vdd.n4072 vdd.n4064 0.0196151
R18398 vdd.n4085 vdd.n4057 0.0196151
R18399 vdd.n5530 vdd.n5522 0.0196151
R18400 vdd.n5543 vdd.n5515 0.0196151
R18401 vdd.n4135 vdd.n4102 0.0196151
R18402 vdd.n4181 vdd.n4148 0.0196151
R18403 vdd.n4278 vdd.n4245 0.0196151
R18404 vdd.n4324 vdd.n4291 0.0196151
R18405 vdd.n4370 vdd.n4337 0.0196151
R18406 vdd.n4416 vdd.n4383 0.0196151
R18407 vdd.n4513 vdd.n4480 0.0196151
R18408 vdd.n3662 vdd.n3629 0.0196151
R18409 vdd.n4557 vdd.n4524 0.0196151
R18410 vdd.n4602 vdd.n4569 0.0196151
R18411 vdd.n4652 vdd.n4619 0.0196151
R18412 vdd.n4698 vdd.n4665 0.0196151
R18413 vdd.n4746 vdd.n4713 0.0196151
R18414 vdd.n4458 vdd.n4434 0.0196151
R18415 vdd.n4793 vdd.n4760 0.0196151
R18416 vdd.n4838 vdd.n4805 0.0196151
R18417 vdd.n4884 vdd.n4851 0.0196151
R18418 vdd.n4935 vdd.n4902 0.0196151
R18419 vdd.n4981 vdd.n4948 0.0196151
R18420 vdd.n5029 vdd.n4996 0.0196151
R18421 vdd.n5075 vdd.n5042 0.0196151
R18422 vdd.n5120 vdd.n5087 0.0196151
R18423 vdd.n5170 vdd.n5137 0.0196151
R18424 vdd.n5216 vdd.n5183 0.0196151
R18425 vdd.n5264 vdd.n5231 0.0196151
R18426 vdd.n4223 vdd.n4199 0.0196151
R18427 vdd.n5311 vdd.n5278 0.0196151
R18428 vdd.n5356 vdd.n5323 0.0196151
R18429 vdd.n5406 vdd.n5373 0.0196151
R18430 vdd.n5452 vdd.n5419 0.0196151
R18431 vdd.n5500 vdd.n5467 0.0196151
R18432 vdd.n5623 vdd.n5615 0.0196151
R18433 vdd.n5636 vdd.n5608 0.0196151
R18434 vdd.n5577 vdd.n5569 0.0196151
R18435 vdd.n5590 vdd.n5562 0.0196151
R18436 vdd.n5670 vdd.n5662 0.0196151
R18437 vdd.n5683 vdd.n5655 0.0196151
R18438 vdd.n5718 vdd.n5710 0.0196151
R18439 vdd.n5731 vdd.n5703 0.0196151
R18440 vdd.n5764 vdd.n5756 0.0196151
R18441 vdd.n5777 vdd.n5749 0.0196151
R18442 vdd.n4020 vdd.n4019 0.0196151
R18443 vdd.n4041 vdd.n4040 0.0196151
R18444 vdd.n5906 vdd.n5898 0.0196151
R18445 vdd.n5919 vdd.n5891 0.0196151
R18446 vdd.n5859 vdd.n5851 0.0196151
R18447 vdd.n5872 vdd.n5844 0.0196151
R18448 vdd.n5813 vdd.n5805 0.0196151
R18449 vdd.n5826 vdd.n5798 0.0196151
R18450 vdd.n5953 vdd.n5945 0.0196151
R18451 vdd.n5966 vdd.n5938 0.0196151
R18452 vdd.n6001 vdd.n5993 0.0196151
R18453 vdd.n6014 vdd.n5986 0.0196151
R18454 vdd.n6047 vdd.n6039 0.0196151
R18455 vdd.n6060 vdd.n6032 0.0196151
R18456 vdd.n6141 vdd.n6133 0.0196151
R18457 vdd.n6154 vdd.n6126 0.0196151
R18458 vdd.n6095 vdd.n6087 0.0196151
R18459 vdd.n6108 vdd.n6080 0.0196151
R18460 vdd.n6188 vdd.n6180 0.0196151
R18461 vdd.n6201 vdd.n6173 0.0196151
R18462 vdd.n6236 vdd.n6228 0.0196151
R18463 vdd.n6249 vdd.n6221 0.0196151
R18464 vdd.n6282 vdd.n6274 0.0196151
R18465 vdd.n6295 vdd.n6267 0.0196151
R18466 vdd.n3784 vdd.n3783 0.0196151
R18467 vdd.n3805 vdd.n3804 0.0196151
R18468 vdd.n6377 vdd.n6369 0.0196151
R18469 vdd.n6390 vdd.n6362 0.0196151
R18470 vdd.n6331 vdd.n6323 0.0196151
R18471 vdd.n6344 vdd.n6316 0.0196151
R18472 vdd.n6424 vdd.n6416 0.0196151
R18473 vdd.n6437 vdd.n6409 0.0196151
R18474 vdd.n6472 vdd.n6464 0.0196151
R18475 vdd.n6485 vdd.n6457 0.0196151
R18476 vdd.n6518 vdd.n6510 0.0196151
R18477 vdd.n6531 vdd.n6503 0.0196151
R18478 vdd.n678 vdd.n670 0.0196151
R18479 vdd.n691 vdd.n663 0.0196151
R18480 vdd.n724 vdd.n716 0.0196151
R18481 vdd.n737 vdd.n709 0.0196151
R18482 vdd.n822 vdd.n814 0.0196151
R18483 vdd.n835 vdd.n807 0.0196151
R18484 vdd.n868 vdd.n860 0.0196151
R18485 vdd.n881 vdd.n853 0.0196151
R18486 vdd.n914 vdd.n906 0.0196151
R18487 vdd.n927 vdd.n899 0.0196151
R18488 vdd.n960 vdd.n952 0.0196151
R18489 vdd.n973 vdd.n945 0.0196151
R18490 vdd.n1058 vdd.n1050 0.0196151
R18491 vdd.n1071 vdd.n1043 0.0196151
R18492 vdd.n2516 vdd.n2508 0.0196151
R18493 vdd.n2529 vdd.n2501 0.0196151
R18494 vdd.n1121 vdd.n1088 0.0196151
R18495 vdd.n1167 vdd.n1134 0.0196151
R18496 vdd.n1264 vdd.n1231 0.0196151
R18497 vdd.n1310 vdd.n1277 0.0196151
R18498 vdd.n1356 vdd.n1323 0.0196151
R18499 vdd.n1402 vdd.n1369 0.0196151
R18500 vdd.n1499 vdd.n1466 0.0196151
R18501 vdd.n648 vdd.n615 0.0196151
R18502 vdd.n1543 vdd.n1510 0.0196151
R18503 vdd.n1588 vdd.n1555 0.0196151
R18504 vdd.n1638 vdd.n1605 0.0196151
R18505 vdd.n1684 vdd.n1651 0.0196151
R18506 vdd.n1732 vdd.n1699 0.0196151
R18507 vdd.n1444 vdd.n1420 0.0196151
R18508 vdd.n1779 vdd.n1746 0.0196151
R18509 vdd.n1824 vdd.n1791 0.0196151
R18510 vdd.n1870 vdd.n1837 0.0196151
R18511 vdd.n1921 vdd.n1888 0.0196151
R18512 vdd.n1967 vdd.n1934 0.0196151
R18513 vdd.n2015 vdd.n1982 0.0196151
R18514 vdd.n2061 vdd.n2028 0.0196151
R18515 vdd.n2106 vdd.n2073 0.0196151
R18516 vdd.n2156 vdd.n2123 0.0196151
R18517 vdd.n2202 vdd.n2169 0.0196151
R18518 vdd.n2250 vdd.n2217 0.0196151
R18519 vdd.n1209 vdd.n1185 0.0196151
R18520 vdd.n2297 vdd.n2264 0.0196151
R18521 vdd.n2342 vdd.n2309 0.0196151
R18522 vdd.n2392 vdd.n2359 0.0196151
R18523 vdd.n2438 vdd.n2405 0.0196151
R18524 vdd.n2486 vdd.n2453 0.0196151
R18525 vdd.n2609 vdd.n2601 0.0196151
R18526 vdd.n2622 vdd.n2594 0.0196151
R18527 vdd.n2563 vdd.n2555 0.0196151
R18528 vdd.n2576 vdd.n2548 0.0196151
R18529 vdd.n2656 vdd.n2648 0.0196151
R18530 vdd.n2669 vdd.n2641 0.0196151
R18531 vdd.n2704 vdd.n2696 0.0196151
R18532 vdd.n2717 vdd.n2689 0.0196151
R18533 vdd.n2750 vdd.n2742 0.0196151
R18534 vdd.n2763 vdd.n2735 0.0196151
R18535 vdd.n1006 vdd.n1005 0.0196151
R18536 vdd.n1027 vdd.n1026 0.0196151
R18537 vdd.n2892 vdd.n2884 0.0196151
R18538 vdd.n2905 vdd.n2877 0.0196151
R18539 vdd.n2845 vdd.n2837 0.0196151
R18540 vdd.n2858 vdd.n2830 0.0196151
R18541 vdd.n2799 vdd.n2791 0.0196151
R18542 vdd.n2812 vdd.n2784 0.0196151
R18543 vdd.n2939 vdd.n2931 0.0196151
R18544 vdd.n2952 vdd.n2924 0.0196151
R18545 vdd.n2987 vdd.n2979 0.0196151
R18546 vdd.n3000 vdd.n2972 0.0196151
R18547 vdd.n3033 vdd.n3025 0.0196151
R18548 vdd.n3046 vdd.n3018 0.0196151
R18549 vdd.n3127 vdd.n3119 0.0196151
R18550 vdd.n3140 vdd.n3112 0.0196151
R18551 vdd.n3081 vdd.n3073 0.0196151
R18552 vdd.n3094 vdd.n3066 0.0196151
R18553 vdd.n3174 vdd.n3166 0.0196151
R18554 vdd.n3187 vdd.n3159 0.0196151
R18555 vdd.n3222 vdd.n3214 0.0196151
R18556 vdd.n3235 vdd.n3207 0.0196151
R18557 vdd.n3268 vdd.n3260 0.0196151
R18558 vdd.n3281 vdd.n3253 0.0196151
R18559 vdd.n770 vdd.n769 0.0196151
R18560 vdd.n791 vdd.n790 0.0196151
R18561 vdd.n3363 vdd.n3355 0.0196151
R18562 vdd.n3376 vdd.n3348 0.0196151
R18563 vdd.n3317 vdd.n3309 0.0196151
R18564 vdd.n3330 vdd.n3302 0.0196151
R18565 vdd.n3410 vdd.n3402 0.0196151
R18566 vdd.n3423 vdd.n3395 0.0196151
R18567 vdd.n3458 vdd.n3450 0.0196151
R18568 vdd.n3471 vdd.n3443 0.0196151
R18569 vdd.n3504 vdd.n3496 0.0196151
R18570 vdd.n3517 vdd.n3489 0.0196151
R18571 vdd.n586 vdd.n578 0.0196151
R18572 vdd.n599 vdd.n571 0.0196151
R18573 vdd.n3599 vdd.n3591 0.0196151
R18574 vdd.n3612 vdd.n3584 0.0196151
R18575 vdd.n3553 vdd.n3545 0.0196151
R18576 vdd.n3566 vdd.n3538 0.0196151
R18577 vdd.n6613 vdd.n6605 0.0196151
R18578 vdd.n6626 vdd.n6598 0.0196151
R18579 vdd.n6567 vdd.n6559 0.0196151
R18580 vdd.n6580 vdd.n6552 0.0196151
R18581 vdd.n9627 vdd.n9619 0.0196151
R18582 vdd.n9640 vdd.n9612 0.0196151
R18583 vdd.n9581 vdd.n9573 0.0196151
R18584 vdd.n9594 vdd.n9566 0.0196151
R18585 vdd.n9673 vdd.n9665 0.0196151
R18586 vdd.n9686 vdd.n9658 0.0196151
R18587 vdd.n9719 vdd.n9711 0.0196151
R18588 vdd.n9732 vdd.n9704 0.0196151
R18589 vdd.n9817 vdd.n9809 0.0196151
R18590 vdd.n9830 vdd.n9802 0.0196151
R18591 vdd.n9863 vdd.n9855 0.0196151
R18592 vdd.n9876 vdd.n9848 0.0196151
R18593 vdd.n9909 vdd.n9901 0.0196151
R18594 vdd.n9922 vdd.n9894 0.0196151
R18595 vdd.n9955 vdd.n9947 0.0196151
R18596 vdd.n9968 vdd.n9940 0.0196151
R18597 vdd.n10053 vdd.n10045 0.0196151
R18598 vdd.n10066 vdd.n10038 0.0196151
R18599 vdd.n69 vdd.n61 0.0196151
R18600 vdd.n82 vdd.n54 0.0196151
R18601 vdd.n23 vdd.n15 0.0196151
R18602 vdd.n36 vdd.n8 0.0196151
R18603 vdd.n10099 vdd.n10091 0.0196151
R18604 vdd.n10112 vdd.n10084 0.0196151
R18605 vdd.n10147 vdd.n10139 0.0196151
R18606 vdd.n10160 vdd.n10132 0.0196151
R18607 vdd.n10193 vdd.n10185 0.0196151
R18608 vdd.n10206 vdd.n10178 0.0196151
R18609 vdd.n10001 vdd.n10000 0.0196151
R18610 vdd.n10022 vdd.n10021 0.0196151
R18611 vdd.n10335 vdd.n10327 0.0196151
R18612 vdd.n10348 vdd.n10320 0.0196151
R18613 vdd.n10288 vdd.n10280 0.0196151
R18614 vdd.n10301 vdd.n10273 0.0196151
R18615 vdd.n10242 vdd.n10234 0.0196151
R18616 vdd.n10255 vdd.n10227 0.0196151
R18617 vdd.n10382 vdd.n10374 0.0196151
R18618 vdd.n10395 vdd.n10367 0.0196151
R18619 vdd.n10430 vdd.n10422 0.0196151
R18620 vdd.n10443 vdd.n10415 0.0196151
R18621 vdd.n10476 vdd.n10468 0.0196151
R18622 vdd.n10489 vdd.n10461 0.0196151
R18623 vdd.n10570 vdd.n10562 0.0196151
R18624 vdd.n10583 vdd.n10555 0.0196151
R18625 vdd.n10524 vdd.n10516 0.0196151
R18626 vdd.n10537 vdd.n10509 0.0196151
R18627 vdd.n10617 vdd.n10609 0.0196151
R18628 vdd.n10630 vdd.n10602 0.0196151
R18629 vdd.n10665 vdd.n10657 0.0196151
R18630 vdd.n10678 vdd.n10650 0.0196151
R18631 vdd.n10711 vdd.n10703 0.0196151
R18632 vdd.n10724 vdd.n10696 0.0196151
R18633 vdd.n9765 vdd.n9764 0.0196151
R18634 vdd.n9786 vdd.n9785 0.0196151
R18635 vdd.n10806 vdd.n10798 0.0196151
R18636 vdd.n10819 vdd.n10791 0.0196151
R18637 vdd.n10760 vdd.n10752 0.0196151
R18638 vdd.n10773 vdd.n10745 0.0196151
R18639 vdd.n10853 vdd.n10845 0.0196151
R18640 vdd.n10866 vdd.n10838 0.0196151
R18641 vdd.n10901 vdd.n10893 0.0196151
R18642 vdd.n10914 vdd.n10886 0.0196151
R18643 vdd.n10947 vdd.n10939 0.0196151
R18644 vdd.n10960 vdd.n10932 0.0196151
R18645 vdd.n11011 vdd.n10978 0.0196151
R18646 vdd.n11056 vdd.n11023 0.0196151
R18647 vdd.n11106 vdd.n11073 0.0196151
R18648 vdd.n11152 vdd.n11119 0.0196151
R18649 vdd.n11200 vdd.n11167 0.0196151
R18650 vdd.n456 vdd.n432 0.0196151
R18651 vdd.n11247 vdd.n11214 0.0196151
R18652 vdd.n11292 vdd.n11259 0.0196151
R18653 vdd.n11338 vdd.n11305 0.0196151
R18654 vdd.n11389 vdd.n11356 0.0196151
R18655 vdd.n11435 vdd.n11402 0.0196151
R18656 vdd.n11483 vdd.n11450 0.0196151
R18657 vdd.n11529 vdd.n11496 0.0196151
R18658 vdd.n11574 vdd.n11541 0.0196151
R18659 vdd.n11624 vdd.n11591 0.0196151
R18660 vdd.n11670 vdd.n11637 0.0196151
R18661 vdd.n11718 vdd.n11685 0.0196151
R18662 vdd.n221 vdd.n197 0.0196151
R18663 vdd.n11765 vdd.n11732 0.0196151
R18664 vdd.n11810 vdd.n11777 0.0196151
R18665 vdd.n11860 vdd.n11827 0.0196151
R18666 vdd.n11906 vdd.n11873 0.0196151
R18667 vdd.n11954 vdd.n11921 0.0196151
R18668 vdd.n7485 vdd.n7484 0.0185921
R18669 vdd.n7250 vdd.n7249 0.0185921
R18670 vdd.n7061 vdd.n7059 0.0185921
R18671 vdd.n6825 vdd.n6823 0.0185921
R18672 vdd.n4471 vdd.n4470 0.0185921
R18673 vdd.n4236 vdd.n4235 0.0185921
R18674 vdd.n4047 vdd.n4045 0.0185921
R18675 vdd.n3811 vdd.n3809 0.0185921
R18676 vdd.n1457 vdd.n1456 0.0185921
R18677 vdd.n1222 vdd.n1221 0.0185921
R18678 vdd.n1033 vdd.n1031 0.0185921
R18679 vdd.n797 vdd.n795 0.0185921
R18680 vdd.n10028 vdd.n10026 0.0185921
R18681 vdd.n9792 vdd.n9790 0.0185921
R18682 vdd.n469 vdd.n468 0.0185921
R18683 vdd.n234 vdd.n233 0.0185921
R18684 vdd.n7485 vdd 0.0136579
R18685 vdd.n7250 vdd 0.0136579
R18686 vdd.n4471 vdd 0.0136579
R18687 vdd.n4236 vdd 0.0136579
R18688 vdd.n1457 vdd 0.0136579
R18689 vdd.n1222 vdd 0.0136579
R18690 vdd.n469 vdd 0.0136579
R18691 vdd.n234 vdd 0.0136579
R18692 vdd.n11964 vdd.n11963 0.0130799
R18693 vdd.n11963 vdd.n11962 0.0130799
R18694 vdd.n11967 vdd.n11966 0.0130799
R18695 vdd.n11966 vdd.n11965 0.0130799
R18696 vdd.n11986 vdd.n11985 0.0130799
R18697 vdd.n11985 vdd.n11984 0.0130799
R18698 vdd.n11988 vdd.n11987 0.0130799
R18699 vdd.n11969 vdd.n11968 0.0130799
R18700 vdd.n106 vdd.n95 0.0130799
R18701 vdd.n107 vdd.n106 0.0130799
R18702 vdd.n123 vdd.n99 0.0130799
R18703 vdd.n128 vdd.n99 0.0130799
R18704 vdd.n114 vdd.n108 0.0130799
R18705 vdd.n108 vdd.n105 0.0130799
R18706 vdd.n113 vdd.n109 0.0130799
R18707 vdd.n131 vdd.n130 0.0130799
R18708 vdd.n152 vdd.n141 0.0130799
R18709 vdd.n153 vdd.n152 0.0130799
R18710 vdd.n169 vdd.n145 0.0130799
R18711 vdd.n174 vdd.n145 0.0130799
R18712 vdd.n160 vdd.n154 0.0130799
R18713 vdd.n154 vdd.n151 0.0130799
R18714 vdd.n159 vdd.n155 0.0130799
R18715 vdd.n177 vdd.n176 0.0130799
R18716 vdd.n249 vdd.n238 0.0130799
R18717 vdd.n250 vdd.n249 0.0130799
R18718 vdd.n266 vdd.n242 0.0130799
R18719 vdd.n271 vdd.n242 0.0130799
R18720 vdd.n257 vdd.n251 0.0130799
R18721 vdd.n251 vdd.n248 0.0130799
R18722 vdd.n256 vdd.n252 0.0130799
R18723 vdd.n274 vdd.n273 0.0130799
R18724 vdd.n295 vdd.n284 0.0130799
R18725 vdd.n296 vdd.n295 0.0130799
R18726 vdd.n312 vdd.n288 0.0130799
R18727 vdd.n317 vdd.n288 0.0130799
R18728 vdd.n303 vdd.n297 0.0130799
R18729 vdd.n297 vdd.n294 0.0130799
R18730 vdd.n302 vdd.n298 0.0130799
R18731 vdd.n320 vdd.n319 0.0130799
R18732 vdd.n341 vdd.n330 0.0130799
R18733 vdd.n342 vdd.n341 0.0130799
R18734 vdd.n358 vdd.n334 0.0130799
R18735 vdd.n363 vdd.n334 0.0130799
R18736 vdd.n349 vdd.n343 0.0130799
R18737 vdd.n343 vdd.n340 0.0130799
R18738 vdd.n348 vdd.n344 0.0130799
R18739 vdd.n366 vdd.n365 0.0130799
R18740 vdd.n387 vdd.n376 0.0130799
R18741 vdd.n388 vdd.n387 0.0130799
R18742 vdd.n404 vdd.n380 0.0130799
R18743 vdd.n409 vdd.n380 0.0130799
R18744 vdd.n395 vdd.n389 0.0130799
R18745 vdd.n389 vdd.n386 0.0130799
R18746 vdd.n394 vdd.n390 0.0130799
R18747 vdd.n412 vdd.n411 0.0130799
R18748 vdd.n484 vdd.n473 0.0130799
R18749 vdd.n485 vdd.n484 0.0130799
R18750 vdd.n501 vdd.n477 0.0130799
R18751 vdd.n506 vdd.n477 0.0130799
R18752 vdd.n492 vdd.n486 0.0130799
R18753 vdd.n486 vdd.n483 0.0130799
R18754 vdd.n491 vdd.n487 0.0130799
R18755 vdd.n509 vdd.n508 0.0130799
R18756 vdd.n530 vdd.n519 0.0130799
R18757 vdd.n531 vdd.n530 0.0130799
R18758 vdd.n547 vdd.n523 0.0130799
R18759 vdd.n552 vdd.n523 0.0130799
R18760 vdd.n538 vdd.n532 0.0130799
R18761 vdd.n532 vdd.n529 0.0130799
R18762 vdd.n537 vdd.n533 0.0130799
R18763 vdd.n555 vdd.n554 0.0130799
R18764 vdd.n6694 vdd.n6683 0.0130799
R18765 vdd.n6694 vdd.n6688 0.0130799
R18766 vdd.n6703 vdd.n6697 0.0130799
R18767 vdd.n6697 vdd.n6696 0.0130799
R18768 vdd.n6721 vdd.n6690 0.0130799
R18769 vdd.n6722 vdd.n6721 0.0130799
R18770 vdd.n6717 vdd.n6716 0.0130799
R18771 vdd.n6702 vdd.n6701 0.0130799
R18772 vdd.n6740 vdd.n6729 0.0130799
R18773 vdd.n6740 vdd.n6734 0.0130799
R18774 vdd.n6749 vdd.n6743 0.0130799
R18775 vdd.n6743 vdd.n6742 0.0130799
R18776 vdd.n6767 vdd.n6736 0.0130799
R18777 vdd.n6768 vdd.n6767 0.0130799
R18778 vdd.n6763 vdd.n6762 0.0130799
R18779 vdd.n6748 vdd.n6747 0.0130799
R18780 vdd.n6838 vdd.n6827 0.0130799
R18781 vdd.n6838 vdd.n6832 0.0130799
R18782 vdd.n6847 vdd.n6841 0.0130799
R18783 vdd.n6841 vdd.n6840 0.0130799
R18784 vdd.n6865 vdd.n6834 0.0130799
R18785 vdd.n6866 vdd.n6865 0.0130799
R18786 vdd.n6861 vdd.n6860 0.0130799
R18787 vdd.n6846 vdd.n6845 0.0130799
R18788 vdd.n6884 vdd.n6873 0.0130799
R18789 vdd.n6884 vdd.n6878 0.0130799
R18790 vdd.n6893 vdd.n6887 0.0130799
R18791 vdd.n6887 vdd.n6886 0.0130799
R18792 vdd.n6911 vdd.n6880 0.0130799
R18793 vdd.n6912 vdd.n6911 0.0130799
R18794 vdd.n6907 vdd.n6906 0.0130799
R18795 vdd.n6892 vdd.n6891 0.0130799
R18796 vdd.n6930 vdd.n6919 0.0130799
R18797 vdd.n6930 vdd.n6924 0.0130799
R18798 vdd.n6939 vdd.n6933 0.0130799
R18799 vdd.n6933 vdd.n6932 0.0130799
R18800 vdd.n6957 vdd.n6926 0.0130799
R18801 vdd.n6958 vdd.n6957 0.0130799
R18802 vdd.n6953 vdd.n6952 0.0130799
R18803 vdd.n6938 vdd.n6937 0.0130799
R18804 vdd.n6976 vdd.n6965 0.0130799
R18805 vdd.n6976 vdd.n6970 0.0130799
R18806 vdd.n6985 vdd.n6979 0.0130799
R18807 vdd.n6979 vdd.n6978 0.0130799
R18808 vdd.n7003 vdd.n6972 0.0130799
R18809 vdd.n7004 vdd.n7003 0.0130799
R18810 vdd.n6999 vdd.n6998 0.0130799
R18811 vdd.n6984 vdd.n6983 0.0130799
R18812 vdd.n7074 vdd.n7063 0.0130799
R18813 vdd.n7074 vdd.n7068 0.0130799
R18814 vdd.n7083 vdd.n7077 0.0130799
R18815 vdd.n7077 vdd.n7076 0.0130799
R18816 vdd.n7101 vdd.n7070 0.0130799
R18817 vdd.n7102 vdd.n7101 0.0130799
R18818 vdd.n7097 vdd.n7096 0.0130799
R18819 vdd.n7082 vdd.n7081 0.0130799
R18820 vdd.n8532 vdd.n8521 0.0130799
R18821 vdd.n8532 vdd.n8526 0.0130799
R18822 vdd.n8541 vdd.n8535 0.0130799
R18823 vdd.n8535 vdd.n8534 0.0130799
R18824 vdd.n8559 vdd.n8528 0.0130799
R18825 vdd.n8560 vdd.n8559 0.0130799
R18826 vdd.n8555 vdd.n8554 0.0130799
R18827 vdd.n8540 vdd.n8539 0.0130799
R18828 vdd.n7122 vdd.n7111 0.0130799
R18829 vdd.n7123 vdd.n7122 0.0130799
R18830 vdd.n7139 vdd.n7115 0.0130799
R18831 vdd.n7144 vdd.n7115 0.0130799
R18832 vdd.n7130 vdd.n7124 0.0130799
R18833 vdd.n7124 vdd.n7121 0.0130799
R18834 vdd.n7129 vdd.n7125 0.0130799
R18835 vdd.n7147 vdd.n7146 0.0130799
R18836 vdd.n7168 vdd.n7157 0.0130799
R18837 vdd.n7169 vdd.n7168 0.0130799
R18838 vdd.n7185 vdd.n7161 0.0130799
R18839 vdd.n7190 vdd.n7161 0.0130799
R18840 vdd.n7176 vdd.n7170 0.0130799
R18841 vdd.n7170 vdd.n7167 0.0130799
R18842 vdd.n7175 vdd.n7171 0.0130799
R18843 vdd.n7193 vdd.n7192 0.0130799
R18844 vdd.n7265 vdd.n7254 0.0130799
R18845 vdd.n7266 vdd.n7265 0.0130799
R18846 vdd.n7282 vdd.n7258 0.0130799
R18847 vdd.n7287 vdd.n7258 0.0130799
R18848 vdd.n7273 vdd.n7267 0.0130799
R18849 vdd.n7267 vdd.n7264 0.0130799
R18850 vdd.n7272 vdd.n7268 0.0130799
R18851 vdd.n7290 vdd.n7289 0.0130799
R18852 vdd.n7311 vdd.n7300 0.0130799
R18853 vdd.n7312 vdd.n7311 0.0130799
R18854 vdd.n7328 vdd.n7304 0.0130799
R18855 vdd.n7333 vdd.n7304 0.0130799
R18856 vdd.n7319 vdd.n7313 0.0130799
R18857 vdd.n7313 vdd.n7310 0.0130799
R18858 vdd.n7318 vdd.n7314 0.0130799
R18859 vdd.n7336 vdd.n7335 0.0130799
R18860 vdd.n7357 vdd.n7346 0.0130799
R18861 vdd.n7358 vdd.n7357 0.0130799
R18862 vdd.n7374 vdd.n7350 0.0130799
R18863 vdd.n7379 vdd.n7350 0.0130799
R18864 vdd.n7365 vdd.n7359 0.0130799
R18865 vdd.n7359 vdd.n7356 0.0130799
R18866 vdd.n7364 vdd.n7360 0.0130799
R18867 vdd.n7382 vdd.n7381 0.0130799
R18868 vdd.n7403 vdd.n7392 0.0130799
R18869 vdd.n7404 vdd.n7403 0.0130799
R18870 vdd.n7420 vdd.n7396 0.0130799
R18871 vdd.n7425 vdd.n7396 0.0130799
R18872 vdd.n7411 vdd.n7405 0.0130799
R18873 vdd.n7405 vdd.n7402 0.0130799
R18874 vdd.n7410 vdd.n7406 0.0130799
R18875 vdd.n7428 vdd.n7427 0.0130799
R18876 vdd.n7500 vdd.n7489 0.0130799
R18877 vdd.n7501 vdd.n7500 0.0130799
R18878 vdd.n7517 vdd.n7493 0.0130799
R18879 vdd.n7522 vdd.n7493 0.0130799
R18880 vdd.n7508 vdd.n7502 0.0130799
R18881 vdd.n7502 vdd.n7499 0.0130799
R18882 vdd.n7507 vdd.n7503 0.0130799
R18883 vdd.n7525 vdd.n7524 0.0130799
R18884 vdd.n6649 vdd.n6638 0.0130799
R18885 vdd.n6650 vdd.n6649 0.0130799
R18886 vdd.n6666 vdd.n6642 0.0130799
R18887 vdd.n6671 vdd.n6642 0.0130799
R18888 vdd.n6657 vdd.n6651 0.0130799
R18889 vdd.n6651 vdd.n6648 0.0130799
R18890 vdd.n6656 vdd.n6652 0.0130799
R18891 vdd.n6674 vdd.n6673 0.0130799
R18892 vdd.n7544 vdd.n7533 0.0130799
R18893 vdd.n7545 vdd.n7544 0.0130799
R18894 vdd.n7561 vdd.n7537 0.0130799
R18895 vdd.n7566 vdd.n7537 0.0130799
R18896 vdd.n7552 vdd.n7546 0.0130799
R18897 vdd.n7546 vdd.n7543 0.0130799
R18898 vdd.n7551 vdd.n7547 0.0130799
R18899 vdd.n7569 vdd.n7568 0.0130799
R18900 vdd.n7589 vdd.n7578 0.0130799
R18901 vdd.n7590 vdd.n7589 0.0130799
R18902 vdd.n7606 vdd.n7582 0.0130799
R18903 vdd.n7611 vdd.n7582 0.0130799
R18904 vdd.n7597 vdd.n7591 0.0130799
R18905 vdd.n7591 vdd.n7588 0.0130799
R18906 vdd.n7596 vdd.n7592 0.0130799
R18907 vdd.n7614 vdd.n7613 0.0130799
R18908 vdd.n7639 vdd.n7628 0.0130799
R18909 vdd.n7640 vdd.n7639 0.0130799
R18910 vdd.n7656 vdd.n7632 0.0130799
R18911 vdd.n7661 vdd.n7632 0.0130799
R18912 vdd.n7647 vdd.n7641 0.0130799
R18913 vdd.n7641 vdd.n7638 0.0130799
R18914 vdd.n7646 vdd.n7642 0.0130799
R18915 vdd.n7664 vdd.n7663 0.0130799
R18916 vdd.n7685 vdd.n7674 0.0130799
R18917 vdd.n7686 vdd.n7685 0.0130799
R18918 vdd.n7702 vdd.n7678 0.0130799
R18919 vdd.n7707 vdd.n7678 0.0130799
R18920 vdd.n7693 vdd.n7687 0.0130799
R18921 vdd.n7687 vdd.n7684 0.0130799
R18922 vdd.n7692 vdd.n7688 0.0130799
R18923 vdd.n7710 vdd.n7709 0.0130799
R18924 vdd.n7733 vdd.n7722 0.0130799
R18925 vdd.n7734 vdd.n7733 0.0130799
R18926 vdd.n7750 vdd.n7726 0.0130799
R18927 vdd.n7755 vdd.n7726 0.0130799
R18928 vdd.n7741 vdd.n7735 0.0130799
R18929 vdd.n7735 vdd.n7732 0.0130799
R18930 vdd.n7740 vdd.n7736 0.0130799
R18931 vdd.n7758 vdd.n7757 0.0130799
R18932 vdd.n7451 vdd.n7444 0.0130799
R18933 vdd.n7451 vdd.n7450 0.0130799
R18934 vdd.n7462 vdd.n7447 0.0130799
R18935 vdd.n7467 vdd.n7447 0.0130799
R18936 vdd.n7453 vdd.n7441 0.0130799
R18937 vdd.n7442 vdd.n7441 0.0130799
R18938 vdd.n7440 vdd.n7438 0.0130799
R18939 vdd.n7470 vdd.n7469 0.0130799
R18940 vdd.n7780 vdd.n7769 0.0130799
R18941 vdd.n7781 vdd.n7780 0.0130799
R18942 vdd.n7797 vdd.n7773 0.0130799
R18943 vdd.n7802 vdd.n7773 0.0130799
R18944 vdd.n7788 vdd.n7782 0.0130799
R18945 vdd.n7782 vdd.n7779 0.0130799
R18946 vdd.n7787 vdd.n7783 0.0130799
R18947 vdd.n7805 vdd.n7804 0.0130799
R18948 vdd.n7825 vdd.n7814 0.0130799
R18949 vdd.n7826 vdd.n7825 0.0130799
R18950 vdd.n7842 vdd.n7818 0.0130799
R18951 vdd.n7847 vdd.n7818 0.0130799
R18952 vdd.n7833 vdd.n7827 0.0130799
R18953 vdd.n7827 vdd.n7824 0.0130799
R18954 vdd.n7832 vdd.n7828 0.0130799
R18955 vdd.n7850 vdd.n7849 0.0130799
R18956 vdd.n7871 vdd.n7860 0.0130799
R18957 vdd.n7872 vdd.n7871 0.0130799
R18958 vdd.n7888 vdd.n7864 0.0130799
R18959 vdd.n7893 vdd.n7864 0.0130799
R18960 vdd.n7879 vdd.n7873 0.0130799
R18961 vdd.n7873 vdd.n7870 0.0130799
R18962 vdd.n7878 vdd.n7874 0.0130799
R18963 vdd.n7896 vdd.n7895 0.0130799
R18964 vdd.n7922 vdd.n7911 0.0130799
R18965 vdd.n7923 vdd.n7922 0.0130799
R18966 vdd.n7939 vdd.n7915 0.0130799
R18967 vdd.n7944 vdd.n7915 0.0130799
R18968 vdd.n7930 vdd.n7924 0.0130799
R18969 vdd.n7924 vdd.n7921 0.0130799
R18970 vdd.n7929 vdd.n7925 0.0130799
R18971 vdd.n7947 vdd.n7946 0.0130799
R18972 vdd.n7968 vdd.n7957 0.0130799
R18973 vdd.n7969 vdd.n7968 0.0130799
R18974 vdd.n7985 vdd.n7961 0.0130799
R18975 vdd.n7990 vdd.n7961 0.0130799
R18976 vdd.n7976 vdd.n7970 0.0130799
R18977 vdd.n7970 vdd.n7967 0.0130799
R18978 vdd.n7975 vdd.n7971 0.0130799
R18979 vdd.n7993 vdd.n7992 0.0130799
R18980 vdd.n8016 vdd.n8005 0.0130799
R18981 vdd.n8017 vdd.n8016 0.0130799
R18982 vdd.n8033 vdd.n8009 0.0130799
R18983 vdd.n8038 vdd.n8009 0.0130799
R18984 vdd.n8024 vdd.n8018 0.0130799
R18985 vdd.n8018 vdd.n8015 0.0130799
R18986 vdd.n8023 vdd.n8019 0.0130799
R18987 vdd.n8041 vdd.n8040 0.0130799
R18988 vdd.n8062 vdd.n8051 0.0130799
R18989 vdd.n8063 vdd.n8062 0.0130799
R18990 vdd.n8079 vdd.n8055 0.0130799
R18991 vdd.n8084 vdd.n8055 0.0130799
R18992 vdd.n8070 vdd.n8064 0.0130799
R18993 vdd.n8064 vdd.n8061 0.0130799
R18994 vdd.n8069 vdd.n8065 0.0130799
R18995 vdd.n8087 vdd.n8086 0.0130799
R18996 vdd.n8107 vdd.n8096 0.0130799
R18997 vdd.n8108 vdd.n8107 0.0130799
R18998 vdd.n8124 vdd.n8100 0.0130799
R18999 vdd.n8129 vdd.n8100 0.0130799
R19000 vdd.n8115 vdd.n8109 0.0130799
R19001 vdd.n8109 vdd.n8106 0.0130799
R19002 vdd.n8114 vdd.n8110 0.0130799
R19003 vdd.n8132 vdd.n8131 0.0130799
R19004 vdd.n8157 vdd.n8146 0.0130799
R19005 vdd.n8158 vdd.n8157 0.0130799
R19006 vdd.n8174 vdd.n8150 0.0130799
R19007 vdd.n8179 vdd.n8150 0.0130799
R19008 vdd.n8165 vdd.n8159 0.0130799
R19009 vdd.n8159 vdd.n8156 0.0130799
R19010 vdd.n8164 vdd.n8160 0.0130799
R19011 vdd.n8182 vdd.n8181 0.0130799
R19012 vdd.n8203 vdd.n8192 0.0130799
R19013 vdd.n8204 vdd.n8203 0.0130799
R19014 vdd.n8220 vdd.n8196 0.0130799
R19015 vdd.n8225 vdd.n8196 0.0130799
R19016 vdd.n8211 vdd.n8205 0.0130799
R19017 vdd.n8205 vdd.n8202 0.0130799
R19018 vdd.n8210 vdd.n8206 0.0130799
R19019 vdd.n8228 vdd.n8227 0.0130799
R19020 vdd.n8251 vdd.n8240 0.0130799
R19021 vdd.n8252 vdd.n8251 0.0130799
R19022 vdd.n8268 vdd.n8244 0.0130799
R19023 vdd.n8273 vdd.n8244 0.0130799
R19024 vdd.n8259 vdd.n8253 0.0130799
R19025 vdd.n8253 vdd.n8250 0.0130799
R19026 vdd.n8258 vdd.n8254 0.0130799
R19027 vdd.n8276 vdd.n8275 0.0130799
R19028 vdd.n7216 vdd.n7209 0.0130799
R19029 vdd.n7216 vdd.n7215 0.0130799
R19030 vdd.n7227 vdd.n7212 0.0130799
R19031 vdd.n7232 vdd.n7212 0.0130799
R19032 vdd.n7218 vdd.n7206 0.0130799
R19033 vdd.n7207 vdd.n7206 0.0130799
R19034 vdd.n7205 vdd.n7203 0.0130799
R19035 vdd.n7235 vdd.n7234 0.0130799
R19036 vdd.n8298 vdd.n8287 0.0130799
R19037 vdd.n8299 vdd.n8298 0.0130799
R19038 vdd.n8315 vdd.n8291 0.0130799
R19039 vdd.n8320 vdd.n8291 0.0130799
R19040 vdd.n8306 vdd.n8300 0.0130799
R19041 vdd.n8300 vdd.n8297 0.0130799
R19042 vdd.n8305 vdd.n8301 0.0130799
R19043 vdd.n8323 vdd.n8322 0.0130799
R19044 vdd.n8343 vdd.n8332 0.0130799
R19045 vdd.n8344 vdd.n8343 0.0130799
R19046 vdd.n8360 vdd.n8336 0.0130799
R19047 vdd.n8365 vdd.n8336 0.0130799
R19048 vdd.n8351 vdd.n8345 0.0130799
R19049 vdd.n8345 vdd.n8342 0.0130799
R19050 vdd.n8350 vdd.n8346 0.0130799
R19051 vdd.n8368 vdd.n8367 0.0130799
R19052 vdd.n8393 vdd.n8382 0.0130799
R19053 vdd.n8394 vdd.n8393 0.0130799
R19054 vdd.n8410 vdd.n8386 0.0130799
R19055 vdd.n8415 vdd.n8386 0.0130799
R19056 vdd.n8401 vdd.n8395 0.0130799
R19057 vdd.n8395 vdd.n8392 0.0130799
R19058 vdd.n8400 vdd.n8396 0.0130799
R19059 vdd.n8418 vdd.n8417 0.0130799
R19060 vdd.n8439 vdd.n8428 0.0130799
R19061 vdd.n8440 vdd.n8439 0.0130799
R19062 vdd.n8456 vdd.n8432 0.0130799
R19063 vdd.n8461 vdd.n8432 0.0130799
R19064 vdd.n8447 vdd.n8441 0.0130799
R19065 vdd.n8441 vdd.n8438 0.0130799
R19066 vdd.n8446 vdd.n8442 0.0130799
R19067 vdd.n8464 vdd.n8463 0.0130799
R19068 vdd.n8487 vdd.n8476 0.0130799
R19069 vdd.n8488 vdd.n8487 0.0130799
R19070 vdd.n8504 vdd.n8480 0.0130799
R19071 vdd.n8509 vdd.n8480 0.0130799
R19072 vdd.n8495 vdd.n8489 0.0130799
R19073 vdd.n8489 vdd.n8486 0.0130799
R19074 vdd.n8494 vdd.n8490 0.0130799
R19075 vdd.n8512 vdd.n8511 0.0130799
R19076 vdd.n8625 vdd.n8614 0.0130799
R19077 vdd.n8625 vdd.n8619 0.0130799
R19078 vdd.n8634 vdd.n8628 0.0130799
R19079 vdd.n8628 vdd.n8627 0.0130799
R19080 vdd.n8652 vdd.n8621 0.0130799
R19081 vdd.n8653 vdd.n8652 0.0130799
R19082 vdd.n8648 vdd.n8647 0.0130799
R19083 vdd.n8633 vdd.n8632 0.0130799
R19084 vdd.n8579 vdd.n8568 0.0130799
R19085 vdd.n8579 vdd.n8573 0.0130799
R19086 vdd.n8588 vdd.n8582 0.0130799
R19087 vdd.n8582 vdd.n8581 0.0130799
R19088 vdd.n8606 vdd.n8575 0.0130799
R19089 vdd.n8607 vdd.n8606 0.0130799
R19090 vdd.n8602 vdd.n8601 0.0130799
R19091 vdd.n8587 vdd.n8586 0.0130799
R19092 vdd.n8672 vdd.n8661 0.0130799
R19093 vdd.n8672 vdd.n8666 0.0130799
R19094 vdd.n8681 vdd.n8675 0.0130799
R19095 vdd.n8675 vdd.n8674 0.0130799
R19096 vdd.n8699 vdd.n8668 0.0130799
R19097 vdd.n8700 vdd.n8699 0.0130799
R19098 vdd.n8695 vdd.n8694 0.0130799
R19099 vdd.n8680 vdd.n8679 0.0130799
R19100 vdd.n8720 vdd.n8709 0.0130799
R19101 vdd.n8720 vdd.n8714 0.0130799
R19102 vdd.n8729 vdd.n8723 0.0130799
R19103 vdd.n8723 vdd.n8722 0.0130799
R19104 vdd.n8747 vdd.n8716 0.0130799
R19105 vdd.n8748 vdd.n8747 0.0130799
R19106 vdd.n8743 vdd.n8742 0.0130799
R19107 vdd.n8728 vdd.n8727 0.0130799
R19108 vdd.n8766 vdd.n8755 0.0130799
R19109 vdd.n8766 vdd.n8760 0.0130799
R19110 vdd.n8775 vdd.n8769 0.0130799
R19111 vdd.n8769 vdd.n8768 0.0130799
R19112 vdd.n8793 vdd.n8762 0.0130799
R19113 vdd.n8794 vdd.n8793 0.0130799
R19114 vdd.n8789 vdd.n8788 0.0130799
R19115 vdd.n8774 vdd.n8773 0.0130799
R19116 vdd.n7025 vdd.n7019 0.0130799
R19117 vdd.n7042 vdd.n7025 0.0130799
R19118 vdd.n7030 vdd.n7027 0.0130799
R19119 vdd.n7030 vdd.n7023 0.0130799
R19120 vdd.n7051 vdd.n7050 0.0130799
R19121 vdd.n7051 vdd.n7017 0.0130799
R19122 vdd.n7057 vdd.n7014 0.0130799
R19123 vdd.n7029 vdd.n7028 0.0130799
R19124 vdd.n8908 vdd.n8897 0.0130799
R19125 vdd.n8908 vdd.n8902 0.0130799
R19126 vdd.n8917 vdd.n8911 0.0130799
R19127 vdd.n8911 vdd.n8910 0.0130799
R19128 vdd.n8935 vdd.n8904 0.0130799
R19129 vdd.n8936 vdd.n8935 0.0130799
R19130 vdd.n8931 vdd.n8930 0.0130799
R19131 vdd.n8916 vdd.n8915 0.0130799
R19132 vdd.n8861 vdd.n8850 0.0130799
R19133 vdd.n8861 vdd.n8855 0.0130799
R19134 vdd.n8870 vdd.n8864 0.0130799
R19135 vdd.n8864 vdd.n8863 0.0130799
R19136 vdd.n8888 vdd.n8857 0.0130799
R19137 vdd.n8889 vdd.n8888 0.0130799
R19138 vdd.n8884 vdd.n8883 0.0130799
R19139 vdd.n8869 vdd.n8868 0.0130799
R19140 vdd.n8815 vdd.n8804 0.0130799
R19141 vdd.n8815 vdd.n8809 0.0130799
R19142 vdd.n8824 vdd.n8818 0.0130799
R19143 vdd.n8818 vdd.n8817 0.0130799
R19144 vdd.n8842 vdd.n8811 0.0130799
R19145 vdd.n8843 vdd.n8842 0.0130799
R19146 vdd.n8838 vdd.n8837 0.0130799
R19147 vdd.n8823 vdd.n8822 0.0130799
R19148 vdd.n8955 vdd.n8944 0.0130799
R19149 vdd.n8955 vdd.n8949 0.0130799
R19150 vdd.n8964 vdd.n8958 0.0130799
R19151 vdd.n8958 vdd.n8957 0.0130799
R19152 vdd.n8982 vdd.n8951 0.0130799
R19153 vdd.n8983 vdd.n8982 0.0130799
R19154 vdd.n8978 vdd.n8977 0.0130799
R19155 vdd.n8963 vdd.n8962 0.0130799
R19156 vdd.n9003 vdd.n8992 0.0130799
R19157 vdd.n9003 vdd.n8997 0.0130799
R19158 vdd.n9012 vdd.n9006 0.0130799
R19159 vdd.n9006 vdd.n9005 0.0130799
R19160 vdd.n9030 vdd.n8999 0.0130799
R19161 vdd.n9031 vdd.n9030 0.0130799
R19162 vdd.n9026 vdd.n9025 0.0130799
R19163 vdd.n9011 vdd.n9010 0.0130799
R19164 vdd.n9049 vdd.n9038 0.0130799
R19165 vdd.n9049 vdd.n9043 0.0130799
R19166 vdd.n9058 vdd.n9052 0.0130799
R19167 vdd.n9052 vdd.n9051 0.0130799
R19168 vdd.n9076 vdd.n9045 0.0130799
R19169 vdd.n9077 vdd.n9076 0.0130799
R19170 vdd.n9072 vdd.n9071 0.0130799
R19171 vdd.n9057 vdd.n9056 0.0130799
R19172 vdd.n9143 vdd.n9132 0.0130799
R19173 vdd.n9143 vdd.n9137 0.0130799
R19174 vdd.n9152 vdd.n9146 0.0130799
R19175 vdd.n9146 vdd.n9145 0.0130799
R19176 vdd.n9170 vdd.n9139 0.0130799
R19177 vdd.n9171 vdd.n9170 0.0130799
R19178 vdd.n9166 vdd.n9165 0.0130799
R19179 vdd.n9151 vdd.n9150 0.0130799
R19180 vdd.n9097 vdd.n9086 0.0130799
R19181 vdd.n9097 vdd.n9091 0.0130799
R19182 vdd.n9106 vdd.n9100 0.0130799
R19183 vdd.n9100 vdd.n9099 0.0130799
R19184 vdd.n9124 vdd.n9093 0.0130799
R19185 vdd.n9125 vdd.n9124 0.0130799
R19186 vdd.n9120 vdd.n9119 0.0130799
R19187 vdd.n9105 vdd.n9104 0.0130799
R19188 vdd.n9190 vdd.n9179 0.0130799
R19189 vdd.n9190 vdd.n9184 0.0130799
R19190 vdd.n9199 vdd.n9193 0.0130799
R19191 vdd.n9193 vdd.n9192 0.0130799
R19192 vdd.n9217 vdd.n9186 0.0130799
R19193 vdd.n9218 vdd.n9217 0.0130799
R19194 vdd.n9213 vdd.n9212 0.0130799
R19195 vdd.n9198 vdd.n9197 0.0130799
R19196 vdd.n9238 vdd.n9227 0.0130799
R19197 vdd.n9238 vdd.n9232 0.0130799
R19198 vdd.n9247 vdd.n9241 0.0130799
R19199 vdd.n9241 vdd.n9240 0.0130799
R19200 vdd.n9265 vdd.n9234 0.0130799
R19201 vdd.n9266 vdd.n9265 0.0130799
R19202 vdd.n9261 vdd.n9260 0.0130799
R19203 vdd.n9246 vdd.n9245 0.0130799
R19204 vdd.n9284 vdd.n9273 0.0130799
R19205 vdd.n9284 vdd.n9278 0.0130799
R19206 vdd.n9293 vdd.n9287 0.0130799
R19207 vdd.n9287 vdd.n9286 0.0130799
R19208 vdd.n9311 vdd.n9280 0.0130799
R19209 vdd.n9312 vdd.n9311 0.0130799
R19210 vdd.n9307 vdd.n9306 0.0130799
R19211 vdd.n9292 vdd.n9291 0.0130799
R19212 vdd.n6789 vdd.n6783 0.0130799
R19213 vdd.n6806 vdd.n6789 0.0130799
R19214 vdd.n6794 vdd.n6791 0.0130799
R19215 vdd.n6794 vdd.n6787 0.0130799
R19216 vdd.n6815 vdd.n6814 0.0130799
R19217 vdd.n6815 vdd.n6781 0.0130799
R19218 vdd.n6821 vdd.n6778 0.0130799
R19219 vdd.n6793 vdd.n6792 0.0130799
R19220 vdd.n9379 vdd.n9368 0.0130799
R19221 vdd.n9379 vdd.n9373 0.0130799
R19222 vdd.n9388 vdd.n9382 0.0130799
R19223 vdd.n9382 vdd.n9381 0.0130799
R19224 vdd.n9406 vdd.n9375 0.0130799
R19225 vdd.n9407 vdd.n9406 0.0130799
R19226 vdd.n9402 vdd.n9401 0.0130799
R19227 vdd.n9387 vdd.n9386 0.0130799
R19228 vdd.n9333 vdd.n9322 0.0130799
R19229 vdd.n9333 vdd.n9327 0.0130799
R19230 vdd.n9342 vdd.n9336 0.0130799
R19231 vdd.n9336 vdd.n9335 0.0130799
R19232 vdd.n9360 vdd.n9329 0.0130799
R19233 vdd.n9361 vdd.n9360 0.0130799
R19234 vdd.n9356 vdd.n9355 0.0130799
R19235 vdd.n9341 vdd.n9340 0.0130799
R19236 vdd.n9426 vdd.n9415 0.0130799
R19237 vdd.n9426 vdd.n9420 0.0130799
R19238 vdd.n9435 vdd.n9429 0.0130799
R19239 vdd.n9429 vdd.n9428 0.0130799
R19240 vdd.n9453 vdd.n9422 0.0130799
R19241 vdd.n9454 vdd.n9453 0.0130799
R19242 vdd.n9449 vdd.n9448 0.0130799
R19243 vdd.n9434 vdd.n9433 0.0130799
R19244 vdd.n9474 vdd.n9463 0.0130799
R19245 vdd.n9474 vdd.n9468 0.0130799
R19246 vdd.n9483 vdd.n9477 0.0130799
R19247 vdd.n9477 vdd.n9476 0.0130799
R19248 vdd.n9501 vdd.n9470 0.0130799
R19249 vdd.n9502 vdd.n9501 0.0130799
R19250 vdd.n9497 vdd.n9496 0.0130799
R19251 vdd.n9482 vdd.n9481 0.0130799
R19252 vdd.n9520 vdd.n9509 0.0130799
R19253 vdd.n9520 vdd.n9514 0.0130799
R19254 vdd.n9529 vdd.n9523 0.0130799
R19255 vdd.n9523 vdd.n9522 0.0130799
R19256 vdd.n9547 vdd.n9516 0.0130799
R19257 vdd.n9548 vdd.n9547 0.0130799
R19258 vdd.n9543 vdd.n9542 0.0130799
R19259 vdd.n9528 vdd.n9527 0.0130799
R19260 vdd.n3680 vdd.n3669 0.0130799
R19261 vdd.n3680 vdd.n3674 0.0130799
R19262 vdd.n3689 vdd.n3683 0.0130799
R19263 vdd.n3683 vdd.n3682 0.0130799
R19264 vdd.n3707 vdd.n3676 0.0130799
R19265 vdd.n3708 vdd.n3707 0.0130799
R19266 vdd.n3703 vdd.n3702 0.0130799
R19267 vdd.n3688 vdd.n3687 0.0130799
R19268 vdd.n3726 vdd.n3715 0.0130799
R19269 vdd.n3726 vdd.n3720 0.0130799
R19270 vdd.n3735 vdd.n3729 0.0130799
R19271 vdd.n3729 vdd.n3728 0.0130799
R19272 vdd.n3753 vdd.n3722 0.0130799
R19273 vdd.n3754 vdd.n3753 0.0130799
R19274 vdd.n3749 vdd.n3748 0.0130799
R19275 vdd.n3734 vdd.n3733 0.0130799
R19276 vdd.n3824 vdd.n3813 0.0130799
R19277 vdd.n3824 vdd.n3818 0.0130799
R19278 vdd.n3833 vdd.n3827 0.0130799
R19279 vdd.n3827 vdd.n3826 0.0130799
R19280 vdd.n3851 vdd.n3820 0.0130799
R19281 vdd.n3852 vdd.n3851 0.0130799
R19282 vdd.n3847 vdd.n3846 0.0130799
R19283 vdd.n3832 vdd.n3831 0.0130799
R19284 vdd.n3870 vdd.n3859 0.0130799
R19285 vdd.n3870 vdd.n3864 0.0130799
R19286 vdd.n3879 vdd.n3873 0.0130799
R19287 vdd.n3873 vdd.n3872 0.0130799
R19288 vdd.n3897 vdd.n3866 0.0130799
R19289 vdd.n3898 vdd.n3897 0.0130799
R19290 vdd.n3893 vdd.n3892 0.0130799
R19291 vdd.n3878 vdd.n3877 0.0130799
R19292 vdd.n3916 vdd.n3905 0.0130799
R19293 vdd.n3916 vdd.n3910 0.0130799
R19294 vdd.n3925 vdd.n3919 0.0130799
R19295 vdd.n3919 vdd.n3918 0.0130799
R19296 vdd.n3943 vdd.n3912 0.0130799
R19297 vdd.n3944 vdd.n3943 0.0130799
R19298 vdd.n3939 vdd.n3938 0.0130799
R19299 vdd.n3924 vdd.n3923 0.0130799
R19300 vdd.n3962 vdd.n3951 0.0130799
R19301 vdd.n3962 vdd.n3956 0.0130799
R19302 vdd.n3971 vdd.n3965 0.0130799
R19303 vdd.n3965 vdd.n3964 0.0130799
R19304 vdd.n3989 vdd.n3958 0.0130799
R19305 vdd.n3990 vdd.n3989 0.0130799
R19306 vdd.n3985 vdd.n3984 0.0130799
R19307 vdd.n3970 vdd.n3969 0.0130799
R19308 vdd.n4060 vdd.n4049 0.0130799
R19309 vdd.n4060 vdd.n4054 0.0130799
R19310 vdd.n4069 vdd.n4063 0.0130799
R19311 vdd.n4063 vdd.n4062 0.0130799
R19312 vdd.n4087 vdd.n4056 0.0130799
R19313 vdd.n4088 vdd.n4087 0.0130799
R19314 vdd.n4083 vdd.n4082 0.0130799
R19315 vdd.n4068 vdd.n4067 0.0130799
R19316 vdd.n5518 vdd.n5507 0.0130799
R19317 vdd.n5518 vdd.n5512 0.0130799
R19318 vdd.n5527 vdd.n5521 0.0130799
R19319 vdd.n5521 vdd.n5520 0.0130799
R19320 vdd.n5545 vdd.n5514 0.0130799
R19321 vdd.n5546 vdd.n5545 0.0130799
R19322 vdd.n5541 vdd.n5540 0.0130799
R19323 vdd.n5526 vdd.n5525 0.0130799
R19324 vdd.n4108 vdd.n4097 0.0130799
R19325 vdd.n4109 vdd.n4108 0.0130799
R19326 vdd.n4125 vdd.n4101 0.0130799
R19327 vdd.n4130 vdd.n4101 0.0130799
R19328 vdd.n4116 vdd.n4110 0.0130799
R19329 vdd.n4110 vdd.n4107 0.0130799
R19330 vdd.n4115 vdd.n4111 0.0130799
R19331 vdd.n4133 vdd.n4132 0.0130799
R19332 vdd.n4154 vdd.n4143 0.0130799
R19333 vdd.n4155 vdd.n4154 0.0130799
R19334 vdd.n4171 vdd.n4147 0.0130799
R19335 vdd.n4176 vdd.n4147 0.0130799
R19336 vdd.n4162 vdd.n4156 0.0130799
R19337 vdd.n4156 vdd.n4153 0.0130799
R19338 vdd.n4161 vdd.n4157 0.0130799
R19339 vdd.n4179 vdd.n4178 0.0130799
R19340 vdd.n4251 vdd.n4240 0.0130799
R19341 vdd.n4252 vdd.n4251 0.0130799
R19342 vdd.n4268 vdd.n4244 0.0130799
R19343 vdd.n4273 vdd.n4244 0.0130799
R19344 vdd.n4259 vdd.n4253 0.0130799
R19345 vdd.n4253 vdd.n4250 0.0130799
R19346 vdd.n4258 vdd.n4254 0.0130799
R19347 vdd.n4276 vdd.n4275 0.0130799
R19348 vdd.n4297 vdd.n4286 0.0130799
R19349 vdd.n4298 vdd.n4297 0.0130799
R19350 vdd.n4314 vdd.n4290 0.0130799
R19351 vdd.n4319 vdd.n4290 0.0130799
R19352 vdd.n4305 vdd.n4299 0.0130799
R19353 vdd.n4299 vdd.n4296 0.0130799
R19354 vdd.n4304 vdd.n4300 0.0130799
R19355 vdd.n4322 vdd.n4321 0.0130799
R19356 vdd.n4343 vdd.n4332 0.0130799
R19357 vdd.n4344 vdd.n4343 0.0130799
R19358 vdd.n4360 vdd.n4336 0.0130799
R19359 vdd.n4365 vdd.n4336 0.0130799
R19360 vdd.n4351 vdd.n4345 0.0130799
R19361 vdd.n4345 vdd.n4342 0.0130799
R19362 vdd.n4350 vdd.n4346 0.0130799
R19363 vdd.n4368 vdd.n4367 0.0130799
R19364 vdd.n4389 vdd.n4378 0.0130799
R19365 vdd.n4390 vdd.n4389 0.0130799
R19366 vdd.n4406 vdd.n4382 0.0130799
R19367 vdd.n4411 vdd.n4382 0.0130799
R19368 vdd.n4397 vdd.n4391 0.0130799
R19369 vdd.n4391 vdd.n4388 0.0130799
R19370 vdd.n4396 vdd.n4392 0.0130799
R19371 vdd.n4414 vdd.n4413 0.0130799
R19372 vdd.n4486 vdd.n4475 0.0130799
R19373 vdd.n4487 vdd.n4486 0.0130799
R19374 vdd.n4503 vdd.n4479 0.0130799
R19375 vdd.n4508 vdd.n4479 0.0130799
R19376 vdd.n4494 vdd.n4488 0.0130799
R19377 vdd.n4488 vdd.n4485 0.0130799
R19378 vdd.n4493 vdd.n4489 0.0130799
R19379 vdd.n4511 vdd.n4510 0.0130799
R19380 vdd.n3635 vdd.n3624 0.0130799
R19381 vdd.n3636 vdd.n3635 0.0130799
R19382 vdd.n3652 vdd.n3628 0.0130799
R19383 vdd.n3657 vdd.n3628 0.0130799
R19384 vdd.n3643 vdd.n3637 0.0130799
R19385 vdd.n3637 vdd.n3634 0.0130799
R19386 vdd.n3642 vdd.n3638 0.0130799
R19387 vdd.n3660 vdd.n3659 0.0130799
R19388 vdd.n4530 vdd.n4519 0.0130799
R19389 vdd.n4531 vdd.n4530 0.0130799
R19390 vdd.n4547 vdd.n4523 0.0130799
R19391 vdd.n4552 vdd.n4523 0.0130799
R19392 vdd.n4538 vdd.n4532 0.0130799
R19393 vdd.n4532 vdd.n4529 0.0130799
R19394 vdd.n4537 vdd.n4533 0.0130799
R19395 vdd.n4555 vdd.n4554 0.0130799
R19396 vdd.n4575 vdd.n4564 0.0130799
R19397 vdd.n4576 vdd.n4575 0.0130799
R19398 vdd.n4592 vdd.n4568 0.0130799
R19399 vdd.n4597 vdd.n4568 0.0130799
R19400 vdd.n4583 vdd.n4577 0.0130799
R19401 vdd.n4577 vdd.n4574 0.0130799
R19402 vdd.n4582 vdd.n4578 0.0130799
R19403 vdd.n4600 vdd.n4599 0.0130799
R19404 vdd.n4625 vdd.n4614 0.0130799
R19405 vdd.n4626 vdd.n4625 0.0130799
R19406 vdd.n4642 vdd.n4618 0.0130799
R19407 vdd.n4647 vdd.n4618 0.0130799
R19408 vdd.n4633 vdd.n4627 0.0130799
R19409 vdd.n4627 vdd.n4624 0.0130799
R19410 vdd.n4632 vdd.n4628 0.0130799
R19411 vdd.n4650 vdd.n4649 0.0130799
R19412 vdd.n4671 vdd.n4660 0.0130799
R19413 vdd.n4672 vdd.n4671 0.0130799
R19414 vdd.n4688 vdd.n4664 0.0130799
R19415 vdd.n4693 vdd.n4664 0.0130799
R19416 vdd.n4679 vdd.n4673 0.0130799
R19417 vdd.n4673 vdd.n4670 0.0130799
R19418 vdd.n4678 vdd.n4674 0.0130799
R19419 vdd.n4696 vdd.n4695 0.0130799
R19420 vdd.n4719 vdd.n4708 0.0130799
R19421 vdd.n4720 vdd.n4719 0.0130799
R19422 vdd.n4736 vdd.n4712 0.0130799
R19423 vdd.n4741 vdd.n4712 0.0130799
R19424 vdd.n4727 vdd.n4721 0.0130799
R19425 vdd.n4721 vdd.n4718 0.0130799
R19426 vdd.n4726 vdd.n4722 0.0130799
R19427 vdd.n4744 vdd.n4743 0.0130799
R19428 vdd.n4437 vdd.n4430 0.0130799
R19429 vdd.n4437 vdd.n4436 0.0130799
R19430 vdd.n4448 vdd.n4433 0.0130799
R19431 vdd.n4453 vdd.n4433 0.0130799
R19432 vdd.n4439 vdd.n4427 0.0130799
R19433 vdd.n4428 vdd.n4427 0.0130799
R19434 vdd.n4426 vdd.n4424 0.0130799
R19435 vdd.n4456 vdd.n4455 0.0130799
R19436 vdd.n4766 vdd.n4755 0.0130799
R19437 vdd.n4767 vdd.n4766 0.0130799
R19438 vdd.n4783 vdd.n4759 0.0130799
R19439 vdd.n4788 vdd.n4759 0.0130799
R19440 vdd.n4774 vdd.n4768 0.0130799
R19441 vdd.n4768 vdd.n4765 0.0130799
R19442 vdd.n4773 vdd.n4769 0.0130799
R19443 vdd.n4791 vdd.n4790 0.0130799
R19444 vdd.n4811 vdd.n4800 0.0130799
R19445 vdd.n4812 vdd.n4811 0.0130799
R19446 vdd.n4828 vdd.n4804 0.0130799
R19447 vdd.n4833 vdd.n4804 0.0130799
R19448 vdd.n4819 vdd.n4813 0.0130799
R19449 vdd.n4813 vdd.n4810 0.0130799
R19450 vdd.n4818 vdd.n4814 0.0130799
R19451 vdd.n4836 vdd.n4835 0.0130799
R19452 vdd.n4857 vdd.n4846 0.0130799
R19453 vdd.n4858 vdd.n4857 0.0130799
R19454 vdd.n4874 vdd.n4850 0.0130799
R19455 vdd.n4879 vdd.n4850 0.0130799
R19456 vdd.n4865 vdd.n4859 0.0130799
R19457 vdd.n4859 vdd.n4856 0.0130799
R19458 vdd.n4864 vdd.n4860 0.0130799
R19459 vdd.n4882 vdd.n4881 0.0130799
R19460 vdd.n4908 vdd.n4897 0.0130799
R19461 vdd.n4909 vdd.n4908 0.0130799
R19462 vdd.n4925 vdd.n4901 0.0130799
R19463 vdd.n4930 vdd.n4901 0.0130799
R19464 vdd.n4916 vdd.n4910 0.0130799
R19465 vdd.n4910 vdd.n4907 0.0130799
R19466 vdd.n4915 vdd.n4911 0.0130799
R19467 vdd.n4933 vdd.n4932 0.0130799
R19468 vdd.n4954 vdd.n4943 0.0130799
R19469 vdd.n4955 vdd.n4954 0.0130799
R19470 vdd.n4971 vdd.n4947 0.0130799
R19471 vdd.n4976 vdd.n4947 0.0130799
R19472 vdd.n4962 vdd.n4956 0.0130799
R19473 vdd.n4956 vdd.n4953 0.0130799
R19474 vdd.n4961 vdd.n4957 0.0130799
R19475 vdd.n4979 vdd.n4978 0.0130799
R19476 vdd.n5002 vdd.n4991 0.0130799
R19477 vdd.n5003 vdd.n5002 0.0130799
R19478 vdd.n5019 vdd.n4995 0.0130799
R19479 vdd.n5024 vdd.n4995 0.0130799
R19480 vdd.n5010 vdd.n5004 0.0130799
R19481 vdd.n5004 vdd.n5001 0.0130799
R19482 vdd.n5009 vdd.n5005 0.0130799
R19483 vdd.n5027 vdd.n5026 0.0130799
R19484 vdd.n5048 vdd.n5037 0.0130799
R19485 vdd.n5049 vdd.n5048 0.0130799
R19486 vdd.n5065 vdd.n5041 0.0130799
R19487 vdd.n5070 vdd.n5041 0.0130799
R19488 vdd.n5056 vdd.n5050 0.0130799
R19489 vdd.n5050 vdd.n5047 0.0130799
R19490 vdd.n5055 vdd.n5051 0.0130799
R19491 vdd.n5073 vdd.n5072 0.0130799
R19492 vdd.n5093 vdd.n5082 0.0130799
R19493 vdd.n5094 vdd.n5093 0.0130799
R19494 vdd.n5110 vdd.n5086 0.0130799
R19495 vdd.n5115 vdd.n5086 0.0130799
R19496 vdd.n5101 vdd.n5095 0.0130799
R19497 vdd.n5095 vdd.n5092 0.0130799
R19498 vdd.n5100 vdd.n5096 0.0130799
R19499 vdd.n5118 vdd.n5117 0.0130799
R19500 vdd.n5143 vdd.n5132 0.0130799
R19501 vdd.n5144 vdd.n5143 0.0130799
R19502 vdd.n5160 vdd.n5136 0.0130799
R19503 vdd.n5165 vdd.n5136 0.0130799
R19504 vdd.n5151 vdd.n5145 0.0130799
R19505 vdd.n5145 vdd.n5142 0.0130799
R19506 vdd.n5150 vdd.n5146 0.0130799
R19507 vdd.n5168 vdd.n5167 0.0130799
R19508 vdd.n5189 vdd.n5178 0.0130799
R19509 vdd.n5190 vdd.n5189 0.0130799
R19510 vdd.n5206 vdd.n5182 0.0130799
R19511 vdd.n5211 vdd.n5182 0.0130799
R19512 vdd.n5197 vdd.n5191 0.0130799
R19513 vdd.n5191 vdd.n5188 0.0130799
R19514 vdd.n5196 vdd.n5192 0.0130799
R19515 vdd.n5214 vdd.n5213 0.0130799
R19516 vdd.n5237 vdd.n5226 0.0130799
R19517 vdd.n5238 vdd.n5237 0.0130799
R19518 vdd.n5254 vdd.n5230 0.0130799
R19519 vdd.n5259 vdd.n5230 0.0130799
R19520 vdd.n5245 vdd.n5239 0.0130799
R19521 vdd.n5239 vdd.n5236 0.0130799
R19522 vdd.n5244 vdd.n5240 0.0130799
R19523 vdd.n5262 vdd.n5261 0.0130799
R19524 vdd.n4202 vdd.n4195 0.0130799
R19525 vdd.n4202 vdd.n4201 0.0130799
R19526 vdd.n4213 vdd.n4198 0.0130799
R19527 vdd.n4218 vdd.n4198 0.0130799
R19528 vdd.n4204 vdd.n4192 0.0130799
R19529 vdd.n4193 vdd.n4192 0.0130799
R19530 vdd.n4191 vdd.n4189 0.0130799
R19531 vdd.n4221 vdd.n4220 0.0130799
R19532 vdd.n5284 vdd.n5273 0.0130799
R19533 vdd.n5285 vdd.n5284 0.0130799
R19534 vdd.n5301 vdd.n5277 0.0130799
R19535 vdd.n5306 vdd.n5277 0.0130799
R19536 vdd.n5292 vdd.n5286 0.0130799
R19537 vdd.n5286 vdd.n5283 0.0130799
R19538 vdd.n5291 vdd.n5287 0.0130799
R19539 vdd.n5309 vdd.n5308 0.0130799
R19540 vdd.n5329 vdd.n5318 0.0130799
R19541 vdd.n5330 vdd.n5329 0.0130799
R19542 vdd.n5346 vdd.n5322 0.0130799
R19543 vdd.n5351 vdd.n5322 0.0130799
R19544 vdd.n5337 vdd.n5331 0.0130799
R19545 vdd.n5331 vdd.n5328 0.0130799
R19546 vdd.n5336 vdd.n5332 0.0130799
R19547 vdd.n5354 vdd.n5353 0.0130799
R19548 vdd.n5379 vdd.n5368 0.0130799
R19549 vdd.n5380 vdd.n5379 0.0130799
R19550 vdd.n5396 vdd.n5372 0.0130799
R19551 vdd.n5401 vdd.n5372 0.0130799
R19552 vdd.n5387 vdd.n5381 0.0130799
R19553 vdd.n5381 vdd.n5378 0.0130799
R19554 vdd.n5386 vdd.n5382 0.0130799
R19555 vdd.n5404 vdd.n5403 0.0130799
R19556 vdd.n5425 vdd.n5414 0.0130799
R19557 vdd.n5426 vdd.n5425 0.0130799
R19558 vdd.n5442 vdd.n5418 0.0130799
R19559 vdd.n5447 vdd.n5418 0.0130799
R19560 vdd.n5433 vdd.n5427 0.0130799
R19561 vdd.n5427 vdd.n5424 0.0130799
R19562 vdd.n5432 vdd.n5428 0.0130799
R19563 vdd.n5450 vdd.n5449 0.0130799
R19564 vdd.n5473 vdd.n5462 0.0130799
R19565 vdd.n5474 vdd.n5473 0.0130799
R19566 vdd.n5490 vdd.n5466 0.0130799
R19567 vdd.n5495 vdd.n5466 0.0130799
R19568 vdd.n5481 vdd.n5475 0.0130799
R19569 vdd.n5475 vdd.n5472 0.0130799
R19570 vdd.n5480 vdd.n5476 0.0130799
R19571 vdd.n5498 vdd.n5497 0.0130799
R19572 vdd.n5611 vdd.n5600 0.0130799
R19573 vdd.n5611 vdd.n5605 0.0130799
R19574 vdd.n5620 vdd.n5614 0.0130799
R19575 vdd.n5614 vdd.n5613 0.0130799
R19576 vdd.n5638 vdd.n5607 0.0130799
R19577 vdd.n5639 vdd.n5638 0.0130799
R19578 vdd.n5634 vdd.n5633 0.0130799
R19579 vdd.n5619 vdd.n5618 0.0130799
R19580 vdd.n5565 vdd.n5554 0.0130799
R19581 vdd.n5565 vdd.n5559 0.0130799
R19582 vdd.n5574 vdd.n5568 0.0130799
R19583 vdd.n5568 vdd.n5567 0.0130799
R19584 vdd.n5592 vdd.n5561 0.0130799
R19585 vdd.n5593 vdd.n5592 0.0130799
R19586 vdd.n5588 vdd.n5587 0.0130799
R19587 vdd.n5573 vdd.n5572 0.0130799
R19588 vdd.n5658 vdd.n5647 0.0130799
R19589 vdd.n5658 vdd.n5652 0.0130799
R19590 vdd.n5667 vdd.n5661 0.0130799
R19591 vdd.n5661 vdd.n5660 0.0130799
R19592 vdd.n5685 vdd.n5654 0.0130799
R19593 vdd.n5686 vdd.n5685 0.0130799
R19594 vdd.n5681 vdd.n5680 0.0130799
R19595 vdd.n5666 vdd.n5665 0.0130799
R19596 vdd.n5706 vdd.n5695 0.0130799
R19597 vdd.n5706 vdd.n5700 0.0130799
R19598 vdd.n5715 vdd.n5709 0.0130799
R19599 vdd.n5709 vdd.n5708 0.0130799
R19600 vdd.n5733 vdd.n5702 0.0130799
R19601 vdd.n5734 vdd.n5733 0.0130799
R19602 vdd.n5729 vdd.n5728 0.0130799
R19603 vdd.n5714 vdd.n5713 0.0130799
R19604 vdd.n5752 vdd.n5741 0.0130799
R19605 vdd.n5752 vdd.n5746 0.0130799
R19606 vdd.n5761 vdd.n5755 0.0130799
R19607 vdd.n5755 vdd.n5754 0.0130799
R19608 vdd.n5779 vdd.n5748 0.0130799
R19609 vdd.n5780 vdd.n5779 0.0130799
R19610 vdd.n5775 vdd.n5774 0.0130799
R19611 vdd.n5760 vdd.n5759 0.0130799
R19612 vdd.n4011 vdd.n4005 0.0130799
R19613 vdd.n4028 vdd.n4011 0.0130799
R19614 vdd.n4016 vdd.n4013 0.0130799
R19615 vdd.n4016 vdd.n4009 0.0130799
R19616 vdd.n4037 vdd.n4036 0.0130799
R19617 vdd.n4037 vdd.n4003 0.0130799
R19618 vdd.n4043 vdd.n4000 0.0130799
R19619 vdd.n4015 vdd.n4014 0.0130799
R19620 vdd.n5894 vdd.n5883 0.0130799
R19621 vdd.n5894 vdd.n5888 0.0130799
R19622 vdd.n5903 vdd.n5897 0.0130799
R19623 vdd.n5897 vdd.n5896 0.0130799
R19624 vdd.n5921 vdd.n5890 0.0130799
R19625 vdd.n5922 vdd.n5921 0.0130799
R19626 vdd.n5917 vdd.n5916 0.0130799
R19627 vdd.n5902 vdd.n5901 0.0130799
R19628 vdd.n5847 vdd.n5836 0.0130799
R19629 vdd.n5847 vdd.n5841 0.0130799
R19630 vdd.n5856 vdd.n5850 0.0130799
R19631 vdd.n5850 vdd.n5849 0.0130799
R19632 vdd.n5874 vdd.n5843 0.0130799
R19633 vdd.n5875 vdd.n5874 0.0130799
R19634 vdd.n5870 vdd.n5869 0.0130799
R19635 vdd.n5855 vdd.n5854 0.0130799
R19636 vdd.n5801 vdd.n5790 0.0130799
R19637 vdd.n5801 vdd.n5795 0.0130799
R19638 vdd.n5810 vdd.n5804 0.0130799
R19639 vdd.n5804 vdd.n5803 0.0130799
R19640 vdd.n5828 vdd.n5797 0.0130799
R19641 vdd.n5829 vdd.n5828 0.0130799
R19642 vdd.n5824 vdd.n5823 0.0130799
R19643 vdd.n5809 vdd.n5808 0.0130799
R19644 vdd.n5941 vdd.n5930 0.0130799
R19645 vdd.n5941 vdd.n5935 0.0130799
R19646 vdd.n5950 vdd.n5944 0.0130799
R19647 vdd.n5944 vdd.n5943 0.0130799
R19648 vdd.n5968 vdd.n5937 0.0130799
R19649 vdd.n5969 vdd.n5968 0.0130799
R19650 vdd.n5964 vdd.n5963 0.0130799
R19651 vdd.n5949 vdd.n5948 0.0130799
R19652 vdd.n5989 vdd.n5978 0.0130799
R19653 vdd.n5989 vdd.n5983 0.0130799
R19654 vdd.n5998 vdd.n5992 0.0130799
R19655 vdd.n5992 vdd.n5991 0.0130799
R19656 vdd.n6016 vdd.n5985 0.0130799
R19657 vdd.n6017 vdd.n6016 0.0130799
R19658 vdd.n6012 vdd.n6011 0.0130799
R19659 vdd.n5997 vdd.n5996 0.0130799
R19660 vdd.n6035 vdd.n6024 0.0130799
R19661 vdd.n6035 vdd.n6029 0.0130799
R19662 vdd.n6044 vdd.n6038 0.0130799
R19663 vdd.n6038 vdd.n6037 0.0130799
R19664 vdd.n6062 vdd.n6031 0.0130799
R19665 vdd.n6063 vdd.n6062 0.0130799
R19666 vdd.n6058 vdd.n6057 0.0130799
R19667 vdd.n6043 vdd.n6042 0.0130799
R19668 vdd.n6129 vdd.n6118 0.0130799
R19669 vdd.n6129 vdd.n6123 0.0130799
R19670 vdd.n6138 vdd.n6132 0.0130799
R19671 vdd.n6132 vdd.n6131 0.0130799
R19672 vdd.n6156 vdd.n6125 0.0130799
R19673 vdd.n6157 vdd.n6156 0.0130799
R19674 vdd.n6152 vdd.n6151 0.0130799
R19675 vdd.n6137 vdd.n6136 0.0130799
R19676 vdd.n6083 vdd.n6072 0.0130799
R19677 vdd.n6083 vdd.n6077 0.0130799
R19678 vdd.n6092 vdd.n6086 0.0130799
R19679 vdd.n6086 vdd.n6085 0.0130799
R19680 vdd.n6110 vdd.n6079 0.0130799
R19681 vdd.n6111 vdd.n6110 0.0130799
R19682 vdd.n6106 vdd.n6105 0.0130799
R19683 vdd.n6091 vdd.n6090 0.0130799
R19684 vdd.n6176 vdd.n6165 0.0130799
R19685 vdd.n6176 vdd.n6170 0.0130799
R19686 vdd.n6185 vdd.n6179 0.0130799
R19687 vdd.n6179 vdd.n6178 0.0130799
R19688 vdd.n6203 vdd.n6172 0.0130799
R19689 vdd.n6204 vdd.n6203 0.0130799
R19690 vdd.n6199 vdd.n6198 0.0130799
R19691 vdd.n6184 vdd.n6183 0.0130799
R19692 vdd.n6224 vdd.n6213 0.0130799
R19693 vdd.n6224 vdd.n6218 0.0130799
R19694 vdd.n6233 vdd.n6227 0.0130799
R19695 vdd.n6227 vdd.n6226 0.0130799
R19696 vdd.n6251 vdd.n6220 0.0130799
R19697 vdd.n6252 vdd.n6251 0.0130799
R19698 vdd.n6247 vdd.n6246 0.0130799
R19699 vdd.n6232 vdd.n6231 0.0130799
R19700 vdd.n6270 vdd.n6259 0.0130799
R19701 vdd.n6270 vdd.n6264 0.0130799
R19702 vdd.n6279 vdd.n6273 0.0130799
R19703 vdd.n6273 vdd.n6272 0.0130799
R19704 vdd.n6297 vdd.n6266 0.0130799
R19705 vdd.n6298 vdd.n6297 0.0130799
R19706 vdd.n6293 vdd.n6292 0.0130799
R19707 vdd.n6278 vdd.n6277 0.0130799
R19708 vdd.n3775 vdd.n3769 0.0130799
R19709 vdd.n3792 vdd.n3775 0.0130799
R19710 vdd.n3780 vdd.n3777 0.0130799
R19711 vdd.n3780 vdd.n3773 0.0130799
R19712 vdd.n3801 vdd.n3800 0.0130799
R19713 vdd.n3801 vdd.n3767 0.0130799
R19714 vdd.n3807 vdd.n3764 0.0130799
R19715 vdd.n3779 vdd.n3778 0.0130799
R19716 vdd.n6365 vdd.n6354 0.0130799
R19717 vdd.n6365 vdd.n6359 0.0130799
R19718 vdd.n6374 vdd.n6368 0.0130799
R19719 vdd.n6368 vdd.n6367 0.0130799
R19720 vdd.n6392 vdd.n6361 0.0130799
R19721 vdd.n6393 vdd.n6392 0.0130799
R19722 vdd.n6388 vdd.n6387 0.0130799
R19723 vdd.n6373 vdd.n6372 0.0130799
R19724 vdd.n6319 vdd.n6308 0.0130799
R19725 vdd.n6319 vdd.n6313 0.0130799
R19726 vdd.n6328 vdd.n6322 0.0130799
R19727 vdd.n6322 vdd.n6321 0.0130799
R19728 vdd.n6346 vdd.n6315 0.0130799
R19729 vdd.n6347 vdd.n6346 0.0130799
R19730 vdd.n6342 vdd.n6341 0.0130799
R19731 vdd.n6327 vdd.n6326 0.0130799
R19732 vdd.n6412 vdd.n6401 0.0130799
R19733 vdd.n6412 vdd.n6406 0.0130799
R19734 vdd.n6421 vdd.n6415 0.0130799
R19735 vdd.n6415 vdd.n6414 0.0130799
R19736 vdd.n6439 vdd.n6408 0.0130799
R19737 vdd.n6440 vdd.n6439 0.0130799
R19738 vdd.n6435 vdd.n6434 0.0130799
R19739 vdd.n6420 vdd.n6419 0.0130799
R19740 vdd.n6460 vdd.n6449 0.0130799
R19741 vdd.n6460 vdd.n6454 0.0130799
R19742 vdd.n6469 vdd.n6463 0.0130799
R19743 vdd.n6463 vdd.n6462 0.0130799
R19744 vdd.n6487 vdd.n6456 0.0130799
R19745 vdd.n6488 vdd.n6487 0.0130799
R19746 vdd.n6483 vdd.n6482 0.0130799
R19747 vdd.n6468 vdd.n6467 0.0130799
R19748 vdd.n6506 vdd.n6495 0.0130799
R19749 vdd.n6506 vdd.n6500 0.0130799
R19750 vdd.n6515 vdd.n6509 0.0130799
R19751 vdd.n6509 vdd.n6508 0.0130799
R19752 vdd.n6533 vdd.n6502 0.0130799
R19753 vdd.n6534 vdd.n6533 0.0130799
R19754 vdd.n6529 vdd.n6528 0.0130799
R19755 vdd.n6514 vdd.n6513 0.0130799
R19756 vdd.n666 vdd.n655 0.0130799
R19757 vdd.n666 vdd.n660 0.0130799
R19758 vdd.n675 vdd.n669 0.0130799
R19759 vdd.n669 vdd.n668 0.0130799
R19760 vdd.n693 vdd.n662 0.0130799
R19761 vdd.n694 vdd.n693 0.0130799
R19762 vdd.n689 vdd.n688 0.0130799
R19763 vdd.n674 vdd.n673 0.0130799
R19764 vdd.n712 vdd.n701 0.0130799
R19765 vdd.n712 vdd.n706 0.0130799
R19766 vdd.n721 vdd.n715 0.0130799
R19767 vdd.n715 vdd.n714 0.0130799
R19768 vdd.n739 vdd.n708 0.0130799
R19769 vdd.n740 vdd.n739 0.0130799
R19770 vdd.n735 vdd.n734 0.0130799
R19771 vdd.n720 vdd.n719 0.0130799
R19772 vdd.n810 vdd.n799 0.0130799
R19773 vdd.n810 vdd.n804 0.0130799
R19774 vdd.n819 vdd.n813 0.0130799
R19775 vdd.n813 vdd.n812 0.0130799
R19776 vdd.n837 vdd.n806 0.0130799
R19777 vdd.n838 vdd.n837 0.0130799
R19778 vdd.n833 vdd.n832 0.0130799
R19779 vdd.n818 vdd.n817 0.0130799
R19780 vdd.n856 vdd.n845 0.0130799
R19781 vdd.n856 vdd.n850 0.0130799
R19782 vdd.n865 vdd.n859 0.0130799
R19783 vdd.n859 vdd.n858 0.0130799
R19784 vdd.n883 vdd.n852 0.0130799
R19785 vdd.n884 vdd.n883 0.0130799
R19786 vdd.n879 vdd.n878 0.0130799
R19787 vdd.n864 vdd.n863 0.0130799
R19788 vdd.n902 vdd.n891 0.0130799
R19789 vdd.n902 vdd.n896 0.0130799
R19790 vdd.n911 vdd.n905 0.0130799
R19791 vdd.n905 vdd.n904 0.0130799
R19792 vdd.n929 vdd.n898 0.0130799
R19793 vdd.n930 vdd.n929 0.0130799
R19794 vdd.n925 vdd.n924 0.0130799
R19795 vdd.n910 vdd.n909 0.0130799
R19796 vdd.n948 vdd.n937 0.0130799
R19797 vdd.n948 vdd.n942 0.0130799
R19798 vdd.n957 vdd.n951 0.0130799
R19799 vdd.n951 vdd.n950 0.0130799
R19800 vdd.n975 vdd.n944 0.0130799
R19801 vdd.n976 vdd.n975 0.0130799
R19802 vdd.n971 vdd.n970 0.0130799
R19803 vdd.n956 vdd.n955 0.0130799
R19804 vdd.n1046 vdd.n1035 0.0130799
R19805 vdd.n1046 vdd.n1040 0.0130799
R19806 vdd.n1055 vdd.n1049 0.0130799
R19807 vdd.n1049 vdd.n1048 0.0130799
R19808 vdd.n1073 vdd.n1042 0.0130799
R19809 vdd.n1074 vdd.n1073 0.0130799
R19810 vdd.n1069 vdd.n1068 0.0130799
R19811 vdd.n1054 vdd.n1053 0.0130799
R19812 vdd.n2504 vdd.n2493 0.0130799
R19813 vdd.n2504 vdd.n2498 0.0130799
R19814 vdd.n2513 vdd.n2507 0.0130799
R19815 vdd.n2507 vdd.n2506 0.0130799
R19816 vdd.n2531 vdd.n2500 0.0130799
R19817 vdd.n2532 vdd.n2531 0.0130799
R19818 vdd.n2527 vdd.n2526 0.0130799
R19819 vdd.n2512 vdd.n2511 0.0130799
R19820 vdd.n1094 vdd.n1083 0.0130799
R19821 vdd.n1095 vdd.n1094 0.0130799
R19822 vdd.n1111 vdd.n1087 0.0130799
R19823 vdd.n1116 vdd.n1087 0.0130799
R19824 vdd.n1102 vdd.n1096 0.0130799
R19825 vdd.n1096 vdd.n1093 0.0130799
R19826 vdd.n1101 vdd.n1097 0.0130799
R19827 vdd.n1119 vdd.n1118 0.0130799
R19828 vdd.n1140 vdd.n1129 0.0130799
R19829 vdd.n1141 vdd.n1140 0.0130799
R19830 vdd.n1157 vdd.n1133 0.0130799
R19831 vdd.n1162 vdd.n1133 0.0130799
R19832 vdd.n1148 vdd.n1142 0.0130799
R19833 vdd.n1142 vdd.n1139 0.0130799
R19834 vdd.n1147 vdd.n1143 0.0130799
R19835 vdd.n1165 vdd.n1164 0.0130799
R19836 vdd.n1237 vdd.n1226 0.0130799
R19837 vdd.n1238 vdd.n1237 0.0130799
R19838 vdd.n1254 vdd.n1230 0.0130799
R19839 vdd.n1259 vdd.n1230 0.0130799
R19840 vdd.n1245 vdd.n1239 0.0130799
R19841 vdd.n1239 vdd.n1236 0.0130799
R19842 vdd.n1244 vdd.n1240 0.0130799
R19843 vdd.n1262 vdd.n1261 0.0130799
R19844 vdd.n1283 vdd.n1272 0.0130799
R19845 vdd.n1284 vdd.n1283 0.0130799
R19846 vdd.n1300 vdd.n1276 0.0130799
R19847 vdd.n1305 vdd.n1276 0.0130799
R19848 vdd.n1291 vdd.n1285 0.0130799
R19849 vdd.n1285 vdd.n1282 0.0130799
R19850 vdd.n1290 vdd.n1286 0.0130799
R19851 vdd.n1308 vdd.n1307 0.0130799
R19852 vdd.n1329 vdd.n1318 0.0130799
R19853 vdd.n1330 vdd.n1329 0.0130799
R19854 vdd.n1346 vdd.n1322 0.0130799
R19855 vdd.n1351 vdd.n1322 0.0130799
R19856 vdd.n1337 vdd.n1331 0.0130799
R19857 vdd.n1331 vdd.n1328 0.0130799
R19858 vdd.n1336 vdd.n1332 0.0130799
R19859 vdd.n1354 vdd.n1353 0.0130799
R19860 vdd.n1375 vdd.n1364 0.0130799
R19861 vdd.n1376 vdd.n1375 0.0130799
R19862 vdd.n1392 vdd.n1368 0.0130799
R19863 vdd.n1397 vdd.n1368 0.0130799
R19864 vdd.n1383 vdd.n1377 0.0130799
R19865 vdd.n1377 vdd.n1374 0.0130799
R19866 vdd.n1382 vdd.n1378 0.0130799
R19867 vdd.n1400 vdd.n1399 0.0130799
R19868 vdd.n1472 vdd.n1461 0.0130799
R19869 vdd.n1473 vdd.n1472 0.0130799
R19870 vdd.n1489 vdd.n1465 0.0130799
R19871 vdd.n1494 vdd.n1465 0.0130799
R19872 vdd.n1480 vdd.n1474 0.0130799
R19873 vdd.n1474 vdd.n1471 0.0130799
R19874 vdd.n1479 vdd.n1475 0.0130799
R19875 vdd.n1497 vdd.n1496 0.0130799
R19876 vdd.n621 vdd.n610 0.0130799
R19877 vdd.n622 vdd.n621 0.0130799
R19878 vdd.n638 vdd.n614 0.0130799
R19879 vdd.n643 vdd.n614 0.0130799
R19880 vdd.n629 vdd.n623 0.0130799
R19881 vdd.n623 vdd.n620 0.0130799
R19882 vdd.n628 vdd.n624 0.0130799
R19883 vdd.n646 vdd.n645 0.0130799
R19884 vdd.n1516 vdd.n1505 0.0130799
R19885 vdd.n1517 vdd.n1516 0.0130799
R19886 vdd.n1533 vdd.n1509 0.0130799
R19887 vdd.n1538 vdd.n1509 0.0130799
R19888 vdd.n1524 vdd.n1518 0.0130799
R19889 vdd.n1518 vdd.n1515 0.0130799
R19890 vdd.n1523 vdd.n1519 0.0130799
R19891 vdd.n1541 vdd.n1540 0.0130799
R19892 vdd.n1561 vdd.n1550 0.0130799
R19893 vdd.n1562 vdd.n1561 0.0130799
R19894 vdd.n1578 vdd.n1554 0.0130799
R19895 vdd.n1583 vdd.n1554 0.0130799
R19896 vdd.n1569 vdd.n1563 0.0130799
R19897 vdd.n1563 vdd.n1560 0.0130799
R19898 vdd.n1568 vdd.n1564 0.0130799
R19899 vdd.n1586 vdd.n1585 0.0130799
R19900 vdd.n1611 vdd.n1600 0.0130799
R19901 vdd.n1612 vdd.n1611 0.0130799
R19902 vdd.n1628 vdd.n1604 0.0130799
R19903 vdd.n1633 vdd.n1604 0.0130799
R19904 vdd.n1619 vdd.n1613 0.0130799
R19905 vdd.n1613 vdd.n1610 0.0130799
R19906 vdd.n1618 vdd.n1614 0.0130799
R19907 vdd.n1636 vdd.n1635 0.0130799
R19908 vdd.n1657 vdd.n1646 0.0130799
R19909 vdd.n1658 vdd.n1657 0.0130799
R19910 vdd.n1674 vdd.n1650 0.0130799
R19911 vdd.n1679 vdd.n1650 0.0130799
R19912 vdd.n1665 vdd.n1659 0.0130799
R19913 vdd.n1659 vdd.n1656 0.0130799
R19914 vdd.n1664 vdd.n1660 0.0130799
R19915 vdd.n1682 vdd.n1681 0.0130799
R19916 vdd.n1705 vdd.n1694 0.0130799
R19917 vdd.n1706 vdd.n1705 0.0130799
R19918 vdd.n1722 vdd.n1698 0.0130799
R19919 vdd.n1727 vdd.n1698 0.0130799
R19920 vdd.n1713 vdd.n1707 0.0130799
R19921 vdd.n1707 vdd.n1704 0.0130799
R19922 vdd.n1712 vdd.n1708 0.0130799
R19923 vdd.n1730 vdd.n1729 0.0130799
R19924 vdd.n1423 vdd.n1416 0.0130799
R19925 vdd.n1423 vdd.n1422 0.0130799
R19926 vdd.n1434 vdd.n1419 0.0130799
R19927 vdd.n1439 vdd.n1419 0.0130799
R19928 vdd.n1425 vdd.n1413 0.0130799
R19929 vdd.n1414 vdd.n1413 0.0130799
R19930 vdd.n1412 vdd.n1410 0.0130799
R19931 vdd.n1442 vdd.n1441 0.0130799
R19932 vdd.n1752 vdd.n1741 0.0130799
R19933 vdd.n1753 vdd.n1752 0.0130799
R19934 vdd.n1769 vdd.n1745 0.0130799
R19935 vdd.n1774 vdd.n1745 0.0130799
R19936 vdd.n1760 vdd.n1754 0.0130799
R19937 vdd.n1754 vdd.n1751 0.0130799
R19938 vdd.n1759 vdd.n1755 0.0130799
R19939 vdd.n1777 vdd.n1776 0.0130799
R19940 vdd.n1797 vdd.n1786 0.0130799
R19941 vdd.n1798 vdd.n1797 0.0130799
R19942 vdd.n1814 vdd.n1790 0.0130799
R19943 vdd.n1819 vdd.n1790 0.0130799
R19944 vdd.n1805 vdd.n1799 0.0130799
R19945 vdd.n1799 vdd.n1796 0.0130799
R19946 vdd.n1804 vdd.n1800 0.0130799
R19947 vdd.n1822 vdd.n1821 0.0130799
R19948 vdd.n1843 vdd.n1832 0.0130799
R19949 vdd.n1844 vdd.n1843 0.0130799
R19950 vdd.n1860 vdd.n1836 0.0130799
R19951 vdd.n1865 vdd.n1836 0.0130799
R19952 vdd.n1851 vdd.n1845 0.0130799
R19953 vdd.n1845 vdd.n1842 0.0130799
R19954 vdd.n1850 vdd.n1846 0.0130799
R19955 vdd.n1868 vdd.n1867 0.0130799
R19956 vdd.n1894 vdd.n1883 0.0130799
R19957 vdd.n1895 vdd.n1894 0.0130799
R19958 vdd.n1911 vdd.n1887 0.0130799
R19959 vdd.n1916 vdd.n1887 0.0130799
R19960 vdd.n1902 vdd.n1896 0.0130799
R19961 vdd.n1896 vdd.n1893 0.0130799
R19962 vdd.n1901 vdd.n1897 0.0130799
R19963 vdd.n1919 vdd.n1918 0.0130799
R19964 vdd.n1940 vdd.n1929 0.0130799
R19965 vdd.n1941 vdd.n1940 0.0130799
R19966 vdd.n1957 vdd.n1933 0.0130799
R19967 vdd.n1962 vdd.n1933 0.0130799
R19968 vdd.n1948 vdd.n1942 0.0130799
R19969 vdd.n1942 vdd.n1939 0.0130799
R19970 vdd.n1947 vdd.n1943 0.0130799
R19971 vdd.n1965 vdd.n1964 0.0130799
R19972 vdd.n1988 vdd.n1977 0.0130799
R19973 vdd.n1989 vdd.n1988 0.0130799
R19974 vdd.n2005 vdd.n1981 0.0130799
R19975 vdd.n2010 vdd.n1981 0.0130799
R19976 vdd.n1996 vdd.n1990 0.0130799
R19977 vdd.n1990 vdd.n1987 0.0130799
R19978 vdd.n1995 vdd.n1991 0.0130799
R19979 vdd.n2013 vdd.n2012 0.0130799
R19980 vdd.n2034 vdd.n2023 0.0130799
R19981 vdd.n2035 vdd.n2034 0.0130799
R19982 vdd.n2051 vdd.n2027 0.0130799
R19983 vdd.n2056 vdd.n2027 0.0130799
R19984 vdd.n2042 vdd.n2036 0.0130799
R19985 vdd.n2036 vdd.n2033 0.0130799
R19986 vdd.n2041 vdd.n2037 0.0130799
R19987 vdd.n2059 vdd.n2058 0.0130799
R19988 vdd.n2079 vdd.n2068 0.0130799
R19989 vdd.n2080 vdd.n2079 0.0130799
R19990 vdd.n2096 vdd.n2072 0.0130799
R19991 vdd.n2101 vdd.n2072 0.0130799
R19992 vdd.n2087 vdd.n2081 0.0130799
R19993 vdd.n2081 vdd.n2078 0.0130799
R19994 vdd.n2086 vdd.n2082 0.0130799
R19995 vdd.n2104 vdd.n2103 0.0130799
R19996 vdd.n2129 vdd.n2118 0.0130799
R19997 vdd.n2130 vdd.n2129 0.0130799
R19998 vdd.n2146 vdd.n2122 0.0130799
R19999 vdd.n2151 vdd.n2122 0.0130799
R20000 vdd.n2137 vdd.n2131 0.0130799
R20001 vdd.n2131 vdd.n2128 0.0130799
R20002 vdd.n2136 vdd.n2132 0.0130799
R20003 vdd.n2154 vdd.n2153 0.0130799
R20004 vdd.n2175 vdd.n2164 0.0130799
R20005 vdd.n2176 vdd.n2175 0.0130799
R20006 vdd.n2192 vdd.n2168 0.0130799
R20007 vdd.n2197 vdd.n2168 0.0130799
R20008 vdd.n2183 vdd.n2177 0.0130799
R20009 vdd.n2177 vdd.n2174 0.0130799
R20010 vdd.n2182 vdd.n2178 0.0130799
R20011 vdd.n2200 vdd.n2199 0.0130799
R20012 vdd.n2223 vdd.n2212 0.0130799
R20013 vdd.n2224 vdd.n2223 0.0130799
R20014 vdd.n2240 vdd.n2216 0.0130799
R20015 vdd.n2245 vdd.n2216 0.0130799
R20016 vdd.n2231 vdd.n2225 0.0130799
R20017 vdd.n2225 vdd.n2222 0.0130799
R20018 vdd.n2230 vdd.n2226 0.0130799
R20019 vdd.n2248 vdd.n2247 0.0130799
R20020 vdd.n1188 vdd.n1181 0.0130799
R20021 vdd.n1188 vdd.n1187 0.0130799
R20022 vdd.n1199 vdd.n1184 0.0130799
R20023 vdd.n1204 vdd.n1184 0.0130799
R20024 vdd.n1190 vdd.n1178 0.0130799
R20025 vdd.n1179 vdd.n1178 0.0130799
R20026 vdd.n1177 vdd.n1175 0.0130799
R20027 vdd.n1207 vdd.n1206 0.0130799
R20028 vdd.n2270 vdd.n2259 0.0130799
R20029 vdd.n2271 vdd.n2270 0.0130799
R20030 vdd.n2287 vdd.n2263 0.0130799
R20031 vdd.n2292 vdd.n2263 0.0130799
R20032 vdd.n2278 vdd.n2272 0.0130799
R20033 vdd.n2272 vdd.n2269 0.0130799
R20034 vdd.n2277 vdd.n2273 0.0130799
R20035 vdd.n2295 vdd.n2294 0.0130799
R20036 vdd.n2315 vdd.n2304 0.0130799
R20037 vdd.n2316 vdd.n2315 0.0130799
R20038 vdd.n2332 vdd.n2308 0.0130799
R20039 vdd.n2337 vdd.n2308 0.0130799
R20040 vdd.n2323 vdd.n2317 0.0130799
R20041 vdd.n2317 vdd.n2314 0.0130799
R20042 vdd.n2322 vdd.n2318 0.0130799
R20043 vdd.n2340 vdd.n2339 0.0130799
R20044 vdd.n2365 vdd.n2354 0.0130799
R20045 vdd.n2366 vdd.n2365 0.0130799
R20046 vdd.n2382 vdd.n2358 0.0130799
R20047 vdd.n2387 vdd.n2358 0.0130799
R20048 vdd.n2373 vdd.n2367 0.0130799
R20049 vdd.n2367 vdd.n2364 0.0130799
R20050 vdd.n2372 vdd.n2368 0.0130799
R20051 vdd.n2390 vdd.n2389 0.0130799
R20052 vdd.n2411 vdd.n2400 0.0130799
R20053 vdd.n2412 vdd.n2411 0.0130799
R20054 vdd.n2428 vdd.n2404 0.0130799
R20055 vdd.n2433 vdd.n2404 0.0130799
R20056 vdd.n2419 vdd.n2413 0.0130799
R20057 vdd.n2413 vdd.n2410 0.0130799
R20058 vdd.n2418 vdd.n2414 0.0130799
R20059 vdd.n2436 vdd.n2435 0.0130799
R20060 vdd.n2459 vdd.n2448 0.0130799
R20061 vdd.n2460 vdd.n2459 0.0130799
R20062 vdd.n2476 vdd.n2452 0.0130799
R20063 vdd.n2481 vdd.n2452 0.0130799
R20064 vdd.n2467 vdd.n2461 0.0130799
R20065 vdd.n2461 vdd.n2458 0.0130799
R20066 vdd.n2466 vdd.n2462 0.0130799
R20067 vdd.n2484 vdd.n2483 0.0130799
R20068 vdd.n2597 vdd.n2586 0.0130799
R20069 vdd.n2597 vdd.n2591 0.0130799
R20070 vdd.n2606 vdd.n2600 0.0130799
R20071 vdd.n2600 vdd.n2599 0.0130799
R20072 vdd.n2624 vdd.n2593 0.0130799
R20073 vdd.n2625 vdd.n2624 0.0130799
R20074 vdd.n2620 vdd.n2619 0.0130799
R20075 vdd.n2605 vdd.n2604 0.0130799
R20076 vdd.n2551 vdd.n2540 0.0130799
R20077 vdd.n2551 vdd.n2545 0.0130799
R20078 vdd.n2560 vdd.n2554 0.0130799
R20079 vdd.n2554 vdd.n2553 0.0130799
R20080 vdd.n2578 vdd.n2547 0.0130799
R20081 vdd.n2579 vdd.n2578 0.0130799
R20082 vdd.n2574 vdd.n2573 0.0130799
R20083 vdd.n2559 vdd.n2558 0.0130799
R20084 vdd.n2644 vdd.n2633 0.0130799
R20085 vdd.n2644 vdd.n2638 0.0130799
R20086 vdd.n2653 vdd.n2647 0.0130799
R20087 vdd.n2647 vdd.n2646 0.0130799
R20088 vdd.n2671 vdd.n2640 0.0130799
R20089 vdd.n2672 vdd.n2671 0.0130799
R20090 vdd.n2667 vdd.n2666 0.0130799
R20091 vdd.n2652 vdd.n2651 0.0130799
R20092 vdd.n2692 vdd.n2681 0.0130799
R20093 vdd.n2692 vdd.n2686 0.0130799
R20094 vdd.n2701 vdd.n2695 0.0130799
R20095 vdd.n2695 vdd.n2694 0.0130799
R20096 vdd.n2719 vdd.n2688 0.0130799
R20097 vdd.n2720 vdd.n2719 0.0130799
R20098 vdd.n2715 vdd.n2714 0.0130799
R20099 vdd.n2700 vdd.n2699 0.0130799
R20100 vdd.n2738 vdd.n2727 0.0130799
R20101 vdd.n2738 vdd.n2732 0.0130799
R20102 vdd.n2747 vdd.n2741 0.0130799
R20103 vdd.n2741 vdd.n2740 0.0130799
R20104 vdd.n2765 vdd.n2734 0.0130799
R20105 vdd.n2766 vdd.n2765 0.0130799
R20106 vdd.n2761 vdd.n2760 0.0130799
R20107 vdd.n2746 vdd.n2745 0.0130799
R20108 vdd.n997 vdd.n991 0.0130799
R20109 vdd.n1014 vdd.n997 0.0130799
R20110 vdd.n1002 vdd.n999 0.0130799
R20111 vdd.n1002 vdd.n995 0.0130799
R20112 vdd.n1023 vdd.n1022 0.0130799
R20113 vdd.n1023 vdd.n989 0.0130799
R20114 vdd.n1029 vdd.n986 0.0130799
R20115 vdd.n1001 vdd.n1000 0.0130799
R20116 vdd.n2880 vdd.n2869 0.0130799
R20117 vdd.n2880 vdd.n2874 0.0130799
R20118 vdd.n2889 vdd.n2883 0.0130799
R20119 vdd.n2883 vdd.n2882 0.0130799
R20120 vdd.n2907 vdd.n2876 0.0130799
R20121 vdd.n2908 vdd.n2907 0.0130799
R20122 vdd.n2903 vdd.n2902 0.0130799
R20123 vdd.n2888 vdd.n2887 0.0130799
R20124 vdd.n2833 vdd.n2822 0.0130799
R20125 vdd.n2833 vdd.n2827 0.0130799
R20126 vdd.n2842 vdd.n2836 0.0130799
R20127 vdd.n2836 vdd.n2835 0.0130799
R20128 vdd.n2860 vdd.n2829 0.0130799
R20129 vdd.n2861 vdd.n2860 0.0130799
R20130 vdd.n2856 vdd.n2855 0.0130799
R20131 vdd.n2841 vdd.n2840 0.0130799
R20132 vdd.n2787 vdd.n2776 0.0130799
R20133 vdd.n2787 vdd.n2781 0.0130799
R20134 vdd.n2796 vdd.n2790 0.0130799
R20135 vdd.n2790 vdd.n2789 0.0130799
R20136 vdd.n2814 vdd.n2783 0.0130799
R20137 vdd.n2815 vdd.n2814 0.0130799
R20138 vdd.n2810 vdd.n2809 0.0130799
R20139 vdd.n2795 vdd.n2794 0.0130799
R20140 vdd.n2927 vdd.n2916 0.0130799
R20141 vdd.n2927 vdd.n2921 0.0130799
R20142 vdd.n2936 vdd.n2930 0.0130799
R20143 vdd.n2930 vdd.n2929 0.0130799
R20144 vdd.n2954 vdd.n2923 0.0130799
R20145 vdd.n2955 vdd.n2954 0.0130799
R20146 vdd.n2950 vdd.n2949 0.0130799
R20147 vdd.n2935 vdd.n2934 0.0130799
R20148 vdd.n2975 vdd.n2964 0.0130799
R20149 vdd.n2975 vdd.n2969 0.0130799
R20150 vdd.n2984 vdd.n2978 0.0130799
R20151 vdd.n2978 vdd.n2977 0.0130799
R20152 vdd.n3002 vdd.n2971 0.0130799
R20153 vdd.n3003 vdd.n3002 0.0130799
R20154 vdd.n2998 vdd.n2997 0.0130799
R20155 vdd.n2983 vdd.n2982 0.0130799
R20156 vdd.n3021 vdd.n3010 0.0130799
R20157 vdd.n3021 vdd.n3015 0.0130799
R20158 vdd.n3030 vdd.n3024 0.0130799
R20159 vdd.n3024 vdd.n3023 0.0130799
R20160 vdd.n3048 vdd.n3017 0.0130799
R20161 vdd.n3049 vdd.n3048 0.0130799
R20162 vdd.n3044 vdd.n3043 0.0130799
R20163 vdd.n3029 vdd.n3028 0.0130799
R20164 vdd.n3115 vdd.n3104 0.0130799
R20165 vdd.n3115 vdd.n3109 0.0130799
R20166 vdd.n3124 vdd.n3118 0.0130799
R20167 vdd.n3118 vdd.n3117 0.0130799
R20168 vdd.n3142 vdd.n3111 0.0130799
R20169 vdd.n3143 vdd.n3142 0.0130799
R20170 vdd.n3138 vdd.n3137 0.0130799
R20171 vdd.n3123 vdd.n3122 0.0130799
R20172 vdd.n3069 vdd.n3058 0.0130799
R20173 vdd.n3069 vdd.n3063 0.0130799
R20174 vdd.n3078 vdd.n3072 0.0130799
R20175 vdd.n3072 vdd.n3071 0.0130799
R20176 vdd.n3096 vdd.n3065 0.0130799
R20177 vdd.n3097 vdd.n3096 0.0130799
R20178 vdd.n3092 vdd.n3091 0.0130799
R20179 vdd.n3077 vdd.n3076 0.0130799
R20180 vdd.n3162 vdd.n3151 0.0130799
R20181 vdd.n3162 vdd.n3156 0.0130799
R20182 vdd.n3171 vdd.n3165 0.0130799
R20183 vdd.n3165 vdd.n3164 0.0130799
R20184 vdd.n3189 vdd.n3158 0.0130799
R20185 vdd.n3190 vdd.n3189 0.0130799
R20186 vdd.n3185 vdd.n3184 0.0130799
R20187 vdd.n3170 vdd.n3169 0.0130799
R20188 vdd.n3210 vdd.n3199 0.0130799
R20189 vdd.n3210 vdd.n3204 0.0130799
R20190 vdd.n3219 vdd.n3213 0.0130799
R20191 vdd.n3213 vdd.n3212 0.0130799
R20192 vdd.n3237 vdd.n3206 0.0130799
R20193 vdd.n3238 vdd.n3237 0.0130799
R20194 vdd.n3233 vdd.n3232 0.0130799
R20195 vdd.n3218 vdd.n3217 0.0130799
R20196 vdd.n3256 vdd.n3245 0.0130799
R20197 vdd.n3256 vdd.n3250 0.0130799
R20198 vdd.n3265 vdd.n3259 0.0130799
R20199 vdd.n3259 vdd.n3258 0.0130799
R20200 vdd.n3283 vdd.n3252 0.0130799
R20201 vdd.n3284 vdd.n3283 0.0130799
R20202 vdd.n3279 vdd.n3278 0.0130799
R20203 vdd.n3264 vdd.n3263 0.0130799
R20204 vdd.n761 vdd.n755 0.0130799
R20205 vdd.n778 vdd.n761 0.0130799
R20206 vdd.n766 vdd.n763 0.0130799
R20207 vdd.n766 vdd.n759 0.0130799
R20208 vdd.n787 vdd.n786 0.0130799
R20209 vdd.n787 vdd.n753 0.0130799
R20210 vdd.n793 vdd.n750 0.0130799
R20211 vdd.n765 vdd.n764 0.0130799
R20212 vdd.n3351 vdd.n3340 0.0130799
R20213 vdd.n3351 vdd.n3345 0.0130799
R20214 vdd.n3360 vdd.n3354 0.0130799
R20215 vdd.n3354 vdd.n3353 0.0130799
R20216 vdd.n3378 vdd.n3347 0.0130799
R20217 vdd.n3379 vdd.n3378 0.0130799
R20218 vdd.n3374 vdd.n3373 0.0130799
R20219 vdd.n3359 vdd.n3358 0.0130799
R20220 vdd.n3305 vdd.n3294 0.0130799
R20221 vdd.n3305 vdd.n3299 0.0130799
R20222 vdd.n3314 vdd.n3308 0.0130799
R20223 vdd.n3308 vdd.n3307 0.0130799
R20224 vdd.n3332 vdd.n3301 0.0130799
R20225 vdd.n3333 vdd.n3332 0.0130799
R20226 vdd.n3328 vdd.n3327 0.0130799
R20227 vdd.n3313 vdd.n3312 0.0130799
R20228 vdd.n3398 vdd.n3387 0.0130799
R20229 vdd.n3398 vdd.n3392 0.0130799
R20230 vdd.n3407 vdd.n3401 0.0130799
R20231 vdd.n3401 vdd.n3400 0.0130799
R20232 vdd.n3425 vdd.n3394 0.0130799
R20233 vdd.n3426 vdd.n3425 0.0130799
R20234 vdd.n3421 vdd.n3420 0.0130799
R20235 vdd.n3406 vdd.n3405 0.0130799
R20236 vdd.n3446 vdd.n3435 0.0130799
R20237 vdd.n3446 vdd.n3440 0.0130799
R20238 vdd.n3455 vdd.n3449 0.0130799
R20239 vdd.n3449 vdd.n3448 0.0130799
R20240 vdd.n3473 vdd.n3442 0.0130799
R20241 vdd.n3474 vdd.n3473 0.0130799
R20242 vdd.n3469 vdd.n3468 0.0130799
R20243 vdd.n3454 vdd.n3453 0.0130799
R20244 vdd.n3492 vdd.n3481 0.0130799
R20245 vdd.n3492 vdd.n3486 0.0130799
R20246 vdd.n3501 vdd.n3495 0.0130799
R20247 vdd.n3495 vdd.n3494 0.0130799
R20248 vdd.n3519 vdd.n3488 0.0130799
R20249 vdd.n3520 vdd.n3519 0.0130799
R20250 vdd.n3515 vdd.n3514 0.0130799
R20251 vdd.n3500 vdd.n3499 0.0130799
R20252 vdd.n574 vdd.n563 0.0130799
R20253 vdd.n574 vdd.n568 0.0130799
R20254 vdd.n583 vdd.n577 0.0130799
R20255 vdd.n577 vdd.n576 0.0130799
R20256 vdd.n601 vdd.n570 0.0130799
R20257 vdd.n602 vdd.n601 0.0130799
R20258 vdd.n597 vdd.n596 0.0130799
R20259 vdd.n582 vdd.n581 0.0130799
R20260 vdd.n3587 vdd.n3576 0.0130799
R20261 vdd.n3587 vdd.n3581 0.0130799
R20262 vdd.n3596 vdd.n3590 0.0130799
R20263 vdd.n3590 vdd.n3589 0.0130799
R20264 vdd.n3614 vdd.n3583 0.0130799
R20265 vdd.n3615 vdd.n3614 0.0130799
R20266 vdd.n3610 vdd.n3609 0.0130799
R20267 vdd.n3595 vdd.n3594 0.0130799
R20268 vdd.n3541 vdd.n3530 0.0130799
R20269 vdd.n3541 vdd.n3535 0.0130799
R20270 vdd.n3550 vdd.n3544 0.0130799
R20271 vdd.n3544 vdd.n3543 0.0130799
R20272 vdd.n3568 vdd.n3537 0.0130799
R20273 vdd.n3569 vdd.n3568 0.0130799
R20274 vdd.n3564 vdd.n3563 0.0130799
R20275 vdd.n3549 vdd.n3548 0.0130799
R20276 vdd.n6601 vdd.n6590 0.0130799
R20277 vdd.n6601 vdd.n6595 0.0130799
R20278 vdd.n6610 vdd.n6604 0.0130799
R20279 vdd.n6604 vdd.n6603 0.0130799
R20280 vdd.n6628 vdd.n6597 0.0130799
R20281 vdd.n6629 vdd.n6628 0.0130799
R20282 vdd.n6624 vdd.n6623 0.0130799
R20283 vdd.n6609 vdd.n6608 0.0130799
R20284 vdd.n6555 vdd.n6544 0.0130799
R20285 vdd.n6555 vdd.n6549 0.0130799
R20286 vdd.n6564 vdd.n6558 0.0130799
R20287 vdd.n6558 vdd.n6557 0.0130799
R20288 vdd.n6582 vdd.n6551 0.0130799
R20289 vdd.n6583 vdd.n6582 0.0130799
R20290 vdd.n6578 vdd.n6577 0.0130799
R20291 vdd.n6563 vdd.n6562 0.0130799
R20292 vdd.n9615 vdd.n9604 0.0130799
R20293 vdd.n9615 vdd.n9609 0.0130799
R20294 vdd.n9624 vdd.n9618 0.0130799
R20295 vdd.n9618 vdd.n9617 0.0130799
R20296 vdd.n9642 vdd.n9611 0.0130799
R20297 vdd.n9643 vdd.n9642 0.0130799
R20298 vdd.n9638 vdd.n9637 0.0130799
R20299 vdd.n9623 vdd.n9622 0.0130799
R20300 vdd.n9569 vdd.n9558 0.0130799
R20301 vdd.n9569 vdd.n9563 0.0130799
R20302 vdd.n9578 vdd.n9572 0.0130799
R20303 vdd.n9572 vdd.n9571 0.0130799
R20304 vdd.n9596 vdd.n9565 0.0130799
R20305 vdd.n9597 vdd.n9596 0.0130799
R20306 vdd.n9592 vdd.n9591 0.0130799
R20307 vdd.n9577 vdd.n9576 0.0130799
R20308 vdd.n9661 vdd.n9650 0.0130799
R20309 vdd.n9661 vdd.n9655 0.0130799
R20310 vdd.n9670 vdd.n9664 0.0130799
R20311 vdd.n9664 vdd.n9663 0.0130799
R20312 vdd.n9688 vdd.n9657 0.0130799
R20313 vdd.n9689 vdd.n9688 0.0130799
R20314 vdd.n9684 vdd.n9683 0.0130799
R20315 vdd.n9669 vdd.n9668 0.0130799
R20316 vdd.n9707 vdd.n9696 0.0130799
R20317 vdd.n9707 vdd.n9701 0.0130799
R20318 vdd.n9716 vdd.n9710 0.0130799
R20319 vdd.n9710 vdd.n9709 0.0130799
R20320 vdd.n9734 vdd.n9703 0.0130799
R20321 vdd.n9735 vdd.n9734 0.0130799
R20322 vdd.n9730 vdd.n9729 0.0130799
R20323 vdd.n9715 vdd.n9714 0.0130799
R20324 vdd.n9805 vdd.n9794 0.0130799
R20325 vdd.n9805 vdd.n9799 0.0130799
R20326 vdd.n9814 vdd.n9808 0.0130799
R20327 vdd.n9808 vdd.n9807 0.0130799
R20328 vdd.n9832 vdd.n9801 0.0130799
R20329 vdd.n9833 vdd.n9832 0.0130799
R20330 vdd.n9828 vdd.n9827 0.0130799
R20331 vdd.n9813 vdd.n9812 0.0130799
R20332 vdd.n9851 vdd.n9840 0.0130799
R20333 vdd.n9851 vdd.n9845 0.0130799
R20334 vdd.n9860 vdd.n9854 0.0130799
R20335 vdd.n9854 vdd.n9853 0.0130799
R20336 vdd.n9878 vdd.n9847 0.0130799
R20337 vdd.n9879 vdd.n9878 0.0130799
R20338 vdd.n9874 vdd.n9873 0.0130799
R20339 vdd.n9859 vdd.n9858 0.0130799
R20340 vdd.n9897 vdd.n9886 0.0130799
R20341 vdd.n9897 vdd.n9891 0.0130799
R20342 vdd.n9906 vdd.n9900 0.0130799
R20343 vdd.n9900 vdd.n9899 0.0130799
R20344 vdd.n9924 vdd.n9893 0.0130799
R20345 vdd.n9925 vdd.n9924 0.0130799
R20346 vdd.n9920 vdd.n9919 0.0130799
R20347 vdd.n9905 vdd.n9904 0.0130799
R20348 vdd.n9943 vdd.n9932 0.0130799
R20349 vdd.n9943 vdd.n9937 0.0130799
R20350 vdd.n9952 vdd.n9946 0.0130799
R20351 vdd.n9946 vdd.n9945 0.0130799
R20352 vdd.n9970 vdd.n9939 0.0130799
R20353 vdd.n9971 vdd.n9970 0.0130799
R20354 vdd.n9966 vdd.n9965 0.0130799
R20355 vdd.n9951 vdd.n9950 0.0130799
R20356 vdd.n10041 vdd.n10030 0.0130799
R20357 vdd.n10041 vdd.n10035 0.0130799
R20358 vdd.n10050 vdd.n10044 0.0130799
R20359 vdd.n10044 vdd.n10043 0.0130799
R20360 vdd.n10068 vdd.n10037 0.0130799
R20361 vdd.n10069 vdd.n10068 0.0130799
R20362 vdd.n10064 vdd.n10063 0.0130799
R20363 vdd.n10049 vdd.n10048 0.0130799
R20364 vdd.n57 vdd.n46 0.0130799
R20365 vdd.n57 vdd.n51 0.0130799
R20366 vdd.n66 vdd.n60 0.0130799
R20367 vdd.n60 vdd.n59 0.0130799
R20368 vdd.n84 vdd.n53 0.0130799
R20369 vdd.n85 vdd.n84 0.0130799
R20370 vdd.n80 vdd.n79 0.0130799
R20371 vdd.n65 vdd.n64 0.0130799
R20372 vdd.n11 vdd.n0 0.0130799
R20373 vdd.n11 vdd.n5 0.0130799
R20374 vdd.n20 vdd.n14 0.0130799
R20375 vdd.n14 vdd.n13 0.0130799
R20376 vdd.n38 vdd.n7 0.0130799
R20377 vdd.n39 vdd.n38 0.0130799
R20378 vdd.n34 vdd.n33 0.0130799
R20379 vdd.n19 vdd.n18 0.0130799
R20380 vdd.n10087 vdd.n10076 0.0130799
R20381 vdd.n10087 vdd.n10081 0.0130799
R20382 vdd.n10096 vdd.n10090 0.0130799
R20383 vdd.n10090 vdd.n10089 0.0130799
R20384 vdd.n10114 vdd.n10083 0.0130799
R20385 vdd.n10115 vdd.n10114 0.0130799
R20386 vdd.n10110 vdd.n10109 0.0130799
R20387 vdd.n10095 vdd.n10094 0.0130799
R20388 vdd.n10135 vdd.n10124 0.0130799
R20389 vdd.n10135 vdd.n10129 0.0130799
R20390 vdd.n10144 vdd.n10138 0.0130799
R20391 vdd.n10138 vdd.n10137 0.0130799
R20392 vdd.n10162 vdd.n10131 0.0130799
R20393 vdd.n10163 vdd.n10162 0.0130799
R20394 vdd.n10158 vdd.n10157 0.0130799
R20395 vdd.n10143 vdd.n10142 0.0130799
R20396 vdd.n10181 vdd.n10170 0.0130799
R20397 vdd.n10181 vdd.n10175 0.0130799
R20398 vdd.n10190 vdd.n10184 0.0130799
R20399 vdd.n10184 vdd.n10183 0.0130799
R20400 vdd.n10208 vdd.n10177 0.0130799
R20401 vdd.n10209 vdd.n10208 0.0130799
R20402 vdd.n10204 vdd.n10203 0.0130799
R20403 vdd.n10189 vdd.n10188 0.0130799
R20404 vdd.n9992 vdd.n9986 0.0130799
R20405 vdd.n10009 vdd.n9992 0.0130799
R20406 vdd.n9997 vdd.n9994 0.0130799
R20407 vdd.n9997 vdd.n9990 0.0130799
R20408 vdd.n10018 vdd.n10017 0.0130799
R20409 vdd.n10018 vdd.n9984 0.0130799
R20410 vdd.n10024 vdd.n9981 0.0130799
R20411 vdd.n9996 vdd.n9995 0.0130799
R20412 vdd.n10323 vdd.n10312 0.0130799
R20413 vdd.n10323 vdd.n10317 0.0130799
R20414 vdd.n10332 vdd.n10326 0.0130799
R20415 vdd.n10326 vdd.n10325 0.0130799
R20416 vdd.n10350 vdd.n10319 0.0130799
R20417 vdd.n10351 vdd.n10350 0.0130799
R20418 vdd.n10346 vdd.n10345 0.0130799
R20419 vdd.n10331 vdd.n10330 0.0130799
R20420 vdd.n10276 vdd.n10265 0.0130799
R20421 vdd.n10276 vdd.n10270 0.0130799
R20422 vdd.n10285 vdd.n10279 0.0130799
R20423 vdd.n10279 vdd.n10278 0.0130799
R20424 vdd.n10303 vdd.n10272 0.0130799
R20425 vdd.n10304 vdd.n10303 0.0130799
R20426 vdd.n10299 vdd.n10298 0.0130799
R20427 vdd.n10284 vdd.n10283 0.0130799
R20428 vdd.n10230 vdd.n10219 0.0130799
R20429 vdd.n10230 vdd.n10224 0.0130799
R20430 vdd.n10239 vdd.n10233 0.0130799
R20431 vdd.n10233 vdd.n10232 0.0130799
R20432 vdd.n10257 vdd.n10226 0.0130799
R20433 vdd.n10258 vdd.n10257 0.0130799
R20434 vdd.n10253 vdd.n10252 0.0130799
R20435 vdd.n10238 vdd.n10237 0.0130799
R20436 vdd.n10370 vdd.n10359 0.0130799
R20437 vdd.n10370 vdd.n10364 0.0130799
R20438 vdd.n10379 vdd.n10373 0.0130799
R20439 vdd.n10373 vdd.n10372 0.0130799
R20440 vdd.n10397 vdd.n10366 0.0130799
R20441 vdd.n10398 vdd.n10397 0.0130799
R20442 vdd.n10393 vdd.n10392 0.0130799
R20443 vdd.n10378 vdd.n10377 0.0130799
R20444 vdd.n10418 vdd.n10407 0.0130799
R20445 vdd.n10418 vdd.n10412 0.0130799
R20446 vdd.n10427 vdd.n10421 0.0130799
R20447 vdd.n10421 vdd.n10420 0.0130799
R20448 vdd.n10445 vdd.n10414 0.0130799
R20449 vdd.n10446 vdd.n10445 0.0130799
R20450 vdd.n10441 vdd.n10440 0.0130799
R20451 vdd.n10426 vdd.n10425 0.0130799
R20452 vdd.n10464 vdd.n10453 0.0130799
R20453 vdd.n10464 vdd.n10458 0.0130799
R20454 vdd.n10473 vdd.n10467 0.0130799
R20455 vdd.n10467 vdd.n10466 0.0130799
R20456 vdd.n10491 vdd.n10460 0.0130799
R20457 vdd.n10492 vdd.n10491 0.0130799
R20458 vdd.n10487 vdd.n10486 0.0130799
R20459 vdd.n10472 vdd.n10471 0.0130799
R20460 vdd.n10558 vdd.n10547 0.0130799
R20461 vdd.n10558 vdd.n10552 0.0130799
R20462 vdd.n10567 vdd.n10561 0.0130799
R20463 vdd.n10561 vdd.n10560 0.0130799
R20464 vdd.n10585 vdd.n10554 0.0130799
R20465 vdd.n10586 vdd.n10585 0.0130799
R20466 vdd.n10581 vdd.n10580 0.0130799
R20467 vdd.n10566 vdd.n10565 0.0130799
R20468 vdd.n10512 vdd.n10501 0.0130799
R20469 vdd.n10512 vdd.n10506 0.0130799
R20470 vdd.n10521 vdd.n10515 0.0130799
R20471 vdd.n10515 vdd.n10514 0.0130799
R20472 vdd.n10539 vdd.n10508 0.0130799
R20473 vdd.n10540 vdd.n10539 0.0130799
R20474 vdd.n10535 vdd.n10534 0.0130799
R20475 vdd.n10520 vdd.n10519 0.0130799
R20476 vdd.n10605 vdd.n10594 0.0130799
R20477 vdd.n10605 vdd.n10599 0.0130799
R20478 vdd.n10614 vdd.n10608 0.0130799
R20479 vdd.n10608 vdd.n10607 0.0130799
R20480 vdd.n10632 vdd.n10601 0.0130799
R20481 vdd.n10633 vdd.n10632 0.0130799
R20482 vdd.n10628 vdd.n10627 0.0130799
R20483 vdd.n10613 vdd.n10612 0.0130799
R20484 vdd.n10653 vdd.n10642 0.0130799
R20485 vdd.n10653 vdd.n10647 0.0130799
R20486 vdd.n10662 vdd.n10656 0.0130799
R20487 vdd.n10656 vdd.n10655 0.0130799
R20488 vdd.n10680 vdd.n10649 0.0130799
R20489 vdd.n10681 vdd.n10680 0.0130799
R20490 vdd.n10676 vdd.n10675 0.0130799
R20491 vdd.n10661 vdd.n10660 0.0130799
R20492 vdd.n10699 vdd.n10688 0.0130799
R20493 vdd.n10699 vdd.n10693 0.0130799
R20494 vdd.n10708 vdd.n10702 0.0130799
R20495 vdd.n10702 vdd.n10701 0.0130799
R20496 vdd.n10726 vdd.n10695 0.0130799
R20497 vdd.n10727 vdd.n10726 0.0130799
R20498 vdd.n10722 vdd.n10721 0.0130799
R20499 vdd.n10707 vdd.n10706 0.0130799
R20500 vdd.n9756 vdd.n9750 0.0130799
R20501 vdd.n9773 vdd.n9756 0.0130799
R20502 vdd.n9761 vdd.n9758 0.0130799
R20503 vdd.n9761 vdd.n9754 0.0130799
R20504 vdd.n9782 vdd.n9781 0.0130799
R20505 vdd.n9782 vdd.n9748 0.0130799
R20506 vdd.n9788 vdd.n9745 0.0130799
R20507 vdd.n9760 vdd.n9759 0.0130799
R20508 vdd.n10794 vdd.n10783 0.0130799
R20509 vdd.n10794 vdd.n10788 0.0130799
R20510 vdd.n10803 vdd.n10797 0.0130799
R20511 vdd.n10797 vdd.n10796 0.0130799
R20512 vdd.n10821 vdd.n10790 0.0130799
R20513 vdd.n10822 vdd.n10821 0.0130799
R20514 vdd.n10817 vdd.n10816 0.0130799
R20515 vdd.n10802 vdd.n10801 0.0130799
R20516 vdd.n10748 vdd.n10737 0.0130799
R20517 vdd.n10748 vdd.n10742 0.0130799
R20518 vdd.n10757 vdd.n10751 0.0130799
R20519 vdd.n10751 vdd.n10750 0.0130799
R20520 vdd.n10775 vdd.n10744 0.0130799
R20521 vdd.n10776 vdd.n10775 0.0130799
R20522 vdd.n10771 vdd.n10770 0.0130799
R20523 vdd.n10756 vdd.n10755 0.0130799
R20524 vdd.n10841 vdd.n10830 0.0130799
R20525 vdd.n10841 vdd.n10835 0.0130799
R20526 vdd.n10850 vdd.n10844 0.0130799
R20527 vdd.n10844 vdd.n10843 0.0130799
R20528 vdd.n10868 vdd.n10837 0.0130799
R20529 vdd.n10869 vdd.n10868 0.0130799
R20530 vdd.n10864 vdd.n10863 0.0130799
R20531 vdd.n10849 vdd.n10848 0.0130799
R20532 vdd.n10889 vdd.n10878 0.0130799
R20533 vdd.n10889 vdd.n10883 0.0130799
R20534 vdd.n10898 vdd.n10892 0.0130799
R20535 vdd.n10892 vdd.n10891 0.0130799
R20536 vdd.n10916 vdd.n10885 0.0130799
R20537 vdd.n10917 vdd.n10916 0.0130799
R20538 vdd.n10912 vdd.n10911 0.0130799
R20539 vdd.n10897 vdd.n10896 0.0130799
R20540 vdd.n10935 vdd.n10924 0.0130799
R20541 vdd.n10935 vdd.n10929 0.0130799
R20542 vdd.n10944 vdd.n10938 0.0130799
R20543 vdd.n10938 vdd.n10937 0.0130799
R20544 vdd.n10962 vdd.n10931 0.0130799
R20545 vdd.n10963 vdd.n10962 0.0130799
R20546 vdd.n10958 vdd.n10957 0.0130799
R20547 vdd.n10943 vdd.n10942 0.0130799
R20548 vdd.n10984 vdd.n10973 0.0130799
R20549 vdd.n10985 vdd.n10984 0.0130799
R20550 vdd.n11001 vdd.n10977 0.0130799
R20551 vdd.n11006 vdd.n10977 0.0130799
R20552 vdd.n10992 vdd.n10986 0.0130799
R20553 vdd.n10986 vdd.n10983 0.0130799
R20554 vdd.n10991 vdd.n10987 0.0130799
R20555 vdd.n11009 vdd.n11008 0.0130799
R20556 vdd.n11029 vdd.n11018 0.0130799
R20557 vdd.n11030 vdd.n11029 0.0130799
R20558 vdd.n11046 vdd.n11022 0.0130799
R20559 vdd.n11051 vdd.n11022 0.0130799
R20560 vdd.n11037 vdd.n11031 0.0130799
R20561 vdd.n11031 vdd.n11028 0.0130799
R20562 vdd.n11036 vdd.n11032 0.0130799
R20563 vdd.n11054 vdd.n11053 0.0130799
R20564 vdd.n11079 vdd.n11068 0.0130799
R20565 vdd.n11080 vdd.n11079 0.0130799
R20566 vdd.n11096 vdd.n11072 0.0130799
R20567 vdd.n11101 vdd.n11072 0.0130799
R20568 vdd.n11087 vdd.n11081 0.0130799
R20569 vdd.n11081 vdd.n11078 0.0130799
R20570 vdd.n11086 vdd.n11082 0.0130799
R20571 vdd.n11104 vdd.n11103 0.0130799
R20572 vdd.n11125 vdd.n11114 0.0130799
R20573 vdd.n11126 vdd.n11125 0.0130799
R20574 vdd.n11142 vdd.n11118 0.0130799
R20575 vdd.n11147 vdd.n11118 0.0130799
R20576 vdd.n11133 vdd.n11127 0.0130799
R20577 vdd.n11127 vdd.n11124 0.0130799
R20578 vdd.n11132 vdd.n11128 0.0130799
R20579 vdd.n11150 vdd.n11149 0.0130799
R20580 vdd.n11173 vdd.n11162 0.0130799
R20581 vdd.n11174 vdd.n11173 0.0130799
R20582 vdd.n11190 vdd.n11166 0.0130799
R20583 vdd.n11195 vdd.n11166 0.0130799
R20584 vdd.n11181 vdd.n11175 0.0130799
R20585 vdd.n11175 vdd.n11172 0.0130799
R20586 vdd.n11180 vdd.n11176 0.0130799
R20587 vdd.n11198 vdd.n11197 0.0130799
R20588 vdd.n435 vdd.n428 0.0130799
R20589 vdd.n435 vdd.n434 0.0130799
R20590 vdd.n446 vdd.n431 0.0130799
R20591 vdd.n451 vdd.n431 0.0130799
R20592 vdd.n437 vdd.n425 0.0130799
R20593 vdd.n426 vdd.n425 0.0130799
R20594 vdd.n424 vdd.n422 0.0130799
R20595 vdd.n454 vdd.n453 0.0130799
R20596 vdd.n11220 vdd.n11209 0.0130799
R20597 vdd.n11221 vdd.n11220 0.0130799
R20598 vdd.n11237 vdd.n11213 0.0130799
R20599 vdd.n11242 vdd.n11213 0.0130799
R20600 vdd.n11228 vdd.n11222 0.0130799
R20601 vdd.n11222 vdd.n11219 0.0130799
R20602 vdd.n11227 vdd.n11223 0.0130799
R20603 vdd.n11245 vdd.n11244 0.0130799
R20604 vdd.n11265 vdd.n11254 0.0130799
R20605 vdd.n11266 vdd.n11265 0.0130799
R20606 vdd.n11282 vdd.n11258 0.0130799
R20607 vdd.n11287 vdd.n11258 0.0130799
R20608 vdd.n11273 vdd.n11267 0.0130799
R20609 vdd.n11267 vdd.n11264 0.0130799
R20610 vdd.n11272 vdd.n11268 0.0130799
R20611 vdd.n11290 vdd.n11289 0.0130799
R20612 vdd.n11311 vdd.n11300 0.0130799
R20613 vdd.n11312 vdd.n11311 0.0130799
R20614 vdd.n11328 vdd.n11304 0.0130799
R20615 vdd.n11333 vdd.n11304 0.0130799
R20616 vdd.n11319 vdd.n11313 0.0130799
R20617 vdd.n11313 vdd.n11310 0.0130799
R20618 vdd.n11318 vdd.n11314 0.0130799
R20619 vdd.n11336 vdd.n11335 0.0130799
R20620 vdd.n11362 vdd.n11351 0.0130799
R20621 vdd.n11363 vdd.n11362 0.0130799
R20622 vdd.n11379 vdd.n11355 0.0130799
R20623 vdd.n11384 vdd.n11355 0.0130799
R20624 vdd.n11370 vdd.n11364 0.0130799
R20625 vdd.n11364 vdd.n11361 0.0130799
R20626 vdd.n11369 vdd.n11365 0.0130799
R20627 vdd.n11387 vdd.n11386 0.0130799
R20628 vdd.n11408 vdd.n11397 0.0130799
R20629 vdd.n11409 vdd.n11408 0.0130799
R20630 vdd.n11425 vdd.n11401 0.0130799
R20631 vdd.n11430 vdd.n11401 0.0130799
R20632 vdd.n11416 vdd.n11410 0.0130799
R20633 vdd.n11410 vdd.n11407 0.0130799
R20634 vdd.n11415 vdd.n11411 0.0130799
R20635 vdd.n11433 vdd.n11432 0.0130799
R20636 vdd.n11456 vdd.n11445 0.0130799
R20637 vdd.n11457 vdd.n11456 0.0130799
R20638 vdd.n11473 vdd.n11449 0.0130799
R20639 vdd.n11478 vdd.n11449 0.0130799
R20640 vdd.n11464 vdd.n11458 0.0130799
R20641 vdd.n11458 vdd.n11455 0.0130799
R20642 vdd.n11463 vdd.n11459 0.0130799
R20643 vdd.n11481 vdd.n11480 0.0130799
R20644 vdd.n11502 vdd.n11491 0.0130799
R20645 vdd.n11503 vdd.n11502 0.0130799
R20646 vdd.n11519 vdd.n11495 0.0130799
R20647 vdd.n11524 vdd.n11495 0.0130799
R20648 vdd.n11510 vdd.n11504 0.0130799
R20649 vdd.n11504 vdd.n11501 0.0130799
R20650 vdd.n11509 vdd.n11505 0.0130799
R20651 vdd.n11527 vdd.n11526 0.0130799
R20652 vdd.n11547 vdd.n11536 0.0130799
R20653 vdd.n11548 vdd.n11547 0.0130799
R20654 vdd.n11564 vdd.n11540 0.0130799
R20655 vdd.n11569 vdd.n11540 0.0130799
R20656 vdd.n11555 vdd.n11549 0.0130799
R20657 vdd.n11549 vdd.n11546 0.0130799
R20658 vdd.n11554 vdd.n11550 0.0130799
R20659 vdd.n11572 vdd.n11571 0.0130799
R20660 vdd.n11597 vdd.n11586 0.0130799
R20661 vdd.n11598 vdd.n11597 0.0130799
R20662 vdd.n11614 vdd.n11590 0.0130799
R20663 vdd.n11619 vdd.n11590 0.0130799
R20664 vdd.n11605 vdd.n11599 0.0130799
R20665 vdd.n11599 vdd.n11596 0.0130799
R20666 vdd.n11604 vdd.n11600 0.0130799
R20667 vdd.n11622 vdd.n11621 0.0130799
R20668 vdd.n11643 vdd.n11632 0.0130799
R20669 vdd.n11644 vdd.n11643 0.0130799
R20670 vdd.n11660 vdd.n11636 0.0130799
R20671 vdd.n11665 vdd.n11636 0.0130799
R20672 vdd.n11651 vdd.n11645 0.0130799
R20673 vdd.n11645 vdd.n11642 0.0130799
R20674 vdd.n11650 vdd.n11646 0.0130799
R20675 vdd.n11668 vdd.n11667 0.0130799
R20676 vdd.n11691 vdd.n11680 0.0130799
R20677 vdd.n11692 vdd.n11691 0.0130799
R20678 vdd.n11708 vdd.n11684 0.0130799
R20679 vdd.n11713 vdd.n11684 0.0130799
R20680 vdd.n11699 vdd.n11693 0.0130799
R20681 vdd.n11693 vdd.n11690 0.0130799
R20682 vdd.n11698 vdd.n11694 0.0130799
R20683 vdd.n11716 vdd.n11715 0.0130799
R20684 vdd.n200 vdd.n193 0.0130799
R20685 vdd.n200 vdd.n199 0.0130799
R20686 vdd.n211 vdd.n196 0.0130799
R20687 vdd.n216 vdd.n196 0.0130799
R20688 vdd.n202 vdd.n190 0.0130799
R20689 vdd.n191 vdd.n190 0.0130799
R20690 vdd.n189 vdd.n187 0.0130799
R20691 vdd.n219 vdd.n218 0.0130799
R20692 vdd.n11738 vdd.n11727 0.0130799
R20693 vdd.n11739 vdd.n11738 0.0130799
R20694 vdd.n11755 vdd.n11731 0.0130799
R20695 vdd.n11760 vdd.n11731 0.0130799
R20696 vdd.n11746 vdd.n11740 0.0130799
R20697 vdd.n11740 vdd.n11737 0.0130799
R20698 vdd.n11745 vdd.n11741 0.0130799
R20699 vdd.n11763 vdd.n11762 0.0130799
R20700 vdd.n11783 vdd.n11772 0.0130799
R20701 vdd.n11784 vdd.n11783 0.0130799
R20702 vdd.n11800 vdd.n11776 0.0130799
R20703 vdd.n11805 vdd.n11776 0.0130799
R20704 vdd.n11791 vdd.n11785 0.0130799
R20705 vdd.n11785 vdd.n11782 0.0130799
R20706 vdd.n11790 vdd.n11786 0.0130799
R20707 vdd.n11808 vdd.n11807 0.0130799
R20708 vdd.n11833 vdd.n11822 0.0130799
R20709 vdd.n11834 vdd.n11833 0.0130799
R20710 vdd.n11850 vdd.n11826 0.0130799
R20711 vdd.n11855 vdd.n11826 0.0130799
R20712 vdd.n11841 vdd.n11835 0.0130799
R20713 vdd.n11835 vdd.n11832 0.0130799
R20714 vdd.n11840 vdd.n11836 0.0130799
R20715 vdd.n11858 vdd.n11857 0.0130799
R20716 vdd.n11879 vdd.n11868 0.0130799
R20717 vdd.n11880 vdd.n11879 0.0130799
R20718 vdd.n11896 vdd.n11872 0.0130799
R20719 vdd.n11901 vdd.n11872 0.0130799
R20720 vdd.n11887 vdd.n11881 0.0130799
R20721 vdd.n11881 vdd.n11878 0.0130799
R20722 vdd.n11886 vdd.n11882 0.0130799
R20723 vdd.n11904 vdd.n11903 0.0130799
R20724 vdd.n11927 vdd.n11916 0.0130799
R20725 vdd.n11928 vdd.n11927 0.0130799
R20726 vdd.n11944 vdd.n11920 0.0130799
R20727 vdd.n11949 vdd.n11920 0.0130799
R20728 vdd.n11935 vdd.n11929 0.0130799
R20729 vdd.n11929 vdd.n11926 0.0130799
R20730 vdd.n11934 vdd.n11930 0.0130799
R20731 vdd.n11952 vdd.n11951 0.0130799
R20732 vdd.n7484 vdd.n7437 0.0103684
R20733 vdd.n7249 vdd.n7202 0.0103684
R20734 vdd.n7059 vdd.n7012 0.0103684
R20735 vdd.n6823 vdd.n6776 0.0103684
R20736 vdd.n4470 vdd.n4423 0.0103684
R20737 vdd.n4235 vdd.n4188 0.0103684
R20738 vdd.n4045 vdd.n3998 0.0103684
R20739 vdd.n3809 vdd.n3762 0.0103684
R20740 vdd.n1456 vdd.n1409 0.0103684
R20741 vdd.n1221 vdd.n1174 0.0103684
R20742 vdd.n1031 vdd.n984 0.0103684
R20743 vdd.n795 vdd.n748 0.0103684
R20744 vdd.n10026 vdd.n9979 0.0103684
R20745 vdd.n9790 vdd.n9743 0.0103684
R20746 vdd.n468 vdd.n421 0.0103684
R20747 vdd.n233 vdd.n186 0.0103684
R20748 vdd.n110 vdd.t1047 0.00463816
R20749 vdd.n156 vdd.t7 0.00463816
R20750 vdd.n253 vdd.t1475 0.00463816
R20751 vdd.n299 vdd.t562 0.00463816
R20752 vdd.n345 vdd.t1298 0.00463816
R20753 vdd.n391 vdd.t1485 0.00463816
R20754 vdd.n488 vdd.t209 0.00463816
R20755 vdd.n534 vdd.t375 0.00463816
R20756 vdd.n7126 vdd.t1463 0.00463816
R20757 vdd.n7172 vdd.t1310 0.00463816
R20758 vdd.n7269 vdd.t1049 0.00463816
R20759 vdd.n7315 vdd.t1360 0.00463816
R20760 vdd.n7361 vdd.t593 0.00463816
R20761 vdd.n7407 vdd.t379 0.00463816
R20762 vdd.n7504 vdd.t1326 0.00463816
R20763 vdd.n6653 vdd.t484 0.00463816
R20764 vdd.n7548 vdd.t898 0.00463816
R20765 vdd.n7593 vdd.t166 0.00463816
R20766 vdd.n7643 vdd.t589 0.00463816
R20767 vdd.n7689 vdd.t862 0.00463816
R20768 vdd.n7737 vdd.t1342 0.00463816
R20769 vdd.n7455 vdd.t1154 0.00463816
R20770 vdd.n7784 vdd.t896 0.00463816
R20771 vdd.n7829 vdd.t837 0.00463816
R20772 vdd.n7875 vdd.t1375 0.00463816
R20773 vdd.n7926 vdd.t486 0.00463816
R20774 vdd.n7972 vdd.t872 0.00463816
R20775 vdd.n8020 vdd.t1330 0.00463816
R20776 vdd.n8066 vdd.t36 0.00463816
R20777 vdd.n8111 vdd.t835 0.00463816
R20778 vdd.n8161 vdd.t201 0.00463816
R20779 vdd.n8207 vdd.t973 0.00463816
R20780 vdd.n8255 vdd.t1346 0.00463816
R20781 vdd.n7220 vdd.t1459 0.00463816
R20782 vdd.n8302 vdd.t854 0.00463816
R20783 vdd.n8347 vdd.t56 0.00463816
R20784 vdd.n8397 vdd.t9 0.00463816
R20785 vdd.n8443 vdd.t40 0.00463816
R20786 vdd.n8491 vdd.t211 0.00463816
R20787 vdd.n4112 vdd.t203 0.00463816
R20788 vdd.n4158 vdd.t554 0.00463816
R20789 vdd.n4255 vdd.t1290 0.00463816
R20790 vdd.n4301 vdd.t1316 0.00463816
R20791 vdd.n4347 vdd.t1055 0.00463816
R20792 vdd.n4393 vdd.t570 0.00463816
R20793 vdd.n4490 vdd.t1045 0.00463816
R20794 vdd.n3639 vdd.t560 0.00463816
R20795 vdd.n4534 vdd.t1000 0.00463816
R20796 vdd.n4579 vdd.t174 0.00463816
R20797 vdd.n4629 vdd.t197 0.00463816
R20798 vdd.n4675 vdd.t34 0.00463816
R20799 vdd.n4723 vdd.t1473 0.00463816
R20800 vdd.n4441 vdd.t1457 0.00463816
R20801 vdd.n4770 vdd.t827 0.00463816
R20802 vdd.n4815 vdd.t52 0.00463816
R20803 vdd.n4861 vdd.t1371 0.00463816
R20804 vdd.n4912 vdd.t1487 0.00463816
R20805 vdd.n4958 vdd.t858 0.00463816
R20806 vdd.n5006 vdd.t1300 0.00463816
R20807 vdd.n5052 vdd.t1010 0.00463816
R20808 vdd.n5097 vdd.t50 0.00463816
R20809 vdd.n5147 vdd.t1043 0.00463816
R20810 vdd.n5193 vdd.t942 0.00463816
R20811 vdd.n5241 vdd.t1304 0.00463816
R20812 vdd.n4206 vdd.t1455 0.00463816
R20813 vdd.n5288 vdd.t844 0.00463816
R20814 vdd.n5333 vdd.t172 0.00463816
R20815 vdd.n5383 vdd.t456 0.00463816
R20816 vdd.n5429 vdd.t1012 0.00463816
R20817 vdd.n5477 vdd.t1051 0.00463816
R20818 vdd.n1098 vdd.t3 0.00463816
R20819 vdd.n1144 vdd.t195 0.00463816
R20820 vdd.n1241 vdd.t1308 0.00463816
R20821 vdd.n1287 vdd.t1495 0.00463816
R20822 vdd.n1333 vdd.t1356 0.00463816
R20823 vdd.n1379 vdd.t591 0.00463816
R20824 vdd.n1476 vdd.t385 0.00463816
R20825 vdd.n625 vdd.t552 0.00463816
R20826 vdd.n1520 vdd.t823 0.00463816
R20827 vdd.n1565 vdd.t833 0.00463816
R20828 vdd.n1615 vdd.t466 0.00463816
R20829 vdd.n1661 vdd.t998 0.00463816
R20830 vdd.n1709 vdd.t1493 0.00463816
R20831 vdd.n1427 vdd.t101 0.00463816
R20832 vdd.n1756 vdd.t870 0.00463816
R20833 vdd.n1801 vdd.t170 0.00463816
R20834 vdd.n1847 vdd.t1127 0.00463816
R20835 vdd.n1898 vdd.t1324 0.00463816
R20836 vdd.n1944 vdd.t992 0.00463816
R20837 vdd.n1992 vdd.t371 0.00463816
R20838 vdd.n2038 vdd.t971 0.00463816
R20839 vdd.n2083 vdd.t168 0.00463816
R20840 vdd.n2133 vdd.t1344 0.00463816
R20841 vdd.n2179 vdd.t940 0.00463816
R20842 vdd.n2227 vdd.t1481 0.00463816
R20843 vdd.n1192 vdd.t95 0.00463816
R20844 vdd.n2274 vdd.t900 0.00463816
R20845 vdd.n2319 vdd.t771 0.00463816
R20846 vdd.n2369 vdd.t492 0.00463816
R20847 vdd.n2415 vdd.t975 0.00463816
R20848 vdd.n2463 vdd.t1348 0.00463816
R20849 vdd.n10988 vdd.t821 0.00463816
R20850 vdd.n11033 vdd.t58 0.00463816
R20851 vdd.n11083 vdd.t1499 0.00463816
R20852 vdd.n11129 vdd.t996 0.00463816
R20853 vdd.n11177 vdd.t1294 0.00463816
R20854 vdd.n439 vdd.t579 0.00463816
R20855 vdd.n11224 vdd.t965 0.00463816
R20856 vdd.n11269 vdd.t796 0.00463816
R20857 vdd.n11315 vdd.t1377 0.00463816
R20858 vdd.n11366 vdd.t199 0.00463816
R20859 vdd.n11412 vdd.t850 0.00463816
R20860 vdd.n11460 vdd.t1340 0.00463816
R20861 vdd.n11506 vdd.t811 0.00463816
R20862 vdd.n11551 vdd.t794 0.00463816
R20863 vdd.n11601 vdd.t1286 0.00463816
R20864 vdd.n11647 vdd.t994 0.00463816
R20865 vdd.n11695 vdd.t1338 0.00463816
R20866 vdd.n204 vdd.t577 0.00463816
R20867 vdd.n11742 vdd.t1014 0.00463816
R20868 vdd.n11787 vdd.t792 0.00463816
R20869 vdd.n11837 vdd.t1320 0.00463816
R20870 vdd.n11883 vdd.t813 0.00463816
R20871 vdd.n11931 vdd.t1292 0.00463816
R20872 vdd.t1471 vdd.n11991 0.00442942
R20873 vdd.n11972 vdd.t829 0.00442942
R20874 vdd.t1182 vdd.n100 0.00442942
R20875 vdd.t977 vdd.n146 0.00442942
R20876 vdd.t527 vdd.n243 0.00442942
R20877 vdd.t1238 vdd.n289 0.00442942
R20878 vdd.t156 vdd.n335 0.00442942
R20879 vdd.t959 vdd.n381 0.00442942
R20880 vdd.t336 vdd.n478 0.00442942
R20881 vdd.t122 vdd.n524 0.00442942
R20882 vdd.n6691 vdd.t1288 0.00442942
R20883 vdd.t728 vdd.n6698 0.00442942
R20884 vdd.n6737 vdd.t207 0.00442942
R20885 vdd.t235 vdd.n6744 0.00442942
R20886 vdd.n6835 vdd.t1318 0.00442942
R20887 vdd.t155 vdd.n6842 0.00442942
R20888 vdd.n6881 vdd.t205 0.00442942
R20889 vdd.t413 vdd.n6888 0.00442942
R20890 vdd.n6927 vdd.t558 0.00442942
R20891 vdd.t983 vdd.n6934 0.00442942
R20892 vdd.n6973 vdd.t377 0.00442942
R20893 vdd.t1107 vdd.n6980 0.00442942
R20894 vdd.n7071 vdd.t587 0.00442942
R20895 vdd.t353 vdd.n7078 0.00442942
R20896 vdd.n8529 vdd.t482 0.00442942
R20897 vdd.t634 vdd.n8536 0.00442942
R20898 vdd.t1025 vdd.n7116 0.00442942
R20899 vdd.t979 vdd.n7162 0.00442942
R20900 vdd.t1285 vdd.n7259 0.00442942
R20901 vdd.t536 vdd.n7305 0.00442942
R20902 vdd.t1094 vdd.n7351 0.00442942
R20903 vdd.t1255 vdd.n7397 0.00442942
R20904 vdd.t143 vdd.n7494 0.00442942
R20905 vdd.t1088 vdd.n6643 0.00442942
R20906 vdd.t1263 vdd.n7538 0.00442942
R20907 vdd.t809 vdd.n7583 0.00442942
R20908 vdd.t1226 vdd.n7633 0.00442942
R20909 vdd.t874 vdd.n7679 0.00442942
R20910 vdd.t1078 vdd.n7727 0.00442942
R20911 vdd.t892 vdd.n7448 0.00442942
R20912 vdd.t1506 vdd.n7774 0.00442942
R20913 vdd.t241 vdd.n7819 0.00442942
R20914 vdd.t543 vdd.n7865 0.00442942
R20915 vdd.t306 vdd.n7916 0.00442942
R20916 vdd.t620 vdd.n7962 0.00442942
R20917 vdd.t978 vdd.n8010 0.00442942
R20918 vdd.t22 vdd.n8056 0.00442942
R20919 vdd.t335 vdd.n8101 0.00442942
R20920 vdd.t70 vdd.n8151 0.00442942
R20921 vdd.t1442 vdd.n8197 0.00442942
R20922 vdd.t743 vdd.n8245 0.00442942
R20923 vdd.t277 vdd.n7213 0.00442942
R20924 vdd.t1112 vdd.n8292 0.00442942
R20925 vdd.t343 vdd.n8337 0.00442942
R20926 vdd.t881 vdd.n8387 0.00442942
R20927 vdd.t1149 vdd.n8433 0.00442942
R20928 vdd.t1066 vdd.n8481 0.00442942
R20929 vdd.n8622 vdd.t848 0.00442942
R20930 vdd.t284 vdd.n8629 0.00442942
R20931 vdd.n8576 vdd.t773 0.00442942
R20932 vdd.t412 vdd.n8583 0.00442942
R20933 vdd.n8669 vdd.t1314 0.00442942
R20934 vdd.t1143 vdd.n8676 0.00442942
R20935 vdd.n8717 vdd.t856 0.00442942
R20936 vdd.t658 vdd.n8724 0.00442942
R20937 vdd.n8763 vdd.t1467 0.00442942
R20938 vdd.t1507 vdd.n8770 0.00442942
R20939 vdd.n7054 vdd.t97 0.00442942
R20940 vdd.t1089 vdd.n7034 0.00442942
R20941 vdd.n8905 vdd.t825 0.00442942
R20942 vdd.t66 vdd.n8912 0.00442942
R20943 vdd.n8858 vdd.t765 0.00442942
R20944 vdd.t1195 vdd.n8865 0.00442942
R20945 vdd.n8812 vdd.t1129 0.00442942
R20946 vdd.t264 vdd.n8819 0.00442942
R20947 vdd.n8952 vdd.t458 0.00442942
R20948 vdd.t758 vdd.n8959 0.00442942
R20949 vdd.n9000 vdd.t864 0.00442942
R20950 vdd.t1062 vdd.n9007 0.00442942
R20951 vdd.n9046 vdd.t1477 0.00442942
R20952 vdd.t1108 vdd.n9053 0.00442942
R20953 vdd.n9140 vdd.t1006 0.00442942
R20954 vdd.t64 vdd.n9147 0.00442942
R20955 vdd.n9094 vdd.t430 0.00442942
R20956 vdd.t1024 vdd.n9101 0.00442942
R20957 vdd.n9187 vdd.t566 0.00442942
R20958 vdd.t1270 vdd.n9194 0.00442942
R20959 vdd.n9235 vdd.t42 0.00442942
R20960 vdd.t675 vdd.n9242 0.00442942
R20961 vdd.n9281 vdd.t1302 0.00442942
R20962 vdd.t547 vdd.n9288 0.00442942
R20963 vdd.n6818 vdd.t89 0.00442942
R20964 vdd.t1362 vdd.n6798 0.00442942
R20965 vdd.n9376 vdd.t988 0.00442942
R20966 vdd.t523 vdd.n9383 0.00442942
R20967 vdd.n9330 vdd.t627 0.00442942
R20968 vdd.t1031 vdd.n9337 0.00442942
R20969 vdd.n9423 vdd.t601 0.00442942
R20970 vdd.t428 vdd.n9430 0.00442942
R20971 vdd.n9471 vdd.t860 0.00442942
R20972 vdd.t1191 vdd.n9478 0.00442942
R20973 vdd.n9517 vdd.t1041 0.00442942
R20974 vdd.t76 vdd.n9524 0.00442942
R20975 vdd.n3677 vdd.t1483 0.00442942
R20976 vdd.t441 vdd.n3684 0.00442942
R20977 vdd.n3723 vdd.t464 0.00442942
R20978 vdd.t234 vdd.n3730 0.00442942
R20979 vdd.n3821 vdd.t599 0.00442942
R20980 vdd.t503 vdd.n3828 0.00442942
R20981 vdd.n3867 vdd.t460 0.00442942
R20982 vdd.t136 vdd.n3874 0.00442942
R20983 vdd.n3913 vdd.t1057 0.00442942
R20984 vdd.t611 vdd.n3920 0.00442942
R20985 vdd.n3959 vdd.t603 0.00442942
R20986 vdd.t802 vdd.n3966 0.00442942
R20987 vdd.n4057 vdd.t468 0.00442942
R20988 vdd.t473 vdd.n4064 0.00442942
R20989 vdd.n5515 vdd.t556 0.00442942
R20990 vdd.t327 vdd.n5522 0.00442942
R20991 vdd.t440 vdd.n4102 0.00442942
R20992 vdd.t477 vdd.n4148 0.00442942
R20993 vdd.t114 vdd.n4245 0.00442942
R20994 vdd.t810 vdd.n4291 0.00442942
R20995 vdd.t1427 vdd.n4337 0.00442942
R20996 vdd.t1225 vdd.n4383 0.00442942
R20997 vdd.t951 vdd.n4480 0.00442942
R20998 vdd.t230 vdd.n3629 0.00442942
R20999 vdd.t1148 vdd.n4524 0.00442942
R21000 vdd.t145 vdd.n4569 0.00442942
R21001 vdd.t1178 vdd.n4619 0.00442942
R21002 vdd.t670 vdd.n4665 0.00442942
R21003 vdd.t1032 vdd.n4713 0.00442942
R21004 vdd.t455 vdd.n4434 0.00442942
R21005 vdd.t72 vdd.n4760 0.00442942
R21006 vdd.t1256 vdd.n4805 0.00442942
R21007 vdd.t411 vdd.n4851 0.00442942
R21008 vdd.t1090 vdd.n4902 0.00442942
R21009 vdd.t1165 vdd.n4948 0.00442942
R21010 vdd.t308 vdd.n4996 0.00442942
R21011 vdd.t1412 vdd.n5042 0.00442942
R21012 vdd.t607 vdd.n5087 0.00442942
R21013 vdd.t191 vdd.n5137 0.00442942
R21014 vdd.t1278 vdd.n5183 0.00442942
R21015 vdd.t537 vdd.n5231 0.00442942
R21016 vdd.t1067 vdd.n4199 0.00442942
R21017 vdd.t888 vdd.n5278 0.00442942
R21018 vdd.t660 vdd.n5323 0.00442942
R21019 vdd.t63 vdd.n5373 0.00442942
R21020 vdd.t1411 vdd.n5419 0.00442942
R21021 vdd.t269 vdd.n5467 0.00442942
R21022 vdd.n5608 vdd.t906 0.00442942
R21023 vdd.t716 vdd.n5615 0.00442942
R21024 vdd.n5562 vdd.t164 0.00442942
R21025 vdd.t1237 vdd.n5569 0.00442942
R21026 vdd.n5655 vdd.t595 0.00442942
R21027 vdd.t144 vdd.n5662 0.00442942
R21028 vdd.n5703 vdd.t990 0.00442942
R21029 vdd.t924 vdd.n5710 0.00442942
R21030 vdd.n5749 vdd.t13 0.00442942
R21031 vdd.t424 vdd.n5756 0.00442942
R21032 vdd.n4040 vdd.t99 0.00442942
R21033 vdd.t1422 vdd.n4020 0.00442942
R21034 vdd.n5891 vdd.t866 0.00442942
R21035 vdd.t23 vdd.n5898 0.00442942
R21036 vdd.n5844 vdd.t767 0.00442942
R21037 vdd.t786 vdd.n5851 0.00442942
R21038 vdd.n5798 vdd.t1373 0.00442942
R21039 vdd.t928 vdd.n5805 0.00442942
R21040 vdd.n5938 vdd.t1479 0.00442942
R21041 vdd.t679 vdd.n5945 0.00442942
R21042 vdd.n5986 vdd.t1002 0.00442942
R21043 vdd.t1258 vdd.n5993 0.00442942
R21044 vdd.n6032 vdd.t1489 0.00442942
R21045 vdd.t429 vdd.n6039 0.00442942
R21046 vdd.n6126 vdd.t969 0.00442942
R21047 vdd.t305 vdd.n6133 0.00442942
R21048 vdd.n6080 vdd.t434 0.00442942
R21049 vdd.t671 vdd.n6087 0.00442942
R21050 vdd.n6173 vdd.t1336 0.00442942
R21051 vdd.t387 vdd.n6180 0.00442942
R21052 vdd.n6221 vdd.t32 0.00442942
R21053 vdd.t246 vdd.n6228 0.00442942
R21054 vdd.n6267 vdd.t496 0.00442942
R21055 vdd.t1026 vdd.n6274 0.00442942
R21056 vdd.n3804 vdd.t93 0.00442942
R21057 vdd.t724 vdd.n3784 0.00442942
R21058 vdd.n6362 vdd.t868 0.00442942
R21059 vdd.t20 vdd.n6369 0.00442942
R21060 vdd.n6316 vdd.t432 0.00442942
R21061 vdd.t331 vdd.n6323 0.00442942
R21062 vdd.n6409 vdd.t1053 0.00442942
R21063 vdd.t615 vdd.n6416 0.00442942
R21064 vdd.n6457 vdd.t894 0.00442942
R21065 vdd.t1367 vdd.n6464 0.00442942
R21066 vdd.n6503 vdd.t564 0.00442942
R21067 vdd.t314 vdd.n6510 0.00442942
R21068 vdd.n663 vdd.t1465 0.00442942
R21069 vdd.t695 vdd.n670 0.00442942
R21070 vdd.n709 vdd.t1501 0.00442942
R21071 vdd.t1406 vdd.n716 0.00442942
R21072 vdd.n807 vdd.t1358 0.00442942
R21073 vdd.t1202 vdd.n814 0.00442942
R21074 vdd.n853 vdd.t1497 0.00442942
R21075 vdd.t1383 vdd.n860 0.00442942
R21076 vdd.n899 vdd.t1312 0.00442942
R21077 vdd.t361 vdd.n906 0.00442942
R21078 vdd.n945 vdd.t462 0.00442942
R21079 vdd.t236 vdd.n952 0.00442942
R21080 vdd.n1043 vdd.t1469 0.00442942
R21081 vdd.t1259 vdd.n1050 0.00442942
R21082 vdd.n2501 vdd.t381 0.00442942
R21083 vdd.t1213 vdd.n2508 0.00442942
R21084 vdd.t947 vdd.n1088 0.00442942
R21085 vdd.t747 vdd.n1134 0.00442942
R21086 vdd.t86 vdd.n1231 0.00442942
R21087 vdd.t157 vdd.n1277 0.00442942
R21088 vdd.t65 vdd.n1323 0.00442942
R21089 vdd.t920 vdd.n1369 0.00442942
R21090 vdd.t1447 vdd.n1466 0.00442942
R21091 vdd.t893 vdd.n615 0.00442942
R21092 vdd.t1142 vdd.n1510 0.00442942
R21093 vdd.t1121 vdd.n1555 0.00442942
R21094 vdd.t1033 vdd.n1605 0.00442942
R21095 vdd.t309 vdd.n1651 0.00442942
R21096 vdd.t1018 vdd.n1699 0.00442942
R21097 vdd.t1443 vdd.n1420 0.00442942
R21098 vdd.t683 vdd.n1746 0.00442942
R21099 vdd.t132 vdd.n1791 0.00442942
R21100 vdd.t657 vdd.n1837 0.00442942
R21101 vdd.t1283 vdd.n1888 0.00442942
R21102 vdd.t391 vdd.n1934 0.00442942
R21103 vdd.t268 vdd.n1982 0.00442942
R21104 vdd.t1220 vdd.n2028 0.00442942
R21105 vdd.t226 vdd.n2073 0.00442942
R21106 vdd.t110 vdd.n2123 0.00442942
R21107 vdd.t1131 vdd.n2169 0.00442942
R21108 vdd.t1119 vdd.n2217 0.00442942
R21109 vdd.t1163 vdd.n1185 0.00442942
R21110 vdd.t929 vdd.n2264 0.00442942
R21111 vdd.t516 vdd.n2309 0.00442942
R21112 vdd.t103 vdd.n2359 0.00442942
R21113 vdd.t606 vdd.n2405 0.00442942
R21114 vdd.t1423 vdd.n2453 0.00442942
R21115 vdd.n2594 vdd.t815 0.00442942
R21116 vdd.t423 vdd.n2601 0.00442942
R21117 vdd.n2548 vdd.t769 0.00442942
R21118 vdd.t1027 vdd.n2555 0.00442942
R21119 vdd.n2641 vdd.t1350 0.00442942
R21120 vdd.t916 vdd.n2648 0.00442942
R21121 vdd.n2689 vdd.t1016 0.00442942
R21122 vdd.t717 vdd.n2696 0.00442942
R21123 vdd.n2735 vdd.t494 0.00442942
R21124 vdd.t392 vdd.n2742 0.00442942
R21125 vdd.n1026 vdd.t91 0.00442942
R21126 vdd.t1230 vdd.n1006 0.00442942
R21127 vdd.n2877 vdd.t44 0.00442942
R21128 vdd.t445 vdd.n2884 0.00442942
R21129 vdd.n2830 vdd.t438 0.00442942
R21130 vdd.t1106 vdd.n2837 0.00442942
R21131 vdd.n2784 vdd.t1125 0.00442942
R21132 vdd.t729 vdd.n2791 0.00442942
R21133 vdd.n2924 vdd.t11 0.00442942
R21134 vdd.t605 vdd.n2931 0.00442942
R21135 vdd.n2972 vdd.t38 0.00442942
R21136 vdd.t1221 vdd.n2979 0.00442942
R21137 vdd.n3018 vdd.t1296 0.00442942
R21138 vdd.t1434 vdd.n3025 0.00442942
R21139 vdd.n3112 vdd.t852 0.00442942
R21140 vdd.t1156 vdd.n3119 0.00442942
R21141 vdd.n3066 vdd.t790 0.00442942
R21142 vdd.t21 vdd.n3073 0.00442942
R21143 vdd.n3159 vdd.t373 0.00442942
R21144 vdd.t245 vdd.n3166 0.00442942
R21145 vdd.n3207 vdd.t967 0.00442942
R21146 vdd.t1282 vdd.n3214 0.00442942
R21147 vdd.n3253 vdd.t1328 0.00442942
R21148 vdd.t798 vdd.n3260 0.00442942
R21149 vdd.n790 vdd.t87 0.00442942
R21150 vdd.t1410 vdd.n770 0.00442942
R21151 vdd.n3348 vdd.t819 0.00442942
R21152 vdd.t1203 vdd.n3355 0.00442942
R21153 vdd.n3302 vdd.t436 0.00442942
R21154 vdd.t310 vdd.n3309 0.00442942
R21155 vdd.n3395 vdd.t1332 0.00442942
R21156 vdd.t1124 vdd.n3402 0.00442942
R21157 vdd.n3443 vdd.t904 0.00442942
R21158 vdd.t1061 vdd.n3450 0.00442942
R21159 vdd.n3489 vdd.t488 0.00442942
R21160 vdd.t1123 vdd.n3496 0.00442942
R21161 vdd.n571 vdd.t30 0.00442942
R21162 vdd.t748 vdd.n578 0.00442942
R21163 vdd.n3584 vdd.t24 0.00442942
R21164 vdd.t1382 vdd.n3591 0.00442942
R21165 vdd.n3538 vdd.t986 0.00442942
R21166 vdd.t1150 vdd.n3545 0.00442942
R21167 vdd.n6598 vdd.t28 0.00442942
R21168 vdd.t1095 vdd.n6605 0.00442942
R21169 vdd.n6552 vdd.t1186 0.00442942
R21170 vdd.t1243 vdd.n6559 0.00442942
R21171 vdd.n9612 vdd.t26 0.00442942
R21172 vdd.t706 vdd.n9619 0.00442942
R21173 vdd.n9566 vdd.t984 0.00442942
R21174 vdd.t237 vdd.n9573 0.00442942
R21175 vdd.n9658 vdd.t1354 0.00442942
R21176 vdd.t1514 vdd.n9665 0.00442942
R21177 vdd.n9704 vdd.t1322 0.00442942
R21178 vdd.t71 vdd.n9711 0.00442942
R21179 vdd.n9802 vdd.t478 0.00442942
R21180 vdd.t360 vdd.n9809 0.00442942
R21181 vdd.n9848 vdd.t1059 0.00442942
R21182 vdd.t1284 vdd.n9855 0.00442942
R21183 vdd.n9894 vdd.t15 0.00442942
R21184 vdd.t1023 vdd.n9901 0.00442942
R21185 vdd.n9940 vdd.t490 0.00442942
R21186 vdd.t960 vdd.n9947 0.00442942
R21187 vdd.n10038 vdd.t1334 0.00442942
R21188 vdd.t548 vdd.n10045 0.00442942
R21189 vdd.n54 vdd.t1008 0.00442942
R21190 vdd.t422 vdd.n61 0.00442942
R21191 vdd.n8 vdd.t839 0.00442942
R21192 vdd.t260 vdd.n15 0.00442942
R21193 vdd.n10084 vdd.t568 0.00442942
R21194 vdd.t1164 vdd.n10091 0.00442942
R21195 vdd.n10132 vdd.t908 0.00442942
R21196 vdd.t1438 vdd.n10139 0.00442942
R21197 vdd.n10178 vdd.t597 0.00442942
R21198 vdd.t418 vdd.n10185 0.00442942
R21199 vdd.n10021 vdd.t575 0.00442942
R21200 vdd.t694 vdd.n10001 0.00442942
R21201 vdd.n10320 vdd.t938 0.00442942
R21202 vdd.t702 vdd.n10327 0.00442942
R21203 vdd.n10273 vdd.t54 0.00442942
R21204 vdd.t502 vdd.n10280 0.00442942
R21205 vdd.n10227 vdd.t1379 0.00442942
R21206 vdd.t659 vdd.n10234 0.00442942
R21207 vdd.n10367 vdd.t383 0.00442942
R21208 vdd.t1138 vdd.n10374 0.00442942
R21209 vdd.n10415 vdd.t846 0.00442942
R21210 vdd.t1454 vdd.n10422 0.00442942
R21211 vdd.n10461 vdd.t1306 0.00442942
R21212 vdd.t1257 vdd.n10468 0.00442942
R21213 vdd.n10555 vdd.t1004 0.00442942
R21214 vdd.t1366 vdd.n10562 0.00442942
R21215 vdd.n10509 vdd.t775 0.00442942
R21216 vdd.t1102 vdd.n10516 0.00442942
R21217 vdd.n10602 vdd.t1491 0.00442942
R21218 vdd.t1019 vdd.n10609 0.00442942
R21219 vdd.n10650 vdd.t817 0.00442942
R21220 vdd.t253 vdd.n10657 0.00442942
R21221 vdd.n10696 vdd.t1352 0.00442942
R21222 vdd.t292 vdd.n10703 0.00442942
R21223 vdd.n9785 vdd.t1461 0.00442942
R21224 vdd.t964 vdd.n9765 0.00442942
R21225 vdd.n10791 vdd.t902 0.00442942
R21226 vdd.t742 vdd.n10798 0.00442942
R21227 vdd.n10745 vdd.t629 0.00442942
R21228 vdd.t1247 vdd.n10752 0.00442942
R21229 vdd.n10838 vdd.t480 0.00442942
R21230 vdd.t417 vdd.n10845 0.00442942
R21231 vdd.n10886 vdd.t936 0.00442942
R21232 vdd.t285 vdd.n10893 0.00442942
R21233 vdd.n10932 vdd.t5 0.00442942
R21234 vdd.t690 vdd.n10939 0.00442942
R21235 vdd.t498 vdd.n10978 0.00442942
R21236 vdd.t1251 vdd.n11023 0.00442942
R21237 vdd.t538 vdd.n11073 0.00442942
R21238 vdd.t539 vdd.n11119 0.00442942
R21239 vdd.t216 vdd.n11167 0.00442942
R21240 vdd.t1122 vdd.n432 0.00442942
R21241 vdd.t115 vdd.n11214 0.00442942
R21242 vdd.t531 vdd.n11259 0.00442942
R21243 vdd.t1037 vdd.n11305 0.00442942
R21244 vdd.t1147 vdd.n11356 0.00442942
R21245 vdd.t958 vdd.n11402 0.00442942
R21246 vdd.t1242 vdd.n11450 0.00442942
R21247 vdd.t273 vdd.n11496 0.00442942
R21248 vdd.t307 vdd.n11541 0.00442942
R21249 vdd.t535 vdd.n11591 0.00442942
R21250 vdd.t641 vdd.n11637 0.00442942
R21251 vdd.t1120 vdd.n11685 0.00442942
R21252 vdd.t1381 vdd.n197 0.00442942
R21253 vdd.t49 vdd.n11732 0.00442942
R21254 vdd.t1396 vdd.n11777 0.00442942
R21255 vdd.t1271 vdd.n11827 0.00442942
R21256 vdd.t619 vdd.n11873 0.00442942
R21257 vdd.t1071 vdd.n11921 0.00442942
R21258 vdd.n7047 vdd.n7046 0.00100279
R21259 vdd.n6811 vdd.n6810 0.00100279
R21260 vdd.n4033 vdd.n4032 0.00100279
R21261 vdd.n3797 vdd.n3796 0.00100279
R21262 vdd.n1019 vdd.n1018 0.00100279
R21263 vdd.n783 vdd.n782 0.00100279
R21264 vdd.n10014 vdd.n10013 0.00100279
R21265 vdd.n9778 vdd.n9777 0.00100279
R21266 vdd.n7477 vdd.n7476 0.00100279
R21267 vdd.n7242 vdd.n7241 0.00100279
R21268 vdd.n4463 vdd.n4462 0.00100279
R21269 vdd.n4228 vdd.n4227 0.00100279
R21270 vdd.n1449 vdd.n1448 0.00100279
R21271 vdd.n1214 vdd.n1213 0.00100279
R21272 vdd.n461 vdd.n460 0.00100279
R21273 vdd.n226 vdd.n225 0.00100279
R21274 vdd.n7486 vdd.n7485 0.00100001
R21275 vdd.n7251 vdd.n7250 0.00100001
R21276 vdd.n7062 vdd.n7061 0.00100001
R21277 vdd.n6826 vdd.n6825 0.00100001
R21278 vdd.n4472 vdd.n4471 0.00100001
R21279 vdd.n4237 vdd.n4236 0.00100001
R21280 vdd.n4048 vdd.n4047 0.00100001
R21281 vdd.n3812 vdd.n3811 0.00100001
R21282 vdd.n1458 vdd.n1457 0.00100001
R21283 vdd.n1223 vdd.n1222 0.00100001
R21284 vdd.n1034 vdd.n1033 0.00100001
R21285 vdd.n798 vdd.n797 0.00100001
R21286 vdd.n10029 vdd.n10028 0.00100001
R21287 vdd.n9793 vdd.n9792 0.00100001
R21288 vdd.n470 vdd.n469 0.00100001
R21289 vdd.n235 vdd.n234 0.00100001
R21290 vdd.n6681 vdd.n6680 0.000501408
R21291 vdd.n7621 vdd.n7620 0.000501408
R21292 vdd.n7622 vdd.n7575 0.000501408
R21293 vdd.n7671 vdd.n7670 0.000501408
R21294 vdd.n7532 vdd.n7531 0.000501408
R21295 vdd.n7765 vdd.n7764 0.000501408
R21296 vdd.n7435 vdd.n7434 0.000501408
R21297 vdd.n7903 vdd.n7902 0.000501408
R21298 vdd.n7857 vdd.n7856 0.000501408
R21299 vdd.n7905 vdd.n7811 0.000501408
R21300 vdd.n7954 vdd.n7953 0.000501408
R21301 vdd.n7389 vdd.n7388 0.000501408
R21302 vdd.n8048 vdd.n8047 0.000501408
R21303 vdd.n7343 vdd.n7342 0.000501408
R21304 vdd.n8139 vdd.n8138 0.000501408
R21305 vdd.n8140 vdd.n8093 0.000501408
R21306 vdd.n8189 vdd.n8188 0.000501408
R21307 vdd.n7297 vdd.n7296 0.000501408
R21308 vdd.n8283 vdd.n8282 0.000501408
R21309 vdd.n7200 vdd.n7199 0.000501408
R21310 vdd.n8375 vdd.n8374 0.000501408
R21311 vdd.n8376 vdd.n8329 0.000501408
R21312 vdd.n8425 vdd.n8424 0.000501408
R21313 vdd.n7154 vdd.n7153 0.000501408
R21314 vdd.n8519 vdd.n8518 0.000501408
R21315 vdd.n8566 vdd.n8563 0.000501408
R21316 vdd.n8613 vdd.n8610 0.000501408
R21317 vdd.n8657 vdd.n8656 0.000501408
R21318 vdd.n8706 vdd.n8703 0.000501408
R21319 vdd.n7108 vdd.n7105 0.000501408
R21320 vdd.n8800 vdd.n8797 0.000501408
R21321 vdd.n7010 vdd.n7007 0.000501408
R21322 vdd.n8849 vdd.n8846 0.000501408
R21323 vdd.n8895 vdd.n8892 0.000501408
R21324 vdd.n8940 vdd.n8939 0.000501408
R21325 vdd.n8989 vdd.n8986 0.000501408
R21326 vdd.n6964 vdd.n6961 0.000501408
R21327 vdd.n9083 vdd.n9080 0.000501408
R21328 vdd.n6918 vdd.n6915 0.000501408
R21329 vdd.n9131 vdd.n9128 0.000501408
R21330 vdd.n9175 vdd.n9174 0.000501408
R21331 vdd.n9224 vdd.n9221 0.000501408
R21332 vdd.n6872 vdd.n6869 0.000501408
R21333 vdd.n9318 vdd.n9315 0.000501408
R21334 vdd.n6774 vdd.n6771 0.000501408
R21335 vdd.n9367 vdd.n9364 0.000501408
R21336 vdd.n9411 vdd.n9410 0.000501408
R21337 vdd.n9460 vdd.n9457 0.000501408
R21338 vdd.n6728 vdd.n6725 0.000501408
R21339 vdd.n9554 vdd.n9551 0.000501408
R21340 vdd.n3667 vdd.n3666 0.000501408
R21341 vdd.n4607 vdd.n4606 0.000501408
R21342 vdd.n4608 vdd.n4561 0.000501408
R21343 vdd.n4657 vdd.n4656 0.000501408
R21344 vdd.n4518 vdd.n4517 0.000501408
R21345 vdd.n4751 vdd.n4750 0.000501408
R21346 vdd.n4421 vdd.n4420 0.000501408
R21347 vdd.n4889 vdd.n4888 0.000501408
R21348 vdd.n4843 vdd.n4842 0.000501408
R21349 vdd.n4891 vdd.n4797 0.000501408
R21350 vdd.n4940 vdd.n4939 0.000501408
R21351 vdd.n4375 vdd.n4374 0.000501408
R21352 vdd.n5034 vdd.n5033 0.000501408
R21353 vdd.n4329 vdd.n4328 0.000501408
R21354 vdd.n5125 vdd.n5124 0.000501408
R21355 vdd.n5126 vdd.n5079 0.000501408
R21356 vdd.n5175 vdd.n5174 0.000501408
R21357 vdd.n4283 vdd.n4282 0.000501408
R21358 vdd.n5269 vdd.n5268 0.000501408
R21359 vdd.n4186 vdd.n4185 0.000501408
R21360 vdd.n5361 vdd.n5360 0.000501408
R21361 vdd.n5362 vdd.n5315 0.000501408
R21362 vdd.n5411 vdd.n5410 0.000501408
R21363 vdd.n4140 vdd.n4139 0.000501408
R21364 vdd.n5505 vdd.n5504 0.000501408
R21365 vdd.n5552 vdd.n5549 0.000501408
R21366 vdd.n5599 vdd.n5596 0.000501408
R21367 vdd.n5643 vdd.n5642 0.000501408
R21368 vdd.n5692 vdd.n5689 0.000501408
R21369 vdd.n4094 vdd.n4091 0.000501408
R21370 vdd.n5786 vdd.n5783 0.000501408
R21371 vdd.n3996 vdd.n3993 0.000501408
R21372 vdd.n5835 vdd.n5832 0.000501408
R21373 vdd.n5881 vdd.n5878 0.000501408
R21374 vdd.n5926 vdd.n5925 0.000501408
R21375 vdd.n5975 vdd.n5972 0.000501408
R21376 vdd.n3950 vdd.n3947 0.000501408
R21377 vdd.n6069 vdd.n6066 0.000501408
R21378 vdd.n3904 vdd.n3901 0.000501408
R21379 vdd.n6117 vdd.n6114 0.000501408
R21380 vdd.n6161 vdd.n6160 0.000501408
R21381 vdd.n6210 vdd.n6207 0.000501408
R21382 vdd.n3858 vdd.n3855 0.000501408
R21383 vdd.n6304 vdd.n6301 0.000501408
R21384 vdd.n3760 vdd.n3757 0.000501408
R21385 vdd.n6353 vdd.n6350 0.000501408
R21386 vdd.n6397 vdd.n6396 0.000501408
R21387 vdd.n6446 vdd.n6443 0.000501408
R21388 vdd.n3714 vdd.n3711 0.000501408
R21389 vdd.n6540 vdd.n6537 0.000501408
R21390 vdd.n653 vdd.n652 0.000501408
R21391 vdd.n1593 vdd.n1592 0.000501408
R21392 vdd.n1594 vdd.n1547 0.000501408
R21393 vdd.n1643 vdd.n1642 0.000501408
R21394 vdd.n1504 vdd.n1503 0.000501408
R21395 vdd.n1737 vdd.n1736 0.000501408
R21396 vdd.n1407 vdd.n1406 0.000501408
R21397 vdd.n1875 vdd.n1874 0.000501408
R21398 vdd.n1829 vdd.n1828 0.000501408
R21399 vdd.n1877 vdd.n1783 0.000501408
R21400 vdd.n1926 vdd.n1925 0.000501408
R21401 vdd.n1361 vdd.n1360 0.000501408
R21402 vdd.n2020 vdd.n2019 0.000501408
R21403 vdd.n1315 vdd.n1314 0.000501408
R21404 vdd.n2111 vdd.n2110 0.000501408
R21405 vdd.n2112 vdd.n2065 0.000501408
R21406 vdd.n2161 vdd.n2160 0.000501408
R21407 vdd.n1269 vdd.n1268 0.000501408
R21408 vdd.n2255 vdd.n2254 0.000501408
R21409 vdd.n1172 vdd.n1171 0.000501408
R21410 vdd.n2347 vdd.n2346 0.000501408
R21411 vdd.n2348 vdd.n2301 0.000501408
R21412 vdd.n2397 vdd.n2396 0.000501408
R21413 vdd.n1126 vdd.n1125 0.000501408
R21414 vdd.n2491 vdd.n2490 0.000501408
R21415 vdd.n2538 vdd.n2535 0.000501408
R21416 vdd.n2585 vdd.n2582 0.000501408
R21417 vdd.n2629 vdd.n2628 0.000501408
R21418 vdd.n2678 vdd.n2675 0.000501408
R21419 vdd.n1080 vdd.n1077 0.000501408
R21420 vdd.n2772 vdd.n2769 0.000501408
R21421 vdd.n982 vdd.n979 0.000501408
R21422 vdd.n2821 vdd.n2818 0.000501408
R21423 vdd.n2867 vdd.n2864 0.000501408
R21424 vdd.n2912 vdd.n2911 0.000501408
R21425 vdd.n2961 vdd.n2958 0.000501408
R21426 vdd.n936 vdd.n933 0.000501408
R21427 vdd.n3055 vdd.n3052 0.000501408
R21428 vdd.n890 vdd.n887 0.000501408
R21429 vdd.n3103 vdd.n3100 0.000501408
R21430 vdd.n3147 vdd.n3146 0.000501408
R21431 vdd.n3196 vdd.n3193 0.000501408
R21432 vdd.n844 vdd.n841 0.000501408
R21433 vdd.n3290 vdd.n3287 0.000501408
R21434 vdd.n746 vdd.n743 0.000501408
R21435 vdd.n3339 vdd.n3336 0.000501408
R21436 vdd.n3383 vdd.n3382 0.000501408
R21437 vdd.n3432 vdd.n3429 0.000501408
R21438 vdd.n700 vdd.n697 0.000501408
R21439 vdd.n3526 vdd.n3523 0.000501408
R21440 vdd.n9601 vdd.n9600 0.000501408
R21441 vdd.n9647 vdd.n9646 0.000501408
R21442 vdd.n6587 vdd.n6586 0.000501408
R21443 vdd.n6633 vdd.n6632 0.000501408
R21444 vdd.n3573 vdd.n3572 0.000501408
R21445 vdd.n3619 vdd.n3618 0.000501408
R21446 vdd.n45 vdd.n42 0.000501408
R21447 vdd.n89 vdd.n88 0.000501408
R21448 vdd.n10121 vdd.n10118 0.000501408
R21449 vdd.n10075 vdd.n10072 0.000501408
R21450 vdd.n10215 vdd.n10212 0.000501408
R21451 vdd.n9977 vdd.n9974 0.000501408
R21452 vdd.n10264 vdd.n10261 0.000501408
R21453 vdd.n10310 vdd.n10307 0.000501408
R21454 vdd.n10355 vdd.n10354 0.000501408
R21455 vdd.n10404 vdd.n10401 0.000501408
R21456 vdd.n9931 vdd.n9928 0.000501408
R21457 vdd.n10498 vdd.n10495 0.000501408
R21458 vdd.n9885 vdd.n9882 0.000501408
R21459 vdd.n10546 vdd.n10543 0.000501408
R21460 vdd.n10590 vdd.n10589 0.000501408
R21461 vdd.n10639 vdd.n10636 0.000501408
R21462 vdd.n9839 vdd.n9836 0.000501408
R21463 vdd.n10733 vdd.n10730 0.000501408
R21464 vdd.n9741 vdd.n9738 0.000501408
R21465 vdd.n10782 vdd.n10779 0.000501408
R21466 vdd.n10826 vdd.n10825 0.000501408
R21467 vdd.n10875 vdd.n10872 0.000501408
R21468 vdd.n9695 vdd.n9692 0.000501408
R21469 vdd.n10969 vdd.n10966 0.000501408
R21470 vdd.n562 vdd.n561 0.000501408
R21471 vdd.n11061 vdd.n11060 0.000501408
R21472 vdd.n11062 vdd.n11015 0.000501408
R21473 vdd.n11111 vdd.n11110 0.000501408
R21474 vdd.n516 vdd.n515 0.000501408
R21475 vdd.n11205 vdd.n11204 0.000501408
R21476 vdd.n419 vdd.n418 0.000501408
R21477 vdd.n11343 vdd.n11342 0.000501408
R21478 vdd.n11297 vdd.n11296 0.000501408
R21479 vdd.n11345 vdd.n11251 0.000501408
R21480 vdd.n11394 vdd.n11393 0.000501408
R21481 vdd.n373 vdd.n372 0.000501408
R21482 vdd.n11488 vdd.n11487 0.000501408
R21483 vdd.n327 vdd.n326 0.000501408
R21484 vdd.n11579 vdd.n11578 0.000501408
R21485 vdd.n11580 vdd.n11533 0.000501408
R21486 vdd.n11629 vdd.n11628 0.000501408
R21487 vdd.n281 vdd.n280 0.000501408
R21488 vdd.n11723 vdd.n11722 0.000501408
R21489 vdd.n184 vdd.n183 0.000501408
R21490 vdd.n11815 vdd.n11814 0.000501408
R21491 vdd.n11816 vdd.n11769 0.000501408
R21492 vdd.n11865 vdd.n11864 0.000501408
R21493 vdd.n138 vdd.n137 0.000501408
R21494 vdd.n11959 vdd.n11958 0.000501408
R21495 vdd.n12007 vdd.n12004 0.000501408
R21496 vss.n6064 vss.n5973 25903.6
R21497 vss.n13077 vss.n2119 24224
R21498 vss.n9670 vss.n5972 21784
R21499 vss.n13921 vss.n13920 18761
R21500 vss.n8510 vss.n6555 18761
R21501 vss.n5363 vss.n3611 18761
R21502 vss.n12100 vss.n12099 18761
R21503 vss.n13921 vss.n18 18099.8
R21504 vss.n7324 vss.n6555 18099.8
R21505 vss.n3611 vss.n2767 18099.8
R21506 vss.n12099 vss.n2145 18099.8
R21507 vss.n14221 vss.n14176 16848
R21508 vss.n9898 vss.n9897 16848
R21509 vss.n14731 vss.n14730 15248
R21510 vss.n14684 vss.n193 15248
R21511 vss.n14536 vss.n14535 15248
R21512 vss.n14489 vss.n252 15248
R21513 vss.n14341 vss.n14340 15248
R21514 vss.n14294 vss.n311 15248
R21515 vss.n14222 vss.n14221 15248
R21516 vss.n9953 vss.n9952 15248
R21517 vss.n9950 vss.n9949 15248
R21518 vss.n9947 vss.n9946 15248
R21519 vss.n9944 vss.n9943 15248
R21520 vss.n9941 vss.n9940 15248
R21521 vss.n9938 vss.n9937 15248
R21522 vss.n9935 vss.n9934 15248
R21523 vss.n9818 vss.n9817 15248
R21524 vss.n9815 vss.n9814 15248
R21525 vss.n9812 vss.n9811 15248
R21526 vss.n9809 vss.n9808 15248
R21527 vss.n9806 vss.n9805 15248
R21528 vss.n9803 vss.n2739 15248
R21529 vss.n9899 vss.n9898 15248
R21530 vss.n9385 vss.n9384 15248
R21531 vss.n9388 vss.n9387 15248
R21532 vss.n9391 vss.n9390 15248
R21533 vss.n9394 vss.n9393 15248
R21534 vss.n9397 vss.n9396 15248
R21535 vss.n9491 vss.n9399 15248
R21536 vss.n9489 vss.n9488 15248
R21537 vss.n8949 vss.n8948 15248
R21538 vss.n8902 vss.n7539 15248
R21539 vss.n8830 vss.n8829 15248
R21540 vss.n8783 vss.n7682 15248
R21541 vss.n8711 vss.n7298 15248
R21542 vss.n9007 vss.n7299 15248
R21543 vss.n13264 vss.n13263 15248
R21544 vss.n13261 vss.n13260 15248
R21545 vss.n13258 vss.n13257 15248
R21546 vss.n13255 vss.n13254 15248
R21547 vss.n13252 vss.n13251 15248
R21548 vss.n13942 vss.n611 15248
R21549 vss.n13940 vss.n13939 15248
R21550 vss.n12993 vss.n12992 15248
R21551 vss.n12990 vss.n12989 15248
R21552 vss.n12987 vss.n12986 15248
R21553 vss.n12984 vss.n12983 15248
R21554 vss.n12981 vss.n12980 15248
R21555 vss.n12978 vss.n12977 15248
R21556 vss.n12975 vss.n2119 15248
R21557 vss.n13136 vss.n13135 15248
R21558 vss.n13133 vss.n13132 15248
R21559 vss.n13130 vss.n13129 15248
R21560 vss.n13127 vss.n13126 15248
R21561 vss.n13124 vss.n13123 15248
R21562 vss.n13121 vss.n13120 15248
R21563 vss.n13118 vss.n13117 15248
R21564 vss.n191 vss.n190 14872
R21565 vss.n14730 vss.n14685 14872
R21566 vss.n250 vss.n193 14872
R21567 vss.n14535 vss.n14490 14872
R21568 vss.n309 vss.n252 14872
R21569 vss.n14340 vss.n14295 14872
R21570 vss.n432 vss.n311 14872
R21571 vss.n9951 vss.n9950 14872
R21572 vss.n9948 vss.n9947 14872
R21573 vss.n9945 vss.n9944 14872
R21574 vss.n9942 vss.n9941 14872
R21575 vss.n9939 vss.n9938 14872
R21576 vss.n9936 vss.n9935 14872
R21577 vss.n2935 vss.n2934 14872
R21578 vss.n9817 vss.n9816 14872
R21579 vss.n9814 vss.n9813 14872
R21580 vss.n9811 vss.n9810 14872
R21581 vss.n9808 vss.n9807 14872
R21582 vss.n9805 vss.n9804 14872
R21583 vss.n9900 vss.n2739 14872
R21584 vss.n9387 vss.n9386 14872
R21585 vss.n9390 vss.n9389 14872
R21586 vss.n9393 vss.n9392 14872
R21587 vss.n9396 vss.n9395 14872
R21588 vss.n9399 vss.n9398 14872
R21589 vss.n9490 vss.n9489 14872
R21590 vss.n9487 vss.n5972 14872
R21591 vss.n7537 vss.n7536 14872
R21592 vss.n8948 vss.n8903 14872
R21593 vss.n7680 vss.n7539 14872
R21594 vss.n8829 vss.n8784 14872
R21595 vss.n8710 vss.n7682 14872
R21596 vss.n9008 vss.n7298 14872
R21597 vss.n13262 vss.n13261 14872
R21598 vss.n13259 vss.n13258 14872
R21599 vss.n13256 vss.n13255 14872
R21600 vss.n13253 vss.n13252 14872
R21601 vss.n13250 vss.n611 14872
R21602 vss.n13941 vss.n13940 14872
R21603 vss.n2305 vss.n2304 14872
R21604 vss.n12992 vss.n12991 14872
R21605 vss.n12989 vss.n12988 14872
R21606 vss.n12986 vss.n12985 14872
R21607 vss.n12983 vss.n12982 14872
R21608 vss.n12980 vss.n12979 14872
R21609 vss.n12977 vss.n12976 14872
R21610 vss.n13134 vss.n13133 14872
R21611 vss.n13131 vss.n13130 14872
R21612 vss.n13128 vss.n13127 14872
R21613 vss.n13125 vss.n13124 14872
R21614 vss.n13122 vss.n13121 14872
R21615 vss.n13119 vss.n13118 14872
R21616 vss.n9932 vss.n9931 14493.4
R21617 vss.n13937 vss.n13936 14493.4
R21618 vss.n9933 vss.n9932 13800
R21619 vss.n13938 vss.n13937 13800
R21620 vss.n13116 vss.n13115 13800
R21621 vss.n9954 vss.n9953 12952
R21622 vss.n9384 vss.n9383 12952
R21623 vss.n13265 vss.n13264 12952
R21624 vss.n13137 vss.n13136 12952
R21625 vss.n9670 vss.n9669 11556.6
R21626 vss.n14176 vss.n433 11376
R21627 vss.n9897 vss.n9896 11376
R21628 vss.n13056 vss.n2145 10957.3
R21629 vss.n14783 vss.n18 10957.3
R21630 vss.n9875 vss.n2767 10957.3
R21631 vss.n8986 vss.n7324 10957.3
R21632 vss.n190 vss.n18 10512
R21633 vss.n2934 vss.n2767 10512
R21634 vss.n7536 vss.n7324 10512
R21635 vss.n2304 vss.n2145 10512
R21636 vss.n8010 vss.n7299 9960
R21637 vss.n8122 vss.n7267 9648.25
R21638 vss.n5643 vss.n5642 8543.71
R21639 vss.n9049 vss.n9048 8543.71
R21640 vss.n13923 vss.n13922 8543.71
R21641 vss.n12098 vss.n11850 8543.71
R21642 vss.n9931 vss.n2708 7207.83
R21643 vss.n13936 vss.n13934 7207.83
R21644 vss.n5641 vss.n5640 6926.6
R21645 vss.n5639 vss.n5638 6926.6
R21646 vss.n5637 vss.n5636 6926.6
R21647 vss.n5635 vss.n5634 6926.6
R21648 vss.n5633 vss.n5632 6926.6
R21649 vss.n9047 vss.n9046 6926.6
R21650 vss.n9045 vss.n9044 6926.6
R21651 vss.n9043 vss.n9042 6926.6
R21652 vss.n9041 vss.n9040 6926.6
R21653 vss.n9039 vss.n9038 6926.6
R21654 vss.n13925 vss.n13924 6926.6
R21655 vss.n13927 vss.n13926 6926.6
R21656 vss.n13929 vss.n13928 6926.6
R21657 vss.n13931 vss.n13930 6926.6
R21658 vss.n13933 vss.n13932 6926.6
R21659 vss.n12035 vss.n10614 6926.6
R21660 vss.n12590 vss.n12589 6926.6
R21661 vss.n12588 vss.n12587 6926.6
R21662 vss.n12770 vss.n10321 6926.6
R21663 vss.n12769 vss.n12768 6926.6
R21664 vss.n8220 vss.n8219 6336
R21665 vss.n481 vss.n433 5848
R21666 vss.n9896 vss.n2743 5848
R21667 vss.n14061 vss.n495 5501.82
R21668 vss.n14061 vss.n14060 5365.58
R21669 vss.n8220 vss.n8010 5288
R21670 vss.n9669 vss.n9668 5056.22
R21671 vss.n13936 vss.n659 4856.95
R21672 vss.n9931 vss.n2707 4856.95
R21673 vss.n9669 vss.n5973 4549.42
R21674 vss.n11155 vss.n10433 4548.38
R21675 vss.n11155 vss.n11083 4548.38
R21676 vss.n11098 vss.n11080 4548.38
R21677 vss.n11080 vss.n10430 4548.38
R21678 vss.n11174 vss.n10436 4548.38
R21679 vss.n11174 vss.n11158 4548.38
R21680 vss.n11351 vss.n11047 4548.38
R21681 vss.n11351 vss.n10429 4548.38
R21682 vss.n11205 vss.n10439 4548.38
R21683 vss.n11205 vss.n11178 4548.38
R21684 vss.n11193 vss.n11175 4548.38
R21685 vss.n11175 vss.n10428 4548.38
R21686 vss.n11236 vss.n10442 4548.38
R21687 vss.n11236 vss.n11209 4548.38
R21688 vss.n11224 vss.n11206 4548.38
R21689 vss.n11206 vss.n10427 4548.38
R21690 vss.n11266 vss.n10445 4548.38
R21691 vss.n11266 vss.n11240 4548.38
R21692 vss.n11252 vss.n11237 4548.38
R21693 vss.n11237 vss.n10426 4548.38
R21694 vss.n11297 vss.n10448 4548.38
R21695 vss.n11297 vss.n11270 4548.38
R21696 vss.n11285 vss.n11267 4548.38
R21697 vss.n11267 vss.n10425 4548.38
R21698 vss.n11327 vss.n10451 4548.38
R21699 vss.n11327 vss.n11301 4548.38
R21700 vss.n11313 vss.n11298 4548.38
R21701 vss.n11298 vss.n10424 4548.38
R21702 vss.n3324 vss.n2603 4548.38
R21703 vss.n3335 vss.n3324 4548.38
R21704 vss.n3323 vss.n3314 4548.38
R21705 vss.n3314 vss.n2599 4548.38
R21706 vss.n4305 vss.n2606 4548.38
R21707 vss.n4305 vss.n3339 4548.38
R21708 vss.n4294 vss.n3336 4548.38
R21709 vss.n4294 vss.n2598 4548.38
R21710 vss.n4229 vss.n2609 4548.38
R21711 vss.n4229 vss.n3343 4548.38
R21712 vss.n4218 vss.n3340 4548.38
R21713 vss.n4218 vss.n2597 4548.38
R21714 vss.n3660 vss.n2612 4548.38
R21715 vss.n3660 vss.n3347 4548.38
R21716 vss.n3649 vss.n3344 4548.38
R21717 vss.n3649 vss.n2596 4548.38
R21718 vss.n3962 vss.n2615 4548.38
R21719 vss.n3962 vss.n3351 4548.38
R21720 vss.n3951 vss.n3348 4548.38
R21721 vss.n3951 vss.n2595 4548.38
R21722 vss.n3440 vss.n2618 4548.38
R21723 vss.n3440 vss.n3355 4548.38
R21724 vss.n3429 vss.n3352 4548.38
R21725 vss.n3429 vss.n2594 4548.38
R21726 vss.n3359 vss.n2621 4548.38
R21727 vss.n5857 vss.n3359 4548.38
R21728 vss.n3366 vss.n3356 4548.38
R21729 vss.n3366 vss.n2593 4548.38
R21730 vss.n9998 vss.n2624 4548.38
R21731 vss.n5881 vss.n2624 4548.38
R21732 vss.n5867 vss.n5858 4548.38
R21733 vss.n5867 vss.n2592 4548.38
R21734 vss.n2234 vss.n2196 4548.38
R21735 vss.n2230 vss.n2196 4548.38
R21736 vss.n2218 vss.n2199 4548.38
R21737 vss.n2222 vss.n2199 4548.38
R21738 vss.n12397 vss.n2192 4548.38
R21739 vss.n12393 vss.n2192 4548.38
R21740 vss.n12381 vss.n2195 4548.38
R21741 vss.n12385 vss.n2195 4548.38
R21742 vss.n12526 vss.n2188 4548.38
R21743 vss.n12522 vss.n2188 4548.38
R21744 vss.n12510 vss.n2191 4548.38
R21745 vss.n12514 vss.n2191 4548.38
R21746 vss.n10293 vss.n2184 4548.38
R21747 vss.n10289 vss.n2184 4548.38
R21748 vss.n10277 vss.n2187 4548.38
R21749 vss.n10281 vss.n2187 4548.38
R21750 vss.n10215 vss.n2180 4548.38
R21751 vss.n10211 vss.n2180 4548.38
R21752 vss.n10199 vss.n2183 4548.38
R21753 vss.n10203 vss.n2183 4548.38
R21754 vss.n2473 vss.n2176 4548.38
R21755 vss.n2469 vss.n2176 4548.38
R21756 vss.n2457 vss.n2179 4548.38
R21757 vss.n2461 vss.n2179 4548.38
R21758 vss.n2552 vss.n2172 4548.38
R21759 vss.n2548 vss.n2172 4548.38
R21760 vss.n2536 vss.n2175 4548.38
R21761 vss.n2540 vss.n2175 4548.38
R21762 vss.n7427 vss.n7403 4548.38
R21763 vss.n7430 vss.n7427 4548.38
R21764 vss.n8984 vss.n7406 4548.38
R21765 vss.n7419 vss.n7406 4548.38
R21766 vss.n7461 vss.n7399 4548.38
R21767 vss.n7464 vss.n7461 4548.38
R21768 vss.n7448 vss.n7402 4548.38
R21769 vss.n7448 vss.n7445 4548.38
R21770 vss.n7615 vss.n7395 4548.38
R21771 vss.n7618 vss.n7615 4548.38
R21772 vss.n7602 vss.n7398 4548.38
R21773 vss.n7602 vss.n7599 4548.38
R21774 vss.n7650 vss.n7391 4548.38
R21775 vss.n7653 vss.n7650 4548.38
R21776 vss.n7637 vss.n7394 4548.38
R21777 vss.n7637 vss.n7634 4548.38
R21778 vss.n7758 vss.n7387 4548.38
R21779 vss.n7761 vss.n7758 4548.38
R21780 vss.n7745 vss.n7390 4548.38
R21781 vss.n7745 vss.n7742 4548.38
R21782 vss.n7837 vss.n7383 4548.38
R21783 vss.n7840 vss.n7837 4548.38
R21784 vss.n7824 vss.n7386 4548.38
R21785 vss.n7824 vss.n7821 4548.38
R21786 vss.n7979 vss.n7379 4548.38
R21787 vss.n7982 vss.n7979 4548.38
R21788 vss.n7966 vss.n7382 4548.38
R21789 vss.n7966 vss.n7963 4548.38
R21790 vss.n7364 vss.n7348 4548.38
R21791 vss.n7365 vss.n7364 4548.38
R21792 vss.n7378 vss.n7341 4548.38
R21793 vss.n7354 vss.n7341 4548.38
R21794 vss.n14041 vss.n500 4548.38
R21795 vss.n14041 vss.n513 4548.38
R21796 vss.n509 vss.n503 4548.38
R21797 vss.n14058 vss.n503 4548.38
R21798 vss.n968 vss.n934 4548.38
R21799 vss.n942 vss.n934 4548.38
R21800 vss.n950 vss.n949 4548.38
R21801 vss.n950 vss.n931 4548.38
R21802 vss.n1495 vss.n971 4548.38
R21803 vss.n1495 vss.n1494 4548.38
R21804 vss.n1508 vss.n1507 4548.38
R21805 vss.n1508 vss.n930 4548.38
R21806 vss.n1578 vss.n974 4548.38
R21807 vss.n1578 vss.n1577 4548.38
R21808 vss.n1591 vss.n1590 4548.38
R21809 vss.n1591 vss.n929 4548.38
R21810 vss.n1415 vss.n977 4548.38
R21811 vss.n1415 vss.n1414 4548.38
R21812 vss.n1428 vss.n1427 4548.38
R21813 vss.n1428 vss.n928 4548.38
R21814 vss.n1283 vss.n980 4548.38
R21815 vss.n1283 vss.n1282 4548.38
R21816 vss.n1296 vss.n1295 4548.38
R21817 vss.n1296 vss.n927 4548.38
R21818 vss.n1022 vss.n983 4548.38
R21819 vss.n1022 vss.n1021 4548.38
R21820 vss.n1035 vss.n1034 4548.38
R21821 vss.n1035 vss.n926 4548.38
R21822 vss.n13208 vss.n986 4548.38
R21823 vss.n994 vss.n986 4548.38
R21824 vss.n1002 vss.n1001 4548.38
R21825 vss.n1002 vss.n925 4548.38
R21826 vss.n401 vss.n64 4548.38
R21827 vss.n401 vss.n71 4548.38
R21828 vss.n394 vss.n61 4548.38
R21829 vss.n394 vss.n74 4548.38
R21830 vss.n278 vss.n57 4548.38
R21831 vss.n278 vss.n77 4548.38
R21832 vss.n271 vss.n54 4548.38
R21833 vss.n271 vss.n80 4548.38
R21834 vss.n14435 vss.n53 4548.38
R21835 vss.n14435 vss.n81 4548.38
R21836 vss.n14428 vss.n50 4548.38
R21837 vss.n14428 vss.n84 4548.38
R21838 vss.n219 vss.n49 4548.38
R21839 vss.n219 vss.n85 4548.38
R21840 vss.n212 vss.n46 4548.38
R21841 vss.n212 vss.n88 4548.38
R21842 vss.n14630 vss.n45 4548.38
R21843 vss.n14630 vss.n89 4548.38
R21844 vss.n14623 vss.n42 4548.38
R21845 vss.n14623 vss.n92 4548.38
R21846 vss.n142 vss.n41 4548.38
R21847 vss.n142 vss.n93 4548.38
R21848 vss.n135 vss.n38 4548.38
R21849 vss.n135 vss.n96 4548.38
R21850 vss.n112 vss.n37 4548.38
R21851 vss.n112 vss.n97 4548.38
R21852 vss.n100 vss.n34 4548.38
R21853 vss.n14771 vss.n100 4548.38
R21854 vss.n14781 vss.n14780 4548.38
R21855 vss.n14780 vss.n67 4548.38
R21856 vss.n369 vss.n76 4548.38
R21857 vss.n369 vss.n58 4548.38
R21858 vss.n9857 vss.n2822 4548.38
R21859 vss.n2832 vss.n2822 4548.38
R21860 vss.n9872 vss.n2825 4548.38
R21861 vss.n9872 vss.n2826 4548.38
R21862 vss.n2865 vss.n2818 4548.38
R21863 vss.n2861 vss.n2818 4548.38
R21864 vss.n2849 vss.n2821 4548.38
R21865 vss.n2853 vss.n2821 4548.38
R21866 vss.n4996 vss.n2814 4548.38
R21867 vss.n4992 vss.n2814 4548.38
R21868 vss.n4980 vss.n2817 4548.38
R21869 vss.n4984 vss.n2817 4548.38
R21870 vss.n5073 vss.n2810 4548.38
R21871 vss.n5069 vss.n2810 4548.38
R21872 vss.n5057 vss.n2813 4548.38
R21873 vss.n5061 vss.n2813 4548.38
R21874 vss.n5198 vss.n2806 4548.38
R21875 vss.n5194 vss.n2806 4548.38
R21876 vss.n5182 vss.n2809 4548.38
R21877 vss.n5186 vss.n2809 4548.38
R21878 vss.n3099 vss.n2802 4548.38
R21879 vss.n3095 vss.n2802 4548.38
R21880 vss.n3083 vss.n2805 4548.38
R21881 vss.n3087 vss.n2805 4548.38
R21882 vss.n3179 vss.n2798 4548.38
R21883 vss.n3175 vss.n2798 4548.38
R21884 vss.n3163 vss.n2801 4548.38
R21885 vss.n3167 vss.n2801 4548.38
R21886 vss.n3256 vss.n2794 4548.38
R21887 vss.n3252 vss.n2794 4548.38
R21888 vss.n3240 vss.n2797 4548.38
R21889 vss.n3244 vss.n2797 4548.38
R21890 vss.n6257 vss.n6226 4548.38
R21891 vss.n6257 vss.n6225 4548.38
R21892 vss.n6244 vss.n6221 4548.38
R21893 vss.n6231 vss.n6221 4548.38
R21894 vss.n6295 vss.n6263 4548.38
R21895 vss.n6295 vss.n6262 4548.38
R21896 vss.n6282 vss.n6258 4548.38
R21897 vss.n6269 vss.n6258 4548.38
R21898 vss.n7108 vss.n6300 4548.38
R21899 vss.n7102 vss.n6300 4548.38
R21900 vss.n7118 vss.n6296 4548.38
R21901 vss.n7114 vss.n6296 4548.38
R21902 vss.n6610 vss.n6305 4548.38
R21903 vss.n6604 vss.n6305 4548.38
R21904 vss.n6620 vss.n6301 4548.38
R21905 vss.n6616 vss.n6301 4548.38
R21906 vss.n6919 vss.n6310 4548.38
R21907 vss.n6913 vss.n6310 4548.38
R21908 vss.n6929 vss.n6306 4548.38
R21909 vss.n6925 vss.n6306 4548.38
R21910 vss.n6383 vss.n6315 4548.38
R21911 vss.n6377 vss.n6315 4548.38
R21912 vss.n6393 vss.n6311 4548.38
R21913 vss.n6389 vss.n6311 4548.38
R21914 vss.n9286 vss.n6321 4548.38
R21915 vss.n9286 vss.n6320 4548.38
R21916 vss.n9273 vss.n6316 4548.38
R21917 vss.n9260 vss.n6316 4548.38
R21918 vss.n9316 vss.n9306 4548.38
R21919 vss.n9316 vss.n9303 4548.38
R21920 vss.n9295 vss.n9287 4548.38
R21921 vss.n9294 vss.n9287 4548.38
R21922 vss.n13047 vss.n2200 4548.38
R21923 vss.n13051 vss.n2200 4548.38
R21924 vss.n13032 vss.n2161 4548.38
R21925 vss.n13028 vss.n2161 4548.38
R21926 vss.n11343 vss.n11328 4548.38
R21927 vss.n11328 vss.n10452 4548.38
R21928 vss.n12670 vss.n10455 4548.38
R21929 vss.n11333 vss.n10455 4548.38
R21930 vss.n12767 vss.n2071 4186.8
R21931 vss.n13138 vss.n13137 4137.66
R21932 vss.n13265 vss.n728 4137.66
R21933 vss.n9383 vss.n9382 4137.66
R21934 vss.n9955 vss.n9954 4137.66
R21935 vss.n10000 vss.n2591 4121.92
R21936 vss.n13113 vss.n2072 4066.11
R21937 vss.n13077 vss.n13076 4051.68
R21938 vss.n9672 vss.n5970 3977.25
R21939 vss.n11091 vss.n11077 3789.35
R21940 vss.n11077 vss.n11076 3789.35
R21941 vss.n11089 vss.n11082 3789.35
R21942 vss.n11082 vss.n11081 3789.35
R21943 vss.n11097 vss.n11079 3789.35
R21944 vss.n11079 vss.n11078 3789.35
R21945 vss.n11161 vss.n11073 3789.35
R21946 vss.n11073 vss.n11072 3789.35
R21947 vss.n11166 vss.n11157 3789.35
R21948 vss.n11157 vss.n11156 3789.35
R21949 vss.n11162 vss.n11075 3789.35
R21950 vss.n11075 vss.n11074 3789.35
R21951 vss.n11186 vss.n11069 3789.35
R21952 vss.n11069 vss.n11068 3789.35
R21953 vss.n11184 vss.n11177 3789.35
R21954 vss.n11177 vss.n11176 3789.35
R21955 vss.n11192 vss.n11071 3789.35
R21956 vss.n11071 vss.n11070 3789.35
R21957 vss.n11217 vss.n11065 3789.35
R21958 vss.n11065 vss.n11064 3789.35
R21959 vss.n11215 vss.n11208 3789.35
R21960 vss.n11208 vss.n11207 3789.35
R21961 vss.n11223 vss.n11067 3789.35
R21962 vss.n11067 vss.n11066 3789.35
R21963 vss.n11243 vss.n11061 3789.35
R21964 vss.n11061 vss.n11060 3789.35
R21965 vss.n11257 vss.n11239 3789.35
R21966 vss.n11239 vss.n11238 3789.35
R21967 vss.n11244 vss.n11063 3789.35
R21968 vss.n11063 vss.n11062 3789.35
R21969 vss.n11278 vss.n11057 3789.35
R21970 vss.n11057 vss.n11056 3789.35
R21971 vss.n11276 vss.n11269 3789.35
R21972 vss.n11269 vss.n11268 3789.35
R21973 vss.n11284 vss.n11059 3789.35
R21974 vss.n11059 vss.n11058 3789.35
R21975 vss.n11304 vss.n11053 3789.35
R21976 vss.n11053 vss.n11052 3789.35
R21977 vss.n11318 vss.n11300 3789.35
R21978 vss.n11300 vss.n11299 3789.35
R21979 vss.n11305 vss.n11055 3789.35
R21980 vss.n11055 vss.n11054 3789.35
R21981 vss.n3331 vss.n3325 3789.35
R21982 vss.n3331 vss.n3330 3789.35
R21983 vss.n5886 vss.n5884 3789.35
R21984 vss.n5886 vss.n5885 3789.35
R21985 vss.n3317 vss.n3312 3789.35
R21986 vss.n3317 vss.n3316 3789.35
R21987 vss.n4311 vss.n4309 3789.35
R21988 vss.n4311 vss.n4310 3789.35
R21989 vss.n4318 vss.n4316 3789.35
R21990 vss.n4318 vss.n4317 3789.35
R21991 vss.n4300 vss.n4298 3789.35
R21992 vss.n4300 vss.n4299 3789.35
R21993 vss.n4235 vss.n4233 3789.35
R21994 vss.n4235 vss.n4234 3789.35
R21995 vss.n4242 vss.n4240 3789.35
R21996 vss.n4242 vss.n4241 3789.35
R21997 vss.n4224 vss.n4222 3789.35
R21998 vss.n4224 vss.n4223 3789.35
R21999 vss.n3666 vss.n3664 3789.35
R22000 vss.n3666 vss.n3665 3789.35
R22001 vss.n3673 vss.n3671 3789.35
R22002 vss.n3673 vss.n3672 3789.35
R22003 vss.n3655 vss.n3653 3789.35
R22004 vss.n3655 vss.n3654 3789.35
R22005 vss.n3968 vss.n3966 3789.35
R22006 vss.n3968 vss.n3967 3789.35
R22007 vss.n3975 vss.n3973 3789.35
R22008 vss.n3975 vss.n3974 3789.35
R22009 vss.n3957 vss.n3955 3789.35
R22010 vss.n3957 vss.n3956 3789.35
R22011 vss.n3446 vss.n3444 3789.35
R22012 vss.n3446 vss.n3445 3789.35
R22013 vss.n3453 vss.n3451 3789.35
R22014 vss.n3453 vss.n3452 3789.35
R22015 vss.n3435 vss.n3433 3789.35
R22016 vss.n3435 vss.n3434 3789.35
R22017 vss.n5853 vss.n3360 3789.35
R22018 vss.n5853 vss.n5852 3789.35
R22019 vss.n3379 vss.n3377 3789.35
R22020 vss.n3379 vss.n3378 3789.35
R22021 vss.n3372 vss.n3370 3789.35
R22022 vss.n3372 vss.n3371 3789.35
R22023 vss.n5865 vss.n5864 3789.35
R22024 vss.n5864 vss.n2625 3789.35
R22025 vss.n5862 vss.n5861 3789.35
R22026 vss.n5861 vss.n5860 3789.35
R22027 vss.n5873 vss.n5871 3789.35
R22028 vss.n5873 vss.n5872 3789.35
R22029 vss.n2235 vss.n2164 3789.35
R22030 vss.n2229 vss.n2164 3789.35
R22031 vss.n2207 vss.n2197 3789.35
R22032 vss.n2210 vss.n2197 3789.35
R22033 vss.n2217 vss.n2198 3789.35
R22034 vss.n2223 vss.n2198 3789.35
R22035 vss.n12398 vss.n2165 3789.35
R22036 vss.n12392 vss.n2165 3789.35
R22037 vss.n12370 vss.n2193 3789.35
R22038 vss.n12373 vss.n2193 3789.35
R22039 vss.n12380 vss.n2194 3789.35
R22040 vss.n12386 vss.n2194 3789.35
R22041 vss.n12527 vss.n2166 3789.35
R22042 vss.n12521 vss.n2166 3789.35
R22043 vss.n12499 vss.n2189 3789.35
R22044 vss.n12502 vss.n2189 3789.35
R22045 vss.n12509 vss.n2190 3789.35
R22046 vss.n12515 vss.n2190 3789.35
R22047 vss.n10294 vss.n2167 3789.35
R22048 vss.n10288 vss.n2167 3789.35
R22049 vss.n10266 vss.n2185 3789.35
R22050 vss.n10269 vss.n2185 3789.35
R22051 vss.n10276 vss.n2186 3789.35
R22052 vss.n10282 vss.n2186 3789.35
R22053 vss.n10216 vss.n2168 3789.35
R22054 vss.n10210 vss.n2168 3789.35
R22055 vss.n10188 vss.n2181 3789.35
R22056 vss.n10191 vss.n2181 3789.35
R22057 vss.n10198 vss.n2182 3789.35
R22058 vss.n10204 vss.n2182 3789.35
R22059 vss.n2474 vss.n2169 3789.35
R22060 vss.n2468 vss.n2169 3789.35
R22061 vss.n2446 vss.n2177 3789.35
R22062 vss.n2449 vss.n2177 3789.35
R22063 vss.n2456 vss.n2178 3789.35
R22064 vss.n2462 vss.n2178 3789.35
R22065 vss.n2553 vss.n2170 3789.35
R22066 vss.n2547 vss.n2170 3789.35
R22067 vss.n2525 vss.n2173 3789.35
R22068 vss.n2528 vss.n2173 3789.35
R22069 vss.n2535 vss.n2174 3789.35
R22070 vss.n2541 vss.n2174 3789.35
R22071 vss.n7432 vss.n7413 3789.35
R22072 vss.n7432 vss.n7431 3789.35
R22073 vss.n7415 vss.n7414 3789.35
R22074 vss.n7416 vss.n7415 3789.35
R22075 vss.n7420 vss.n7407 3789.35
R22076 vss.n7421 vss.n7420 3789.35
R22077 vss.n7466 vss.n7439 3789.35
R22078 vss.n7466 vss.n7465 3789.35
R22079 vss.n7442 vss.n7441 3789.35
R22080 vss.n7442 vss.n7440 3789.35
R22081 vss.n7454 vss.n7446 3789.35
R22082 vss.n7455 vss.n7454 3789.35
R22083 vss.n7620 vss.n7593 3789.35
R22084 vss.n7620 vss.n7619 3789.35
R22085 vss.n7596 vss.n7595 3789.35
R22086 vss.n7596 vss.n7594 3789.35
R22087 vss.n7608 vss.n7600 3789.35
R22088 vss.n7609 vss.n7608 3789.35
R22089 vss.n7655 vss.n7628 3789.35
R22090 vss.n7655 vss.n7654 3789.35
R22091 vss.n7631 vss.n7630 3789.35
R22092 vss.n7631 vss.n7629 3789.35
R22093 vss.n7643 vss.n7635 3789.35
R22094 vss.n7644 vss.n7643 3789.35
R22095 vss.n7763 vss.n7736 3789.35
R22096 vss.n7763 vss.n7762 3789.35
R22097 vss.n7739 vss.n7738 3789.35
R22098 vss.n7739 vss.n7737 3789.35
R22099 vss.n7751 vss.n7743 3789.35
R22100 vss.n7752 vss.n7751 3789.35
R22101 vss.n7842 vss.n7815 3789.35
R22102 vss.n7842 vss.n7841 3789.35
R22103 vss.n7818 vss.n7817 3789.35
R22104 vss.n7818 vss.n7816 3789.35
R22105 vss.n7830 vss.n7822 3789.35
R22106 vss.n7831 vss.n7830 3789.35
R22107 vss.n7984 vss.n7957 3789.35
R22108 vss.n7984 vss.n7983 3789.35
R22109 vss.n7960 vss.n7959 3789.35
R22110 vss.n7960 vss.n7958 3789.35
R22111 vss.n7972 vss.n7964 3789.35
R22112 vss.n7973 vss.n7972 3789.35
R22113 vss.n7370 vss.n7369 3789.35
R22114 vss.n7369 vss.n7349 3789.35
R22115 vss.n7351 vss.n7347 3789.35
R22116 vss.n7359 vss.n7351 3789.35
R22117 vss.n7352 vss.n7342 3789.35
R22118 vss.n7353 vss.n7352 3789.35
R22119 vss.n14046 vss.n14045 3789.35
R22120 vss.n14046 vss.n514 3789.35
R22121 vss.n14037 vss.n14036 3789.35
R22122 vss.n14037 vss.n510 3789.35
R22123 vss.n14054 vss.n504 3789.35
R22124 vss.n14054 vss.n14053 3789.35
R22125 vss.n941 vss.n940 3789.35
R22126 vss.n940 vss.n935 3789.35
R22127 vss.n962 vss.n960 3789.35
R22128 vss.n962 vss.n961 3789.35
R22129 vss.n955 vss.n947 3789.35
R22130 vss.n955 vss.n954 3789.35
R22131 vss.n1500 vss.n1492 3789.35
R22132 vss.n1500 vss.n1499 3789.35
R22133 vss.n1520 vss.n1518 3789.35
R22134 vss.n1520 vss.n1519 3789.35
R22135 vss.n1513 vss.n1505 3789.35
R22136 vss.n1513 vss.n1512 3789.35
R22137 vss.n1583 vss.n1575 3789.35
R22138 vss.n1583 vss.n1582 3789.35
R22139 vss.n1603 vss.n1601 3789.35
R22140 vss.n1603 vss.n1602 3789.35
R22141 vss.n1596 vss.n1588 3789.35
R22142 vss.n1596 vss.n1595 3789.35
R22143 vss.n1420 vss.n1412 3789.35
R22144 vss.n1420 vss.n1419 3789.35
R22145 vss.n1440 vss.n1438 3789.35
R22146 vss.n1440 vss.n1439 3789.35
R22147 vss.n1433 vss.n1425 3789.35
R22148 vss.n1433 vss.n1432 3789.35
R22149 vss.n1288 vss.n1280 3789.35
R22150 vss.n1288 vss.n1287 3789.35
R22151 vss.n1308 vss.n1306 3789.35
R22152 vss.n1308 vss.n1307 3789.35
R22153 vss.n1301 vss.n1293 3789.35
R22154 vss.n1301 vss.n1300 3789.35
R22155 vss.n1027 vss.n1019 3789.35
R22156 vss.n1027 vss.n1026 3789.35
R22157 vss.n1047 vss.n1045 3789.35
R22158 vss.n1047 vss.n1046 3789.35
R22159 vss.n1040 vss.n1032 3789.35
R22160 vss.n1040 vss.n1039 3789.35
R22161 vss.n993 vss.n992 3789.35
R22162 vss.n992 vss.n987 3789.35
R22163 vss.n1014 vss.n1012 3789.35
R22164 vss.n1014 vss.n1013 3789.35
R22165 vss.n1007 vss.n999 3789.35
R22166 vss.n1007 vss.n1006 3789.35
R22167 vss.n407 vss.n405 3789.35
R22168 vss.n407 vss.n406 3789.35
R22169 vss.n385 vss.n383 3789.35
R22170 vss.n385 vss.n384 3789.35
R22171 vss.n389 vss.n387 3789.35
R22172 vss.n389 vss.n388 3789.35
R22173 vss.n284 vss.n282 3789.35
R22174 vss.n284 vss.n283 3789.35
R22175 vss.n262 vss.n260 3789.35
R22176 vss.n262 vss.n261 3789.35
R22177 vss.n266 vss.n264 3789.35
R22178 vss.n266 vss.n265 3789.35
R22179 vss.n14441 vss.n14439 3789.35
R22180 vss.n14441 vss.n14440 3789.35
R22181 vss.n14419 vss.n14417 3789.35
R22182 vss.n14419 vss.n14418 3789.35
R22183 vss.n14423 vss.n14421 3789.35
R22184 vss.n14423 vss.n14422 3789.35
R22185 vss.n225 vss.n223 3789.35
R22186 vss.n225 vss.n224 3789.35
R22187 vss.n203 vss.n201 3789.35
R22188 vss.n203 vss.n202 3789.35
R22189 vss.n207 vss.n205 3789.35
R22190 vss.n207 vss.n206 3789.35
R22191 vss.n14636 vss.n14634 3789.35
R22192 vss.n14636 vss.n14635 3789.35
R22193 vss.n14614 vss.n14612 3789.35
R22194 vss.n14614 vss.n14613 3789.35
R22195 vss.n14618 vss.n14616 3789.35
R22196 vss.n14618 vss.n14617 3789.35
R22197 vss.n148 vss.n146 3789.35
R22198 vss.n148 vss.n147 3789.35
R22199 vss.n126 vss.n124 3789.35
R22200 vss.n126 vss.n125 3789.35
R22201 vss.n130 vss.n128 3789.35
R22202 vss.n130 vss.n129 3789.35
R22203 vss.n118 vss.n116 3789.35
R22204 vss.n118 vss.n117 3789.35
R22205 vss.n107 vss.n105 3789.35
R22206 vss.n107 vss.n106 3789.35
R22207 vss.n14767 vss.n14766 3789.35
R22208 vss.n14767 vss.n101 3789.35
R22209 vss.n14775 vss.n65 3789.35
R22210 vss.n14775 vss.n14774 3789.35
R22211 vss.n363 vss.n362 3789.35
R22212 vss.n363 vss.n70 3789.35
R22213 vss.n367 vss.n365 3789.35
R22214 vss.n367 vss.n366 3789.35
R22215 vss.n9858 vss.n2785 3789.35
R22216 vss.n2831 vss.n2785 3789.35
R22217 vss.n9856 vss.n2823 3789.35
R22218 vss.n9866 vss.n2823 3789.35
R22219 vss.n9850 vss.n2824 3789.35
R22220 vss.n2830 vss.n2824 3789.35
R22221 vss.n2866 vss.n2786 3789.35
R22222 vss.n2860 vss.n2786 3789.35
R22223 vss.n2838 vss.n2819 3789.35
R22224 vss.n2841 vss.n2819 3789.35
R22225 vss.n2848 vss.n2820 3789.35
R22226 vss.n2854 vss.n2820 3789.35
R22227 vss.n4997 vss.n2787 3789.35
R22228 vss.n4991 vss.n2787 3789.35
R22229 vss.n4969 vss.n2815 3789.35
R22230 vss.n4972 vss.n2815 3789.35
R22231 vss.n4979 vss.n2816 3789.35
R22232 vss.n4985 vss.n2816 3789.35
R22233 vss.n5074 vss.n2788 3789.35
R22234 vss.n5068 vss.n2788 3789.35
R22235 vss.n5046 vss.n2811 3789.35
R22236 vss.n5049 vss.n2811 3789.35
R22237 vss.n5056 vss.n2812 3789.35
R22238 vss.n5062 vss.n2812 3789.35
R22239 vss.n5199 vss.n2789 3789.35
R22240 vss.n5193 vss.n2789 3789.35
R22241 vss.n5171 vss.n2807 3789.35
R22242 vss.n5174 vss.n2807 3789.35
R22243 vss.n5181 vss.n2808 3789.35
R22244 vss.n5187 vss.n2808 3789.35
R22245 vss.n3100 vss.n2790 3789.35
R22246 vss.n3094 vss.n2790 3789.35
R22247 vss.n3072 vss.n2803 3789.35
R22248 vss.n3075 vss.n2803 3789.35
R22249 vss.n3082 vss.n2804 3789.35
R22250 vss.n3088 vss.n2804 3789.35
R22251 vss.n3180 vss.n2791 3789.35
R22252 vss.n3174 vss.n2791 3789.35
R22253 vss.n3152 vss.n2799 3789.35
R22254 vss.n3155 vss.n2799 3789.35
R22255 vss.n3162 vss.n2800 3789.35
R22256 vss.n3168 vss.n2800 3789.35
R22257 vss.n3257 vss.n2792 3789.35
R22258 vss.n3251 vss.n2792 3789.35
R22259 vss.n3229 vss.n2795 3789.35
R22260 vss.n3232 vss.n2795 3789.35
R22261 vss.n3239 vss.n2796 3789.35
R22262 vss.n3245 vss.n2796 3789.35
R22263 vss.n6235 vss.n6224 3789.35
R22264 vss.n6229 vss.n6224 3789.35
R22265 vss.n6241 vss.n6223 3789.35
R22266 vss.n6251 vss.n6223 3789.35
R22267 vss.n6243 vss.n6222 3789.35
R22268 vss.n6230 vss.n6222 3789.35
R22269 vss.n6273 vss.n6261 3789.35
R22270 vss.n6267 vss.n6261 3789.35
R22271 vss.n6279 vss.n6260 3789.35
R22272 vss.n6289 vss.n6260 3789.35
R22273 vss.n6281 vss.n6259 3789.35
R22274 vss.n6268 vss.n6259 3789.35
R22275 vss.n7098 vss.n6299 3789.35
R22276 vss.n7109 vss.n6299 3789.35
R22277 vss.n7121 vss.n6298 3789.35
R22278 vss.n7111 vss.n6298 3789.35
R22279 vss.n7119 vss.n6297 3789.35
R22280 vss.n7113 vss.n6297 3789.35
R22281 vss.n6600 vss.n6304 3789.35
R22282 vss.n6611 vss.n6304 3789.35
R22283 vss.n6623 vss.n6303 3789.35
R22284 vss.n6613 vss.n6303 3789.35
R22285 vss.n6621 vss.n6302 3789.35
R22286 vss.n6615 vss.n6302 3789.35
R22287 vss.n6909 vss.n6309 3789.35
R22288 vss.n6920 vss.n6309 3789.35
R22289 vss.n6932 vss.n6308 3789.35
R22290 vss.n6922 vss.n6308 3789.35
R22291 vss.n6930 vss.n6307 3789.35
R22292 vss.n6924 vss.n6307 3789.35
R22293 vss.n6373 vss.n6314 3789.35
R22294 vss.n6384 vss.n6314 3789.35
R22295 vss.n6396 vss.n6313 3789.35
R22296 vss.n6386 vss.n6313 3789.35
R22297 vss.n6394 vss.n6312 3789.35
R22298 vss.n6388 vss.n6312 3789.35
R22299 vss.n9264 vss.n6319 3789.35
R22300 vss.n9258 vss.n6319 3789.35
R22301 vss.n9270 vss.n6318 3789.35
R22302 vss.n9280 vss.n6318 3789.35
R22303 vss.n9272 vss.n6317 3789.35
R22304 vss.n9259 vss.n6317 3789.35
R22305 vss.n9308 vss.n9302 3789.35
R22306 vss.n9305 vss.n9302 3789.35
R22307 vss.n9317 vss.n6217 3789.35
R22308 vss.n9317 vss.n6218 3789.35
R22309 vss.n9301 vss.n9288 3789.35
R22310 vss.n9301 vss.n9290 3789.35
R22311 vss.n13053 vss.n2201 3789.35
R22312 vss.n13053 vss.n13052 3789.35
R22313 vss.n13043 vss.n2163 3789.35
R22314 vss.n13034 vss.n2163 3789.35
R22315 vss.n13024 vss.n2162 3789.35
R22316 vss.n13033 vss.n2162 3789.35
R22317 vss.n11350 vss.n11329 3789.35
R22318 vss.n11350 vss.n11349 3789.35
R22319 vss.n11338 vss.n11051 3789.35
R22320 vss.n11051 vss.n11050 3789.35
R22321 vss.n11332 vss.n11049 3789.35
R22322 vss.n11049 vss.n10456 3789.35
R22323 vss.n9671 vss.n9670 3624
R22324 vss.n482 vss.n481 3479.54
R22325 vss.n9720 vss.n2743 3479.54
R22326 vss.n9704 vss.n9703 3404.02
R22327 vss.n14063 vss.n14062 3385.58
R22328 vss.n9604 vss.n498 3056.88
R22329 vss.n9930 vss.n2706 3021.03
R22330 vss.n13935 vss.n494 3021.03
R22331 vss.n13113 vss.n13112 2820.86
R22332 vss.n9672 vss.n9671 2618.67
R22333 vss.n13115 vss.n13114 2602
R22334 vss.n14060 vss.n498 2563.49
R22335 vss.n2600 vss.n2591 2458.67
R22336 vss.n9671 vss.n5971 2458.67
R22337 vss.n9931 vss.n9930 2440.41
R22338 vss.n13936 vss.n13935 2440.41
R22339 vss.n9932 vss.n2706 2289.76
R22340 vss.n13937 vss.n494 2289.76
R22341 vss.t257 vss.n7332 2269.4
R22342 vss.t257 vss.n499 2269.4
R22343 vss.n14059 vss.t242 2269.4
R22344 vss.n14051 vss.t242 2269.4
R22345 vss.n9873 vss.n2784 2257.36
R22346 vss.n13139 vss.n2047 2172.79
R22347 vss.n13140 vss.n13139 2172.79
R22348 vss.n10408 vss.n10394 2172.79
R22349 vss.n10408 vss.n10393 2172.79
R22350 vss.n12653 vss.n12652 2172.79
R22351 vss.n12654 vss.n12653 2172.79
R22352 vss.n12641 vss.n12635 2172.79
R22353 vss.n12642 vss.n12635 2172.79
R22354 vss.n11137 vss.n11136 2172.79
R22355 vss.n11138 vss.n11137 2172.79
R22356 vss.n11125 vss.n11119 2172.79
R22357 vss.n11126 vss.n11119 2172.79
R22358 vss.n12677 vss.n10389 2172.79
R22359 vss.n12676 vss.n10389 2172.79
R22360 vss.n12685 vss.n10382 2172.79
R22361 vss.n12689 vss.n10382 2172.79
R22362 vss.n11427 vss.n11420 2172.79
R22363 vss.n11426 vss.n11420 2172.79
R22364 vss.n11435 vss.n11413 2172.79
R22365 vss.n11439 vss.n11413 2172.79
R22366 vss.n11380 vss.n11373 2172.79
R22367 vss.n11379 vss.n11373 2172.79
R22368 vss.n11388 vss.n11366 2172.79
R22369 vss.n11392 vss.n11366 2172.79
R22370 vss.n10955 vss.n10948 2172.79
R22371 vss.n10954 vss.n10948 2172.79
R22372 vss.n10963 vss.n10941 2172.79
R22373 vss.n10967 vss.n10941 2172.79
R22374 vss.n10792 vss.n10785 2172.79
R22375 vss.n10791 vss.n10785 2172.79
R22376 vss.n10800 vss.n10778 2172.79
R22377 vss.n10804 vss.n10778 2172.79
R22378 vss.n10748 vss.n10741 2172.79
R22379 vss.n10747 vss.n10741 2172.79
R22380 vss.n10756 vss.n10734 2172.79
R22381 vss.n10760 vss.n10734 2172.79
R22382 vss.n11574 vss.n11567 2172.79
R22383 vss.n11573 vss.n11567 2172.79
R22384 vss.n11582 vss.n11560 2172.79
R22385 vss.n11586 vss.n11560 2172.79
R22386 vss.n10571 vss.n10564 2172.79
R22387 vss.n10570 vss.n10564 2172.79
R22388 vss.n10579 vss.n10557 2172.79
R22389 vss.n10583 vss.n10557 2172.79
R22390 vss.n10527 vss.n10520 2172.79
R22391 vss.n10526 vss.n10520 2172.79
R22392 vss.n10535 vss.n10513 2172.79
R22393 vss.n10539 vss.n10513 2172.79
R22394 vss.n11948 vss.n11941 2172.79
R22395 vss.n11947 vss.n11941 2172.79
R22396 vss.n11956 vss.n11934 2172.79
R22397 vss.n11960 vss.n11934 2172.79
R22398 vss.n12096 vss.n11851 2172.79
R22399 vss.n12096 vss.n11852 2172.79
R22400 vss.n12064 vss.n11903 2172.79
R22401 vss.n12063 vss.n11903 2172.79
R22402 vss.n12046 vss.n11980 2172.79
R22403 vss.n12047 vss.n12046 2172.79
R22404 vss.n11911 vss.n11910 2172.79
R22405 vss.n11910 vss.n11909 2172.79
R22406 vss.n12037 vss.n12034 2172.79
R22407 vss.n12038 vss.n12037 2172.79
R22408 vss.n12024 vss.n11990 2172.79
R22409 vss.n12023 vss.n11990 2172.79
R22410 vss.n12601 vss.n10606 2172.79
R22411 vss.n12602 vss.n12601 2172.79
R22412 vss.n11999 vss.n11998 2172.79
R22413 vss.n11998 vss.n11997 2172.79
R22414 vss.n12592 vss.n10613 2172.79
R22415 vss.n12593 vss.n12592 2172.79
R22416 vss.n10669 vss.n10644 2172.79
R22417 vss.n10669 vss.n10643 2172.79
R22418 vss.n11611 vss.n10623 2172.79
R22419 vss.n11611 vss.n10624 2172.79
R22420 vss.n10672 vss.n10640 2172.79
R22421 vss.n10642 vss.n10640 2172.79
R22422 vss.n11622 vss.n10616 2172.79
R22423 vss.n11622 vss.n10617 2172.79
R22424 vss.n10856 vss.n10831 2172.79
R22425 vss.n10856 vss.n10830 2172.79
R22426 vss.n11530 vss.n10872 2172.79
R22427 vss.n11531 vss.n11530 2172.79
R22428 vss.n10861 vss.n10826 2172.79
R22429 vss.n10862 vss.n10826 2172.79
R22430 vss.n11521 vss.n11519 2172.79
R22431 vss.n11522 vss.n11521 2172.79
R22432 vss.n11509 vss.n10882 2172.79
R22433 vss.n11508 vss.n10882 2172.79
R22434 vss.n11481 vss.n10898 2172.79
R22435 vss.n11482 vss.n11481 2172.79
R22436 vss.n10890 vss.n10889 2172.79
R22437 vss.n10889 vss.n10888 2172.79
R22438 vss.n11472 vss.n11471 2172.79
R22439 vss.n11473 vss.n11472 2172.79
R22440 vss.n11461 vss.n10908 2172.79
R22441 vss.n11460 vss.n10908 2172.79
R22442 vss.n12754 vss.n10330 2172.79
R22443 vss.n12754 vss.n10331 2172.79
R22444 vss.n10919 vss.n10918 2172.79
R22445 vss.n10918 vss.n10917 2172.79
R22446 vss.n12765 vss.n10323 2172.79
R22447 vss.n12765 vss.n10324 2172.79
R22448 vss.n12729 vss.n10352 2172.79
R22449 vss.n12728 vss.n10352 2172.79
R22450 vss.n12711 vss.n12709 2172.79
R22451 vss.n12712 vss.n12711 2172.79
R22452 vss.n10360 vss.n10359 2172.79
R22453 vss.n10359 vss.n10358 2172.79
R22454 vss.n13111 vss.n2073 2172.79
R22455 vss.n13111 vss.n2074 2172.79
R22456 vss.n13094 vss.n2095 2172.79
R22457 vss.n13095 vss.n13094 2172.79
R22458 vss.n12924 vss.n10082 2172.79
R22459 vss.n12925 vss.n10082 2172.79
R22460 vss.n12941 vss.n10061 2172.79
R22461 vss.n10061 vss.n10059 2172.79
R22462 vss.n12997 vss.n2255 2172.79
R22463 vss.n12998 vss.n2255 2172.79
R22464 vss.n13010 vss.n13007 2172.79
R22465 vss.n13009 vss.n13007 2172.79
R22466 vss.n2302 vss.n2259 2172.79
R22467 vss.n2302 vss.n2260 2172.79
R22468 vss.n2285 vss.n2284 2172.79
R22469 vss.n2286 vss.n2285 2172.79
R22470 vss.n13075 vss.n2120 2172.79
R22471 vss.n13075 vss.n2121 2172.79
R22472 vss.n13058 vss.n2142 2172.79
R22473 vss.n13059 vss.n13058 2172.79
R22474 vss.n14157 vss.n456 2172.79
R22475 vss.n14158 vss.n456 2172.79
R22476 vss.n14174 vss.n434 2172.79
R22477 vss.n14174 vss.n435 2172.79
R22478 vss.n657 vss.n614 2172.79
R22479 vss.n657 vss.n615 2172.79
R22480 vss.n634 vss.n631 2172.79
R22481 vss.n633 vss.n631 2172.79
R22482 vss.n2017 vss.n2016 2172.79
R22483 vss.n2018 vss.n2017 2172.79
R22484 vss.n2005 vss.n1999 2172.79
R22485 vss.n2006 vss.n1999 2172.79
R22486 vss.n1082 vss.n1081 2172.79
R22487 vss.n1083 vss.n1082 2172.79
R22488 vss.n1070 vss.n1064 2172.79
R22489 vss.n1071 vss.n1064 2172.79
R22490 vss.n1343 vss.n1342 2172.79
R22491 vss.n1344 vss.n1343 2172.79
R22492 vss.n1331 vss.n1325 2172.79
R22493 vss.n1332 vss.n1325 2172.79
R22494 vss.n1475 vss.n1474 2172.79
R22495 vss.n1476 vss.n1475 2172.79
R22496 vss.n1463 vss.n1457 2172.79
R22497 vss.n1464 vss.n1457 2172.79
R22498 vss.n1638 vss.n1637 2172.79
R22499 vss.n1639 vss.n1638 2172.79
R22500 vss.n1626 vss.n1620 2172.79
R22501 vss.n1627 vss.n1620 2172.79
R22502 vss.n1556 vss.n1554 2172.79
R22503 vss.n1557 vss.n1556 2172.79
R22504 vss.n1543 vss.n1537 2172.79
R22505 vss.n1544 vss.n1537 2172.79
R22506 vss.n905 vss.n904 2172.79
R22507 vss.n906 vss.n905 2172.79
R22508 vss.n917 vss.n876 2172.79
R22509 vss.n917 vss.n875 2172.79
R22510 vss.n861 vss.n860 2172.79
R22511 vss.n862 vss.n861 2172.79
R22512 vss.n873 vss.n835 2172.79
R22513 vss.n873 vss.n834 2172.79
R22514 vss.n13944 vss.n610 2172.79
R22515 vss.n13945 vss.n13944 2172.79
R22516 vss.n832 vss.n818 2172.79
R22517 vss.n832 vss.n817 2172.79
R22518 vss.n13226 vss.n13225 2172.79
R22519 vss.n13227 vss.n13226 2172.79
R22520 vss.n13214 vss.n808 2172.79
R22521 vss.n13215 vss.n808 2172.79
R22522 vss.n1685 vss.n1684 2172.79
R22523 vss.n1686 vss.n1685 2172.79
R22524 vss.n1673 vss.n1667 2172.79
R22525 vss.n1674 vss.n1667 2172.79
R22526 vss.n1390 vss.n1389 2172.79
R22527 vss.n1391 vss.n1390 2172.79
R22528 vss.n1378 vss.n1372 2172.79
R22529 vss.n1379 vss.n1372 2172.79
R22530 vss.n1191 vss.n1190 2172.79
R22531 vss.n1192 vss.n1191 2172.79
R22532 vss.n1179 vss.n1173 2172.79
R22533 vss.n1180 vss.n1173 2172.79
R22534 vss.n1127 vss.n1126 2172.79
R22535 vss.n1128 vss.n1127 2172.79
R22536 vss.n1115 vss.n1109 2172.79
R22537 vss.n1116 vss.n1109 2172.79
R22538 vss.n13180 vss.n13173 2172.79
R22539 vss.n13179 vss.n13173 2172.79
R22540 vss.n13190 vss.n13189 2172.79
R22541 vss.n13191 vss.n13190 2172.79
R22542 vss.n188 vss.n173 2172.79
R22543 vss.n188 vss.n174 2172.79
R22544 vss.n14785 vss.n15 2172.79
R22545 vss.n17 vss.n15 2172.79
R22546 vss.n14728 vss.n14686 2172.79
R22547 vss.n14728 vss.n14687 2172.79
R22548 vss.n14711 vss.n14710 2172.79
R22549 vss.n14712 vss.n14711 2172.79
R22550 vss.n14586 vss.n14579 2172.79
R22551 vss.n14587 vss.n14579 2172.79
R22552 vss.n14599 vss.n14596 2172.79
R22553 vss.n14598 vss.n14596 2172.79
R22554 vss.n14533 vss.n14491 2172.79
R22555 vss.n14533 vss.n14492 2172.79
R22556 vss.n14516 vss.n14515 2172.79
R22557 vss.n14517 vss.n14516 2172.79
R22558 vss.n14391 vss.n14384 2172.79
R22559 vss.n14392 vss.n14384 2172.79
R22560 vss.n14404 vss.n14401 2172.79
R22561 vss.n14403 vss.n14401 2172.79
R22562 vss.n14338 vss.n14296 2172.79
R22563 vss.n14338 vss.n14297 2172.79
R22564 vss.n14321 vss.n14320 2172.79
R22565 vss.n14322 vss.n14321 2172.79
R22566 vss.n338 vss.n331 2172.79
R22567 vss.n339 vss.n331 2172.79
R22568 vss.n351 vss.n348 2172.79
R22569 vss.n350 vss.n348 2172.79
R22570 vss.n14219 vss.n14177 2172.79
R22571 vss.n14219 vss.n14178 2172.79
R22572 vss.n14202 vss.n14201 2172.79
R22573 vss.n14203 vss.n14202 2172.79
R22574 vss.n14117 vss.n14110 2172.79
R22575 vss.n14118 vss.n14110 2172.79
R22576 vss.n14130 vss.n14127 2172.79
R22577 vss.n14129 vss.n14127 2172.79
R22578 vss.n14226 vss.n428 2172.79
R22579 vss.n14227 vss.n428 2172.79
R22580 vss.n14239 vss.n14236 2172.79
R22581 vss.n14238 vss.n14236 2172.79
R22582 vss.n14292 vss.n312 2172.79
R22583 vss.n14292 vss.n313 2172.79
R22584 vss.n14275 vss.n14274 2172.79
R22585 vss.n14276 vss.n14275 2172.79
R22586 vss.n14345 vss.n305 2172.79
R22587 vss.n14346 vss.n305 2172.79
R22588 vss.n14358 vss.n14355 2172.79
R22589 vss.n14357 vss.n14355 2172.79
R22590 vss.n14487 vss.n253 2172.79
R22591 vss.n14487 vss.n254 2172.79
R22592 vss.n14470 vss.n14469 2172.79
R22593 vss.n14471 vss.n14470 2172.79
R22594 vss.n14540 vss.n246 2172.79
R22595 vss.n14541 vss.n246 2172.79
R22596 vss.n14553 vss.n14550 2172.79
R22597 vss.n14552 vss.n14550 2172.79
R22598 vss.n14682 vss.n194 2172.79
R22599 vss.n14682 vss.n195 2172.79
R22600 vss.n14665 vss.n14664 2172.79
R22601 vss.n14666 vss.n14665 2172.79
R22602 vss.n14735 vss.n169 2172.79
R22603 vss.n14736 vss.n169 2172.79
R22604 vss.n14748 vss.n14745 2172.79
R22605 vss.n14747 vss.n14745 2172.79
R22606 vss.n14153 vss.n460 2172.79
R22607 vss.n460 vss.n459 2172.79
R22608 vss.n13581 vss.n13566 2172.79
R22609 vss.n13581 vss.n13567 2172.79
R22610 vss.n13607 vss.n13545 2172.79
R22611 vss.n13607 vss.n13546 2172.79
R22612 vss.n13590 vss.n13587 2172.79
R22613 vss.n13591 vss.n13587 2172.79
R22614 vss.n13919 vss.n13302 2172.79
R22615 vss.n13907 vss.n13324 2172.79
R22616 vss.n13908 vss.n13324 2172.79
R22617 vss.n13304 vss.n13302 2172.79
R22618 vss.n13875 vss.n13343 2172.79
R22619 vss.n13876 vss.n13343 2172.79
R22620 vss.n13896 vss.n13326 2172.79
R22621 vss.n13896 vss.n13327 2172.79
R22622 vss.n13871 vss.n13344 2172.79
R22623 vss.n13852 vss.n13363 2172.79
R22624 vss.n13853 vss.n13363 2172.79
R22625 vss.n13346 vss.n13344 2172.79
R22626 vss.n13821 vss.n13384 2172.79
R22627 vss.n13822 vss.n13384 2172.79
R22628 vss.n13842 vss.n13365 2172.79
R22629 vss.n13842 vss.n13366 2172.79
R22630 vss.n13817 vss.n13385 2172.79
R22631 vss.n13802 vss.n13404 2172.79
R22632 vss.n13803 vss.n13404 2172.79
R22633 vss.n13387 vss.n13385 2172.79
R22634 vss.n13770 vss.n13423 2172.79
R22635 vss.n13771 vss.n13423 2172.79
R22636 vss.n13791 vss.n13406 2172.79
R22637 vss.n13791 vss.n13407 2172.79
R22638 vss.n13766 vss.n13424 2172.79
R22639 vss.n13747 vss.n13443 2172.79
R22640 vss.n13748 vss.n13443 2172.79
R22641 vss.n13426 vss.n13424 2172.79
R22642 vss.n13716 vss.n13464 2172.79
R22643 vss.n13717 vss.n13464 2172.79
R22644 vss.n13737 vss.n13445 2172.79
R22645 vss.n13737 vss.n13446 2172.79
R22646 vss.n13712 vss.n13465 2172.79
R22647 vss.n13697 vss.n13484 2172.79
R22648 vss.n13698 vss.n13484 2172.79
R22649 vss.n13467 vss.n13465 2172.79
R22650 vss.n13665 vss.n13503 2172.79
R22651 vss.n13666 vss.n13503 2172.79
R22652 vss.n13686 vss.n13486 2172.79
R22653 vss.n13686 vss.n13487 2172.79
R22654 vss.n13661 vss.n13504 2172.79
R22655 vss.n13642 vss.n13523 2172.79
R22656 vss.n13643 vss.n13523 2172.79
R22657 vss.n13506 vss.n13504 2172.79
R22658 vss.n13611 vss.n13544 2172.79
R22659 vss.n13612 vss.n13544 2172.79
R22660 vss.n13632 vss.n13525 2172.79
R22661 vss.n13632 vss.n13526 2172.79
R22662 vss.n14006 vss.n532 2172.79
R22663 vss.n14005 vss.n532 2172.79
R22664 vss.n14014 vss.n525 2172.79
R22665 vss.n14018 vss.n525 2172.79
R22666 vss.n14000 vss.n537 2172.79
R22667 vss.n14000 vss.n538 2172.79
R22668 vss.n677 vss.n660 2172.79
R22669 vss.n677 vss.n661 2172.79
R22670 vss.n13971 vss.n571 2172.79
R22671 vss.n13970 vss.n571 2172.79
R22672 vss.n13979 vss.n564 2172.79
R22673 vss.n13983 vss.n564 2172.79
R22674 vss.n13965 vss.n576 2172.79
R22675 vss.n13965 vss.n577 2172.79
R22676 vss.n777 vss.n776 2172.79
R22677 vss.n776 vss.n763 2172.79
R22678 vss.n13248 vss.n743 2172.79
R22679 vss.n13248 vss.n744 2172.79
R22680 vss.n783 vss.n780 2172.79
R22681 vss.n787 vss.n780 2172.79
R22682 vss.n1730 vss.n1726 2172.79
R22683 vss.n1731 vss.n1726 2172.79
R22684 vss.n1748 vss.n1747 2172.79
R22685 vss.n1747 vss.n1707 2172.79
R22686 vss.n1783 vss.n1758 2172.79
R22687 vss.n1782 vss.n1758 2172.79
R22688 vss.n1791 vss.n1751 2172.79
R22689 vss.n1795 vss.n1751 2172.79
R22690 vss.n1777 vss.n1762 2172.79
R22691 vss.n1777 vss.n1763 2172.79
R22692 vss.n1819 vss.n1818 2172.79
R22693 vss.n1818 vss.n1264 2172.79
R22694 vss.n1830 vss.n1233 2172.79
R22695 vss.n1233 vss.n1232 2172.79
R22696 vss.n1822 vss.n1248 2172.79
R22697 vss.n1262 vss.n1248 2172.79
R22698 vss.n1834 vss.n1230 2172.79
R22699 vss.n1835 vss.n1230 2172.79
R22700 vss.n1852 vss.n1851 2172.79
R22701 vss.n1851 vss.n1211 2172.79
R22702 vss.n1887 vss.n1862 2172.79
R22703 vss.n1886 vss.n1862 2172.79
R22704 vss.n1895 vss.n1855 2172.79
R22705 vss.n1899 vss.n1855 2172.79
R22706 vss.n1881 vss.n1866 2172.79
R22707 vss.n1881 vss.n1867 2172.79
R22708 vss.n1923 vss.n1922 2172.79
R22709 vss.n1922 vss.n1146 2172.79
R22710 vss.n1958 vss.n1933 2172.79
R22711 vss.n1957 vss.n1933 2172.79
R22712 vss.n1966 vss.n1926 2172.79
R22713 vss.n1970 vss.n1926 2172.79
R22714 vss.n1952 vss.n1937 2172.79
R22715 vss.n1952 vss.n1938 2172.79
R22716 vss.n13300 vss.n690 2172.79
R22717 vss.n13300 vss.n691 2172.79
R22718 vss.n13270 vss.n724 2172.79
R22719 vss.n13269 vss.n724 2172.79
R22720 vss.n13278 vss.n717 2172.79
R22721 vss.n13282 vss.n717 2172.79
R22722 vss.n9607 vss.n9600 2172.79
R22723 vss.n9608 vss.n9600 2172.79
R22724 vss.n9620 vss.n9617 2172.79
R22725 vss.n9619 vss.n9617 2172.79
R22726 vss.n7534 vss.n7491 2172.79
R22727 vss.n7534 vss.n7492 2172.79
R22728 vss.n7517 vss.n7516 2172.79
R22729 vss.n7518 vss.n7517 2172.79
R22730 vss.n8946 vss.n8904 2172.79
R22731 vss.n8946 vss.n8905 2172.79
R22732 vss.n8929 vss.n8928 2172.79
R22733 vss.n8930 vss.n8929 2172.79
R22734 vss.n7566 vss.n7559 2172.79
R22735 vss.n7567 vss.n7559 2172.79
R22736 vss.n7579 vss.n7576 2172.79
R22737 vss.n7578 vss.n7576 2172.79
R22738 vss.n8827 vss.n8785 2172.79
R22739 vss.n8827 vss.n8786 2172.79
R22740 vss.n8810 vss.n8809 2172.79
R22741 vss.n8811 vss.n8810 2172.79
R22742 vss.n7709 vss.n7702 2172.79
R22743 vss.n7710 vss.n7702 2172.79
R22744 vss.n7722 vss.n7719 2172.79
R22745 vss.n7721 vss.n7719 2172.79
R22746 vss.n7789 vss.n7782 2172.79
R22747 vss.n7790 vss.n7782 2172.79
R22748 vss.n7802 vss.n7799 2172.79
R22749 vss.n7801 vss.n7799 2172.79
R22750 vss.n7930 vss.n7923 2172.79
R22751 vss.n7931 vss.n7923 2172.79
R22752 vss.n7943 vss.n7940 2172.79
R22753 vss.n7942 vss.n7940 2172.79
R22754 vss.n8217 vss.n8175 2172.79
R22755 vss.n8217 vss.n8176 2172.79
R22756 vss.n8200 vss.n8199 2172.79
R22757 vss.n8201 vss.n8200 2172.79
R22758 vss.n8224 vss.n8006 2172.79
R22759 vss.n8225 vss.n8006 2172.79
R22760 vss.n8237 vss.n8234 2172.79
R22761 vss.n8236 vss.n8234 2172.79
R22762 vss.n9005 vss.n7300 2172.79
R22763 vss.n9005 vss.n7301 2172.79
R22764 vss.n8988 vss.n7322 2172.79
R22765 vss.n8989 vss.n8988 2172.79
R22766 vss.n8715 vss.n7863 2172.79
R22767 vss.n8716 vss.n7863 2172.79
R22768 vss.n8728 vss.n8725 2172.79
R22769 vss.n8727 vss.n8725 2172.79
R22770 vss.n8781 vss.n7683 2172.79
R22771 vss.n8781 vss.n7684 2172.79
R22772 vss.n8764 vss.n8763 2172.79
R22773 vss.n8765 vss.n8764 2172.79
R22774 vss.n8834 vss.n7676 2172.79
R22775 vss.n8835 vss.n7676 2172.79
R22776 vss.n8847 vss.n8844 2172.79
R22777 vss.n8846 vss.n8844 2172.79
R22778 vss.n8900 vss.n7540 2172.79
R22779 vss.n8900 vss.n7541 2172.79
R22780 vss.n8883 vss.n8882 2172.79
R22781 vss.n8884 vss.n8883 2172.79
R22782 vss.n8953 vss.n7487 2172.79
R22783 vss.n8954 vss.n7487 2172.79
R22784 vss.n8966 vss.n8963 2172.79
R22785 vss.n8965 vss.n8963 2172.79
R22786 vss.n8081 vss.n8077 2172.79
R22787 vss.n8082 vss.n8077 2172.79
R22788 vss.n8098 vss.n8053 2172.79
R22789 vss.n8098 vss.n8054 2172.79
R22790 vss.n9353 vss.n9352 2172.79
R22791 vss.n9354 vss.n9353 2172.79
R22792 vss.n9341 vss.n9334 2172.79
R22793 vss.n9342 vss.n9334 2172.79
R22794 vss.n6357 vss.n6356 2172.79
R22795 vss.n6358 vss.n6357 2172.79
R22796 vss.n6345 vss.n6338 2172.79
R22797 vss.n6346 vss.n6338 2172.79
R22798 vss.n6435 vss.n6434 2172.79
R22799 vss.n6436 vss.n6435 2172.79
R22800 vss.n6423 vss.n6416 2172.79
R22801 vss.n6424 vss.n6416 2172.79
R22802 vss.n6971 vss.n6970 2172.79
R22803 vss.n6972 vss.n6971 2172.79
R22804 vss.n6959 vss.n6952 2172.79
R22805 vss.n6960 vss.n6952 2172.79
R22806 vss.n6662 vss.n6661 2172.79
R22807 vss.n6663 vss.n6662 2172.79
R22808 vss.n6650 vss.n6643 2172.79
R22809 vss.n6651 vss.n6643 2172.79
R22810 vss.n7160 vss.n7159 2172.79
R22811 vss.n7161 vss.n7160 2172.79
R22812 vss.n7148 vss.n7141 2172.79
R22813 vss.n7149 vss.n7141 2172.79
R22814 vss.n9443 vss.n9400 2172.79
R22815 vss.n9443 vss.n9401 2172.79
R22816 vss.n9421 vss.n9417 2172.79
R22817 vss.n9420 vss.n9417 2172.79
R22818 vss.n6042 vss.n6040 2172.79
R22819 vss.n6043 vss.n6042 2172.79
R22820 vss.n6029 vss.n6022 2172.79
R22821 vss.n6030 vss.n6022 2172.79
R22822 vss.n9485 vss.n9445 2172.79
R22823 vss.n9485 vss.n9446 2172.79
R22824 vss.n9466 vss.n9461 2172.79
R22825 vss.n9465 vss.n9461 2172.79
R22826 vss.n9493 vss.n6167 2172.79
R22827 vss.n9494 vss.n9493 2172.79
R22828 vss.n6156 vss.n6149 2172.79
R22829 vss.n6157 vss.n6149 2172.79
R22830 vss.n7211 vss.n7210 2172.79
R22831 vss.n7212 vss.n7211 2172.79
R22832 vss.n7199 vss.n7192 2172.79
R22833 vss.n7200 vss.n7192 2172.79
R22834 vss.n6706 vss.n6705 2172.79
R22835 vss.n6707 vss.n6706 2172.79
R22836 vss.n6694 vss.n6687 2172.79
R22837 vss.n6695 vss.n6687 2172.79
R22838 vss.n7020 vss.n7019 2172.79
R22839 vss.n7021 vss.n7020 2172.79
R22840 vss.n7008 vss.n7001 2172.79
R22841 vss.n7009 vss.n7001 2172.79
R22842 vss.n6480 vss.n6479 2172.79
R22843 vss.n6481 vss.n6480 2172.79
R22844 vss.n6468 vss.n6461 2172.79
R22845 vss.n6469 vss.n6461 2172.79
R22846 vss.n9183 vss.n9182 2172.79
R22847 vss.n9184 vss.n9183 2172.79
R22848 vss.n9171 vss.n9164 2172.79
R22849 vss.n9172 vss.n9164 2172.79
R22850 vss.n9381 vss.n6185 2172.79
R22851 vss.n9381 vss.n6186 2172.79
R22852 vss.n6206 vss.n6202 2172.79
R22853 vss.n6205 vss.n6202 2172.79
R22854 vss.n8050 vss.n8011 2172.79
R22855 vss.n8035 vss.n8034 2172.79
R22856 vss.n8036 vss.n8035 2172.79
R22857 vss.n8013 vss.n8011 2172.79
R22858 vss.n9667 vss.n5974 2172.79
R22859 vss.n9667 vss.n5975 2172.79
R22860 vss.n9650 vss.n5996 2172.79
R22861 vss.n9651 vss.n9650 2172.79
R22862 vss.n8151 vss.n8124 2172.79
R22863 vss.n8136 vss.n8132 2172.79
R22864 vss.n8140 vss.n8132 2172.79
R22865 vss.n8151 vss.n5999 2172.79
R22866 vss.n8155 vss.n8121 2172.79
R22867 vss.n8172 vss.n8100 2172.79
R22868 vss.n8172 vss.n8101 2172.79
R22869 vss.n8156 vss.n8121 2172.79
R22870 vss.n9036 vss.n7268 2172.79
R22871 vss.n9036 vss.n7269 2172.79
R22872 vss.n9019 vss.n7290 2172.79
R22873 vss.n9020 vss.n9019 2172.79
R22874 vss.n8281 vss.n7900 2172.79
R22875 vss.n8281 vss.n7901 2172.79
R22876 vss.n9010 vss.n7297 2172.79
R22877 vss.n9011 vss.n9010 2172.79
R22878 vss.n8285 vss.n7899 2172.79
R22879 vss.n8286 vss.n7899 2172.79
R22880 vss.n8302 vss.n7878 2172.79
R22881 vss.n8302 vss.n7879 2172.79
R22882 vss.n8691 vss.n8318 2172.79
R22883 vss.n8692 vss.n8318 2172.79
R22884 vss.n8708 vss.n7867 2172.79
R22885 vss.n8708 vss.n7868 2172.79
R22886 vss.n8325 vss.n8324 2172.79
R22887 vss.n8326 vss.n8325 2172.79
R22888 vss.n8675 vss.n8345 2172.79
R22889 vss.n8348 vss.n8345 2172.79
R22890 vss.n8650 vss.n8363 2172.79
R22891 vss.n8649 vss.n8363 2172.79
R22892 vss.n8666 vss.n8665 2172.79
R22893 vss.n8667 vss.n8666 2172.79
R22894 vss.n8370 vss.n8369 2172.79
R22895 vss.n8371 vss.n8370 2172.79
R22896 vss.n8632 vss.n8395 2172.79
R22897 vss.n8398 vss.n8395 2172.79
R22898 vss.n8606 vss.n8416 2172.79
R22899 vss.n8605 vss.n8416 2172.79
R22900 vss.n8623 vss.n8621 2172.79
R22901 vss.n8624 vss.n8623 2172.79
R22902 vss.n8423 vss.n8422 2172.79
R22903 vss.n8424 vss.n8423 2172.79
R22904 vss.n8588 vss.n8443 2172.79
R22905 vss.n8446 vss.n8443 2172.79
R22906 vss.n8563 vss.n8461 2172.79
R22907 vss.n8562 vss.n8461 2172.79
R22908 vss.n8579 vss.n8578 2172.79
R22909 vss.n8580 vss.n8579 2172.79
R22910 vss.n8468 vss.n8467 2172.79
R22911 vss.n8469 vss.n8468 2172.79
R22912 vss.n8545 vss.n8493 2172.79
R22913 vss.n8496 vss.n8493 2172.79
R22914 vss.n8523 vss.n8509 2172.79
R22915 vss.n8536 vss.n8534 2172.79
R22916 vss.n8537 vss.n8536 2172.79
R22917 vss.n8524 vss.n8509 2172.79
R22918 vss.n9555 vss.n6072 2172.79
R22919 vss.n9554 vss.n6072 2172.79
R22920 vss.n9563 vss.n6065 2172.79
R22921 vss.n9567 vss.n6065 2172.79
R22922 vss.n9549 vss.n6077 2172.79
R22923 vss.n9549 vss.n6078 2172.79
R22924 vss.n7265 vss.n7248 2172.79
R22925 vss.n7265 vss.n7249 2172.79
R22926 vss.n9520 vss.n6111 2172.79
R22927 vss.n9519 vss.n6111 2172.79
R22928 vss.n9528 vss.n6104 2172.79
R22929 vss.n9532 vss.n6104 2172.79
R22930 vss.n9514 vss.n6116 2172.79
R22931 vss.n9514 vss.n6117 2172.79
R22932 vss.n7246 vss.n6575 2172.79
R22933 vss.n7246 vss.n6576 2172.79
R22934 vss.n6762 vss.n6749 2172.79
R22935 vss.n6749 vss.n6748 2172.79
R22936 vss.n7234 vss.n6581 2172.79
R22937 vss.n7234 vss.n6582 2172.79
R22938 vss.n6766 vss.n6746 2172.79
R22939 vss.n6767 vss.n6746 2172.79
R22940 vss.n6784 vss.n6783 2172.79
R22941 vss.n6783 vss.n6727 2172.79
R22942 vss.n7065 vss.n6794 2172.79
R22943 vss.n7064 vss.n6794 2172.79
R22944 vss.n7073 vss.n6787 2172.79
R22945 vss.n7077 vss.n6787 2172.79
R22946 vss.n7059 vss.n6798 2172.79
R22947 vss.n7059 vss.n6799 2172.79
R22948 vss.n6826 vss.n6825 2172.79
R22949 vss.n6825 vss.n6818 2172.79
R22950 vss.n6895 vss.n6848 2172.79
R22951 vss.n6896 vss.n6848 2172.79
R22952 vss.n7043 vss.n6827 2172.79
R22953 vss.n7043 vss.n6828 2172.79
R22954 vss.n6891 vss.n6849 2172.79
R22955 vss.n6891 vss.n6850 2172.79
R22956 vss.n6877 vss.n6876 2172.79
R22957 vss.n6876 vss.n6869 2172.79
R22958 vss.n9228 vss.n6505 2172.79
R22959 vss.n9227 vss.n6505 2172.79
R22960 vss.n9236 vss.n6498 2172.79
R22961 vss.n9240 vss.n6498 2172.79
R22962 vss.n9222 vss.n6509 2172.79
R22963 vss.n9222 vss.n6510 2172.79
R22964 vss.n6566 vss.n6557 2172.79
R22965 vss.n6566 vss.n6559 2172.79
R22966 vss.n9080 vss.n9067 2172.79
R22967 vss.n9067 vss.n9066 2172.79
R22968 vss.n9206 vss.n6528 2172.79
R22969 vss.n9206 vss.n6529 2172.79
R22970 vss.n9086 vss.n9061 2172.79
R22971 vss.n9085 vss.n9061 2172.79
R22972 vss.n9097 vss.n9096 2172.79
R22973 vss.n9096 vss.n9052 2172.79
R22974 vss.n9121 vss.n9119 2172.79
R22975 vss.n9122 vss.n9119 2172.79
R22976 vss.n9138 vss.n9098 2172.79
R22977 vss.n9138 vss.n9099 2172.79
R22978 vss.n5957 vss.n5951 2172.79
R22979 vss.n5958 vss.n5951 2172.79
R22980 vss.n9674 vss.n5967 2172.79
R22981 vss.n5969 vss.n5967 2172.79
R22982 vss.n9894 vss.n2744 2172.79
R22983 vss.n9894 vss.n2745 2172.79
R22984 vss.n9877 vss.n2766 2172.79
R22985 vss.n9878 vss.n9877 2172.79
R22986 vss.n9707 vss.n9699 2172.79
R22987 vss.n9708 vss.n9699 2172.79
R22988 vss.n9721 vss.n9717 2172.79
R22989 vss.n9719 vss.n9717 2172.79
R22990 vss.n3285 vss.n3277 2172.79
R22991 vss.n3286 vss.n3277 2172.79
R22992 vss.n3299 vss.n3294 2172.79
R22993 vss.n3298 vss.n3294 2172.79
R22994 vss.n2578 vss.n2572 2172.79
R22995 vss.n2579 vss.n2572 2172.79
R22996 vss.n10002 vss.n2588 2172.79
R22997 vss.n2590 vss.n2588 2172.79
R22998 vss.n5922 vss.n5921 2172.79
R22999 vss.n5923 vss.n5922 2172.79
R23000 vss.n5910 vss.n5903 2172.79
R23001 vss.n5911 vss.n5903 2172.79
R23002 vss.n9761 vss.n9760 2172.79
R23003 vss.n9776 vss.n9750 2172.79
R23004 vss.n9780 vss.n9750 2172.79
R23005 vss.n9767 vss.n9760 2172.79
R23006 vss.n3201 vss.n3200 2172.79
R23007 vss.n3216 vss.n3190 2172.79
R23008 vss.n3220 vss.n3190 2172.79
R23009 vss.n3207 vss.n3200 2172.79
R23010 vss.n9801 vss.n2993 2172.79
R23011 vss.n3018 vss.n3012 2172.79
R23012 vss.n3022 vss.n3012 2172.79
R23013 vss.n2995 vss.n2993 2172.79
R23014 vss.n5231 vss.n5230 2172.79
R23015 vss.n5246 vss.n5220 2172.79
R23016 vss.n5250 vss.n5220 2172.79
R23017 vss.n5237 vss.n5230 2172.79
R23018 vss.n3044 vss.n3043 2172.79
R23019 vss.n3059 vss.n3033 2172.79
R23020 vss.n3063 vss.n3033 2172.79
R23021 vss.n3050 vss.n3043 2172.79
R23022 vss.n5101 vss.n5100 2172.79
R23023 vss.n5116 vss.n5090 2172.79
R23024 vss.n5120 vss.n5090 2172.79
R23025 vss.n5107 vss.n5100 2172.79
R23026 vss.n5290 vss.n5289 2172.79
R23027 vss.n5305 vss.n5279 2172.79
R23028 vss.n5309 vss.n5279 2172.79
R23029 vss.n5296 vss.n5289 2172.79
R23030 vss.n5018 vss.n5017 2172.79
R23031 vss.n5033 vss.n5007 2172.79
R23032 vss.n5037 vss.n5007 2172.79
R23033 vss.n5024 vss.n5017 2172.79
R23034 vss.n4899 vss.n4898 2172.79
R23035 vss.n4914 vss.n4888 2172.79
R23036 vss.n4918 vss.n4888 2172.79
R23037 vss.n4905 vss.n4898 2172.79
R23038 vss.n9928 vss.n2709 2172.79
R23039 vss.n9928 vss.n2710 2172.79
R23040 vss.n9911 vss.n2731 2172.79
R23041 vss.n9912 vss.n9911 2172.79
R23042 vss.n4665 vss.n4637 2172.79
R23043 vss.n4665 vss.n4638 2172.79
R23044 vss.n9902 vss.n2738 2172.79
R23045 vss.n9903 vss.n9902 2172.79
R23046 vss.n5630 vss.n4628 2172.79
R23047 vss.n5630 vss.n4629 2172.79
R23048 vss.n5613 vss.n4683 2172.79
R23049 vss.n5614 vss.n5613 2172.79
R23050 vss.n5588 vss.n4698 2172.79
R23051 vss.n5587 vss.n4698 2172.79
R23052 vss.n5604 vss.n5603 2172.79
R23053 vss.n5605 vss.n5604 2172.79
R23054 vss.n4705 vss.n4704 2172.79
R23055 vss.n4706 vss.n4705 2172.79
R23056 vss.n5570 vss.n4723 2172.79
R23057 vss.n4726 vss.n4723 2172.79
R23058 vss.n5545 vss.n4741 2172.79
R23059 vss.n5544 vss.n4741 2172.79
R23060 vss.n5561 vss.n5560 2172.79
R23061 vss.n5562 vss.n5561 2172.79
R23062 vss.n4748 vss.n4747 2172.79
R23063 vss.n4749 vss.n4748 2172.79
R23064 vss.n5527 vss.n4766 2172.79
R23065 vss.n4769 vss.n4766 2172.79
R23066 vss.n5502 vss.n4784 2172.79
R23067 vss.n5501 vss.n4784 2172.79
R23068 vss.n5518 vss.n5517 2172.79
R23069 vss.n5519 vss.n5518 2172.79
R23070 vss.n4791 vss.n4790 2172.79
R23071 vss.n4792 vss.n4791 2172.79
R23072 vss.n5484 vss.n4809 2172.79
R23073 vss.n4812 vss.n4809 2172.79
R23074 vss.n5459 vss.n4827 2172.79
R23075 vss.n5458 vss.n4827 2172.79
R23076 vss.n5475 vss.n5474 2172.79
R23077 vss.n5476 vss.n5475 2172.79
R23078 vss.n4834 vss.n4833 2172.79
R23079 vss.n4835 vss.n4834 2172.79
R23080 vss.n5441 vss.n4852 2172.79
R23081 vss.n4855 vss.n4852 2172.79
R23082 vss.n5416 vss.n4870 2172.79
R23083 vss.n5415 vss.n4870 2172.79
R23084 vss.n5432 vss.n5431 2172.79
R23085 vss.n5433 vss.n5432 2172.79
R23086 vss.n4877 vss.n4876 2172.79
R23087 vss.n4878 vss.n4877 2172.79
R23088 vss.n5398 vss.n5346 2172.79
R23089 vss.n5349 vss.n5346 2172.79
R23090 vss.n5376 vss.n5362 2172.79
R23091 vss.n5389 vss.n5387 2172.79
R23092 vss.n5390 vss.n5389 2172.79
R23093 vss.n5377 vss.n5362 2172.79
R23094 vss.n9820 vss.n2888 2172.79
R23095 vss.n9835 vss.n2878 2172.79
R23096 vss.n9839 vss.n2878 2172.79
R23097 vss.n9826 vss.n2888 2172.79
R23098 vss.n2978 vss.n2936 2172.79
R23099 vss.n2961 vss.n2955 2172.79
R23100 vss.n2965 vss.n2955 2172.79
R23101 vss.n2938 vss.n2936 2172.79
R23102 vss.n2932 vss.n2889 2172.79
R23103 vss.n2914 vss.n2908 2172.79
R23104 vss.n2918 vss.n2908 2172.79
R23105 vss.n2891 vss.n2889 2172.79
R23106 vss.n4940 vss.n4939 2172.79
R23107 vss.n4955 vss.n4929 2172.79
R23108 vss.n4959 vss.n4929 2172.79
R23109 vss.n4946 vss.n4939 2172.79
R23110 vss.n5142 vss.n5141 2172.79
R23111 vss.n5157 vss.n5131 2172.79
R23112 vss.n5161 vss.n5131 2172.79
R23113 vss.n5148 vss.n5141 2172.79
R23114 vss.n3123 vss.n3121 2172.79
R23115 vss.n3138 vss.n3111 2172.79
R23116 vss.n3142 vss.n3111 2172.79
R23117 vss.n3129 vss.n3121 2172.79
R23118 vss.n4484 vss.n4476 2172.79
R23119 vss.n4483 vss.n4476 2172.79
R23120 vss.n4492 vss.n4469 2172.79
R23121 vss.n4496 vss.n4469 2172.79
R23122 vss.n4392 vss.n4384 2172.79
R23123 vss.n4391 vss.n4384 2172.79
R23124 vss.n4400 vss.n4377 2172.79
R23125 vss.n4404 vss.n4377 2172.79
R23126 vss.n4344 vss.n4336 2172.79
R23127 vss.n4343 vss.n4336 2172.79
R23128 vss.n4352 vss.n4329 2172.79
R23129 vss.n4356 vss.n4329 2172.79
R23130 vss.n3744 vss.n3736 2172.79
R23131 vss.n3743 vss.n3736 2172.79
R23132 vss.n3752 vss.n3729 2172.79
R23133 vss.n3756 vss.n3729 2172.79
R23134 vss.n4046 vss.n4038 2172.79
R23135 vss.n4045 vss.n4038 2172.79
R23136 vss.n4054 vss.n4031 2172.79
R23137 vss.n4058 vss.n4031 2172.79
R23138 vss.n3699 vss.n3691 2172.79
R23139 vss.n3698 vss.n3691 2172.79
R23140 vss.n3707 vss.n3684 2172.79
R23141 vss.n3711 vss.n3684 2172.79
R23142 vss.n4100 vss.n4092 2172.79
R23143 vss.n4099 vss.n4092 2172.79
R23144 vss.n4108 vss.n4085 2172.79
R23145 vss.n4112 vss.n4085 2172.79
R23146 vss.n3524 vss.n3516 2172.79
R23147 vss.n3523 vss.n3516 2172.79
R23148 vss.n3532 vss.n3509 2172.79
R23149 vss.n3536 vss.n3509 2172.79
R23150 vss.n3479 vss.n3471 2172.79
R23151 vss.n3478 vss.n3471 2172.79
R23152 vss.n3487 vss.n3464 2172.79
R23153 vss.n3491 vss.n3464 2172.79
R23154 vss.n5767 vss.n5759 2172.79
R23155 vss.n5766 vss.n5759 2172.79
R23156 vss.n5775 vss.n5752 2172.79
R23157 vss.n5779 vss.n5752 2172.79
R23158 vss.n4534 vss.n4445 2172.79
R23159 vss.n4445 vss.n4444 2172.79
R23160 vss.n4526 vss.n4511 2172.79
R23161 vss.n4525 vss.n4511 2172.79
R23162 vss.n4538 vss.n4442 2172.79
R23163 vss.n4539 vss.n4442 2172.79
R23164 vss.n4556 vss.n4555 2172.79
R23165 vss.n4555 vss.n4423 2172.79
R23166 vss.n4591 vss.n4566 2172.79
R23167 vss.n4590 vss.n4566 2172.79
R23168 vss.n4599 vss.n4559 2172.79
R23169 vss.n4603 vss.n4559 2172.79
R23170 vss.n4585 vss.n4570 2172.79
R23171 vss.n4585 vss.n4571 2172.79
R23172 vss.n4626 vss.n3631 2172.79
R23173 vss.n4626 vss.n3632 2172.79
R23174 vss.n4188 vss.n3780 2172.79
R23175 vss.n4187 vss.n3780 2172.79
R23176 vss.n4196 vss.n3773 2172.79
R23177 vss.n4200 vss.n3773 2172.79
R23178 vss.n4182 vss.n3784 2172.79
R23179 vss.n4182 vss.n3785 2172.79
R23180 vss.n3826 vss.n3825 2172.79
R23181 vss.n3825 vss.n3812 2172.79
R23182 vss.n4153 vss.n3836 2172.79
R23183 vss.n4152 vss.n3836 2172.79
R23184 vss.n4161 vss.n3829 2172.79
R23185 vss.n4165 vss.n3829 2172.79
R23186 vss.n4147 vss.n3840 2172.79
R23187 vss.n4147 vss.n3841 2172.79
R23188 vss.n3869 vss.n3868 2172.79
R23189 vss.n3868 vss.n3861 2172.79
R23190 vss.n3938 vss.n3891 2172.79
R23191 vss.n3939 vss.n3891 2172.79
R23192 vss.n4133 vss.n3870 2172.79
R23193 vss.n4133 vss.n3871 2172.79
R23194 vss.n3934 vss.n3892 2172.79
R23195 vss.n3934 vss.n3893 2172.79
R23196 vss.n3920 vss.n3919 2172.79
R23197 vss.n3919 vss.n3912 2172.79
R23198 vss.n5820 vss.n3559 2172.79
R23199 vss.n5819 vss.n3559 2172.79
R23200 vss.n5828 vss.n3552 2172.79
R23201 vss.n5832 vss.n3552 2172.79
R23202 vss.n5814 vss.n3563 2172.79
R23203 vss.n5814 vss.n3564 2172.79
R23204 vss.n3622 vss.n3613 2172.79
R23205 vss.n3622 vss.n3615 2172.79
R23206 vss.n5674 vss.n5661 2172.79
R23207 vss.n5661 vss.n5660 2172.79
R23208 vss.n5800 vss.n3584 2172.79
R23209 vss.n5800 vss.n3585 2172.79
R23210 vss.n5680 vss.n5655 2172.79
R23211 vss.n5679 vss.n5655 2172.79
R23212 vss.n5691 vss.n5690 2172.79
R23213 vss.n5690 vss.n5646 2172.79
R23214 vss.n5715 vss.n5713 2172.79
R23215 vss.n5716 vss.n5713 2172.79
R23216 vss.n5732 vss.n5692 2172.79
R23217 vss.n5732 vss.n5693 2172.79
R23218 vss.n9971 vss.n9963 2172.79
R23219 vss.n9970 vss.n9963 2172.79
R23220 vss.n9979 vss.n9956 2172.79
R23221 vss.n9983 vss.n9956 2172.79
R23222 vss.n2664 vss.n2661 2172.79
R23223 vss.n2665 vss.n2661 2172.79
R23224 vss.n2683 vss.n2640 2172.79
R23225 vss.n2683 vss.n2641 2172.79
R23226 vss.n3404 vss.n3396 2172.79
R23227 vss.n3403 vss.n3396 2172.79
R23228 vss.n3412 vss.n3389 2172.79
R23229 vss.n3416 vss.n3389 2172.79
R23230 vss.n4001 vss.n3993 2172.79
R23231 vss.n4000 vss.n3993 2172.79
R23232 vss.n4009 vss.n3986 2172.79
R23233 vss.n4013 vss.n3986 2172.79
R23234 vss.n4268 vss.n4260 2172.79
R23235 vss.n4267 vss.n4260 2172.79
R23236 vss.n4276 vss.n4253 2172.79
R23237 vss.n4280 vss.n4253 2172.79
R23238 vss.n14064 vss.n493 2172.79
R23239 vss.n14079 vss.n483 2172.79
R23240 vss.n14083 vss.n483 2172.79
R23241 vss.n14070 vss.n493 2172.79
R23242 vss.n10119 vss.n10118 2172.79
R23243 vss.n10134 vss.n10108 2172.79
R23244 vss.n10138 vss.n10108 2172.79
R23245 vss.n10125 vss.n10118 2172.79
R23246 vss.n12877 vss.n12876 2172.79
R23247 vss.n12892 vss.n12866 2172.79
R23248 vss.n12896 vss.n12866 2172.79
R23249 vss.n12883 vss.n12876 2172.79
R23250 vss.n10160 vss.n10159 2172.79
R23251 vss.n10175 vss.n10149 2172.79
R23252 vss.n10179 vss.n10149 2172.79
R23253 vss.n10166 vss.n10159 2172.79
R23254 vss.n12426 vss.n12425 2172.79
R23255 vss.n12441 vss.n12415 2172.79
R23256 vss.n12445 vss.n12415 2172.79
R23257 vss.n12432 vss.n12425 2172.79
R23258 vss.n11755 vss.n11754 2172.79
R23259 vss.n11770 vss.n11744 2172.79
R23260 vss.n11774 vss.n11744 2172.79
R23261 vss.n11761 vss.n11754 2172.79
R23262 vss.n12471 vss.n12470 2172.79
R23263 vss.n12486 vss.n12460 2172.79
R23264 vss.n12490 vss.n12460 2172.79
R23265 vss.n12477 vss.n12470 2172.79
R23266 vss.n2348 vss.n2306 2172.79
R23267 vss.n2331 vss.n2325 2172.79
R23268 vss.n2335 vss.n2325 2172.79
R23269 vss.n2308 vss.n2306 2172.79
R23270 vss.n12296 vss.n12295 2172.79
R23271 vss.n12311 vss.n12285 2172.79
R23272 vss.n12315 vss.n12285 2172.79
R23273 vss.n12302 vss.n12295 2172.79
R23274 vss.n12341 vss.n12340 2172.79
R23275 vss.n12356 vss.n12330 2172.79
R23276 vss.n12360 vss.n12330 2172.79
R23277 vss.n12347 vss.n12340 2172.79
R23278 vss.n10237 vss.n10236 2172.79
R23279 vss.n10252 vss.n10226 2172.79
R23280 vss.n10256 vss.n10226 2172.79
R23281 vss.n10243 vss.n10236 2172.79
R23282 vss.n2417 vss.n2416 2172.79
R23283 vss.n2432 vss.n2406 2172.79
R23284 vss.n2436 vss.n2406 2172.79
R23285 vss.n2423 vss.n2416 2172.79
R23286 vss.n12973 vss.n2366 2172.79
R23287 vss.n2391 vss.n2385 2172.79
R23288 vss.n2395 vss.n2385 2172.79
R23289 vss.n2368 vss.n2366 2172.79
R23290 vss.n10045 vss.n10031 2172.79
R23291 vss.n10046 vss.n10031 2172.79
R23292 vss.n12944 vss.n10055 2172.79
R23293 vss.n10057 vss.n10055 2172.79
R23294 vss.n10040 vss.n10036 2172.79
R23295 vss.n13079 vss.n2115 2172.79
R23296 vss.n2118 vss.n2115 2172.79
R23297 vss.n10040 vss.n10037 2172.79
R23298 vss.n2497 vss.n2495 2172.79
R23299 vss.n2512 vss.n2485 2172.79
R23300 vss.n2516 vss.n2485 2172.79
R23301 vss.n2503 vss.n2495 2172.79
R23302 vss.n12102 vss.n11849 2172.79
R23303 vss.n12121 vss.n11830 2172.79
R23304 vss.n11830 vss.n11827 2172.79
R23305 vss.n12103 vss.n11849 2172.79
R23306 vss.n12151 vss.n11809 2172.79
R23307 vss.n11809 vss.n11808 2172.79
R23308 vss.n12130 vss.n12124 2172.79
R23309 vss.n12134 vss.n12124 2172.79
R23310 vss.n12155 vss.n11805 2172.79
R23311 vss.n12174 vss.n11789 2172.79
R23312 vss.n11789 vss.n11787 2172.79
R23313 vss.n12156 vss.n11805 2172.79
R23314 vss.n12253 vss.n12188 2172.79
R23315 vss.n12253 vss.n12186 2172.79
R23316 vss.n12267 vss.n12177 2172.79
R23317 vss.n12271 vss.n12177 2172.79
R23318 vss.n12249 vss.n12189 2172.79
R23319 vss.n12235 vss.n12208 2172.79
R23320 vss.n12236 vss.n12208 2172.79
R23321 vss.n12191 vss.n12189 2172.79
R23322 vss.n12547 vss.n11721 2172.79
R23323 vss.n11721 vss.n11720 2172.79
R23324 vss.n12225 vss.n12210 2172.79
R23325 vss.n12225 vss.n12211 2172.79
R23326 vss.n12551 vss.n11718 2172.79
R23327 vss.n12570 vss.n11702 2172.79
R23328 vss.n11702 vss.n11700 2172.79
R23329 vss.n12552 vss.n11718 2172.79
R23330 vss.n12585 vss.n11624 2172.79
R23331 vss.n12585 vss.n11625 2172.79
R23332 vss.n12573 vss.n11698 2172.79
R23333 vss.n12574 vss.n12573 2172.79
R23334 vss.n11684 vss.n11640 2172.79
R23335 vss.n11670 vss.n11659 2172.79
R23336 vss.n11671 vss.n11659 2172.79
R23337 vss.n11642 vss.n11640 2172.79
R23338 vss.n12833 vss.n10320 2172.79
R23339 vss.n12833 vss.n10318 2172.79
R23340 vss.n12847 vss.n10309 2172.79
R23341 vss.n12851 vss.n10309 2172.79
R23342 vss.n12829 vss.n12771 2172.79
R23343 vss.n12817 vss.n12790 2172.79
R23344 vss.n12818 vss.n12790 2172.79
R23345 vss.n12773 vss.n12771 2172.79
R23346 vss.n12920 vss.n10086 2172.79
R23347 vss.n10086 vss.n10085 2172.79
R23348 vss.n12807 vss.n12792 2172.79
R23349 vss.n12807 vss.n12793 2172.79
R23350 vss.n11881 vss.n11879 2172.79
R23351 vss.n11882 vss.n11879 2172.79
R23352 vss.n12085 vss.n11858 2172.79
R23353 vss.n12085 vss.n11859 2172.79
R23354 vss.n10483 vss.n10476 2172.79
R23355 vss.n10482 vss.n10476 2172.79
R23356 vss.n10491 vss.n10469 2172.79
R23357 vss.n10495 vss.n10469 2172.79
R23358 vss.n10704 vss.n10697 2172.79
R23359 vss.n10703 vss.n10697 2172.79
R23360 vss.n10712 vss.n10690 2172.79
R23361 vss.n10716 vss.n10690 2172.79
R23362 vss.n11018 vss.n11011 2172.79
R23363 vss.n11017 vss.n11011 2172.79
R23364 vss.n11026 vss.n11004 2172.79
R23365 vss.n11030 vss.n11004 2172.79
R23366 vss.n14051 vss.n512 2054.26
R23367 vss.n13054 vss.n2160 1971.02
R23368 vss.n13114 vss.n2071 1911.25
R23369 vss.n8986 vss.n7332 1870.35
R23370 vss.n8219 vss.n8218 1726.34
R23371 vss.n5642 vss.n5641 1719.18
R23372 vss.n5640 vss.n5639 1719.18
R23373 vss.n5638 vss.n5637 1719.18
R23374 vss.n5636 vss.n5635 1719.18
R23375 vss.n5634 vss.n5633 1719.18
R23376 vss.n5632 vss.n2708 1719.18
R23377 vss.n9048 vss.n9047 1719.18
R23378 vss.n9046 vss.n9045 1719.18
R23379 vss.n9044 vss.n9043 1719.18
R23380 vss.n9042 vss.n9041 1719.18
R23381 vss.n9040 vss.n9039 1719.18
R23382 vss.n9038 vss.n7267 1719.18
R23383 vss.n13924 vss.n13923 1719.18
R23384 vss.n13926 vss.n13925 1719.18
R23385 vss.n13928 vss.n13927 1719.18
R23386 vss.n13930 vss.n13929 1719.18
R23387 vss.n13932 vss.n13931 1719.18
R23388 vss.n13934 vss.n13933 1719.18
R23389 vss.n12035 vss.n11850 1719.18
R23390 vss.n12590 vss.n10614 1719.18
R23391 vss.n12589 vss.n12588 1719.18
R23392 vss.n12587 vss.n10321 1719.18
R23393 vss.n12770 vss.n12769 1719.18
R23394 vss.n12768 vss.n12767 1719.18
R23395 vss.n10001 vss.n10000 1696.62
R23396 vss.n9673 vss.n9672 1569.44
R23397 vss.n12710 vss.n2071 1482.59
R23398 vss.n9703 vss.n2706 1457.22
R23399 vss.n14062 vss.n14061 1438.73
R23400 vss.n14060 vss.n499 1224.92
R23401 vss.n14060 vss.n14059 1224.92
R23402 vss.n14062 vss.n494 1144.63
R23403 vss.n3269 vss.n2743 1122.88
R23404 vss.n481 vss.n442 1122.88
R23405 vss.n10398 vss.n10394 1118.26
R23406 vss.n10403 vss.n10398 1118.26
R23407 vss.n10403 vss.n2040 1118.26
R23408 vss.n13144 vss.n2040 1118.26
R23409 vss.n13144 vss.n2041 1118.26
R23410 vss.n13140 vss.n2041 1118.26
R23411 vss.n10401 vss.n10393 1118.26
R23412 vss.n10402 vss.n10401 1118.26
R23413 vss.n10402 vss.n2035 1118.26
R23414 vss.n13145 vss.n2035 1118.26
R23415 vss.n13145 vss.n2036 1118.26
R23416 vss.n2047 vss.n2036 1118.26
R23417 vss.n12641 vss.n12632 1118.26
R23418 vss.n12645 vss.n12632 1118.26
R23419 vss.n12645 vss.n12629 1118.26
R23420 vss.n12658 vss.n12629 1118.26
R23421 vss.n12658 vss.n12630 1118.26
R23422 vss.n12654 vss.n12630 1118.26
R23423 vss.n12643 vss.n12642 1118.26
R23424 vss.n12644 vss.n12643 1118.26
R23425 vss.n12644 vss.n12624 1118.26
R23426 vss.n12659 vss.n12624 1118.26
R23427 vss.n12659 vss.n12625 1118.26
R23428 vss.n12652 vss.n12625 1118.26
R23429 vss.n11125 vss.n11116 1118.26
R23430 vss.n11129 vss.n11116 1118.26
R23431 vss.n11129 vss.n11113 1118.26
R23432 vss.n11142 vss.n11113 1118.26
R23433 vss.n11142 vss.n11114 1118.26
R23434 vss.n11138 vss.n11114 1118.26
R23435 vss.n11127 vss.n11126 1118.26
R23436 vss.n11128 vss.n11127 1118.26
R23437 vss.n11128 vss.n11108 1118.26
R23438 vss.n11143 vss.n11108 1118.26
R23439 vss.n11143 vss.n11109 1118.26
R23440 vss.n11136 vss.n11109 1118.26
R23441 vss.n12678 vss.n12677 1118.26
R23442 vss.n12679 vss.n12678 1118.26
R23443 vss.n12679 vss.n10377 1118.26
R23444 vss.n12693 vss.n10377 1118.26
R23445 vss.n12693 vss.n10378 1118.26
R23446 vss.n12685 vss.n10378 1118.26
R23447 vss.n12676 vss.n10384 1118.26
R23448 vss.n12680 vss.n10384 1118.26
R23449 vss.n12680 vss.n10386 1118.26
R23450 vss.n10386 vss.n10380 1118.26
R23451 vss.n12690 vss.n10380 1118.26
R23452 vss.n12690 vss.n12689 1118.26
R23453 vss.n11428 vss.n11427 1118.26
R23454 vss.n11429 vss.n11428 1118.26
R23455 vss.n11429 vss.n11408 1118.26
R23456 vss.n11443 vss.n11408 1118.26
R23457 vss.n11443 vss.n11409 1118.26
R23458 vss.n11435 vss.n11409 1118.26
R23459 vss.n11426 vss.n11415 1118.26
R23460 vss.n11430 vss.n11415 1118.26
R23461 vss.n11430 vss.n11417 1118.26
R23462 vss.n11417 vss.n11411 1118.26
R23463 vss.n11440 vss.n11411 1118.26
R23464 vss.n11440 vss.n11439 1118.26
R23465 vss.n11381 vss.n11380 1118.26
R23466 vss.n11382 vss.n11381 1118.26
R23467 vss.n11382 vss.n11361 1118.26
R23468 vss.n11396 vss.n11361 1118.26
R23469 vss.n11396 vss.n11362 1118.26
R23470 vss.n11388 vss.n11362 1118.26
R23471 vss.n11379 vss.n11368 1118.26
R23472 vss.n11383 vss.n11368 1118.26
R23473 vss.n11383 vss.n11370 1118.26
R23474 vss.n11370 vss.n11364 1118.26
R23475 vss.n11393 vss.n11364 1118.26
R23476 vss.n11393 vss.n11392 1118.26
R23477 vss.n10956 vss.n10955 1118.26
R23478 vss.n10957 vss.n10956 1118.26
R23479 vss.n10957 vss.n10936 1118.26
R23480 vss.n10971 vss.n10936 1118.26
R23481 vss.n10971 vss.n10937 1118.26
R23482 vss.n10963 vss.n10937 1118.26
R23483 vss.n10954 vss.n10943 1118.26
R23484 vss.n10958 vss.n10943 1118.26
R23485 vss.n10958 vss.n10945 1118.26
R23486 vss.n10945 vss.n10939 1118.26
R23487 vss.n10968 vss.n10939 1118.26
R23488 vss.n10968 vss.n10967 1118.26
R23489 vss.n10793 vss.n10792 1118.26
R23490 vss.n10794 vss.n10793 1118.26
R23491 vss.n10794 vss.n10773 1118.26
R23492 vss.n10808 vss.n10773 1118.26
R23493 vss.n10808 vss.n10774 1118.26
R23494 vss.n10800 vss.n10774 1118.26
R23495 vss.n10791 vss.n10780 1118.26
R23496 vss.n10795 vss.n10780 1118.26
R23497 vss.n10795 vss.n10782 1118.26
R23498 vss.n10782 vss.n10776 1118.26
R23499 vss.n10805 vss.n10776 1118.26
R23500 vss.n10805 vss.n10804 1118.26
R23501 vss.n10749 vss.n10748 1118.26
R23502 vss.n10750 vss.n10749 1118.26
R23503 vss.n10750 vss.n10729 1118.26
R23504 vss.n10764 vss.n10729 1118.26
R23505 vss.n10764 vss.n10730 1118.26
R23506 vss.n10756 vss.n10730 1118.26
R23507 vss.n10747 vss.n10736 1118.26
R23508 vss.n10751 vss.n10736 1118.26
R23509 vss.n10751 vss.n10738 1118.26
R23510 vss.n10738 vss.n10732 1118.26
R23511 vss.n10761 vss.n10732 1118.26
R23512 vss.n10761 vss.n10760 1118.26
R23513 vss.n11575 vss.n11574 1118.26
R23514 vss.n11576 vss.n11575 1118.26
R23515 vss.n11576 vss.n11555 1118.26
R23516 vss.n11590 vss.n11555 1118.26
R23517 vss.n11590 vss.n11556 1118.26
R23518 vss.n11582 vss.n11556 1118.26
R23519 vss.n11573 vss.n11562 1118.26
R23520 vss.n11577 vss.n11562 1118.26
R23521 vss.n11577 vss.n11564 1118.26
R23522 vss.n11564 vss.n11558 1118.26
R23523 vss.n11587 vss.n11558 1118.26
R23524 vss.n11587 vss.n11586 1118.26
R23525 vss.n10572 vss.n10571 1118.26
R23526 vss.n10573 vss.n10572 1118.26
R23527 vss.n10573 vss.n10552 1118.26
R23528 vss.n10587 vss.n10552 1118.26
R23529 vss.n10587 vss.n10553 1118.26
R23530 vss.n10579 vss.n10553 1118.26
R23531 vss.n10570 vss.n10559 1118.26
R23532 vss.n10574 vss.n10559 1118.26
R23533 vss.n10574 vss.n10561 1118.26
R23534 vss.n10561 vss.n10555 1118.26
R23535 vss.n10584 vss.n10555 1118.26
R23536 vss.n10584 vss.n10583 1118.26
R23537 vss.n10528 vss.n10527 1118.26
R23538 vss.n10529 vss.n10528 1118.26
R23539 vss.n10529 vss.n10508 1118.26
R23540 vss.n10543 vss.n10508 1118.26
R23541 vss.n10543 vss.n10509 1118.26
R23542 vss.n10535 vss.n10509 1118.26
R23543 vss.n10526 vss.n10515 1118.26
R23544 vss.n10530 vss.n10515 1118.26
R23545 vss.n10530 vss.n10517 1118.26
R23546 vss.n10517 vss.n10511 1118.26
R23547 vss.n10540 vss.n10511 1118.26
R23548 vss.n10540 vss.n10539 1118.26
R23549 vss.n11949 vss.n11948 1118.26
R23550 vss.n11950 vss.n11949 1118.26
R23551 vss.n11950 vss.n11929 1118.26
R23552 vss.n11964 vss.n11929 1118.26
R23553 vss.n11964 vss.n11930 1118.26
R23554 vss.n11956 vss.n11930 1118.26
R23555 vss.n11947 vss.n11936 1118.26
R23556 vss.n11951 vss.n11936 1118.26
R23557 vss.n11951 vss.n11938 1118.26
R23558 vss.n11938 vss.n11932 1118.26
R23559 vss.n11961 vss.n11932 1118.26
R23560 vss.n11961 vss.n11960 1118.26
R23561 vss.n12064 vss.n11899 1118.26
R23562 vss.n12068 vss.n11899 1118.26
R23563 vss.n12068 vss.n11856 1118.26
R23564 vss.n12091 vss.n11856 1118.26
R23565 vss.n12091 vss.n12090 1118.26
R23566 vss.n12090 vss.n11852 1118.26
R23567 vss.n12063 vss.n11896 1118.26
R23568 vss.n12069 vss.n11896 1118.26
R23569 vss.n12070 vss.n12069 1118.26
R23570 vss.n12071 vss.n12070 1118.26
R23571 vss.n12071 vss.n11857 1118.26
R23572 vss.n11857 vss.n11851 1118.26
R23573 vss.n11911 vss.n11905 1118.26
R23574 vss.n12053 vss.n11905 1118.26
R23575 vss.n12053 vss.n12052 1118.26
R23576 vss.n12052 vss.n12051 1118.26
R23577 vss.n12051 vss.n11916 1118.26
R23578 vss.n12047 vss.n11916 1118.26
R23579 vss.n11909 vss.n11904 1118.26
R23580 vss.n11974 vss.n11904 1118.26
R23581 vss.n11975 vss.n11974 1118.26
R23582 vss.n11976 vss.n11975 1118.26
R23583 vss.n11976 vss.n11921 1118.26
R23584 vss.n11980 vss.n11921 1118.26
R23585 vss.n12024 vss.n11986 1118.26
R23586 vss.n12028 vss.n11986 1118.26
R23587 vss.n12029 vss.n12028 1118.26
R23588 vss.n12030 vss.n12029 1118.26
R23589 vss.n12030 vss.n11982 1118.26
R23590 vss.n12038 vss.n11982 1118.26
R23591 vss.n12023 vss.n12011 1118.26
R23592 vss.n12019 vss.n12011 1118.26
R23593 vss.n12019 vss.n12018 1118.26
R23594 vss.n12018 vss.n12017 1118.26
R23595 vss.n12017 vss.n11981 1118.26
R23596 vss.n12034 vss.n11981 1118.26
R23597 vss.n11999 vss.n11993 1118.26
R23598 vss.n12001 vss.n11993 1118.26
R23599 vss.n12001 vss.n10599 1118.26
R23600 vss.n12606 vss.n10599 1118.26
R23601 vss.n12606 vss.n10600 1118.26
R23602 vss.n12602 vss.n10600 1118.26
R23603 vss.n11997 vss.n11992 1118.26
R23604 vss.n11992 vss.n11991 1118.26
R23605 vss.n11991 vss.n10594 1118.26
R23606 vss.n12607 vss.n10594 1118.26
R23607 vss.n12607 vss.n10595 1118.26
R23608 vss.n10606 vss.n10595 1118.26
R23609 vss.n10648 vss.n10644 1118.26
R23610 vss.n10664 vss.n10648 1118.26
R23611 vss.n10664 vss.n10663 1118.26
R23612 vss.n10663 vss.n10662 1118.26
R23613 vss.n10662 vss.n10608 1118.26
R23614 vss.n12593 vss.n10608 1118.26
R23615 vss.n10653 vss.n10643 1118.26
R23616 vss.n10654 vss.n10653 1118.26
R23617 vss.n10654 vss.n10649 1118.26
R23618 vss.n10656 vss.n10649 1118.26
R23619 vss.n10656 vss.n10607 1118.26
R23620 vss.n10613 vss.n10607 1118.26
R23621 vss.n10672 vss.n10636 1118.26
R23622 vss.n10676 vss.n10636 1118.26
R23623 vss.n10676 vss.n10628 1118.26
R23624 vss.n11606 vss.n10628 1118.26
R23625 vss.n11606 vss.n11605 1118.26
R23626 vss.n11605 vss.n10624 1118.26
R23627 vss.n10642 vss.n10632 1118.26
R23628 vss.n10677 vss.n10632 1118.26
R23629 vss.n10677 vss.n10629 1118.26
R23630 vss.n11601 vss.n10629 1118.26
R23631 vss.n11602 vss.n11601 1118.26
R23632 vss.n11602 vss.n10623 1118.26
R23633 vss.n10834 vss.n10831 1118.26
R23634 vss.n10851 vss.n10834 1118.26
R23635 vss.n10851 vss.n10621 1118.26
R23636 vss.n11617 vss.n10621 1118.26
R23637 vss.n11617 vss.n11616 1118.26
R23638 vss.n11616 vss.n10617 1118.26
R23639 vss.n10838 vss.n10830 1118.26
R23640 vss.n10850 vss.n10838 1118.26
R23641 vss.n10850 vss.n10839 1118.26
R23642 vss.n10846 vss.n10839 1118.26
R23643 vss.n10846 vss.n10622 1118.26
R23644 vss.n10622 vss.n10616 1118.26
R23645 vss.n10861 vss.n10823 1118.26
R23646 vss.n10865 vss.n10823 1118.26
R23647 vss.n10865 vss.n10820 1118.26
R23648 vss.n11535 vss.n10820 1118.26
R23649 vss.n11535 vss.n10821 1118.26
R23650 vss.n11531 vss.n10821 1118.26
R23651 vss.n10863 vss.n10862 1118.26
R23652 vss.n10864 vss.n10863 1118.26
R23653 vss.n10864 vss.n10815 1118.26
R23654 vss.n11536 vss.n10815 1118.26
R23655 vss.n11536 vss.n10816 1118.26
R23656 vss.n10872 vss.n10816 1118.26
R23657 vss.n11509 vss.n10878 1118.26
R23658 vss.n11513 vss.n10878 1118.26
R23659 vss.n11514 vss.n11513 1118.26
R23660 vss.n11515 vss.n11514 1118.26
R23661 vss.n11515 vss.n10874 1118.26
R23662 vss.n11522 vss.n10874 1118.26
R23663 vss.n11508 vss.n11498 1118.26
R23664 vss.n11504 vss.n11498 1118.26
R23665 vss.n11504 vss.n11503 1118.26
R23666 vss.n11503 vss.n11502 1118.26
R23667 vss.n11502 vss.n10873 1118.26
R23668 vss.n11519 vss.n10873 1118.26
R23669 vss.n10890 vss.n10884 1118.26
R23670 vss.n11488 vss.n10884 1118.26
R23671 vss.n11488 vss.n11487 1118.26
R23672 vss.n11487 vss.n11486 1118.26
R23673 vss.n11486 vss.n10895 1118.26
R23674 vss.n11482 vss.n10895 1118.26
R23675 vss.n10888 vss.n10883 1118.26
R23676 vss.n10980 vss.n10883 1118.26
R23677 vss.n10981 vss.n10980 1118.26
R23678 vss.n10985 vss.n10981 1118.26
R23679 vss.n10985 vss.n10984 1118.26
R23680 vss.n10984 vss.n10898 1118.26
R23681 vss.n11461 vss.n10904 1118.26
R23682 vss.n11465 vss.n10904 1118.26
R23683 vss.n11466 vss.n11465 1118.26
R23684 vss.n11467 vss.n11466 1118.26
R23685 vss.n11467 vss.n10900 1118.26
R23686 vss.n11473 vss.n10900 1118.26
R23687 vss.n11460 vss.n10931 1118.26
R23688 vss.n11456 vss.n10931 1118.26
R23689 vss.n11456 vss.n11455 1118.26
R23690 vss.n11455 vss.n11454 1118.26
R23691 vss.n11454 vss.n10899 1118.26
R23692 vss.n11471 vss.n10899 1118.26
R23693 vss.n10919 vss.n10913 1118.26
R23694 vss.n10921 vss.n10913 1118.26
R23695 vss.n10921 vss.n10335 1118.26
R23696 vss.n12749 vss.n10335 1118.26
R23697 vss.n12749 vss.n12748 1118.26
R23698 vss.n12748 vss.n10331 1118.26
R23699 vss.n10917 vss.n10912 1118.26
R23700 vss.n10912 vss.n10911 1118.26
R23701 vss.n10911 vss.n10336 1118.26
R23702 vss.n12744 vss.n10336 1118.26
R23703 vss.n12745 vss.n12744 1118.26
R23704 vss.n12745 vss.n10330 1118.26
R23705 vss.n12729 vss.n10348 1118.26
R23706 vss.n12733 vss.n10348 1118.26
R23707 vss.n12733 vss.n10328 1118.26
R23708 vss.n12760 vss.n10328 1118.26
R23709 vss.n12760 vss.n12759 1118.26
R23710 vss.n12759 vss.n10324 1118.26
R23711 vss.n12728 vss.n10345 1118.26
R23712 vss.n12734 vss.n10345 1118.26
R23713 vss.n12735 vss.n12734 1118.26
R23714 vss.n12736 vss.n12735 1118.26
R23715 vss.n12736 vss.n10329 1118.26
R23716 vss.n10329 vss.n10323 1118.26
R23717 vss.n10360 vss.n10354 1118.26
R23718 vss.n12718 vss.n10354 1118.26
R23719 vss.n12718 vss.n12717 1118.26
R23720 vss.n12717 vss.n12716 1118.26
R23721 vss.n12716 vss.n10365 1118.26
R23722 vss.n12712 vss.n10365 1118.26
R23723 vss.n10358 vss.n10353 1118.26
R23724 vss.n12703 vss.n10353 1118.26
R23725 vss.n12704 vss.n12703 1118.26
R23726 vss.n12705 vss.n12704 1118.26
R23727 vss.n12705 vss.n10370 1118.26
R23728 vss.n12709 vss.n10370 1118.26
R23729 vss.n2083 vss.n2073 1118.26
R23730 vss.n13105 vss.n2083 1118.26
R23731 vss.n13105 vss.n2084 1118.26
R23732 vss.n13101 vss.n2084 1118.26
R23733 vss.n13101 vss.n2089 1118.26
R23734 vss.n2095 vss.n2089 1118.26
R23735 vss.n2078 vss.n2074 1118.26
R23736 vss.n13106 vss.n2078 1118.26
R23737 vss.n13106 vss.n2079 1118.26
R23738 vss.n2090 vss.n2079 1118.26
R23739 vss.n2091 vss.n2090 1118.26
R23740 vss.n13095 vss.n2091 1118.26
R23741 vss.n12924 vss.n10076 1118.26
R23742 vss.n12930 vss.n10076 1118.26
R23743 vss.n12930 vss.n10072 1118.26
R23744 vss.n12934 vss.n10072 1118.26
R23745 vss.n12934 vss.n10060 1118.26
R23746 vss.n12941 vss.n10060 1118.26
R23747 vss.n12925 vss.n10078 1118.26
R23748 vss.n12929 vss.n10078 1118.26
R23749 vss.n12929 vss.n10068 1118.26
R23750 vss.n12935 vss.n10068 1118.26
R23751 vss.n12935 vss.n10070 1118.26
R23752 vss.n10070 vss.n10059 1118.26
R23753 vss.n12997 vss.n2252 1118.26
R23754 vss.n13001 vss.n2252 1118.26
R23755 vss.n13001 vss.n2249 1118.26
R23756 vss.n13014 vss.n2249 1118.26
R23757 vss.n13014 vss.n2250 1118.26
R23758 vss.n13010 vss.n2250 1118.26
R23759 vss.n12999 vss.n12998 1118.26
R23760 vss.n13000 vss.n12999 1118.26
R23761 vss.n13000 vss.n2244 1118.26
R23762 vss.n13015 vss.n2244 1118.26
R23763 vss.n13015 vss.n2245 1118.26
R23764 vss.n13009 vss.n2245 1118.26
R23765 vss.n2272 vss.n2259 1118.26
R23766 vss.n2296 vss.n2272 1118.26
R23767 vss.n2296 vss.n2273 1118.26
R23768 vss.n2292 vss.n2273 1118.26
R23769 vss.n2292 vss.n2278 1118.26
R23770 vss.n2284 vss.n2278 1118.26
R23771 vss.n2267 vss.n2260 1118.26
R23772 vss.n2297 vss.n2267 1118.26
R23773 vss.n2297 vss.n2268 1118.26
R23774 vss.n2279 vss.n2268 1118.26
R23775 vss.n2280 vss.n2279 1118.26
R23776 vss.n2286 vss.n2280 1118.26
R23777 vss.n2130 vss.n2120 1118.26
R23778 vss.n13069 vss.n2130 1118.26
R23779 vss.n13069 vss.n2131 1118.26
R23780 vss.n13065 vss.n2131 1118.26
R23781 vss.n13065 vss.n2136 1118.26
R23782 vss.n2142 vss.n2136 1118.26
R23783 vss.n2125 vss.n2121 1118.26
R23784 vss.n13070 vss.n2125 1118.26
R23785 vss.n13070 vss.n2126 1118.26
R23786 vss.n2137 vss.n2126 1118.26
R23787 vss.n2138 vss.n2137 1118.26
R23788 vss.n13059 vss.n2138 1118.26
R23789 vss.n14157 vss.n450 1118.26
R23790 vss.n14163 vss.n450 1118.26
R23791 vss.n14163 vss.n443 1118.26
R23792 vss.n14168 vss.n443 1118.26
R23793 vss.n14168 vss.n446 1118.26
R23794 vss.n446 vss.n434 1118.26
R23795 vss.n14158 vss.n452 1118.26
R23796 vss.n14162 vss.n452 1118.26
R23797 vss.n14162 vss.n439 1118.26
R23798 vss.n14169 vss.n439 1118.26
R23799 vss.n14169 vss.n440 1118.26
R23800 vss.n440 vss.n435 1118.26
R23801 vss.n634 vss.n627 1118.26
R23802 vss.n638 vss.n627 1118.26
R23803 vss.n638 vss.n619 1118.26
R23804 vss.n652 vss.n619 1118.26
R23805 vss.n652 vss.n651 1118.26
R23806 vss.n651 vss.n615 1118.26
R23807 vss.n633 vss.n623 1118.26
R23808 vss.n639 vss.n623 1118.26
R23809 vss.n639 vss.n620 1118.26
R23810 vss.n647 vss.n620 1118.26
R23811 vss.n648 vss.n647 1118.26
R23812 vss.n648 vss.n614 1118.26
R23813 vss.n2005 vss.n1996 1118.26
R23814 vss.n2009 vss.n1996 1118.26
R23815 vss.n2009 vss.n1993 1118.26
R23816 vss.n2022 vss.n1993 1118.26
R23817 vss.n2022 vss.n1994 1118.26
R23818 vss.n2018 vss.n1994 1118.26
R23819 vss.n2007 vss.n2006 1118.26
R23820 vss.n2008 vss.n2007 1118.26
R23821 vss.n2008 vss.n1988 1118.26
R23822 vss.n2023 vss.n1988 1118.26
R23823 vss.n2023 vss.n1989 1118.26
R23824 vss.n2016 vss.n1989 1118.26
R23825 vss.n1070 vss.n1061 1118.26
R23826 vss.n1074 vss.n1061 1118.26
R23827 vss.n1074 vss.n1058 1118.26
R23828 vss.n1087 vss.n1058 1118.26
R23829 vss.n1087 vss.n1059 1118.26
R23830 vss.n1083 vss.n1059 1118.26
R23831 vss.n1072 vss.n1071 1118.26
R23832 vss.n1073 vss.n1072 1118.26
R23833 vss.n1073 vss.n1053 1118.26
R23834 vss.n1088 vss.n1053 1118.26
R23835 vss.n1088 vss.n1054 1118.26
R23836 vss.n1081 vss.n1054 1118.26
R23837 vss.n1331 vss.n1322 1118.26
R23838 vss.n1335 vss.n1322 1118.26
R23839 vss.n1335 vss.n1319 1118.26
R23840 vss.n1348 vss.n1319 1118.26
R23841 vss.n1348 vss.n1320 1118.26
R23842 vss.n1344 vss.n1320 1118.26
R23843 vss.n1333 vss.n1332 1118.26
R23844 vss.n1334 vss.n1333 1118.26
R23845 vss.n1334 vss.n1314 1118.26
R23846 vss.n1349 vss.n1314 1118.26
R23847 vss.n1349 vss.n1315 1118.26
R23848 vss.n1342 vss.n1315 1118.26
R23849 vss.n1463 vss.n1454 1118.26
R23850 vss.n1467 vss.n1454 1118.26
R23851 vss.n1467 vss.n1451 1118.26
R23852 vss.n1480 vss.n1451 1118.26
R23853 vss.n1480 vss.n1452 1118.26
R23854 vss.n1476 vss.n1452 1118.26
R23855 vss.n1465 vss.n1464 1118.26
R23856 vss.n1466 vss.n1465 1118.26
R23857 vss.n1466 vss.n1446 1118.26
R23858 vss.n1481 vss.n1446 1118.26
R23859 vss.n1481 vss.n1447 1118.26
R23860 vss.n1474 vss.n1447 1118.26
R23861 vss.n1626 vss.n1617 1118.26
R23862 vss.n1630 vss.n1617 1118.26
R23863 vss.n1630 vss.n1614 1118.26
R23864 vss.n1643 vss.n1614 1118.26
R23865 vss.n1643 vss.n1615 1118.26
R23866 vss.n1639 vss.n1615 1118.26
R23867 vss.n1628 vss.n1627 1118.26
R23868 vss.n1629 vss.n1628 1118.26
R23869 vss.n1629 vss.n1609 1118.26
R23870 vss.n1644 vss.n1609 1118.26
R23871 vss.n1644 vss.n1610 1118.26
R23872 vss.n1637 vss.n1610 1118.26
R23873 vss.n1543 vss.n1534 1118.26
R23874 vss.n1547 vss.n1534 1118.26
R23875 vss.n1547 vss.n1531 1118.26
R23876 vss.n1561 vss.n1531 1118.26
R23877 vss.n1561 vss.n1532 1118.26
R23878 vss.n1557 vss.n1532 1118.26
R23879 vss.n1545 vss.n1544 1118.26
R23880 vss.n1546 vss.n1545 1118.26
R23881 vss.n1546 vss.n1526 1118.26
R23882 vss.n1562 vss.n1526 1118.26
R23883 vss.n1562 vss.n1527 1118.26
R23884 vss.n1554 vss.n1527 1118.26
R23885 vss.n880 vss.n876 1118.26
R23886 vss.n912 vss.n880 1118.26
R23887 vss.n912 vss.n911 1118.26
R23888 vss.n911 vss.n910 1118.26
R23889 vss.n910 vss.n883 1118.26
R23890 vss.n906 vss.n883 1118.26
R23891 vss.n895 vss.n875 1118.26
R23892 vss.n898 vss.n895 1118.26
R23893 vss.n899 vss.n898 1118.26
R23894 vss.n900 vss.n899 1118.26
R23895 vss.n900 vss.n888 1118.26
R23896 vss.n904 vss.n888 1118.26
R23897 vss.n839 vss.n835 1118.26
R23898 vss.n868 vss.n839 1118.26
R23899 vss.n868 vss.n867 1118.26
R23900 vss.n867 vss.n866 1118.26
R23901 vss.n866 vss.n843 1118.26
R23902 vss.n862 vss.n843 1118.26
R23903 vss.n851 vss.n834 1118.26
R23904 vss.n854 vss.n851 1118.26
R23905 vss.n855 vss.n854 1118.26
R23906 vss.n856 vss.n855 1118.26
R23907 vss.n856 vss.n848 1118.26
R23908 vss.n860 vss.n848 1118.26
R23909 vss.n822 vss.n818 1118.26
R23910 vss.n827 vss.n822 1118.26
R23911 vss.n827 vss.n603 1118.26
R23912 vss.n13949 vss.n603 1118.26
R23913 vss.n13949 vss.n604 1118.26
R23914 vss.n13945 vss.n604 1118.26
R23915 vss.n825 vss.n817 1118.26
R23916 vss.n826 vss.n825 1118.26
R23917 vss.n826 vss.n598 1118.26
R23918 vss.n13950 vss.n598 1118.26
R23919 vss.n13950 vss.n599 1118.26
R23920 vss.n610 vss.n599 1118.26
R23921 vss.n13214 vss.n805 1118.26
R23922 vss.n13218 vss.n805 1118.26
R23923 vss.n13218 vss.n802 1118.26
R23924 vss.n13231 vss.n802 1118.26
R23925 vss.n13231 vss.n803 1118.26
R23926 vss.n13227 vss.n803 1118.26
R23927 vss.n13216 vss.n13215 1118.26
R23928 vss.n13217 vss.n13216 1118.26
R23929 vss.n13217 vss.n797 1118.26
R23930 vss.n13232 vss.n797 1118.26
R23931 vss.n13232 vss.n798 1118.26
R23932 vss.n13225 vss.n798 1118.26
R23933 vss.n1673 vss.n1664 1118.26
R23934 vss.n1677 vss.n1664 1118.26
R23935 vss.n1677 vss.n1661 1118.26
R23936 vss.n1690 vss.n1661 1118.26
R23937 vss.n1690 vss.n1662 1118.26
R23938 vss.n1686 vss.n1662 1118.26
R23939 vss.n1675 vss.n1674 1118.26
R23940 vss.n1676 vss.n1675 1118.26
R23941 vss.n1676 vss.n1656 1118.26
R23942 vss.n1691 vss.n1656 1118.26
R23943 vss.n1691 vss.n1657 1118.26
R23944 vss.n1684 vss.n1657 1118.26
R23945 vss.n1378 vss.n1369 1118.26
R23946 vss.n1382 vss.n1369 1118.26
R23947 vss.n1382 vss.n1366 1118.26
R23948 vss.n1395 vss.n1366 1118.26
R23949 vss.n1395 vss.n1367 1118.26
R23950 vss.n1391 vss.n1367 1118.26
R23951 vss.n1380 vss.n1379 1118.26
R23952 vss.n1381 vss.n1380 1118.26
R23953 vss.n1381 vss.n1361 1118.26
R23954 vss.n1396 vss.n1361 1118.26
R23955 vss.n1396 vss.n1362 1118.26
R23956 vss.n1389 vss.n1362 1118.26
R23957 vss.n1179 vss.n1170 1118.26
R23958 vss.n1183 vss.n1170 1118.26
R23959 vss.n1183 vss.n1167 1118.26
R23960 vss.n1196 vss.n1167 1118.26
R23961 vss.n1196 vss.n1168 1118.26
R23962 vss.n1192 vss.n1168 1118.26
R23963 vss.n1181 vss.n1180 1118.26
R23964 vss.n1182 vss.n1181 1118.26
R23965 vss.n1182 vss.n1162 1118.26
R23966 vss.n1197 vss.n1162 1118.26
R23967 vss.n1197 vss.n1163 1118.26
R23968 vss.n1190 vss.n1163 1118.26
R23969 vss.n1115 vss.n1106 1118.26
R23970 vss.n1119 vss.n1106 1118.26
R23971 vss.n1119 vss.n1103 1118.26
R23972 vss.n1132 vss.n1103 1118.26
R23973 vss.n1132 vss.n1104 1118.26
R23974 vss.n1128 vss.n1104 1118.26
R23975 vss.n1117 vss.n1116 1118.26
R23976 vss.n1118 vss.n1117 1118.26
R23977 vss.n1118 vss.n1098 1118.26
R23978 vss.n1133 vss.n1098 1118.26
R23979 vss.n1133 vss.n1099 1118.26
R23980 vss.n1126 vss.n1099 1118.26
R23981 vss.n13181 vss.n13180 1118.26
R23982 vss.n13182 vss.n13181 1118.26
R23983 vss.n13182 vss.n13162 1118.26
R23984 vss.n13197 vss.n13162 1118.26
R23985 vss.n13197 vss.n13163 1118.26
R23986 vss.n13189 vss.n13163 1118.26
R23987 vss.n13179 vss.n13168 1118.26
R23988 vss.n13183 vss.n13168 1118.26
R23989 vss.n13183 vss.n13170 1118.26
R23990 vss.n13170 vss.n13165 1118.26
R23991 vss.n13166 vss.n13165 1118.26
R23992 vss.n13191 vss.n13166 1118.26
R23993 vss.n177 vss.n173 1118.26
R23994 vss.n181 vss.n177 1118.26
R23995 vss.n181 vss.n9 1118.26
R23996 vss.n14789 vss.n9 1118.26
R23997 vss.n14789 vss.n10 1118.26
R23998 vss.n14785 vss.n10 1118.26
R23999 vss.n178 vss.n174 1118.26
R24000 vss.n179 vss.n178 1118.26
R24001 vss.n179 vss.n4 1118.26
R24002 vss.n14790 vss.n4 1118.26
R24003 vss.n14790 vss.n5 1118.26
R24004 vss.n17 vss.n5 1118.26
R24005 vss.n14698 vss.n14686 1118.26
R24006 vss.n14722 vss.n14698 1118.26
R24007 vss.n14722 vss.n14699 1118.26
R24008 vss.n14718 vss.n14699 1118.26
R24009 vss.n14718 vss.n14704 1118.26
R24010 vss.n14710 vss.n14704 1118.26
R24011 vss.n14693 vss.n14687 1118.26
R24012 vss.n14723 vss.n14693 1118.26
R24013 vss.n14723 vss.n14694 1118.26
R24014 vss.n14705 vss.n14694 1118.26
R24015 vss.n14706 vss.n14705 1118.26
R24016 vss.n14712 vss.n14706 1118.26
R24017 vss.n14586 vss.n14576 1118.26
R24018 vss.n14590 vss.n14576 1118.26
R24019 vss.n14590 vss.n14573 1118.26
R24020 vss.n14603 vss.n14573 1118.26
R24021 vss.n14603 vss.n14574 1118.26
R24022 vss.n14599 vss.n14574 1118.26
R24023 vss.n14588 vss.n14587 1118.26
R24024 vss.n14589 vss.n14588 1118.26
R24025 vss.n14589 vss.n14568 1118.26
R24026 vss.n14604 vss.n14568 1118.26
R24027 vss.n14604 vss.n14569 1118.26
R24028 vss.n14598 vss.n14569 1118.26
R24029 vss.n14503 vss.n14491 1118.26
R24030 vss.n14527 vss.n14503 1118.26
R24031 vss.n14527 vss.n14504 1118.26
R24032 vss.n14523 vss.n14504 1118.26
R24033 vss.n14523 vss.n14509 1118.26
R24034 vss.n14515 vss.n14509 1118.26
R24035 vss.n14498 vss.n14492 1118.26
R24036 vss.n14528 vss.n14498 1118.26
R24037 vss.n14528 vss.n14499 1118.26
R24038 vss.n14510 vss.n14499 1118.26
R24039 vss.n14511 vss.n14510 1118.26
R24040 vss.n14517 vss.n14511 1118.26
R24041 vss.n14391 vss.n14381 1118.26
R24042 vss.n14395 vss.n14381 1118.26
R24043 vss.n14395 vss.n14378 1118.26
R24044 vss.n14408 vss.n14378 1118.26
R24045 vss.n14408 vss.n14379 1118.26
R24046 vss.n14404 vss.n14379 1118.26
R24047 vss.n14393 vss.n14392 1118.26
R24048 vss.n14394 vss.n14393 1118.26
R24049 vss.n14394 vss.n14373 1118.26
R24050 vss.n14409 vss.n14373 1118.26
R24051 vss.n14409 vss.n14374 1118.26
R24052 vss.n14403 vss.n14374 1118.26
R24053 vss.n14308 vss.n14296 1118.26
R24054 vss.n14332 vss.n14308 1118.26
R24055 vss.n14332 vss.n14309 1118.26
R24056 vss.n14328 vss.n14309 1118.26
R24057 vss.n14328 vss.n14314 1118.26
R24058 vss.n14320 vss.n14314 1118.26
R24059 vss.n14303 vss.n14297 1118.26
R24060 vss.n14333 vss.n14303 1118.26
R24061 vss.n14333 vss.n14304 1118.26
R24062 vss.n14315 vss.n14304 1118.26
R24063 vss.n14316 vss.n14315 1118.26
R24064 vss.n14322 vss.n14316 1118.26
R24065 vss.n338 vss.n328 1118.26
R24066 vss.n342 vss.n328 1118.26
R24067 vss.n342 vss.n325 1118.26
R24068 vss.n355 vss.n325 1118.26
R24069 vss.n355 vss.n326 1118.26
R24070 vss.n351 vss.n326 1118.26
R24071 vss.n340 vss.n339 1118.26
R24072 vss.n341 vss.n340 1118.26
R24073 vss.n341 vss.n320 1118.26
R24074 vss.n356 vss.n320 1118.26
R24075 vss.n356 vss.n321 1118.26
R24076 vss.n350 vss.n321 1118.26
R24077 vss.n14189 vss.n14177 1118.26
R24078 vss.n14213 vss.n14189 1118.26
R24079 vss.n14213 vss.n14190 1118.26
R24080 vss.n14209 vss.n14190 1118.26
R24081 vss.n14209 vss.n14195 1118.26
R24082 vss.n14201 vss.n14195 1118.26
R24083 vss.n14184 vss.n14178 1118.26
R24084 vss.n14214 vss.n14184 1118.26
R24085 vss.n14214 vss.n14185 1118.26
R24086 vss.n14196 vss.n14185 1118.26
R24087 vss.n14197 vss.n14196 1118.26
R24088 vss.n14203 vss.n14197 1118.26
R24089 vss.n14117 vss.n14107 1118.26
R24090 vss.n14121 vss.n14107 1118.26
R24091 vss.n14121 vss.n14104 1118.26
R24092 vss.n14134 vss.n14104 1118.26
R24093 vss.n14134 vss.n14105 1118.26
R24094 vss.n14130 vss.n14105 1118.26
R24095 vss.n14119 vss.n14118 1118.26
R24096 vss.n14120 vss.n14119 1118.26
R24097 vss.n14120 vss.n14099 1118.26
R24098 vss.n14135 vss.n14099 1118.26
R24099 vss.n14135 vss.n14100 1118.26
R24100 vss.n14129 vss.n14100 1118.26
R24101 vss.n14226 vss.n425 1118.26
R24102 vss.n14230 vss.n425 1118.26
R24103 vss.n14230 vss.n422 1118.26
R24104 vss.n14243 vss.n422 1118.26
R24105 vss.n14243 vss.n423 1118.26
R24106 vss.n14239 vss.n423 1118.26
R24107 vss.n14228 vss.n14227 1118.26
R24108 vss.n14229 vss.n14228 1118.26
R24109 vss.n14229 vss.n417 1118.26
R24110 vss.n14244 vss.n417 1118.26
R24111 vss.n14244 vss.n418 1118.26
R24112 vss.n14238 vss.n418 1118.26
R24113 vss.n14262 vss.n312 1118.26
R24114 vss.n14286 vss.n14262 1118.26
R24115 vss.n14286 vss.n14263 1118.26
R24116 vss.n14282 vss.n14263 1118.26
R24117 vss.n14282 vss.n14268 1118.26
R24118 vss.n14274 vss.n14268 1118.26
R24119 vss.n14257 vss.n313 1118.26
R24120 vss.n14287 vss.n14257 1118.26
R24121 vss.n14287 vss.n14258 1118.26
R24122 vss.n14269 vss.n14258 1118.26
R24123 vss.n14270 vss.n14269 1118.26
R24124 vss.n14276 vss.n14270 1118.26
R24125 vss.n14345 vss.n302 1118.26
R24126 vss.n14349 vss.n302 1118.26
R24127 vss.n14349 vss.n299 1118.26
R24128 vss.n14362 vss.n299 1118.26
R24129 vss.n14362 vss.n300 1118.26
R24130 vss.n14358 vss.n300 1118.26
R24131 vss.n14347 vss.n14346 1118.26
R24132 vss.n14348 vss.n14347 1118.26
R24133 vss.n14348 vss.n294 1118.26
R24134 vss.n14363 vss.n294 1118.26
R24135 vss.n14363 vss.n295 1118.26
R24136 vss.n14357 vss.n295 1118.26
R24137 vss.n14457 vss.n253 1118.26
R24138 vss.n14481 vss.n14457 1118.26
R24139 vss.n14481 vss.n14458 1118.26
R24140 vss.n14477 vss.n14458 1118.26
R24141 vss.n14477 vss.n14463 1118.26
R24142 vss.n14469 vss.n14463 1118.26
R24143 vss.n14452 vss.n254 1118.26
R24144 vss.n14482 vss.n14452 1118.26
R24145 vss.n14482 vss.n14453 1118.26
R24146 vss.n14464 vss.n14453 1118.26
R24147 vss.n14465 vss.n14464 1118.26
R24148 vss.n14471 vss.n14465 1118.26
R24149 vss.n14540 vss.n243 1118.26
R24150 vss.n14544 vss.n243 1118.26
R24151 vss.n14544 vss.n240 1118.26
R24152 vss.n14557 vss.n240 1118.26
R24153 vss.n14557 vss.n241 1118.26
R24154 vss.n14553 vss.n241 1118.26
R24155 vss.n14542 vss.n14541 1118.26
R24156 vss.n14543 vss.n14542 1118.26
R24157 vss.n14543 vss.n235 1118.26
R24158 vss.n14558 vss.n235 1118.26
R24159 vss.n14558 vss.n236 1118.26
R24160 vss.n14552 vss.n236 1118.26
R24161 vss.n14652 vss.n194 1118.26
R24162 vss.n14676 vss.n14652 1118.26
R24163 vss.n14676 vss.n14653 1118.26
R24164 vss.n14672 vss.n14653 1118.26
R24165 vss.n14672 vss.n14658 1118.26
R24166 vss.n14664 vss.n14658 1118.26
R24167 vss.n14647 vss.n195 1118.26
R24168 vss.n14677 vss.n14647 1118.26
R24169 vss.n14677 vss.n14648 1118.26
R24170 vss.n14659 vss.n14648 1118.26
R24171 vss.n14660 vss.n14659 1118.26
R24172 vss.n14666 vss.n14660 1118.26
R24173 vss.n14735 vss.n166 1118.26
R24174 vss.n14739 vss.n166 1118.26
R24175 vss.n14739 vss.n163 1118.26
R24176 vss.n14752 vss.n163 1118.26
R24177 vss.n14752 vss.n164 1118.26
R24178 vss.n14748 vss.n164 1118.26
R24179 vss.n14737 vss.n14736 1118.26
R24180 vss.n14738 vss.n14737 1118.26
R24181 vss.n14738 vss.n158 1118.26
R24182 vss.n14753 vss.n158 1118.26
R24183 vss.n14753 vss.n159 1118.26
R24184 vss.n14747 vss.n159 1118.26
R24185 vss.n14153 vss.n461 1118.26
R24186 vss.n14149 vss.n461 1118.26
R24187 vss.n14149 vss.n465 1118.26
R24188 vss.n13574 vss.n465 1118.26
R24189 vss.n13574 vss.n13570 1118.26
R24190 vss.n13570 vss.n13566 1118.26
R24191 vss.n468 vss.n459 1118.26
R24192 vss.n14148 vss.n468 1118.26
R24193 vss.n14148 vss.n469 1118.26
R24194 vss.n13572 vss.n469 1118.26
R24195 vss.n13572 vss.n13571 1118.26
R24196 vss.n13571 vss.n13567 1118.26
R24197 vss.n13558 vss.n13545 1118.26
R24198 vss.n13601 vss.n13558 1118.26
R24199 vss.n13601 vss.n13559 1118.26
R24200 vss.n13597 vss.n13559 1118.26
R24201 vss.n13597 vss.n13564 1118.26
R24202 vss.n13590 vss.n13564 1118.26
R24203 vss.n13553 vss.n13546 1118.26
R24204 vss.n13602 vss.n13553 1118.26
R24205 vss.n13602 vss.n13554 1118.26
R24206 vss.n13565 vss.n13554 1118.26
R24207 vss.n13584 vss.n13565 1118.26
R24208 vss.n13591 vss.n13584 1118.26
R24209 vss.n13919 vss.n13305 1118.26
R24210 vss.n13915 vss.n13305 1118.26
R24211 vss.n13915 vss.n13309 1118.26
R24212 vss.n13902 vss.n13309 1118.26
R24213 vss.n13902 vss.n13900 1118.26
R24214 vss.n13907 vss.n13900 1118.26
R24215 vss.n13312 vss.n13304 1118.26
R24216 vss.n13914 vss.n13312 1118.26
R24217 vss.n13914 vss.n13313 1118.26
R24218 vss.n13910 vss.n13313 1118.26
R24219 vss.n13910 vss.n13909 1118.26
R24220 vss.n13909 vss.n13908 1118.26
R24221 vss.n13875 vss.n13335 1118.26
R24222 vss.n13881 vss.n13335 1118.26
R24223 vss.n13881 vss.n13332 1118.26
R24224 vss.n13886 vss.n13332 1118.26
R24225 vss.n13887 vss.n13886 1118.26
R24226 vss.n13887 vss.n13326 1118.26
R24227 vss.n13876 vss.n13339 1118.26
R24228 vss.n13880 vss.n13339 1118.26
R24229 vss.n13880 vss.n13331 1118.26
R24230 vss.n13891 vss.n13331 1118.26
R24231 vss.n13891 vss.n13890 1118.26
R24232 vss.n13890 vss.n13327 1118.26
R24233 vss.n13871 vss.n13347 1118.26
R24234 vss.n13867 vss.n13347 1118.26
R24235 vss.n13867 vss.n13351 1118.26
R24236 vss.n13847 vss.n13351 1118.26
R24237 vss.n13847 vss.n13845 1118.26
R24238 vss.n13852 vss.n13845 1118.26
R24239 vss.n13354 vss.n13346 1118.26
R24240 vss.n13866 vss.n13354 1118.26
R24241 vss.n13866 vss.n13355 1118.26
R24242 vss.n13855 vss.n13355 1118.26
R24243 vss.n13855 vss.n13854 1118.26
R24244 vss.n13854 vss.n13853 1118.26
R24245 vss.n13821 vss.n13376 1118.26
R24246 vss.n13827 vss.n13376 1118.26
R24247 vss.n13827 vss.n13373 1118.26
R24248 vss.n13832 vss.n13373 1118.26
R24249 vss.n13833 vss.n13832 1118.26
R24250 vss.n13833 vss.n13365 1118.26
R24251 vss.n13822 vss.n13380 1118.26
R24252 vss.n13826 vss.n13380 1118.26
R24253 vss.n13826 vss.n13372 1118.26
R24254 vss.n13837 vss.n13372 1118.26
R24255 vss.n13837 vss.n13836 1118.26
R24256 vss.n13836 vss.n13366 1118.26
R24257 vss.n13817 vss.n13388 1118.26
R24258 vss.n13813 vss.n13388 1118.26
R24259 vss.n13813 vss.n13392 1118.26
R24260 vss.n13797 vss.n13392 1118.26
R24261 vss.n13797 vss.n13795 1118.26
R24262 vss.n13802 vss.n13795 1118.26
R24263 vss.n13395 vss.n13387 1118.26
R24264 vss.n13812 vss.n13395 1118.26
R24265 vss.n13812 vss.n13396 1118.26
R24266 vss.n13805 vss.n13396 1118.26
R24267 vss.n13805 vss.n13804 1118.26
R24268 vss.n13804 vss.n13803 1118.26
R24269 vss.n13770 vss.n13415 1118.26
R24270 vss.n13776 vss.n13415 1118.26
R24271 vss.n13776 vss.n13412 1118.26
R24272 vss.n13781 vss.n13412 1118.26
R24273 vss.n13782 vss.n13781 1118.26
R24274 vss.n13782 vss.n13406 1118.26
R24275 vss.n13771 vss.n13419 1118.26
R24276 vss.n13775 vss.n13419 1118.26
R24277 vss.n13775 vss.n13411 1118.26
R24278 vss.n13786 vss.n13411 1118.26
R24279 vss.n13786 vss.n13785 1118.26
R24280 vss.n13785 vss.n13407 1118.26
R24281 vss.n13766 vss.n13427 1118.26
R24282 vss.n13762 vss.n13427 1118.26
R24283 vss.n13762 vss.n13431 1118.26
R24284 vss.n13742 vss.n13431 1118.26
R24285 vss.n13742 vss.n13740 1118.26
R24286 vss.n13747 vss.n13740 1118.26
R24287 vss.n13434 vss.n13426 1118.26
R24288 vss.n13761 vss.n13434 1118.26
R24289 vss.n13761 vss.n13435 1118.26
R24290 vss.n13750 vss.n13435 1118.26
R24291 vss.n13750 vss.n13749 1118.26
R24292 vss.n13749 vss.n13748 1118.26
R24293 vss.n13716 vss.n13456 1118.26
R24294 vss.n13722 vss.n13456 1118.26
R24295 vss.n13722 vss.n13453 1118.26
R24296 vss.n13727 vss.n13453 1118.26
R24297 vss.n13728 vss.n13727 1118.26
R24298 vss.n13728 vss.n13445 1118.26
R24299 vss.n13717 vss.n13460 1118.26
R24300 vss.n13721 vss.n13460 1118.26
R24301 vss.n13721 vss.n13452 1118.26
R24302 vss.n13732 vss.n13452 1118.26
R24303 vss.n13732 vss.n13731 1118.26
R24304 vss.n13731 vss.n13446 1118.26
R24305 vss.n13712 vss.n13468 1118.26
R24306 vss.n13708 vss.n13468 1118.26
R24307 vss.n13708 vss.n13472 1118.26
R24308 vss.n13692 vss.n13472 1118.26
R24309 vss.n13692 vss.n13690 1118.26
R24310 vss.n13697 vss.n13690 1118.26
R24311 vss.n13475 vss.n13467 1118.26
R24312 vss.n13707 vss.n13475 1118.26
R24313 vss.n13707 vss.n13476 1118.26
R24314 vss.n13700 vss.n13476 1118.26
R24315 vss.n13700 vss.n13699 1118.26
R24316 vss.n13699 vss.n13698 1118.26
R24317 vss.n13665 vss.n13495 1118.26
R24318 vss.n13671 vss.n13495 1118.26
R24319 vss.n13671 vss.n13492 1118.26
R24320 vss.n13676 vss.n13492 1118.26
R24321 vss.n13677 vss.n13676 1118.26
R24322 vss.n13677 vss.n13486 1118.26
R24323 vss.n13666 vss.n13499 1118.26
R24324 vss.n13670 vss.n13499 1118.26
R24325 vss.n13670 vss.n13491 1118.26
R24326 vss.n13681 vss.n13491 1118.26
R24327 vss.n13681 vss.n13680 1118.26
R24328 vss.n13680 vss.n13487 1118.26
R24329 vss.n13661 vss.n13507 1118.26
R24330 vss.n13657 vss.n13507 1118.26
R24331 vss.n13657 vss.n13511 1118.26
R24332 vss.n13637 vss.n13511 1118.26
R24333 vss.n13637 vss.n13635 1118.26
R24334 vss.n13642 vss.n13635 1118.26
R24335 vss.n13514 vss.n13506 1118.26
R24336 vss.n13656 vss.n13514 1118.26
R24337 vss.n13656 vss.n13515 1118.26
R24338 vss.n13645 vss.n13515 1118.26
R24339 vss.n13645 vss.n13644 1118.26
R24340 vss.n13644 vss.n13643 1118.26
R24341 vss.n13611 vss.n13536 1118.26
R24342 vss.n13617 vss.n13536 1118.26
R24343 vss.n13617 vss.n13533 1118.26
R24344 vss.n13622 vss.n13533 1118.26
R24345 vss.n13623 vss.n13622 1118.26
R24346 vss.n13623 vss.n13525 1118.26
R24347 vss.n13612 vss.n13540 1118.26
R24348 vss.n13616 vss.n13540 1118.26
R24349 vss.n13616 vss.n13532 1118.26
R24350 vss.n13627 vss.n13532 1118.26
R24351 vss.n13627 vss.n13626 1118.26
R24352 vss.n13626 vss.n13526 1118.26
R24353 vss.n14007 vss.n14006 1118.26
R24354 vss.n14008 vss.n14007 1118.26
R24355 vss.n14008 vss.n520 1118.26
R24356 vss.n14022 vss.n520 1118.26
R24357 vss.n14022 vss.n521 1118.26
R24358 vss.n14014 vss.n521 1118.26
R24359 vss.n14005 vss.n527 1118.26
R24360 vss.n14009 vss.n527 1118.26
R24361 vss.n14009 vss.n529 1118.26
R24362 vss.n529 vss.n523 1118.26
R24363 vss.n14019 vss.n523 1118.26
R24364 vss.n14019 vss.n14018 1118.26
R24365 vss.n547 vss.n537 1118.26
R24366 vss.n13994 vss.n547 1118.26
R24367 vss.n13994 vss.n548 1118.26
R24368 vss.n671 vss.n548 1118.26
R24369 vss.n671 vss.n670 1118.26
R24370 vss.n670 vss.n660 1118.26
R24371 vss.n542 vss.n538 1118.26
R24372 vss.n13995 vss.n542 1118.26
R24373 vss.n13995 vss.n543 1118.26
R24374 vss.n672 vss.n543 1118.26
R24375 vss.n672 vss.n665 1118.26
R24376 vss.n665 vss.n661 1118.26
R24377 vss.n13972 vss.n13971 1118.26
R24378 vss.n13973 vss.n13972 1118.26
R24379 vss.n13973 vss.n559 1118.26
R24380 vss.n13987 vss.n559 1118.26
R24381 vss.n13987 vss.n560 1118.26
R24382 vss.n13979 vss.n560 1118.26
R24383 vss.n13970 vss.n566 1118.26
R24384 vss.n13974 vss.n566 1118.26
R24385 vss.n13974 vss.n568 1118.26
R24386 vss.n568 vss.n562 1118.26
R24387 vss.n13984 vss.n562 1118.26
R24388 vss.n13984 vss.n13983 1118.26
R24389 vss.n586 vss.n576 1118.26
R24390 vss.n13959 vss.n586 1118.26
R24391 vss.n13959 vss.n587 1118.26
R24392 vss.n770 vss.n587 1118.26
R24393 vss.n770 vss.n764 1118.26
R24394 vss.n777 vss.n764 1118.26
R24395 vss.n581 vss.n577 1118.26
R24396 vss.n13960 vss.n581 1118.26
R24397 vss.n13960 vss.n582 1118.26
R24398 vss.n771 vss.n582 1118.26
R24399 vss.n771 vss.n769 1118.26
R24400 vss.n769 vss.n763 1118.26
R24401 vss.n753 vss.n743 1118.26
R24402 vss.n13242 vss.n753 1118.26
R24403 vss.n13242 vss.n754 1118.26
R24404 vss.n791 vss.n754 1118.26
R24405 vss.n791 vss.n759 1118.26
R24406 vss.n783 vss.n759 1118.26
R24407 vss.n748 vss.n744 1118.26
R24408 vss.n13243 vss.n748 1118.26
R24409 vss.n13243 vss.n749 1118.26
R24410 vss.n760 vss.n749 1118.26
R24411 vss.n788 vss.n760 1118.26
R24412 vss.n788 vss.n787 1118.26
R24413 vss.n1730 vss.n1720 1118.26
R24414 vss.n1736 vss.n1720 1118.26
R24415 vss.n1736 vss.n1716 1118.26
R24416 vss.n1741 vss.n1716 1118.26
R24417 vss.n1741 vss.n1708 1118.26
R24418 vss.n1748 vss.n1708 1118.26
R24419 vss.n1731 vss.n1722 1118.26
R24420 vss.n1735 vss.n1722 1118.26
R24421 vss.n1735 vss.n1712 1118.26
R24422 vss.n1742 vss.n1712 1118.26
R24423 vss.n1742 vss.n1714 1118.26
R24424 vss.n1714 vss.n1707 1118.26
R24425 vss.n1784 vss.n1783 1118.26
R24426 vss.n1785 vss.n1784 1118.26
R24427 vss.n1785 vss.n1701 1118.26
R24428 vss.n1799 vss.n1701 1118.26
R24429 vss.n1799 vss.n1702 1118.26
R24430 vss.n1791 vss.n1702 1118.26
R24431 vss.n1782 vss.n1753 1118.26
R24432 vss.n1786 vss.n1753 1118.26
R24433 vss.n1786 vss.n1755 1118.26
R24434 vss.n1755 vss.n1704 1118.26
R24435 vss.n1796 vss.n1704 1118.26
R24436 vss.n1796 vss.n1795 1118.26
R24437 vss.n1770 vss.n1762 1118.26
R24438 vss.n1771 vss.n1770 1118.26
R24439 vss.n1771 vss.n1273 1118.26
R24440 vss.n1812 vss.n1273 1118.26
R24441 vss.n1812 vss.n1265 1118.26
R24442 vss.n1819 vss.n1265 1118.26
R24443 vss.n1767 vss.n1763 1118.26
R24444 vss.n1772 vss.n1767 1118.26
R24445 vss.n1772 vss.n1269 1118.26
R24446 vss.n1813 vss.n1269 1118.26
R24447 vss.n1813 vss.n1271 1118.26
R24448 vss.n1271 vss.n1264 1118.26
R24449 vss.n1830 vss.n1829 1118.26
R24450 vss.n1829 vss.n1828 1118.26
R24451 vss.n1828 vss.n1236 1118.26
R24452 vss.n1826 vss.n1236 1118.26
R24453 vss.n1826 vss.n1244 1118.26
R24454 vss.n1822 vss.n1244 1118.26
R24455 vss.n1238 vss.n1232 1118.26
R24456 vss.n1239 vss.n1238 1118.26
R24457 vss.n1241 vss.n1239 1118.26
R24458 vss.n1242 vss.n1241 1118.26
R24459 vss.n1250 vss.n1242 1118.26
R24460 vss.n1262 vss.n1250 1118.26
R24461 vss.n1834 vss.n1224 1118.26
R24462 vss.n1840 vss.n1224 1118.26
R24463 vss.n1840 vss.n1220 1118.26
R24464 vss.n1845 vss.n1220 1118.26
R24465 vss.n1845 vss.n1212 1118.26
R24466 vss.n1852 vss.n1212 1118.26
R24467 vss.n1835 vss.n1226 1118.26
R24468 vss.n1839 vss.n1226 1118.26
R24469 vss.n1839 vss.n1216 1118.26
R24470 vss.n1846 vss.n1216 1118.26
R24471 vss.n1846 vss.n1218 1118.26
R24472 vss.n1218 vss.n1211 1118.26
R24473 vss.n1888 vss.n1887 1118.26
R24474 vss.n1889 vss.n1888 1118.26
R24475 vss.n1889 vss.n1205 1118.26
R24476 vss.n1903 vss.n1205 1118.26
R24477 vss.n1903 vss.n1206 1118.26
R24478 vss.n1895 vss.n1206 1118.26
R24479 vss.n1886 vss.n1857 1118.26
R24480 vss.n1890 vss.n1857 1118.26
R24481 vss.n1890 vss.n1859 1118.26
R24482 vss.n1859 vss.n1208 1118.26
R24483 vss.n1900 vss.n1208 1118.26
R24484 vss.n1900 vss.n1899 1118.26
R24485 vss.n1874 vss.n1866 1118.26
R24486 vss.n1875 vss.n1874 1118.26
R24487 vss.n1875 vss.n1155 1118.26
R24488 vss.n1916 vss.n1155 1118.26
R24489 vss.n1916 vss.n1147 1118.26
R24490 vss.n1923 vss.n1147 1118.26
R24491 vss.n1871 vss.n1867 1118.26
R24492 vss.n1876 vss.n1871 1118.26
R24493 vss.n1876 vss.n1151 1118.26
R24494 vss.n1917 vss.n1151 1118.26
R24495 vss.n1917 vss.n1153 1118.26
R24496 vss.n1153 vss.n1146 1118.26
R24497 vss.n1959 vss.n1958 1118.26
R24498 vss.n1960 vss.n1959 1118.26
R24499 vss.n1960 vss.n1140 1118.26
R24500 vss.n1974 vss.n1140 1118.26
R24501 vss.n1974 vss.n1141 1118.26
R24502 vss.n1966 vss.n1141 1118.26
R24503 vss.n1957 vss.n1928 1118.26
R24504 vss.n1961 vss.n1928 1118.26
R24505 vss.n1961 vss.n1930 1118.26
R24506 vss.n1930 vss.n1143 1118.26
R24507 vss.n1971 vss.n1143 1118.26
R24508 vss.n1971 vss.n1970 1118.26
R24509 vss.n1945 vss.n1937 1118.26
R24510 vss.n1946 vss.n1945 1118.26
R24511 vss.n1946 vss.n699 1118.26
R24512 vss.n13294 vss.n699 1118.26
R24513 vss.n13294 vss.n701 1118.26
R24514 vss.n701 vss.n690 1118.26
R24515 vss.n1942 vss.n1938 1118.26
R24516 vss.n1947 vss.n1942 1118.26
R24517 vss.n1947 vss.n695 1118.26
R24518 vss.n13295 vss.n695 1118.26
R24519 vss.n13295 vss.n696 1118.26
R24520 vss.n696 vss.n691 1118.26
R24521 vss.n13271 vss.n13270 1118.26
R24522 vss.n13272 vss.n13271 1118.26
R24523 vss.n13272 vss.n710 1118.26
R24524 vss.n13286 vss.n710 1118.26
R24525 vss.n13286 vss.n711 1118.26
R24526 vss.n13278 vss.n711 1118.26
R24527 vss.n13269 vss.n719 1118.26
R24528 vss.n13273 vss.n719 1118.26
R24529 vss.n13273 vss.n721 1118.26
R24530 vss.n721 vss.n713 1118.26
R24531 vss.n13283 vss.n713 1118.26
R24532 vss.n13283 vss.n13282 1118.26
R24533 vss.n9607 vss.n9597 1118.26
R24534 vss.n9611 vss.n9597 1118.26
R24535 vss.n9611 vss.n9594 1118.26
R24536 vss.n9624 vss.n9594 1118.26
R24537 vss.n9624 vss.n9595 1118.26
R24538 vss.n9620 vss.n9595 1118.26
R24539 vss.n9609 vss.n9608 1118.26
R24540 vss.n9610 vss.n9609 1118.26
R24541 vss.n9610 vss.n9589 1118.26
R24542 vss.n9625 vss.n9589 1118.26
R24543 vss.n9625 vss.n9590 1118.26
R24544 vss.n9619 vss.n9590 1118.26
R24545 vss.n7504 vss.n7491 1118.26
R24546 vss.n7528 vss.n7504 1118.26
R24547 vss.n7528 vss.n7505 1118.26
R24548 vss.n7524 vss.n7505 1118.26
R24549 vss.n7524 vss.n7510 1118.26
R24550 vss.n7516 vss.n7510 1118.26
R24551 vss.n7499 vss.n7492 1118.26
R24552 vss.n7529 vss.n7499 1118.26
R24553 vss.n7529 vss.n7500 1118.26
R24554 vss.n7511 vss.n7500 1118.26
R24555 vss.n7512 vss.n7511 1118.26
R24556 vss.n7518 vss.n7512 1118.26
R24557 vss.n8916 vss.n8904 1118.26
R24558 vss.n8940 vss.n8916 1118.26
R24559 vss.n8940 vss.n8917 1118.26
R24560 vss.n8936 vss.n8917 1118.26
R24561 vss.n8936 vss.n8922 1118.26
R24562 vss.n8928 vss.n8922 1118.26
R24563 vss.n8911 vss.n8905 1118.26
R24564 vss.n8941 vss.n8911 1118.26
R24565 vss.n8941 vss.n8912 1118.26
R24566 vss.n8923 vss.n8912 1118.26
R24567 vss.n8924 vss.n8923 1118.26
R24568 vss.n8930 vss.n8924 1118.26
R24569 vss.n7566 vss.n7556 1118.26
R24570 vss.n7570 vss.n7556 1118.26
R24571 vss.n7570 vss.n7553 1118.26
R24572 vss.n7583 vss.n7553 1118.26
R24573 vss.n7583 vss.n7554 1118.26
R24574 vss.n7579 vss.n7554 1118.26
R24575 vss.n7568 vss.n7567 1118.26
R24576 vss.n7569 vss.n7568 1118.26
R24577 vss.n7569 vss.n7548 1118.26
R24578 vss.n7584 vss.n7548 1118.26
R24579 vss.n7584 vss.n7549 1118.26
R24580 vss.n7578 vss.n7549 1118.26
R24581 vss.n8797 vss.n8785 1118.26
R24582 vss.n8821 vss.n8797 1118.26
R24583 vss.n8821 vss.n8798 1118.26
R24584 vss.n8817 vss.n8798 1118.26
R24585 vss.n8817 vss.n8803 1118.26
R24586 vss.n8809 vss.n8803 1118.26
R24587 vss.n8792 vss.n8786 1118.26
R24588 vss.n8822 vss.n8792 1118.26
R24589 vss.n8822 vss.n8793 1118.26
R24590 vss.n8804 vss.n8793 1118.26
R24591 vss.n8805 vss.n8804 1118.26
R24592 vss.n8811 vss.n8805 1118.26
R24593 vss.n7709 vss.n7699 1118.26
R24594 vss.n7713 vss.n7699 1118.26
R24595 vss.n7713 vss.n7696 1118.26
R24596 vss.n7726 vss.n7696 1118.26
R24597 vss.n7726 vss.n7697 1118.26
R24598 vss.n7722 vss.n7697 1118.26
R24599 vss.n7711 vss.n7710 1118.26
R24600 vss.n7712 vss.n7711 1118.26
R24601 vss.n7712 vss.n7691 1118.26
R24602 vss.n7727 vss.n7691 1118.26
R24603 vss.n7727 vss.n7692 1118.26
R24604 vss.n7721 vss.n7692 1118.26
R24605 vss.n7789 vss.n7779 1118.26
R24606 vss.n7793 vss.n7779 1118.26
R24607 vss.n7793 vss.n7776 1118.26
R24608 vss.n7806 vss.n7776 1118.26
R24609 vss.n7806 vss.n7777 1118.26
R24610 vss.n7802 vss.n7777 1118.26
R24611 vss.n7791 vss.n7790 1118.26
R24612 vss.n7792 vss.n7791 1118.26
R24613 vss.n7792 vss.n7771 1118.26
R24614 vss.n7807 vss.n7771 1118.26
R24615 vss.n7807 vss.n7772 1118.26
R24616 vss.n7801 vss.n7772 1118.26
R24617 vss.n7930 vss.n7920 1118.26
R24618 vss.n7934 vss.n7920 1118.26
R24619 vss.n7934 vss.n7917 1118.26
R24620 vss.n7947 vss.n7917 1118.26
R24621 vss.n7947 vss.n7918 1118.26
R24622 vss.n7943 vss.n7918 1118.26
R24623 vss.n7932 vss.n7931 1118.26
R24624 vss.n7933 vss.n7932 1118.26
R24625 vss.n7933 vss.n7912 1118.26
R24626 vss.n7948 vss.n7912 1118.26
R24627 vss.n7948 vss.n7913 1118.26
R24628 vss.n7942 vss.n7913 1118.26
R24629 vss.n8187 vss.n8175 1118.26
R24630 vss.n8211 vss.n8187 1118.26
R24631 vss.n8211 vss.n8188 1118.26
R24632 vss.n8207 vss.n8188 1118.26
R24633 vss.n8207 vss.n8193 1118.26
R24634 vss.n8199 vss.n8193 1118.26
R24635 vss.n8182 vss.n8176 1118.26
R24636 vss.n8212 vss.n8182 1118.26
R24637 vss.n8212 vss.n8183 1118.26
R24638 vss.n8194 vss.n8183 1118.26
R24639 vss.n8195 vss.n8194 1118.26
R24640 vss.n8201 vss.n8195 1118.26
R24641 vss.n8224 vss.n8003 1118.26
R24642 vss.n8228 vss.n8003 1118.26
R24643 vss.n8228 vss.n8000 1118.26
R24644 vss.n8241 vss.n8000 1118.26
R24645 vss.n8241 vss.n8001 1118.26
R24646 vss.n8237 vss.n8001 1118.26
R24647 vss.n8226 vss.n8225 1118.26
R24648 vss.n8227 vss.n8226 1118.26
R24649 vss.n8227 vss.n7995 1118.26
R24650 vss.n8242 vss.n7995 1118.26
R24651 vss.n8242 vss.n7996 1118.26
R24652 vss.n8236 vss.n7996 1118.26
R24653 vss.n7310 vss.n7300 1118.26
R24654 vss.n8999 vss.n7310 1118.26
R24655 vss.n8999 vss.n7311 1118.26
R24656 vss.n8995 vss.n7311 1118.26
R24657 vss.n8995 vss.n7316 1118.26
R24658 vss.n7322 vss.n7316 1118.26
R24659 vss.n7305 vss.n7301 1118.26
R24660 vss.n9000 vss.n7305 1118.26
R24661 vss.n9000 vss.n7306 1118.26
R24662 vss.n7317 vss.n7306 1118.26
R24663 vss.n7318 vss.n7317 1118.26
R24664 vss.n8989 vss.n7318 1118.26
R24665 vss.n8715 vss.n7860 1118.26
R24666 vss.n8719 vss.n7860 1118.26
R24667 vss.n8719 vss.n7857 1118.26
R24668 vss.n8732 vss.n7857 1118.26
R24669 vss.n8732 vss.n7858 1118.26
R24670 vss.n8728 vss.n7858 1118.26
R24671 vss.n8717 vss.n8716 1118.26
R24672 vss.n8718 vss.n8717 1118.26
R24673 vss.n8718 vss.n7852 1118.26
R24674 vss.n8733 vss.n7852 1118.26
R24675 vss.n8733 vss.n7853 1118.26
R24676 vss.n8727 vss.n7853 1118.26
R24677 vss.n8751 vss.n7683 1118.26
R24678 vss.n8775 vss.n8751 1118.26
R24679 vss.n8775 vss.n8752 1118.26
R24680 vss.n8771 vss.n8752 1118.26
R24681 vss.n8771 vss.n8757 1118.26
R24682 vss.n8763 vss.n8757 1118.26
R24683 vss.n8746 vss.n7684 1118.26
R24684 vss.n8776 vss.n8746 1118.26
R24685 vss.n8776 vss.n8747 1118.26
R24686 vss.n8758 vss.n8747 1118.26
R24687 vss.n8759 vss.n8758 1118.26
R24688 vss.n8765 vss.n8759 1118.26
R24689 vss.n8834 vss.n7673 1118.26
R24690 vss.n8838 vss.n7673 1118.26
R24691 vss.n8838 vss.n7670 1118.26
R24692 vss.n8851 vss.n7670 1118.26
R24693 vss.n8851 vss.n7671 1118.26
R24694 vss.n8847 vss.n7671 1118.26
R24695 vss.n8836 vss.n8835 1118.26
R24696 vss.n8837 vss.n8836 1118.26
R24697 vss.n8837 vss.n7665 1118.26
R24698 vss.n8852 vss.n7665 1118.26
R24699 vss.n8852 vss.n7666 1118.26
R24700 vss.n8846 vss.n7666 1118.26
R24701 vss.n8870 vss.n7540 1118.26
R24702 vss.n8894 vss.n8870 1118.26
R24703 vss.n8894 vss.n8871 1118.26
R24704 vss.n8890 vss.n8871 1118.26
R24705 vss.n8890 vss.n8876 1118.26
R24706 vss.n8882 vss.n8876 1118.26
R24707 vss.n8865 vss.n7541 1118.26
R24708 vss.n8895 vss.n8865 1118.26
R24709 vss.n8895 vss.n8866 1118.26
R24710 vss.n8877 vss.n8866 1118.26
R24711 vss.n8878 vss.n8877 1118.26
R24712 vss.n8884 vss.n8878 1118.26
R24713 vss.n8953 vss.n7484 1118.26
R24714 vss.n8957 vss.n7484 1118.26
R24715 vss.n8957 vss.n7481 1118.26
R24716 vss.n8970 vss.n7481 1118.26
R24717 vss.n8970 vss.n7482 1118.26
R24718 vss.n8966 vss.n7482 1118.26
R24719 vss.n8955 vss.n8954 1118.26
R24720 vss.n8956 vss.n8955 1118.26
R24721 vss.n8956 vss.n7476 1118.26
R24722 vss.n8971 vss.n7476 1118.26
R24723 vss.n8971 vss.n7477 1118.26
R24724 vss.n8965 vss.n7477 1118.26
R24725 vss.n8081 vss.n8071 1118.26
R24726 vss.n8087 vss.n8071 1118.26
R24727 vss.n8087 vss.n8065 1118.26
R24728 vss.n8092 vss.n8065 1118.26
R24729 vss.n8092 vss.n8067 1118.26
R24730 vss.n8067 vss.n8053 1118.26
R24731 vss.n8082 vss.n8073 1118.26
R24732 vss.n8086 vss.n8073 1118.26
R24733 vss.n8086 vss.n8061 1118.26
R24734 vss.n8093 vss.n8061 1118.26
R24735 vss.n8093 vss.n8062 1118.26
R24736 vss.n8062 vss.n8054 1118.26
R24737 vss.n9341 vss.n9331 1118.26
R24738 vss.n9345 vss.n9331 1118.26
R24739 vss.n9345 vss.n9328 1118.26
R24740 vss.n9358 vss.n9328 1118.26
R24741 vss.n9358 vss.n9329 1118.26
R24742 vss.n9354 vss.n9329 1118.26
R24743 vss.n9343 vss.n9342 1118.26
R24744 vss.n9344 vss.n9343 1118.26
R24745 vss.n9344 vss.n9323 1118.26
R24746 vss.n9359 vss.n9323 1118.26
R24747 vss.n9359 vss.n9324 1118.26
R24748 vss.n9352 vss.n9324 1118.26
R24749 vss.n6345 vss.n6335 1118.26
R24750 vss.n6349 vss.n6335 1118.26
R24751 vss.n6349 vss.n6332 1118.26
R24752 vss.n6362 vss.n6332 1118.26
R24753 vss.n6362 vss.n6333 1118.26
R24754 vss.n6358 vss.n6333 1118.26
R24755 vss.n6347 vss.n6346 1118.26
R24756 vss.n6348 vss.n6347 1118.26
R24757 vss.n6348 vss.n6327 1118.26
R24758 vss.n6363 vss.n6327 1118.26
R24759 vss.n6363 vss.n6328 1118.26
R24760 vss.n6356 vss.n6328 1118.26
R24761 vss.n6423 vss.n6413 1118.26
R24762 vss.n6427 vss.n6413 1118.26
R24763 vss.n6427 vss.n6410 1118.26
R24764 vss.n6440 vss.n6410 1118.26
R24765 vss.n6440 vss.n6411 1118.26
R24766 vss.n6436 vss.n6411 1118.26
R24767 vss.n6425 vss.n6424 1118.26
R24768 vss.n6426 vss.n6425 1118.26
R24769 vss.n6426 vss.n6405 1118.26
R24770 vss.n6441 vss.n6405 1118.26
R24771 vss.n6441 vss.n6406 1118.26
R24772 vss.n6434 vss.n6406 1118.26
R24773 vss.n6959 vss.n6949 1118.26
R24774 vss.n6963 vss.n6949 1118.26
R24775 vss.n6963 vss.n6946 1118.26
R24776 vss.n6976 vss.n6946 1118.26
R24777 vss.n6976 vss.n6947 1118.26
R24778 vss.n6972 vss.n6947 1118.26
R24779 vss.n6961 vss.n6960 1118.26
R24780 vss.n6962 vss.n6961 1118.26
R24781 vss.n6962 vss.n6941 1118.26
R24782 vss.n6977 vss.n6941 1118.26
R24783 vss.n6977 vss.n6942 1118.26
R24784 vss.n6970 vss.n6942 1118.26
R24785 vss.n6650 vss.n6640 1118.26
R24786 vss.n6654 vss.n6640 1118.26
R24787 vss.n6654 vss.n6637 1118.26
R24788 vss.n6667 vss.n6637 1118.26
R24789 vss.n6667 vss.n6638 1118.26
R24790 vss.n6663 vss.n6638 1118.26
R24791 vss.n6652 vss.n6651 1118.26
R24792 vss.n6653 vss.n6652 1118.26
R24793 vss.n6653 vss.n6632 1118.26
R24794 vss.n6668 vss.n6632 1118.26
R24795 vss.n6668 vss.n6633 1118.26
R24796 vss.n6661 vss.n6633 1118.26
R24797 vss.n7148 vss.n7138 1118.26
R24798 vss.n7152 vss.n7138 1118.26
R24799 vss.n7152 vss.n7135 1118.26
R24800 vss.n7165 vss.n7135 1118.26
R24801 vss.n7165 vss.n7136 1118.26
R24802 vss.n7161 vss.n7136 1118.26
R24803 vss.n7150 vss.n7149 1118.26
R24804 vss.n7151 vss.n7150 1118.26
R24805 vss.n7151 vss.n7130 1118.26
R24806 vss.n7166 vss.n7130 1118.26
R24807 vss.n7166 vss.n7131 1118.26
R24808 vss.n7159 vss.n7131 1118.26
R24809 vss.n9421 vss.n9413 1118.26
R24810 vss.n9425 vss.n9413 1118.26
R24811 vss.n9425 vss.n9405 1118.26
R24812 vss.n9438 vss.n9405 1118.26
R24813 vss.n9438 vss.n9437 1118.26
R24814 vss.n9437 vss.n9401 1118.26
R24815 vss.n9420 vss.n9409 1118.26
R24816 vss.n9426 vss.n9409 1118.26
R24817 vss.n9426 vss.n9406 1118.26
R24818 vss.n9433 vss.n9406 1118.26
R24819 vss.n9434 vss.n9433 1118.26
R24820 vss.n9434 vss.n9400 1118.26
R24821 vss.n6029 vss.n6019 1118.26
R24822 vss.n6033 vss.n6019 1118.26
R24823 vss.n6033 vss.n6016 1118.26
R24824 vss.n6047 vss.n6016 1118.26
R24825 vss.n6047 vss.n6017 1118.26
R24826 vss.n6043 vss.n6017 1118.26
R24827 vss.n6031 vss.n6030 1118.26
R24828 vss.n6032 vss.n6031 1118.26
R24829 vss.n6032 vss.n6011 1118.26
R24830 vss.n6048 vss.n6011 1118.26
R24831 vss.n6048 vss.n6012 1118.26
R24832 vss.n6040 vss.n6012 1118.26
R24833 vss.n9466 vss.n9457 1118.26
R24834 vss.n9470 vss.n9457 1118.26
R24835 vss.n9470 vss.n9450 1118.26
R24836 vss.n9480 vss.n9450 1118.26
R24837 vss.n9480 vss.n9479 1118.26
R24838 vss.n9479 vss.n9446 1118.26
R24839 vss.n9465 vss.n9453 1118.26
R24840 vss.n9471 vss.n9453 1118.26
R24841 vss.n9472 vss.n9471 1118.26
R24842 vss.n9475 vss.n9472 1118.26
R24843 vss.n9476 vss.n9475 1118.26
R24844 vss.n9476 vss.n9445 1118.26
R24845 vss.n6156 vss.n6146 1118.26
R24846 vss.n6160 vss.n6146 1118.26
R24847 vss.n6160 vss.n6143 1118.26
R24848 vss.n9498 vss.n6143 1118.26
R24849 vss.n9498 vss.n6144 1118.26
R24850 vss.n9494 vss.n6144 1118.26
R24851 vss.n6158 vss.n6157 1118.26
R24852 vss.n6159 vss.n6158 1118.26
R24853 vss.n6159 vss.n6138 1118.26
R24854 vss.n9499 vss.n6138 1118.26
R24855 vss.n9499 vss.n6139 1118.26
R24856 vss.n6167 vss.n6139 1118.26
R24857 vss.n7199 vss.n7189 1118.26
R24858 vss.n7203 vss.n7189 1118.26
R24859 vss.n7203 vss.n7186 1118.26
R24860 vss.n7216 vss.n7186 1118.26
R24861 vss.n7216 vss.n7187 1118.26
R24862 vss.n7212 vss.n7187 1118.26
R24863 vss.n7201 vss.n7200 1118.26
R24864 vss.n7202 vss.n7201 1118.26
R24865 vss.n7202 vss.n7181 1118.26
R24866 vss.n7217 vss.n7181 1118.26
R24867 vss.n7217 vss.n7182 1118.26
R24868 vss.n7210 vss.n7182 1118.26
R24869 vss.n6694 vss.n6684 1118.26
R24870 vss.n6698 vss.n6684 1118.26
R24871 vss.n6698 vss.n6681 1118.26
R24872 vss.n6711 vss.n6681 1118.26
R24873 vss.n6711 vss.n6682 1118.26
R24874 vss.n6707 vss.n6682 1118.26
R24875 vss.n6696 vss.n6695 1118.26
R24876 vss.n6697 vss.n6696 1118.26
R24877 vss.n6697 vss.n6676 1118.26
R24878 vss.n6712 vss.n6676 1118.26
R24879 vss.n6712 vss.n6677 1118.26
R24880 vss.n6705 vss.n6677 1118.26
R24881 vss.n7008 vss.n6998 1118.26
R24882 vss.n7012 vss.n6998 1118.26
R24883 vss.n7012 vss.n6995 1118.26
R24884 vss.n7025 vss.n6995 1118.26
R24885 vss.n7025 vss.n6996 1118.26
R24886 vss.n7021 vss.n6996 1118.26
R24887 vss.n7010 vss.n7009 1118.26
R24888 vss.n7011 vss.n7010 1118.26
R24889 vss.n7011 vss.n6990 1118.26
R24890 vss.n7026 vss.n6990 1118.26
R24891 vss.n7026 vss.n6991 1118.26
R24892 vss.n7019 vss.n6991 1118.26
R24893 vss.n6468 vss.n6458 1118.26
R24894 vss.n6472 vss.n6458 1118.26
R24895 vss.n6472 vss.n6455 1118.26
R24896 vss.n6485 vss.n6455 1118.26
R24897 vss.n6485 vss.n6456 1118.26
R24898 vss.n6481 vss.n6456 1118.26
R24899 vss.n6470 vss.n6469 1118.26
R24900 vss.n6471 vss.n6470 1118.26
R24901 vss.n6471 vss.n6450 1118.26
R24902 vss.n6486 vss.n6450 1118.26
R24903 vss.n6486 vss.n6451 1118.26
R24904 vss.n6479 vss.n6451 1118.26
R24905 vss.n9171 vss.n9161 1118.26
R24906 vss.n9175 vss.n9161 1118.26
R24907 vss.n9175 vss.n9158 1118.26
R24908 vss.n9188 vss.n9158 1118.26
R24909 vss.n9188 vss.n9159 1118.26
R24910 vss.n9184 vss.n9159 1118.26
R24911 vss.n9173 vss.n9172 1118.26
R24912 vss.n9174 vss.n9173 1118.26
R24913 vss.n9174 vss.n9153 1118.26
R24914 vss.n9189 vss.n9153 1118.26
R24915 vss.n9189 vss.n9154 1118.26
R24916 vss.n9182 vss.n9154 1118.26
R24917 vss.n6206 vss.n6198 1118.26
R24918 vss.n6210 vss.n6198 1118.26
R24919 vss.n6210 vss.n6190 1118.26
R24920 vss.n9376 vss.n6190 1118.26
R24921 vss.n9376 vss.n9375 1118.26
R24922 vss.n9375 vss.n6186 1118.26
R24923 vss.n6205 vss.n6194 1118.26
R24924 vss.n6211 vss.n6194 1118.26
R24925 vss.n6211 vss.n6191 1118.26
R24926 vss.n9371 vss.n6191 1118.26
R24927 vss.n9372 vss.n9371 1118.26
R24928 vss.n9372 vss.n6185 1118.26
R24929 vss.n8050 vss.n8014 1118.26
R24930 vss.n8046 vss.n8014 1118.26
R24931 vss.n8046 vss.n8018 1118.26
R24932 vss.n8030 vss.n8018 1118.26
R24933 vss.n8030 vss.n8029 1118.26
R24934 vss.n8034 vss.n8029 1118.26
R24935 vss.n8021 vss.n8013 1118.26
R24936 vss.n8045 vss.n8021 1118.26
R24937 vss.n8045 vss.n8041 1118.26
R24938 vss.n8041 vss.n8040 1118.26
R24939 vss.n8040 vss.n8024 1118.26
R24940 vss.n8036 vss.n8024 1118.26
R24941 vss.n5984 vss.n5974 1118.26
R24942 vss.n9661 vss.n5984 1118.26
R24943 vss.n9661 vss.n5985 1118.26
R24944 vss.n9657 vss.n5985 1118.26
R24945 vss.n9657 vss.n5990 1118.26
R24946 vss.n5996 vss.n5990 1118.26
R24947 vss.n5979 vss.n5975 1118.26
R24948 vss.n9662 vss.n5979 1118.26
R24949 vss.n9662 vss.n5980 1118.26
R24950 vss.n5991 vss.n5980 1118.26
R24951 vss.n5992 vss.n5991 1118.26
R24952 vss.n9651 vss.n5992 1118.26
R24953 vss.n8124 vss.n5997 1118.26
R24954 vss.n8145 vss.n5997 1118.26
R24955 vss.n8145 vss.n8144 1118.26
R24956 vss.n8144 vss.n8143 1118.26
R24957 vss.n8143 vss.n8127 1118.26
R24958 vss.n8136 vss.n8127 1118.26
R24959 vss.n9645 vss.n5999 1118.26
R24960 vss.n9645 vss.n9644 1118.26
R24961 vss.n9644 vss.n6000 1118.26
R24962 vss.n8142 vss.n6000 1118.26
R24963 vss.n8142 vss.n8141 1118.26
R24964 vss.n8141 vss.n8140 1118.26
R24965 vss.n8155 vss.n8115 1118.26
R24966 vss.n8161 vss.n8115 1118.26
R24967 vss.n8161 vss.n8109 1118.26
R24968 vss.n8166 vss.n8109 1118.26
R24969 vss.n8166 vss.n8111 1118.26
R24970 vss.n8111 vss.n8100 1118.26
R24971 vss.n8156 vss.n8117 1118.26
R24972 vss.n8160 vss.n8117 1118.26
R24973 vss.n8160 vss.n8105 1118.26
R24974 vss.n8167 vss.n8105 1118.26
R24975 vss.n8167 vss.n8106 1118.26
R24976 vss.n8106 vss.n8101 1118.26
R24977 vss.n7278 vss.n7268 1118.26
R24978 vss.n9030 vss.n7278 1118.26
R24979 vss.n9030 vss.n7279 1118.26
R24980 vss.n9026 vss.n7279 1118.26
R24981 vss.n9026 vss.n7284 1118.26
R24982 vss.n7290 vss.n7284 1118.26
R24983 vss.n7273 vss.n7269 1118.26
R24984 vss.n9031 vss.n7273 1118.26
R24985 vss.n9031 vss.n7274 1118.26
R24986 vss.n7285 vss.n7274 1118.26
R24987 vss.n7286 vss.n7285 1118.26
R24988 vss.n9020 vss.n7286 1118.26
R24989 vss.n8266 vss.n7900 1118.26
R24990 vss.n8275 vss.n8266 1118.26
R24991 vss.n8275 vss.n8267 1118.26
R24992 vss.n8271 vss.n8267 1118.26
R24993 vss.n8271 vss.n7291 1118.26
R24994 vss.n7297 vss.n7291 1118.26
R24995 vss.n8260 vss.n7901 1118.26
R24996 vss.n8276 vss.n8260 1118.26
R24997 vss.n8276 vss.n8262 1118.26
R24998 vss.n8262 vss.n8261 1118.26
R24999 vss.n8261 vss.n7292 1118.26
R25000 vss.n9011 vss.n7292 1118.26
R25001 vss.n8285 vss.n7893 1118.26
R25002 vss.n8291 vss.n7893 1118.26
R25003 vss.n8291 vss.n7887 1118.26
R25004 vss.n8296 vss.n7887 1118.26
R25005 vss.n8296 vss.n7889 1118.26
R25006 vss.n7889 vss.n7878 1118.26
R25007 vss.n8286 vss.n7895 1118.26
R25008 vss.n8290 vss.n7895 1118.26
R25009 vss.n8290 vss.n7883 1118.26
R25010 vss.n8297 vss.n7883 1118.26
R25011 vss.n8297 vss.n7884 1118.26
R25012 vss.n7884 vss.n7879 1118.26
R25013 vss.n8691 vss.n8312 1118.26
R25014 vss.n8697 vss.n8312 1118.26
R25015 vss.n8697 vss.n8306 1118.26
R25016 vss.n8702 vss.n8306 1118.26
R25017 vss.n8702 vss.n8308 1118.26
R25018 vss.n8308 vss.n7867 1118.26
R25019 vss.n8692 vss.n8314 1118.26
R25020 vss.n8696 vss.n8314 1118.26
R25021 vss.n8696 vss.n7875 1118.26
R25022 vss.n8703 vss.n7875 1118.26
R25023 vss.n8703 vss.n7876 1118.26
R25024 vss.n7876 vss.n7868 1118.26
R25025 vss.n8324 vss.n8319 1118.26
R25026 vss.n8339 vss.n8319 1118.26
R25027 vss.n8339 vss.n8336 1118.26
R25028 vss.n8679 vss.n8336 1118.26
R25029 vss.n8679 vss.n8337 1118.26
R25030 vss.n8675 vss.n8337 1118.26
R25031 vss.n8326 vss.n8320 1118.26
R25032 vss.n8682 vss.n8320 1118.26
R25033 vss.n8682 vss.n8681 1118.26
R25034 vss.n8681 vss.n8680 1118.26
R25035 vss.n8680 vss.n8332 1118.26
R25036 vss.n8348 vss.n8332 1118.26
R25037 vss.n8650 vss.n8358 1118.26
R25038 vss.n8658 vss.n8358 1118.26
R25039 vss.n8658 vss.n8359 1118.26
R25040 vss.n8654 vss.n8359 1118.26
R25041 vss.n8654 vss.n8349 1118.26
R25042 vss.n8665 vss.n8349 1118.26
R25043 vss.n8649 vss.n8354 1118.26
R25044 vss.n8659 vss.n8354 1118.26
R25045 vss.n8660 vss.n8659 1118.26
R25046 vss.n8661 vss.n8660 1118.26
R25047 vss.n8661 vss.n8350 1118.26
R25048 vss.n8667 vss.n8350 1118.26
R25049 vss.n8369 vss.n8364 1118.26
R25050 vss.n8389 vss.n8364 1118.26
R25051 vss.n8389 vss.n8386 1118.26
R25052 vss.n8636 vss.n8386 1118.26
R25053 vss.n8636 vss.n8387 1118.26
R25054 vss.n8632 vss.n8387 1118.26
R25055 vss.n8371 vss.n8365 1118.26
R25056 vss.n8639 vss.n8365 1118.26
R25057 vss.n8639 vss.n8638 1118.26
R25058 vss.n8638 vss.n8637 1118.26
R25059 vss.n8637 vss.n8382 1118.26
R25060 vss.n8398 vss.n8382 1118.26
R25061 vss.n8606 vss.n8411 1118.26
R25062 vss.n8614 vss.n8411 1118.26
R25063 vss.n8614 vss.n8412 1118.26
R25064 vss.n8610 vss.n8412 1118.26
R25065 vss.n8610 vss.n8399 1118.26
R25066 vss.n8621 vss.n8399 1118.26
R25067 vss.n8605 vss.n8407 1118.26
R25068 vss.n8615 vss.n8407 1118.26
R25069 vss.n8616 vss.n8615 1118.26
R25070 vss.n8617 vss.n8616 1118.26
R25071 vss.n8617 vss.n8400 1118.26
R25072 vss.n8624 vss.n8400 1118.26
R25073 vss.n8422 vss.n8417 1118.26
R25074 vss.n8437 vss.n8417 1118.26
R25075 vss.n8437 vss.n8434 1118.26
R25076 vss.n8592 vss.n8434 1118.26
R25077 vss.n8592 vss.n8435 1118.26
R25078 vss.n8588 vss.n8435 1118.26
R25079 vss.n8424 vss.n8418 1118.26
R25080 vss.n8595 vss.n8418 1118.26
R25081 vss.n8595 vss.n8594 1118.26
R25082 vss.n8594 vss.n8593 1118.26
R25083 vss.n8593 vss.n8430 1118.26
R25084 vss.n8446 vss.n8430 1118.26
R25085 vss.n8563 vss.n8456 1118.26
R25086 vss.n8571 vss.n8456 1118.26
R25087 vss.n8571 vss.n8457 1118.26
R25088 vss.n8567 vss.n8457 1118.26
R25089 vss.n8567 vss.n8447 1118.26
R25090 vss.n8578 vss.n8447 1118.26
R25091 vss.n8562 vss.n8452 1118.26
R25092 vss.n8572 vss.n8452 1118.26
R25093 vss.n8573 vss.n8572 1118.26
R25094 vss.n8574 vss.n8573 1118.26
R25095 vss.n8574 vss.n8448 1118.26
R25096 vss.n8580 vss.n8448 1118.26
R25097 vss.n8467 vss.n8462 1118.26
R25098 vss.n8487 vss.n8462 1118.26
R25099 vss.n8487 vss.n8484 1118.26
R25100 vss.n8549 vss.n8484 1118.26
R25101 vss.n8549 vss.n8485 1118.26
R25102 vss.n8545 vss.n8485 1118.26
R25103 vss.n8469 vss.n8463 1118.26
R25104 vss.n8552 vss.n8463 1118.26
R25105 vss.n8552 vss.n8551 1118.26
R25106 vss.n8551 vss.n8550 1118.26
R25107 vss.n8550 vss.n8480 1118.26
R25108 vss.n8496 vss.n8480 1118.26
R25109 vss.n8523 vss.n8513 1118.26
R25110 vss.n8519 vss.n8513 1118.26
R25111 vss.n8519 vss.n8518 1118.26
R25112 vss.n8518 vss.n8517 1118.26
R25113 vss.n8517 vss.n8497 1118.26
R25114 vss.n8534 vss.n8497 1118.26
R25115 vss.n8524 vss.n8505 1118.26
R25116 vss.n8528 vss.n8505 1118.26
R25117 vss.n8529 vss.n8528 1118.26
R25118 vss.n8530 vss.n8529 1118.26
R25119 vss.n8530 vss.n8498 1118.26
R25120 vss.n8537 vss.n8498 1118.26
R25121 vss.n9556 vss.n9555 1118.26
R25122 vss.n9557 vss.n9556 1118.26
R25123 vss.n9557 vss.n6059 1118.26
R25124 vss.n9571 vss.n6059 1118.26
R25125 vss.n9571 vss.n6060 1118.26
R25126 vss.n9563 vss.n6060 1118.26
R25127 vss.n9554 vss.n6067 1118.26
R25128 vss.n9558 vss.n6067 1118.26
R25129 vss.n9558 vss.n6069 1118.26
R25130 vss.n6069 vss.n6062 1118.26
R25131 vss.n9568 vss.n6062 1118.26
R25132 vss.n9568 vss.n9567 1118.26
R25133 vss.n6087 vss.n6077 1118.26
R25134 vss.n9543 vss.n6087 1118.26
R25135 vss.n9543 vss.n6088 1118.26
R25136 vss.n7259 vss.n6088 1118.26
R25137 vss.n7259 vss.n7258 1118.26
R25138 vss.n7258 vss.n7248 1118.26
R25139 vss.n6082 vss.n6078 1118.26
R25140 vss.n9544 vss.n6082 1118.26
R25141 vss.n9544 vss.n6083 1118.26
R25142 vss.n7260 vss.n6083 1118.26
R25143 vss.n7260 vss.n7253 1118.26
R25144 vss.n7253 vss.n7249 1118.26
R25145 vss.n9521 vss.n9520 1118.26
R25146 vss.n9522 vss.n9521 1118.26
R25147 vss.n9522 vss.n6099 1118.26
R25148 vss.n9536 vss.n6099 1118.26
R25149 vss.n9536 vss.n6100 1118.26
R25150 vss.n9528 vss.n6100 1118.26
R25151 vss.n9519 vss.n6106 1118.26
R25152 vss.n9523 vss.n6106 1118.26
R25153 vss.n9523 vss.n6108 1118.26
R25154 vss.n6108 vss.n6102 1118.26
R25155 vss.n9533 vss.n6102 1118.26
R25156 vss.n9533 vss.n9532 1118.26
R25157 vss.n6126 vss.n6116 1118.26
R25158 vss.n9508 vss.n6126 1118.26
R25159 vss.n9508 vss.n6127 1118.26
R25160 vss.n7240 vss.n6127 1118.26
R25161 vss.n7240 vss.n7239 1118.26
R25162 vss.n7239 vss.n6575 1118.26
R25163 vss.n6121 vss.n6117 1118.26
R25164 vss.n9509 vss.n6121 1118.26
R25165 vss.n9509 vss.n6122 1118.26
R25166 vss.n7241 vss.n6122 1118.26
R25167 vss.n7241 vss.n6580 1118.26
R25168 vss.n6580 vss.n6576 1118.26
R25169 vss.n6762 vss.n6761 1118.26
R25170 vss.n6761 vss.n6760 1118.26
R25171 vss.n6760 vss.n6590 1118.26
R25172 vss.n7228 vss.n6590 1118.26
R25173 vss.n7228 vss.n6592 1118.26
R25174 vss.n6592 vss.n6581 1118.26
R25175 vss.n6752 vss.n6748 1118.26
R25176 vss.n6759 vss.n6752 1118.26
R25177 vss.n6759 vss.n6586 1118.26
R25178 vss.n7229 vss.n6586 1118.26
R25179 vss.n7229 vss.n6587 1118.26
R25180 vss.n6587 vss.n6582 1118.26
R25181 vss.n6766 vss.n6740 1118.26
R25182 vss.n6772 vss.n6740 1118.26
R25183 vss.n6772 vss.n6736 1118.26
R25184 vss.n6777 vss.n6736 1118.26
R25185 vss.n6777 vss.n6728 1118.26
R25186 vss.n6784 vss.n6728 1118.26
R25187 vss.n6767 vss.n6742 1118.26
R25188 vss.n6771 vss.n6742 1118.26
R25189 vss.n6771 vss.n6732 1118.26
R25190 vss.n6778 vss.n6732 1118.26
R25191 vss.n6778 vss.n6734 1118.26
R25192 vss.n6734 vss.n6727 1118.26
R25193 vss.n7066 vss.n7065 1118.26
R25194 vss.n7067 vss.n7066 1118.26
R25195 vss.n7067 vss.n6721 1118.26
R25196 vss.n7081 vss.n6721 1118.26
R25197 vss.n7081 vss.n6722 1118.26
R25198 vss.n7073 vss.n6722 1118.26
R25199 vss.n7064 vss.n6789 1118.26
R25200 vss.n7068 vss.n6789 1118.26
R25201 vss.n7068 vss.n6791 1118.26
R25202 vss.n6791 vss.n6724 1118.26
R25203 vss.n7078 vss.n6724 1118.26
R25204 vss.n7078 vss.n7077 1118.26
R25205 vss.n6808 vss.n6798 1118.26
R25206 vss.n7053 vss.n6808 1118.26
R25207 vss.n7053 vss.n6809 1118.26
R25208 vss.n7047 vss.n6809 1118.26
R25209 vss.n7047 vss.n6814 1118.26
R25210 vss.n6826 vss.n6814 1118.26
R25211 vss.n6803 vss.n6799 1118.26
R25212 vss.n7054 vss.n6803 1118.26
R25213 vss.n7054 vss.n6804 1118.26
R25214 vss.n6815 vss.n6804 1118.26
R25215 vss.n6817 vss.n6815 1118.26
R25216 vss.n6818 vss.n6817 1118.26
R25217 vss.n6895 vss.n6842 1118.26
R25218 vss.n6901 vss.n6842 1118.26
R25219 vss.n6901 vss.n6836 1118.26
R25220 vss.n7037 vss.n6836 1118.26
R25221 vss.n7037 vss.n6838 1118.26
R25222 vss.n6838 vss.n6827 1118.26
R25223 vss.n6896 vss.n6844 1118.26
R25224 vss.n6900 vss.n6844 1118.26
R25225 vss.n6900 vss.n6832 1118.26
R25226 vss.n7038 vss.n6832 1118.26
R25227 vss.n7038 vss.n6833 1118.26
R25228 vss.n6833 vss.n6828 1118.26
R25229 vss.n6859 vss.n6849 1118.26
R25230 vss.n6885 vss.n6859 1118.26
R25231 vss.n6885 vss.n6860 1118.26
R25232 vss.n6881 vss.n6860 1118.26
R25233 vss.n6881 vss.n6865 1118.26
R25234 vss.n6877 vss.n6865 1118.26
R25235 vss.n6854 vss.n6850 1118.26
R25236 vss.n6886 vss.n6854 1118.26
R25237 vss.n6886 vss.n6855 1118.26
R25238 vss.n6866 vss.n6855 1118.26
R25239 vss.n6868 vss.n6866 1118.26
R25240 vss.n6869 vss.n6868 1118.26
R25241 vss.n9229 vss.n9228 1118.26
R25242 vss.n9230 vss.n9229 1118.26
R25243 vss.n9230 vss.n6493 1118.26
R25244 vss.n9244 vss.n6493 1118.26
R25245 vss.n9244 vss.n6494 1118.26
R25246 vss.n9236 vss.n6494 1118.26
R25247 vss.n9227 vss.n6500 1118.26
R25248 vss.n9231 vss.n6500 1118.26
R25249 vss.n9231 vss.n6502 1118.26
R25250 vss.n6502 vss.n6496 1118.26
R25251 vss.n9241 vss.n6496 1118.26
R25252 vss.n9241 vss.n9240 1118.26
R25253 vss.n6519 vss.n6509 1118.26
R25254 vss.n9216 vss.n6519 1118.26
R25255 vss.n9216 vss.n6520 1118.26
R25256 vss.n9210 vss.n6520 1118.26
R25257 vss.n9210 vss.n6525 1118.26
R25258 vss.n6557 vss.n6525 1118.26
R25259 vss.n6514 vss.n6510 1118.26
R25260 vss.n9217 vss.n6514 1118.26
R25261 vss.n9217 vss.n6515 1118.26
R25262 vss.n6526 vss.n6515 1118.26
R25263 vss.n6558 vss.n6526 1118.26
R25264 vss.n6559 vss.n6558 1118.26
R25265 vss.n9080 vss.n9079 1118.26
R25266 vss.n9079 vss.n9078 1118.26
R25267 vss.n9078 vss.n6537 1118.26
R25268 vss.n9200 vss.n6537 1118.26
R25269 vss.n9200 vss.n6539 1118.26
R25270 vss.n6539 vss.n6528 1118.26
R25271 vss.n9070 vss.n9066 1118.26
R25272 vss.n9077 vss.n9070 1118.26
R25273 vss.n9077 vss.n6533 1118.26
R25274 vss.n9201 vss.n6533 1118.26
R25275 vss.n9201 vss.n6534 1118.26
R25276 vss.n6534 vss.n6529 1118.26
R25277 vss.n9087 vss.n9086 1118.26
R25278 vss.n9088 vss.n9087 1118.26
R25279 vss.n9088 vss.n6550 1118.26
R25280 vss.n9142 vss.n6550 1118.26
R25281 vss.n9142 vss.n6551 1118.26
R25282 vss.n9097 vss.n6551 1118.26
R25283 vss.n9085 vss.n9056 1118.26
R25284 vss.n9089 vss.n9056 1118.26
R25285 vss.n9089 vss.n9058 1118.26
R25286 vss.n9058 vss.n6553 1118.26
R25287 vss.n9051 vss.n6553 1118.26
R25288 vss.n9052 vss.n9051 1118.26
R25289 vss.n9121 vss.n9113 1118.26
R25290 vss.n9127 vss.n9113 1118.26
R25291 vss.n9127 vss.n9107 1118.26
R25292 vss.n9132 vss.n9107 1118.26
R25293 vss.n9132 vss.n9109 1118.26
R25294 vss.n9109 vss.n9098 1118.26
R25295 vss.n9122 vss.n9115 1118.26
R25296 vss.n9126 vss.n9115 1118.26
R25297 vss.n9126 vss.n9103 1118.26
R25298 vss.n9133 vss.n9103 1118.26
R25299 vss.n9133 vss.n9104 1118.26
R25300 vss.n9104 vss.n9099 1118.26
R25301 vss.n5957 vss.n5948 1118.26
R25302 vss.n5961 vss.n5948 1118.26
R25303 vss.n5961 vss.n5945 1118.26
R25304 vss.n9678 vss.n5945 1118.26
R25305 vss.n9678 vss.n5946 1118.26
R25306 vss.n9674 vss.n5946 1118.26
R25307 vss.n5959 vss.n5958 1118.26
R25308 vss.n5960 vss.n5959 1118.26
R25309 vss.n5960 vss.n5940 1118.26
R25310 vss.n9679 vss.n5940 1118.26
R25311 vss.n9679 vss.n5941 1118.26
R25312 vss.n5969 vss.n5941 1118.26
R25313 vss.n2754 vss.n2744 1118.26
R25314 vss.n9888 vss.n2754 1118.26
R25315 vss.n9888 vss.n2755 1118.26
R25316 vss.n9884 vss.n2755 1118.26
R25317 vss.n9884 vss.n2760 1118.26
R25318 vss.n2766 vss.n2760 1118.26
R25319 vss.n2749 vss.n2745 1118.26
R25320 vss.n9889 vss.n2749 1118.26
R25321 vss.n9889 vss.n2750 1118.26
R25322 vss.n2761 vss.n2750 1118.26
R25323 vss.n2762 vss.n2761 1118.26
R25324 vss.n9878 vss.n2762 1118.26
R25325 vss.n9707 vss.n9696 1118.26
R25326 vss.n9711 vss.n9696 1118.26
R25327 vss.n9711 vss.n9693 1118.26
R25328 vss.n9725 vss.n9693 1118.26
R25329 vss.n9725 vss.n9694 1118.26
R25330 vss.n9721 vss.n9694 1118.26
R25331 vss.n9709 vss.n9708 1118.26
R25332 vss.n9710 vss.n9709 1118.26
R25333 vss.n9710 vss.n9688 1118.26
R25334 vss.n9726 vss.n9688 1118.26
R25335 vss.n9726 vss.n9689 1118.26
R25336 vss.n9719 vss.n9689 1118.26
R25337 vss.n3285 vss.n3274 1118.26
R25338 vss.n3289 vss.n3274 1118.26
R25339 vss.n3289 vss.n3271 1118.26
R25340 vss.n3303 vss.n3271 1118.26
R25341 vss.n3303 vss.n3272 1118.26
R25342 vss.n3299 vss.n3272 1118.26
R25343 vss.n3287 vss.n3286 1118.26
R25344 vss.n3288 vss.n3287 1118.26
R25345 vss.n3288 vss.n3266 1118.26
R25346 vss.n3304 vss.n3266 1118.26
R25347 vss.n3304 vss.n3267 1118.26
R25348 vss.n3298 vss.n3267 1118.26
R25349 vss.n2578 vss.n2569 1118.26
R25350 vss.n2582 vss.n2569 1118.26
R25351 vss.n2582 vss.n2566 1118.26
R25352 vss.n10006 vss.n2566 1118.26
R25353 vss.n10006 vss.n2567 1118.26
R25354 vss.n10002 vss.n2567 1118.26
R25355 vss.n2580 vss.n2579 1118.26
R25356 vss.n2581 vss.n2580 1118.26
R25357 vss.n2581 vss.n2561 1118.26
R25358 vss.n10007 vss.n2561 1118.26
R25359 vss.n10007 vss.n2562 1118.26
R25360 vss.n2590 vss.n2562 1118.26
R25361 vss.n5910 vss.n5900 1118.26
R25362 vss.n5914 vss.n5900 1118.26
R25363 vss.n5914 vss.n5897 1118.26
R25364 vss.n5927 vss.n5897 1118.26
R25365 vss.n5927 vss.n5898 1118.26
R25366 vss.n5923 vss.n5898 1118.26
R25367 vss.n5912 vss.n5911 1118.26
R25368 vss.n5913 vss.n5912 1118.26
R25369 vss.n5913 vss.n5892 1118.26
R25370 vss.n5928 vss.n5892 1118.26
R25371 vss.n5928 vss.n5893 1118.26
R25372 vss.n5921 vss.n5893 1118.26
R25373 vss.n9761 vss.n9755 1118.26
R25374 vss.n9770 vss.n9755 1118.26
R25375 vss.n9770 vss.n9753 1118.26
R25376 vss.n9774 vss.n9753 1118.26
R25377 vss.n9775 vss.n9774 1118.26
R25378 vss.n9776 vss.n9775 1118.26
R25379 vss.n9768 vss.n9767 1118.26
R25380 vss.n9769 vss.n9768 1118.26
R25381 vss.n9769 vss.n9747 1118.26
R25382 vss.n9782 vss.n9747 1118.26
R25383 vss.n9782 vss.n9781 1118.26
R25384 vss.n9781 vss.n9780 1118.26
R25385 vss.n3201 vss.n3195 1118.26
R25386 vss.n3210 vss.n3195 1118.26
R25387 vss.n3210 vss.n3193 1118.26
R25388 vss.n3214 vss.n3193 1118.26
R25389 vss.n3215 vss.n3214 1118.26
R25390 vss.n3216 vss.n3215 1118.26
R25391 vss.n3208 vss.n3207 1118.26
R25392 vss.n3209 vss.n3208 1118.26
R25393 vss.n3209 vss.n3187 1118.26
R25394 vss.n3222 vss.n3187 1118.26
R25395 vss.n3222 vss.n3221 1118.26
R25396 vss.n3221 vss.n3220 1118.26
R25397 vss.n9801 vss.n2996 1118.26
R25398 vss.n9797 vss.n2996 1118.26
R25399 vss.n9797 vss.n3000 1118.26
R25400 vss.n3016 vss.n3000 1118.26
R25401 vss.n3017 vss.n3016 1118.26
R25402 vss.n3018 vss.n3017 1118.26
R25403 vss.n3003 vss.n2995 1118.26
R25404 vss.n9796 vss.n3003 1118.26
R25405 vss.n9796 vss.n3004 1118.26
R25406 vss.n3024 vss.n3004 1118.26
R25407 vss.n3024 vss.n3023 1118.26
R25408 vss.n3023 vss.n3022 1118.26
R25409 vss.n5231 vss.n5225 1118.26
R25410 vss.n5240 vss.n5225 1118.26
R25411 vss.n5240 vss.n5223 1118.26
R25412 vss.n5244 vss.n5223 1118.26
R25413 vss.n5245 vss.n5244 1118.26
R25414 vss.n5246 vss.n5245 1118.26
R25415 vss.n5238 vss.n5237 1118.26
R25416 vss.n5239 vss.n5238 1118.26
R25417 vss.n5239 vss.n5217 1118.26
R25418 vss.n5252 vss.n5217 1118.26
R25419 vss.n5252 vss.n5251 1118.26
R25420 vss.n5251 vss.n5250 1118.26
R25421 vss.n3044 vss.n3038 1118.26
R25422 vss.n3053 vss.n3038 1118.26
R25423 vss.n3053 vss.n3036 1118.26
R25424 vss.n3057 vss.n3036 1118.26
R25425 vss.n3058 vss.n3057 1118.26
R25426 vss.n3059 vss.n3058 1118.26
R25427 vss.n3051 vss.n3050 1118.26
R25428 vss.n3052 vss.n3051 1118.26
R25429 vss.n3052 vss.n3030 1118.26
R25430 vss.n3065 vss.n3030 1118.26
R25431 vss.n3065 vss.n3064 1118.26
R25432 vss.n3064 vss.n3063 1118.26
R25433 vss.n5101 vss.n5095 1118.26
R25434 vss.n5110 vss.n5095 1118.26
R25435 vss.n5110 vss.n5093 1118.26
R25436 vss.n5114 vss.n5093 1118.26
R25437 vss.n5115 vss.n5114 1118.26
R25438 vss.n5116 vss.n5115 1118.26
R25439 vss.n5108 vss.n5107 1118.26
R25440 vss.n5109 vss.n5108 1118.26
R25441 vss.n5109 vss.n5087 1118.26
R25442 vss.n5122 vss.n5087 1118.26
R25443 vss.n5122 vss.n5121 1118.26
R25444 vss.n5121 vss.n5120 1118.26
R25445 vss.n5290 vss.n5284 1118.26
R25446 vss.n5299 vss.n5284 1118.26
R25447 vss.n5299 vss.n5282 1118.26
R25448 vss.n5303 vss.n5282 1118.26
R25449 vss.n5304 vss.n5303 1118.26
R25450 vss.n5305 vss.n5304 1118.26
R25451 vss.n5297 vss.n5296 1118.26
R25452 vss.n5298 vss.n5297 1118.26
R25453 vss.n5298 vss.n5276 1118.26
R25454 vss.n5311 vss.n5276 1118.26
R25455 vss.n5311 vss.n5310 1118.26
R25456 vss.n5310 vss.n5309 1118.26
R25457 vss.n5018 vss.n5012 1118.26
R25458 vss.n5027 vss.n5012 1118.26
R25459 vss.n5027 vss.n5010 1118.26
R25460 vss.n5031 vss.n5010 1118.26
R25461 vss.n5032 vss.n5031 1118.26
R25462 vss.n5033 vss.n5032 1118.26
R25463 vss.n5025 vss.n5024 1118.26
R25464 vss.n5026 vss.n5025 1118.26
R25465 vss.n5026 vss.n5004 1118.26
R25466 vss.n5039 vss.n5004 1118.26
R25467 vss.n5039 vss.n5038 1118.26
R25468 vss.n5038 vss.n5037 1118.26
R25469 vss.n4899 vss.n4893 1118.26
R25470 vss.n4908 vss.n4893 1118.26
R25471 vss.n4908 vss.n4891 1118.26
R25472 vss.n4912 vss.n4891 1118.26
R25473 vss.n4913 vss.n4912 1118.26
R25474 vss.n4914 vss.n4913 1118.26
R25475 vss.n4906 vss.n4905 1118.26
R25476 vss.n4907 vss.n4906 1118.26
R25477 vss.n4907 vss.n4885 1118.26
R25478 vss.n4920 vss.n4885 1118.26
R25479 vss.n4920 vss.n4919 1118.26
R25480 vss.n4919 vss.n4918 1118.26
R25481 vss.n2719 vss.n2709 1118.26
R25482 vss.n9922 vss.n2719 1118.26
R25483 vss.n9922 vss.n2720 1118.26
R25484 vss.n9918 vss.n2720 1118.26
R25485 vss.n9918 vss.n2725 1118.26
R25486 vss.n2731 vss.n2725 1118.26
R25487 vss.n2714 vss.n2710 1118.26
R25488 vss.n9923 vss.n2714 1118.26
R25489 vss.n9923 vss.n2715 1118.26
R25490 vss.n2726 vss.n2715 1118.26
R25491 vss.n2727 vss.n2726 1118.26
R25492 vss.n9912 vss.n2727 1118.26
R25493 vss.n4650 vss.n4637 1118.26
R25494 vss.n4659 vss.n4650 1118.26
R25495 vss.n4659 vss.n4651 1118.26
R25496 vss.n4655 vss.n4651 1118.26
R25497 vss.n4655 vss.n2732 1118.26
R25498 vss.n2738 vss.n2732 1118.26
R25499 vss.n4644 vss.n4638 1118.26
R25500 vss.n4660 vss.n4644 1118.26
R25501 vss.n4660 vss.n4646 1118.26
R25502 vss.n4646 vss.n4645 1118.26
R25503 vss.n4645 vss.n2733 1118.26
R25504 vss.n9903 vss.n2733 1118.26
R25505 vss.n4671 vss.n4628 1118.26
R25506 vss.n5624 vss.n4671 1118.26
R25507 vss.n5624 vss.n4672 1118.26
R25508 vss.n5620 vss.n4672 1118.26
R25509 vss.n5620 vss.n4677 1118.26
R25510 vss.n4683 vss.n4677 1118.26
R25511 vss.n4635 vss.n4629 1118.26
R25512 vss.n5625 vss.n4635 1118.26
R25513 vss.n5625 vss.n4636 1118.26
R25514 vss.n4678 vss.n4636 1118.26
R25515 vss.n4679 vss.n4678 1118.26
R25516 vss.n5614 vss.n4679 1118.26
R25517 vss.n5588 vss.n4693 1118.26
R25518 vss.n5596 vss.n4693 1118.26
R25519 vss.n5596 vss.n4694 1118.26
R25520 vss.n5592 vss.n4694 1118.26
R25521 vss.n5592 vss.n4684 1118.26
R25522 vss.n5603 vss.n4684 1118.26
R25523 vss.n5587 vss.n4689 1118.26
R25524 vss.n5597 vss.n4689 1118.26
R25525 vss.n5598 vss.n5597 1118.26
R25526 vss.n5599 vss.n5598 1118.26
R25527 vss.n5599 vss.n4685 1118.26
R25528 vss.n5605 vss.n4685 1118.26
R25529 vss.n4704 vss.n4699 1118.26
R25530 vss.n4717 vss.n4699 1118.26
R25531 vss.n4717 vss.n4714 1118.26
R25532 vss.n5574 vss.n4714 1118.26
R25533 vss.n5574 vss.n4715 1118.26
R25534 vss.n5570 vss.n4715 1118.26
R25535 vss.n4706 vss.n4700 1118.26
R25536 vss.n5577 vss.n4700 1118.26
R25537 vss.n5577 vss.n5576 1118.26
R25538 vss.n5576 vss.n5575 1118.26
R25539 vss.n5575 vss.n4710 1118.26
R25540 vss.n4726 vss.n4710 1118.26
R25541 vss.n5545 vss.n4736 1118.26
R25542 vss.n5553 vss.n4736 1118.26
R25543 vss.n5553 vss.n4737 1118.26
R25544 vss.n5549 vss.n4737 1118.26
R25545 vss.n5549 vss.n4727 1118.26
R25546 vss.n5560 vss.n4727 1118.26
R25547 vss.n5544 vss.n4732 1118.26
R25548 vss.n5554 vss.n4732 1118.26
R25549 vss.n5555 vss.n5554 1118.26
R25550 vss.n5556 vss.n5555 1118.26
R25551 vss.n5556 vss.n4728 1118.26
R25552 vss.n5562 vss.n4728 1118.26
R25553 vss.n4747 vss.n4742 1118.26
R25554 vss.n4760 vss.n4742 1118.26
R25555 vss.n4760 vss.n4757 1118.26
R25556 vss.n5531 vss.n4757 1118.26
R25557 vss.n5531 vss.n4758 1118.26
R25558 vss.n5527 vss.n4758 1118.26
R25559 vss.n4749 vss.n4743 1118.26
R25560 vss.n5534 vss.n4743 1118.26
R25561 vss.n5534 vss.n5533 1118.26
R25562 vss.n5533 vss.n5532 1118.26
R25563 vss.n5532 vss.n4753 1118.26
R25564 vss.n4769 vss.n4753 1118.26
R25565 vss.n5502 vss.n4779 1118.26
R25566 vss.n5510 vss.n4779 1118.26
R25567 vss.n5510 vss.n4780 1118.26
R25568 vss.n5506 vss.n4780 1118.26
R25569 vss.n5506 vss.n4770 1118.26
R25570 vss.n5517 vss.n4770 1118.26
R25571 vss.n5501 vss.n4775 1118.26
R25572 vss.n5511 vss.n4775 1118.26
R25573 vss.n5512 vss.n5511 1118.26
R25574 vss.n5513 vss.n5512 1118.26
R25575 vss.n5513 vss.n4771 1118.26
R25576 vss.n5519 vss.n4771 1118.26
R25577 vss.n4790 vss.n4785 1118.26
R25578 vss.n4803 vss.n4785 1118.26
R25579 vss.n4803 vss.n4800 1118.26
R25580 vss.n5488 vss.n4800 1118.26
R25581 vss.n5488 vss.n4801 1118.26
R25582 vss.n5484 vss.n4801 1118.26
R25583 vss.n4792 vss.n4786 1118.26
R25584 vss.n5491 vss.n4786 1118.26
R25585 vss.n5491 vss.n5490 1118.26
R25586 vss.n5490 vss.n5489 1118.26
R25587 vss.n5489 vss.n4796 1118.26
R25588 vss.n4812 vss.n4796 1118.26
R25589 vss.n5459 vss.n4822 1118.26
R25590 vss.n5467 vss.n4822 1118.26
R25591 vss.n5467 vss.n4823 1118.26
R25592 vss.n5463 vss.n4823 1118.26
R25593 vss.n5463 vss.n4813 1118.26
R25594 vss.n5474 vss.n4813 1118.26
R25595 vss.n5458 vss.n4818 1118.26
R25596 vss.n5468 vss.n4818 1118.26
R25597 vss.n5469 vss.n5468 1118.26
R25598 vss.n5470 vss.n5469 1118.26
R25599 vss.n5470 vss.n4814 1118.26
R25600 vss.n5476 vss.n4814 1118.26
R25601 vss.n4833 vss.n4828 1118.26
R25602 vss.n4846 vss.n4828 1118.26
R25603 vss.n4846 vss.n4843 1118.26
R25604 vss.n5445 vss.n4843 1118.26
R25605 vss.n5445 vss.n4844 1118.26
R25606 vss.n5441 vss.n4844 1118.26
R25607 vss.n4835 vss.n4829 1118.26
R25608 vss.n5448 vss.n4829 1118.26
R25609 vss.n5448 vss.n5447 1118.26
R25610 vss.n5447 vss.n5446 1118.26
R25611 vss.n5446 vss.n4839 1118.26
R25612 vss.n4855 vss.n4839 1118.26
R25613 vss.n5416 vss.n4865 1118.26
R25614 vss.n5424 vss.n4865 1118.26
R25615 vss.n5424 vss.n4866 1118.26
R25616 vss.n5420 vss.n4866 1118.26
R25617 vss.n5420 vss.n4856 1118.26
R25618 vss.n5431 vss.n4856 1118.26
R25619 vss.n5415 vss.n4861 1118.26
R25620 vss.n5425 vss.n4861 1118.26
R25621 vss.n5426 vss.n5425 1118.26
R25622 vss.n5427 vss.n5426 1118.26
R25623 vss.n5427 vss.n4857 1118.26
R25624 vss.n5433 vss.n4857 1118.26
R25625 vss.n4876 vss.n4871 1118.26
R25626 vss.n5340 vss.n4871 1118.26
R25627 vss.n5340 vss.n5337 1118.26
R25628 vss.n5402 vss.n5337 1118.26
R25629 vss.n5402 vss.n5338 1118.26
R25630 vss.n5398 vss.n5338 1118.26
R25631 vss.n4878 vss.n4872 1118.26
R25632 vss.n5405 vss.n4872 1118.26
R25633 vss.n5405 vss.n5404 1118.26
R25634 vss.n5404 vss.n5403 1118.26
R25635 vss.n5403 vss.n5333 1118.26
R25636 vss.n5349 vss.n5333 1118.26
R25637 vss.n5376 vss.n5366 1118.26
R25638 vss.n5372 vss.n5366 1118.26
R25639 vss.n5372 vss.n5371 1118.26
R25640 vss.n5371 vss.n5370 1118.26
R25641 vss.n5370 vss.n5350 1118.26
R25642 vss.n5387 vss.n5350 1118.26
R25643 vss.n5377 vss.n5358 1118.26
R25644 vss.n5381 vss.n5358 1118.26
R25645 vss.n5382 vss.n5381 1118.26
R25646 vss.n5383 vss.n5382 1118.26
R25647 vss.n5383 vss.n5351 1118.26
R25648 vss.n5390 vss.n5351 1118.26
R25649 vss.n9820 vss.n2883 1118.26
R25650 vss.n9829 vss.n2883 1118.26
R25651 vss.n9829 vss.n2881 1118.26
R25652 vss.n9833 vss.n2881 1118.26
R25653 vss.n9834 vss.n9833 1118.26
R25654 vss.n9835 vss.n9834 1118.26
R25655 vss.n9827 vss.n9826 1118.26
R25656 vss.n9828 vss.n9827 1118.26
R25657 vss.n9828 vss.n2875 1118.26
R25658 vss.n9841 vss.n2875 1118.26
R25659 vss.n9841 vss.n9840 1118.26
R25660 vss.n9840 vss.n9839 1118.26
R25661 vss.n2978 vss.n2939 1118.26
R25662 vss.n2974 vss.n2939 1118.26
R25663 vss.n2974 vss.n2943 1118.26
R25664 vss.n2959 vss.n2943 1118.26
R25665 vss.n2960 vss.n2959 1118.26
R25666 vss.n2961 vss.n2960 1118.26
R25667 vss.n2946 vss.n2938 1118.26
R25668 vss.n2973 vss.n2946 1118.26
R25669 vss.n2973 vss.n2947 1118.26
R25670 vss.n2967 vss.n2947 1118.26
R25671 vss.n2967 vss.n2966 1118.26
R25672 vss.n2966 vss.n2965 1118.26
R25673 vss.n2932 vss.n2892 1118.26
R25674 vss.n2928 vss.n2892 1118.26
R25675 vss.n2928 vss.n2896 1118.26
R25676 vss.n2912 vss.n2896 1118.26
R25677 vss.n2913 vss.n2912 1118.26
R25678 vss.n2914 vss.n2913 1118.26
R25679 vss.n2899 vss.n2891 1118.26
R25680 vss.n2927 vss.n2899 1118.26
R25681 vss.n2927 vss.n2900 1118.26
R25682 vss.n2920 vss.n2900 1118.26
R25683 vss.n2920 vss.n2919 1118.26
R25684 vss.n2919 vss.n2918 1118.26
R25685 vss.n4940 vss.n4934 1118.26
R25686 vss.n4949 vss.n4934 1118.26
R25687 vss.n4949 vss.n4932 1118.26
R25688 vss.n4953 vss.n4932 1118.26
R25689 vss.n4954 vss.n4953 1118.26
R25690 vss.n4955 vss.n4954 1118.26
R25691 vss.n4947 vss.n4946 1118.26
R25692 vss.n4948 vss.n4947 1118.26
R25693 vss.n4948 vss.n4926 1118.26
R25694 vss.n4961 vss.n4926 1118.26
R25695 vss.n4961 vss.n4960 1118.26
R25696 vss.n4960 vss.n4959 1118.26
R25697 vss.n5142 vss.n5136 1118.26
R25698 vss.n5151 vss.n5136 1118.26
R25699 vss.n5151 vss.n5134 1118.26
R25700 vss.n5155 vss.n5134 1118.26
R25701 vss.n5156 vss.n5155 1118.26
R25702 vss.n5157 vss.n5156 1118.26
R25703 vss.n5149 vss.n5148 1118.26
R25704 vss.n5150 vss.n5149 1118.26
R25705 vss.n5150 vss.n5128 1118.26
R25706 vss.n5163 vss.n5128 1118.26
R25707 vss.n5163 vss.n5162 1118.26
R25708 vss.n5162 vss.n5161 1118.26
R25709 vss.n3123 vss.n3116 1118.26
R25710 vss.n3132 vss.n3116 1118.26
R25711 vss.n3132 vss.n3114 1118.26
R25712 vss.n3136 vss.n3114 1118.26
R25713 vss.n3137 vss.n3136 1118.26
R25714 vss.n3138 vss.n3137 1118.26
R25715 vss.n3130 vss.n3129 1118.26
R25716 vss.n3131 vss.n3130 1118.26
R25717 vss.n3131 vss.n3108 1118.26
R25718 vss.n3144 vss.n3108 1118.26
R25719 vss.n3144 vss.n3143 1118.26
R25720 vss.n3143 vss.n3142 1118.26
R25721 vss.n4485 vss.n4484 1118.26
R25722 vss.n4486 vss.n4485 1118.26
R25723 vss.n4486 vss.n4464 1118.26
R25724 vss.n4500 vss.n4464 1118.26
R25725 vss.n4500 vss.n4465 1118.26
R25726 vss.n4492 vss.n4465 1118.26
R25727 vss.n4483 vss.n4471 1118.26
R25728 vss.n4487 vss.n4471 1118.26
R25729 vss.n4487 vss.n4473 1118.26
R25730 vss.n4473 vss.n4467 1118.26
R25731 vss.n4497 vss.n4467 1118.26
R25732 vss.n4497 vss.n4496 1118.26
R25733 vss.n4393 vss.n4392 1118.26
R25734 vss.n4394 vss.n4393 1118.26
R25735 vss.n4394 vss.n4372 1118.26
R25736 vss.n4408 vss.n4372 1118.26
R25737 vss.n4408 vss.n4373 1118.26
R25738 vss.n4400 vss.n4373 1118.26
R25739 vss.n4391 vss.n4379 1118.26
R25740 vss.n4395 vss.n4379 1118.26
R25741 vss.n4395 vss.n4381 1118.26
R25742 vss.n4381 vss.n4375 1118.26
R25743 vss.n4405 vss.n4375 1118.26
R25744 vss.n4405 vss.n4404 1118.26
R25745 vss.n4345 vss.n4344 1118.26
R25746 vss.n4346 vss.n4345 1118.26
R25747 vss.n4346 vss.n4324 1118.26
R25748 vss.n4360 vss.n4324 1118.26
R25749 vss.n4360 vss.n4325 1118.26
R25750 vss.n4352 vss.n4325 1118.26
R25751 vss.n4343 vss.n4331 1118.26
R25752 vss.n4347 vss.n4331 1118.26
R25753 vss.n4347 vss.n4333 1118.26
R25754 vss.n4333 vss.n4327 1118.26
R25755 vss.n4357 vss.n4327 1118.26
R25756 vss.n4357 vss.n4356 1118.26
R25757 vss.n3745 vss.n3744 1118.26
R25758 vss.n3746 vss.n3745 1118.26
R25759 vss.n3746 vss.n3724 1118.26
R25760 vss.n3760 vss.n3724 1118.26
R25761 vss.n3760 vss.n3725 1118.26
R25762 vss.n3752 vss.n3725 1118.26
R25763 vss.n3743 vss.n3731 1118.26
R25764 vss.n3747 vss.n3731 1118.26
R25765 vss.n3747 vss.n3733 1118.26
R25766 vss.n3733 vss.n3727 1118.26
R25767 vss.n3757 vss.n3727 1118.26
R25768 vss.n3757 vss.n3756 1118.26
R25769 vss.n4047 vss.n4046 1118.26
R25770 vss.n4048 vss.n4047 1118.26
R25771 vss.n4048 vss.n4026 1118.26
R25772 vss.n4062 vss.n4026 1118.26
R25773 vss.n4062 vss.n4027 1118.26
R25774 vss.n4054 vss.n4027 1118.26
R25775 vss.n4045 vss.n4033 1118.26
R25776 vss.n4049 vss.n4033 1118.26
R25777 vss.n4049 vss.n4035 1118.26
R25778 vss.n4035 vss.n4029 1118.26
R25779 vss.n4059 vss.n4029 1118.26
R25780 vss.n4059 vss.n4058 1118.26
R25781 vss.n3700 vss.n3699 1118.26
R25782 vss.n3701 vss.n3700 1118.26
R25783 vss.n3701 vss.n3679 1118.26
R25784 vss.n3715 vss.n3679 1118.26
R25785 vss.n3715 vss.n3680 1118.26
R25786 vss.n3707 vss.n3680 1118.26
R25787 vss.n3698 vss.n3686 1118.26
R25788 vss.n3702 vss.n3686 1118.26
R25789 vss.n3702 vss.n3688 1118.26
R25790 vss.n3688 vss.n3682 1118.26
R25791 vss.n3712 vss.n3682 1118.26
R25792 vss.n3712 vss.n3711 1118.26
R25793 vss.n4101 vss.n4100 1118.26
R25794 vss.n4102 vss.n4101 1118.26
R25795 vss.n4102 vss.n4080 1118.26
R25796 vss.n4116 vss.n4080 1118.26
R25797 vss.n4116 vss.n4081 1118.26
R25798 vss.n4108 vss.n4081 1118.26
R25799 vss.n4099 vss.n4087 1118.26
R25800 vss.n4103 vss.n4087 1118.26
R25801 vss.n4103 vss.n4089 1118.26
R25802 vss.n4089 vss.n4083 1118.26
R25803 vss.n4113 vss.n4083 1118.26
R25804 vss.n4113 vss.n4112 1118.26
R25805 vss.n3525 vss.n3524 1118.26
R25806 vss.n3526 vss.n3525 1118.26
R25807 vss.n3526 vss.n3504 1118.26
R25808 vss.n3540 vss.n3504 1118.26
R25809 vss.n3540 vss.n3505 1118.26
R25810 vss.n3532 vss.n3505 1118.26
R25811 vss.n3523 vss.n3511 1118.26
R25812 vss.n3527 vss.n3511 1118.26
R25813 vss.n3527 vss.n3513 1118.26
R25814 vss.n3513 vss.n3507 1118.26
R25815 vss.n3537 vss.n3507 1118.26
R25816 vss.n3537 vss.n3536 1118.26
R25817 vss.n3480 vss.n3479 1118.26
R25818 vss.n3481 vss.n3480 1118.26
R25819 vss.n3481 vss.n3459 1118.26
R25820 vss.n3495 vss.n3459 1118.26
R25821 vss.n3495 vss.n3460 1118.26
R25822 vss.n3487 vss.n3460 1118.26
R25823 vss.n3478 vss.n3466 1118.26
R25824 vss.n3482 vss.n3466 1118.26
R25825 vss.n3482 vss.n3468 1118.26
R25826 vss.n3468 vss.n3462 1118.26
R25827 vss.n3492 vss.n3462 1118.26
R25828 vss.n3492 vss.n3491 1118.26
R25829 vss.n5768 vss.n5767 1118.26
R25830 vss.n5769 vss.n5768 1118.26
R25831 vss.n5769 vss.n5747 1118.26
R25832 vss.n5783 vss.n5747 1118.26
R25833 vss.n5783 vss.n5748 1118.26
R25834 vss.n5775 vss.n5748 1118.26
R25835 vss.n5766 vss.n5754 1118.26
R25836 vss.n5770 vss.n5754 1118.26
R25837 vss.n5770 vss.n5756 1118.26
R25838 vss.n5756 vss.n5750 1118.26
R25839 vss.n5780 vss.n5750 1118.26
R25840 vss.n5780 vss.n5779 1118.26
R25841 vss.n4534 vss.n4533 1118.26
R25842 vss.n4533 vss.n4532 1118.26
R25843 vss.n4532 vss.n4448 1118.26
R25844 vss.n4530 vss.n4448 1118.26
R25845 vss.n4530 vss.n4456 1118.26
R25846 vss.n4526 vss.n4456 1118.26
R25847 vss.n4450 vss.n4444 1118.26
R25848 vss.n4451 vss.n4450 1118.26
R25849 vss.n4453 vss.n4451 1118.26
R25850 vss.n4454 vss.n4453 1118.26
R25851 vss.n4513 vss.n4454 1118.26
R25852 vss.n4525 vss.n4513 1118.26
R25853 vss.n4538 vss.n4436 1118.26
R25854 vss.n4544 vss.n4436 1118.26
R25855 vss.n4544 vss.n4432 1118.26
R25856 vss.n4549 vss.n4432 1118.26
R25857 vss.n4549 vss.n4424 1118.26
R25858 vss.n4556 vss.n4424 1118.26
R25859 vss.n4539 vss.n4438 1118.26
R25860 vss.n4543 vss.n4438 1118.26
R25861 vss.n4543 vss.n4428 1118.26
R25862 vss.n4550 vss.n4428 1118.26
R25863 vss.n4550 vss.n4430 1118.26
R25864 vss.n4430 vss.n4423 1118.26
R25865 vss.n4592 vss.n4591 1118.26
R25866 vss.n4593 vss.n4592 1118.26
R25867 vss.n4593 vss.n4416 1118.26
R25868 vss.n4607 vss.n4416 1118.26
R25869 vss.n4607 vss.n4417 1118.26
R25870 vss.n4599 vss.n4417 1118.26
R25871 vss.n4590 vss.n4561 1118.26
R25872 vss.n4594 vss.n4561 1118.26
R25873 vss.n4594 vss.n4563 1118.26
R25874 vss.n4563 vss.n4419 1118.26
R25875 vss.n4604 vss.n4419 1118.26
R25876 vss.n4604 vss.n4603 1118.26
R25877 vss.n4578 vss.n4570 1118.26
R25878 vss.n4579 vss.n4578 1118.26
R25879 vss.n4579 vss.n3640 1118.26
R25880 vss.n4620 vss.n3640 1118.26
R25881 vss.n4620 vss.n3642 1118.26
R25882 vss.n3642 vss.n3631 1118.26
R25883 vss.n4575 vss.n4571 1118.26
R25884 vss.n4580 vss.n4575 1118.26
R25885 vss.n4580 vss.n3636 1118.26
R25886 vss.n4621 vss.n3636 1118.26
R25887 vss.n4621 vss.n3637 1118.26
R25888 vss.n3637 vss.n3632 1118.26
R25889 vss.n4189 vss.n4188 1118.26
R25890 vss.n4190 vss.n4189 1118.26
R25891 vss.n4190 vss.n3766 1118.26
R25892 vss.n4204 vss.n3766 1118.26
R25893 vss.n4204 vss.n3767 1118.26
R25894 vss.n4196 vss.n3767 1118.26
R25895 vss.n4187 vss.n3775 1118.26
R25896 vss.n4191 vss.n3775 1118.26
R25897 vss.n4191 vss.n3777 1118.26
R25898 vss.n3777 vss.n3769 1118.26
R25899 vss.n4201 vss.n3769 1118.26
R25900 vss.n4201 vss.n4200 1118.26
R25901 vss.n3794 vss.n3784 1118.26
R25902 vss.n4176 vss.n3794 1118.26
R25903 vss.n4176 vss.n3795 1118.26
R25904 vss.n3819 vss.n3795 1118.26
R25905 vss.n3819 vss.n3813 1118.26
R25906 vss.n3826 vss.n3813 1118.26
R25907 vss.n3789 vss.n3785 1118.26
R25908 vss.n4177 vss.n3789 1118.26
R25909 vss.n4177 vss.n3790 1118.26
R25910 vss.n3820 vss.n3790 1118.26
R25911 vss.n3820 vss.n3818 1118.26
R25912 vss.n3818 vss.n3812 1118.26
R25913 vss.n4154 vss.n4153 1118.26
R25914 vss.n4155 vss.n4154 1118.26
R25915 vss.n4155 vss.n3806 1118.26
R25916 vss.n4169 vss.n3806 1118.26
R25917 vss.n4169 vss.n3807 1118.26
R25918 vss.n4161 vss.n3807 1118.26
R25919 vss.n4152 vss.n3831 1118.26
R25920 vss.n4156 vss.n3831 1118.26
R25921 vss.n4156 vss.n3833 1118.26
R25922 vss.n3833 vss.n3809 1118.26
R25923 vss.n4166 vss.n3809 1118.26
R25924 vss.n4166 vss.n4165 1118.26
R25925 vss.n3850 vss.n3840 1118.26
R25926 vss.n4141 vss.n3850 1118.26
R25927 vss.n4141 vss.n3851 1118.26
R25928 vss.n4137 vss.n3851 1118.26
R25929 vss.n4137 vss.n3857 1118.26
R25930 vss.n3869 vss.n3857 1118.26
R25931 vss.n3845 vss.n3841 1118.26
R25932 vss.n4142 vss.n3845 1118.26
R25933 vss.n4142 vss.n3846 1118.26
R25934 vss.n3858 vss.n3846 1118.26
R25935 vss.n3860 vss.n3858 1118.26
R25936 vss.n3861 vss.n3860 1118.26
R25937 vss.n3938 vss.n3885 1118.26
R25938 vss.n3944 vss.n3885 1118.26
R25939 vss.n3944 vss.n3879 1118.26
R25940 vss.n4127 vss.n3879 1118.26
R25941 vss.n4127 vss.n3881 1118.26
R25942 vss.n3881 vss.n3870 1118.26
R25943 vss.n3939 vss.n3887 1118.26
R25944 vss.n3943 vss.n3887 1118.26
R25945 vss.n3943 vss.n3875 1118.26
R25946 vss.n4128 vss.n3875 1118.26
R25947 vss.n4128 vss.n3876 1118.26
R25948 vss.n3876 vss.n3871 1118.26
R25949 vss.n3902 vss.n3892 1118.26
R25950 vss.n3928 vss.n3902 1118.26
R25951 vss.n3928 vss.n3903 1118.26
R25952 vss.n3924 vss.n3903 1118.26
R25953 vss.n3924 vss.n3908 1118.26
R25954 vss.n3920 vss.n3908 1118.26
R25955 vss.n3897 vss.n3893 1118.26
R25956 vss.n3929 vss.n3897 1118.26
R25957 vss.n3929 vss.n3898 1118.26
R25958 vss.n3909 vss.n3898 1118.26
R25959 vss.n3911 vss.n3909 1118.26
R25960 vss.n3912 vss.n3911 1118.26
R25961 vss.n5821 vss.n5820 1118.26
R25962 vss.n5822 vss.n5821 1118.26
R25963 vss.n5822 vss.n3547 1118.26
R25964 vss.n5836 vss.n3547 1118.26
R25965 vss.n5836 vss.n3548 1118.26
R25966 vss.n5828 vss.n3548 1118.26
R25967 vss.n5819 vss.n3554 1118.26
R25968 vss.n5823 vss.n3554 1118.26
R25969 vss.n5823 vss.n3556 1118.26
R25970 vss.n3556 vss.n3550 1118.26
R25971 vss.n5833 vss.n3550 1118.26
R25972 vss.n5833 vss.n5832 1118.26
R25973 vss.n3573 vss.n3563 1118.26
R25974 vss.n5808 vss.n3573 1118.26
R25975 vss.n5808 vss.n3574 1118.26
R25976 vss.n5804 vss.n3574 1118.26
R25977 vss.n5804 vss.n3581 1118.26
R25978 vss.n3613 vss.n3581 1118.26
R25979 vss.n3568 vss.n3564 1118.26
R25980 vss.n5809 vss.n3568 1118.26
R25981 vss.n5809 vss.n3569 1118.26
R25982 vss.n3582 vss.n3569 1118.26
R25983 vss.n3614 vss.n3582 1118.26
R25984 vss.n3615 vss.n3614 1118.26
R25985 vss.n5674 vss.n5673 1118.26
R25986 vss.n5673 vss.n5672 1118.26
R25987 vss.n5672 vss.n3593 1118.26
R25988 vss.n5794 vss.n3593 1118.26
R25989 vss.n5794 vss.n3595 1118.26
R25990 vss.n3595 vss.n3584 1118.26
R25991 vss.n5664 vss.n5660 1118.26
R25992 vss.n5671 vss.n5664 1118.26
R25993 vss.n5671 vss.n3589 1118.26
R25994 vss.n5795 vss.n3589 1118.26
R25995 vss.n5795 vss.n3590 1118.26
R25996 vss.n3590 vss.n3585 1118.26
R25997 vss.n5681 vss.n5680 1118.26
R25998 vss.n5682 vss.n5681 1118.26
R25999 vss.n5682 vss.n3606 1118.26
R26000 vss.n5736 vss.n3606 1118.26
R26001 vss.n5736 vss.n3607 1118.26
R26002 vss.n5691 vss.n3607 1118.26
R26003 vss.n5679 vss.n5650 1118.26
R26004 vss.n5683 vss.n5650 1118.26
R26005 vss.n5683 vss.n5652 1118.26
R26006 vss.n5652 vss.n3609 1118.26
R26007 vss.n5645 vss.n3609 1118.26
R26008 vss.n5646 vss.n5645 1118.26
R26009 vss.n5715 vss.n5707 1118.26
R26010 vss.n5721 vss.n5707 1118.26
R26011 vss.n5721 vss.n5701 1118.26
R26012 vss.n5726 vss.n5701 1118.26
R26013 vss.n5726 vss.n5703 1118.26
R26014 vss.n5703 vss.n5692 1118.26
R26015 vss.n5716 vss.n5709 1118.26
R26016 vss.n5720 vss.n5709 1118.26
R26017 vss.n5720 vss.n5697 1118.26
R26018 vss.n5727 vss.n5697 1118.26
R26019 vss.n5727 vss.n5698 1118.26
R26020 vss.n5698 vss.n5693 1118.26
R26021 vss.n9972 vss.n9971 1118.26
R26022 vss.n9973 vss.n9972 1118.26
R26023 vss.n9973 vss.n2634 1118.26
R26024 vss.n9987 vss.n2634 1118.26
R26025 vss.n9987 vss.n2635 1118.26
R26026 vss.n9979 vss.n2635 1118.26
R26027 vss.n9970 vss.n9958 1118.26
R26028 vss.n9974 vss.n9958 1118.26
R26029 vss.n9974 vss.n9960 1118.26
R26030 vss.n9960 vss.n2637 1118.26
R26031 vss.n9984 vss.n2637 1118.26
R26032 vss.n9984 vss.n9983 1118.26
R26033 vss.n2664 vss.n2655 1118.26
R26034 vss.n2670 vss.n2655 1118.26
R26035 vss.n2670 vss.n2649 1118.26
R26036 vss.n2677 vss.n2649 1118.26
R26037 vss.n2677 vss.n2651 1118.26
R26038 vss.n2651 vss.n2640 1118.26
R26039 vss.n2665 vss.n2657 1118.26
R26040 vss.n2669 vss.n2657 1118.26
R26041 vss.n2669 vss.n2645 1118.26
R26042 vss.n2678 vss.n2645 1118.26
R26043 vss.n2678 vss.n2646 1118.26
R26044 vss.n2646 vss.n2641 1118.26
R26045 vss.n3405 vss.n3404 1118.26
R26046 vss.n3406 vss.n3405 1118.26
R26047 vss.n3406 vss.n3384 1118.26
R26048 vss.n3420 vss.n3384 1118.26
R26049 vss.n3420 vss.n3385 1118.26
R26050 vss.n3412 vss.n3385 1118.26
R26051 vss.n3403 vss.n3391 1118.26
R26052 vss.n3407 vss.n3391 1118.26
R26053 vss.n3407 vss.n3393 1118.26
R26054 vss.n3393 vss.n3387 1118.26
R26055 vss.n3417 vss.n3387 1118.26
R26056 vss.n3417 vss.n3416 1118.26
R26057 vss.n4002 vss.n4001 1118.26
R26058 vss.n4003 vss.n4002 1118.26
R26059 vss.n4003 vss.n3981 1118.26
R26060 vss.n4017 vss.n3981 1118.26
R26061 vss.n4017 vss.n3982 1118.26
R26062 vss.n4009 vss.n3982 1118.26
R26063 vss.n4000 vss.n3988 1118.26
R26064 vss.n4004 vss.n3988 1118.26
R26065 vss.n4004 vss.n3990 1118.26
R26066 vss.n3990 vss.n3984 1118.26
R26067 vss.n4014 vss.n3984 1118.26
R26068 vss.n4014 vss.n4013 1118.26
R26069 vss.n4269 vss.n4268 1118.26
R26070 vss.n4270 vss.n4269 1118.26
R26071 vss.n4270 vss.n4248 1118.26
R26072 vss.n4284 vss.n4248 1118.26
R26073 vss.n4284 vss.n4249 1118.26
R26074 vss.n4276 vss.n4249 1118.26
R26075 vss.n4267 vss.n4255 1118.26
R26076 vss.n4271 vss.n4255 1118.26
R26077 vss.n4271 vss.n4257 1118.26
R26078 vss.n4257 vss.n4251 1118.26
R26079 vss.n4281 vss.n4251 1118.26
R26080 vss.n4281 vss.n4280 1118.26
R26081 vss.n14064 vss.n488 1118.26
R26082 vss.n14073 vss.n488 1118.26
R26083 vss.n14073 vss.n486 1118.26
R26084 vss.n14077 vss.n486 1118.26
R26085 vss.n14078 vss.n14077 1118.26
R26086 vss.n14079 vss.n14078 1118.26
R26087 vss.n14071 vss.n14070 1118.26
R26088 vss.n14072 vss.n14071 1118.26
R26089 vss.n14072 vss.n478 1118.26
R26090 vss.n14085 vss.n478 1118.26
R26091 vss.n14085 vss.n14084 1118.26
R26092 vss.n14084 vss.n14083 1118.26
R26093 vss.n10119 vss.n10113 1118.26
R26094 vss.n10128 vss.n10113 1118.26
R26095 vss.n10128 vss.n10111 1118.26
R26096 vss.n10132 vss.n10111 1118.26
R26097 vss.n10133 vss.n10132 1118.26
R26098 vss.n10134 vss.n10133 1118.26
R26099 vss.n10126 vss.n10125 1118.26
R26100 vss.n10127 vss.n10126 1118.26
R26101 vss.n10127 vss.n10105 1118.26
R26102 vss.n10140 vss.n10105 1118.26
R26103 vss.n10140 vss.n10139 1118.26
R26104 vss.n10139 vss.n10138 1118.26
R26105 vss.n12877 vss.n12871 1118.26
R26106 vss.n12886 vss.n12871 1118.26
R26107 vss.n12886 vss.n12869 1118.26
R26108 vss.n12890 vss.n12869 1118.26
R26109 vss.n12891 vss.n12890 1118.26
R26110 vss.n12892 vss.n12891 1118.26
R26111 vss.n12884 vss.n12883 1118.26
R26112 vss.n12885 vss.n12884 1118.26
R26113 vss.n12885 vss.n12863 1118.26
R26114 vss.n12898 vss.n12863 1118.26
R26115 vss.n12898 vss.n12897 1118.26
R26116 vss.n12897 vss.n12896 1118.26
R26117 vss.n10160 vss.n10154 1118.26
R26118 vss.n10169 vss.n10154 1118.26
R26119 vss.n10169 vss.n10152 1118.26
R26120 vss.n10173 vss.n10152 1118.26
R26121 vss.n10174 vss.n10173 1118.26
R26122 vss.n10175 vss.n10174 1118.26
R26123 vss.n10167 vss.n10166 1118.26
R26124 vss.n10168 vss.n10167 1118.26
R26125 vss.n10168 vss.n10146 1118.26
R26126 vss.n10181 vss.n10146 1118.26
R26127 vss.n10181 vss.n10180 1118.26
R26128 vss.n10180 vss.n10179 1118.26
R26129 vss.n12426 vss.n12420 1118.26
R26130 vss.n12435 vss.n12420 1118.26
R26131 vss.n12435 vss.n12418 1118.26
R26132 vss.n12439 vss.n12418 1118.26
R26133 vss.n12440 vss.n12439 1118.26
R26134 vss.n12441 vss.n12440 1118.26
R26135 vss.n12433 vss.n12432 1118.26
R26136 vss.n12434 vss.n12433 1118.26
R26137 vss.n12434 vss.n12412 1118.26
R26138 vss.n12447 vss.n12412 1118.26
R26139 vss.n12447 vss.n12446 1118.26
R26140 vss.n12446 vss.n12445 1118.26
R26141 vss.n11755 vss.n11749 1118.26
R26142 vss.n11764 vss.n11749 1118.26
R26143 vss.n11764 vss.n11747 1118.26
R26144 vss.n11768 vss.n11747 1118.26
R26145 vss.n11769 vss.n11768 1118.26
R26146 vss.n11770 vss.n11769 1118.26
R26147 vss.n11762 vss.n11761 1118.26
R26148 vss.n11763 vss.n11762 1118.26
R26149 vss.n11763 vss.n11741 1118.26
R26150 vss.n11776 vss.n11741 1118.26
R26151 vss.n11776 vss.n11775 1118.26
R26152 vss.n11775 vss.n11774 1118.26
R26153 vss.n12471 vss.n12465 1118.26
R26154 vss.n12480 vss.n12465 1118.26
R26155 vss.n12480 vss.n12463 1118.26
R26156 vss.n12484 vss.n12463 1118.26
R26157 vss.n12485 vss.n12484 1118.26
R26158 vss.n12486 vss.n12485 1118.26
R26159 vss.n12478 vss.n12477 1118.26
R26160 vss.n12479 vss.n12478 1118.26
R26161 vss.n12479 vss.n12457 1118.26
R26162 vss.n12492 vss.n12457 1118.26
R26163 vss.n12492 vss.n12491 1118.26
R26164 vss.n12491 vss.n12490 1118.26
R26165 vss.n2348 vss.n2309 1118.26
R26166 vss.n2344 vss.n2309 1118.26
R26167 vss.n2344 vss.n2313 1118.26
R26168 vss.n2329 vss.n2313 1118.26
R26169 vss.n2330 vss.n2329 1118.26
R26170 vss.n2331 vss.n2330 1118.26
R26171 vss.n2316 vss.n2308 1118.26
R26172 vss.n2343 vss.n2316 1118.26
R26173 vss.n2343 vss.n2317 1118.26
R26174 vss.n2337 vss.n2317 1118.26
R26175 vss.n2337 vss.n2336 1118.26
R26176 vss.n2336 vss.n2335 1118.26
R26177 vss.n12296 vss.n12290 1118.26
R26178 vss.n12305 vss.n12290 1118.26
R26179 vss.n12305 vss.n12288 1118.26
R26180 vss.n12309 vss.n12288 1118.26
R26181 vss.n12310 vss.n12309 1118.26
R26182 vss.n12311 vss.n12310 1118.26
R26183 vss.n12303 vss.n12302 1118.26
R26184 vss.n12304 vss.n12303 1118.26
R26185 vss.n12304 vss.n12282 1118.26
R26186 vss.n12317 vss.n12282 1118.26
R26187 vss.n12317 vss.n12316 1118.26
R26188 vss.n12316 vss.n12315 1118.26
R26189 vss.n12341 vss.n12335 1118.26
R26190 vss.n12350 vss.n12335 1118.26
R26191 vss.n12350 vss.n12333 1118.26
R26192 vss.n12354 vss.n12333 1118.26
R26193 vss.n12355 vss.n12354 1118.26
R26194 vss.n12356 vss.n12355 1118.26
R26195 vss.n12348 vss.n12347 1118.26
R26196 vss.n12349 vss.n12348 1118.26
R26197 vss.n12349 vss.n12327 1118.26
R26198 vss.n12362 vss.n12327 1118.26
R26199 vss.n12362 vss.n12361 1118.26
R26200 vss.n12361 vss.n12360 1118.26
R26201 vss.n10237 vss.n10231 1118.26
R26202 vss.n10246 vss.n10231 1118.26
R26203 vss.n10246 vss.n10229 1118.26
R26204 vss.n10250 vss.n10229 1118.26
R26205 vss.n10251 vss.n10250 1118.26
R26206 vss.n10252 vss.n10251 1118.26
R26207 vss.n10244 vss.n10243 1118.26
R26208 vss.n10245 vss.n10244 1118.26
R26209 vss.n10245 vss.n10223 1118.26
R26210 vss.n10258 vss.n10223 1118.26
R26211 vss.n10258 vss.n10257 1118.26
R26212 vss.n10257 vss.n10256 1118.26
R26213 vss.n2417 vss.n2411 1118.26
R26214 vss.n2426 vss.n2411 1118.26
R26215 vss.n2426 vss.n2409 1118.26
R26216 vss.n2430 vss.n2409 1118.26
R26217 vss.n2431 vss.n2430 1118.26
R26218 vss.n2432 vss.n2431 1118.26
R26219 vss.n2424 vss.n2423 1118.26
R26220 vss.n2425 vss.n2424 1118.26
R26221 vss.n2425 vss.n2403 1118.26
R26222 vss.n2438 vss.n2403 1118.26
R26223 vss.n2438 vss.n2437 1118.26
R26224 vss.n2437 vss.n2436 1118.26
R26225 vss.n12973 vss.n2369 1118.26
R26226 vss.n12969 vss.n2369 1118.26
R26227 vss.n12969 vss.n2373 1118.26
R26228 vss.n2389 vss.n2373 1118.26
R26229 vss.n2390 vss.n2389 1118.26
R26230 vss.n2391 vss.n2390 1118.26
R26231 vss.n2376 vss.n2368 1118.26
R26232 vss.n12968 vss.n2376 1118.26
R26233 vss.n12968 vss.n2377 1118.26
R26234 vss.n2397 vss.n2377 1118.26
R26235 vss.n2397 vss.n2396 1118.26
R26236 vss.n2396 vss.n2395 1118.26
R26237 vss.n10045 vss.n10028 1118.26
R26238 vss.n10049 vss.n10028 1118.26
R26239 vss.n10049 vss.n10025 1118.26
R26240 vss.n12948 vss.n10025 1118.26
R26241 vss.n12948 vss.n10026 1118.26
R26242 vss.n12944 vss.n10026 1118.26
R26243 vss.n10047 vss.n10046 1118.26
R26244 vss.n10048 vss.n10047 1118.26
R26245 vss.n10048 vss.n10020 1118.26
R26246 vss.n12949 vss.n10020 1118.26
R26247 vss.n12949 vss.n10021 1118.26
R26248 vss.n10057 vss.n10021 1118.26
R26249 vss.n10036 vss.n2096 1118.26
R26250 vss.n2109 vss.n2096 1118.26
R26251 vss.n2109 vss.n2106 1118.26
R26252 vss.n13083 vss.n2106 1118.26
R26253 vss.n13083 vss.n2107 1118.26
R26254 vss.n13079 vss.n2107 1118.26
R26255 vss.n10037 vss.n2097 1118.26
R26256 vss.n13086 vss.n2097 1118.26
R26257 vss.n13086 vss.n13085 1118.26
R26258 vss.n13085 vss.n13084 1118.26
R26259 vss.n13084 vss.n2102 1118.26
R26260 vss.n2118 vss.n2102 1118.26
R26261 vss.n2497 vss.n2490 1118.26
R26262 vss.n2506 vss.n2490 1118.26
R26263 vss.n2506 vss.n2488 1118.26
R26264 vss.n2510 vss.n2488 1118.26
R26265 vss.n2511 vss.n2510 1118.26
R26266 vss.n2512 vss.n2511 1118.26
R26267 vss.n2504 vss.n2503 1118.26
R26268 vss.n2505 vss.n2504 1118.26
R26269 vss.n2505 vss.n2482 1118.26
R26270 vss.n2518 vss.n2482 1118.26
R26271 vss.n2518 vss.n2517 1118.26
R26272 vss.n2517 vss.n2516 1118.26
R26273 vss.n12102 vss.n11843 1118.26
R26274 vss.n12108 vss.n11843 1118.26
R26275 vss.n12108 vss.n11839 1118.26
R26276 vss.n12112 vss.n11839 1118.26
R26277 vss.n12112 vss.n11829 1118.26
R26278 vss.n12121 vss.n11829 1118.26
R26279 vss.n12103 vss.n11845 1118.26
R26280 vss.n12107 vss.n11845 1118.26
R26281 vss.n12107 vss.n11837 1118.26
R26282 vss.n12115 vss.n11837 1118.26
R26283 vss.n12115 vss.n12114 1118.26
R26284 vss.n12114 vss.n11827 1118.26
R26285 vss.n12151 vss.n11810 1118.26
R26286 vss.n12147 vss.n11810 1118.26
R26287 vss.n12147 vss.n11814 1118.26
R26288 vss.n12128 vss.n11814 1118.26
R26289 vss.n12129 vss.n12128 1118.26
R26290 vss.n12130 vss.n12129 1118.26
R26291 vss.n11817 vss.n11808 1118.26
R26292 vss.n12146 vss.n11817 1118.26
R26293 vss.n12146 vss.n11818 1118.26
R26294 vss.n12136 vss.n11818 1118.26
R26295 vss.n12136 vss.n12135 1118.26
R26296 vss.n12135 vss.n12134 1118.26
R26297 vss.n12155 vss.n11799 1118.26
R26298 vss.n12161 vss.n11799 1118.26
R26299 vss.n12161 vss.n11795 1118.26
R26300 vss.n12165 vss.n11795 1118.26
R26301 vss.n12165 vss.n11788 1118.26
R26302 vss.n12174 vss.n11788 1118.26
R26303 vss.n12156 vss.n11801 1118.26
R26304 vss.n12160 vss.n11801 1118.26
R26305 vss.n12160 vss.n11793 1118.26
R26306 vss.n12168 vss.n11793 1118.26
R26307 vss.n12168 vss.n12167 1118.26
R26308 vss.n12167 vss.n11787 1118.26
R26309 vss.n12188 vss.n12182 1118.26
R26310 vss.n12261 vss.n12182 1118.26
R26311 vss.n12261 vss.n12180 1118.26
R26312 vss.n12265 vss.n12180 1118.26
R26313 vss.n12266 vss.n12265 1118.26
R26314 vss.n12267 vss.n12266 1118.26
R26315 vss.n12259 vss.n12186 1118.26
R26316 vss.n12260 vss.n12259 1118.26
R26317 vss.n12260 vss.n11783 1118.26
R26318 vss.n12273 vss.n11783 1118.26
R26319 vss.n12273 vss.n12272 1118.26
R26320 vss.n12272 vss.n12271 1118.26
R26321 vss.n12249 vss.n12192 1118.26
R26322 vss.n12245 vss.n12192 1118.26
R26323 vss.n12245 vss.n12196 1118.26
R26324 vss.n12230 vss.n12196 1118.26
R26325 vss.n12230 vss.n12228 1118.26
R26326 vss.n12235 vss.n12228 1118.26
R26327 vss.n12199 vss.n12191 1118.26
R26328 vss.n12244 vss.n12199 1118.26
R26329 vss.n12244 vss.n12200 1118.26
R26330 vss.n12238 vss.n12200 1118.26
R26331 vss.n12238 vss.n12237 1118.26
R26332 vss.n12237 vss.n12236 1118.26
R26333 vss.n12547 vss.n11722 1118.26
R26334 vss.n12543 vss.n11722 1118.26
R26335 vss.n12543 vss.n11726 1118.26
R26336 vss.n12218 vss.n11726 1118.26
R26337 vss.n12218 vss.n12214 1118.26
R26338 vss.n12214 vss.n12210 1118.26
R26339 vss.n11729 vss.n11720 1118.26
R26340 vss.n12542 vss.n11729 1118.26
R26341 vss.n12542 vss.n11730 1118.26
R26342 vss.n12216 vss.n11730 1118.26
R26343 vss.n12216 vss.n12215 1118.26
R26344 vss.n12215 vss.n12211 1118.26
R26345 vss.n12551 vss.n11712 1118.26
R26346 vss.n12557 vss.n11712 1118.26
R26347 vss.n12557 vss.n11708 1118.26
R26348 vss.n12561 vss.n11708 1118.26
R26349 vss.n12561 vss.n11701 1118.26
R26350 vss.n12570 vss.n11701 1118.26
R26351 vss.n12552 vss.n11714 1118.26
R26352 vss.n12556 vss.n11714 1118.26
R26353 vss.n12556 vss.n11706 1118.26
R26354 vss.n12564 vss.n11706 1118.26
R26355 vss.n12564 vss.n12563 1118.26
R26356 vss.n12563 vss.n11700 1118.26
R26357 vss.n11689 vss.n11624 1118.26
R26358 vss.n11692 vss.n11689 1118.26
R26359 vss.n11693 vss.n11692 1118.26
R26360 vss.n11694 vss.n11693 1118.26
R26361 vss.n11694 vss.n11637 1118.26
R26362 vss.n11698 vss.n11637 1118.26
R26363 vss.n11629 vss.n11625 1118.26
R26364 vss.n12580 vss.n11629 1118.26
R26365 vss.n12580 vss.n12579 1118.26
R26366 vss.n12579 vss.n12578 1118.26
R26367 vss.n12578 vss.n11632 1118.26
R26368 vss.n12574 vss.n11632 1118.26
R26369 vss.n11684 vss.n11643 1118.26
R26370 vss.n11680 vss.n11643 1118.26
R26371 vss.n11680 vss.n11647 1118.26
R26372 vss.n11665 vss.n11647 1118.26
R26373 vss.n11665 vss.n11663 1118.26
R26374 vss.n11670 vss.n11663 1118.26
R26375 vss.n11650 vss.n11642 1118.26
R26376 vss.n11679 vss.n11650 1118.26
R26377 vss.n11679 vss.n11651 1118.26
R26378 vss.n11673 vss.n11651 1118.26
R26379 vss.n11673 vss.n11672 1118.26
R26380 vss.n11672 vss.n11671 1118.26
R26381 vss.n10320 vss.n10314 1118.26
R26382 vss.n12841 vss.n10314 1118.26
R26383 vss.n12841 vss.n10312 1118.26
R26384 vss.n12845 vss.n10312 1118.26
R26385 vss.n12846 vss.n12845 1118.26
R26386 vss.n12847 vss.n12846 1118.26
R26387 vss.n12839 vss.n10318 1118.26
R26388 vss.n12840 vss.n12839 1118.26
R26389 vss.n12840 vss.n10306 1118.26
R26390 vss.n12853 vss.n10306 1118.26
R26391 vss.n12853 vss.n12852 1118.26
R26392 vss.n12852 vss.n12851 1118.26
R26393 vss.n12829 vss.n12774 1118.26
R26394 vss.n12825 vss.n12774 1118.26
R26395 vss.n12825 vss.n12778 1118.26
R26396 vss.n12812 vss.n12778 1118.26
R26397 vss.n12812 vss.n12810 1118.26
R26398 vss.n12817 vss.n12810 1118.26
R26399 vss.n12781 vss.n12773 1118.26
R26400 vss.n12824 vss.n12781 1118.26
R26401 vss.n12824 vss.n12782 1118.26
R26402 vss.n12820 vss.n12782 1118.26
R26403 vss.n12820 vss.n12819 1118.26
R26404 vss.n12819 vss.n12818 1118.26
R26405 vss.n12920 vss.n10087 1118.26
R26406 vss.n12916 vss.n10087 1118.26
R26407 vss.n12916 vss.n10091 1118.26
R26408 vss.n12800 vss.n10091 1118.26
R26409 vss.n12800 vss.n12796 1118.26
R26410 vss.n12796 vss.n12792 1118.26
R26411 vss.n10094 vss.n10085 1118.26
R26412 vss.n12915 vss.n10094 1118.26
R26413 vss.n12915 vss.n10095 1118.26
R26414 vss.n12798 vss.n10095 1118.26
R26415 vss.n12798 vss.n12797 1118.26
R26416 vss.n12797 vss.n12793 1118.26
R26417 vss.n11881 vss.n11873 1118.26
R26418 vss.n11887 vss.n11873 1118.26
R26419 vss.n11887 vss.n11867 1118.26
R26420 vss.n12079 vss.n11867 1118.26
R26421 vss.n12079 vss.n11869 1118.26
R26422 vss.n11869 vss.n11858 1118.26
R26423 vss.n11882 vss.n11875 1118.26
R26424 vss.n11886 vss.n11875 1118.26
R26425 vss.n11886 vss.n11863 1118.26
R26426 vss.n12080 vss.n11863 1118.26
R26427 vss.n12080 vss.n11864 1118.26
R26428 vss.n11864 vss.n11859 1118.26
R26429 vss.n10484 vss.n10483 1118.26
R26430 vss.n10485 vss.n10484 1118.26
R26431 vss.n10485 vss.n10464 1118.26
R26432 vss.n10499 vss.n10464 1118.26
R26433 vss.n10499 vss.n10465 1118.26
R26434 vss.n10491 vss.n10465 1118.26
R26435 vss.n10482 vss.n10471 1118.26
R26436 vss.n10486 vss.n10471 1118.26
R26437 vss.n10486 vss.n10473 1118.26
R26438 vss.n10473 vss.n10467 1118.26
R26439 vss.n10496 vss.n10467 1118.26
R26440 vss.n10496 vss.n10495 1118.26
R26441 vss.n10705 vss.n10704 1118.26
R26442 vss.n10706 vss.n10705 1118.26
R26443 vss.n10706 vss.n10685 1118.26
R26444 vss.n10720 vss.n10685 1118.26
R26445 vss.n10720 vss.n10686 1118.26
R26446 vss.n10712 vss.n10686 1118.26
R26447 vss.n10703 vss.n10692 1118.26
R26448 vss.n10707 vss.n10692 1118.26
R26449 vss.n10707 vss.n10694 1118.26
R26450 vss.n10694 vss.n10688 1118.26
R26451 vss.n10717 vss.n10688 1118.26
R26452 vss.n10717 vss.n10716 1118.26
R26453 vss.n11019 vss.n11018 1118.26
R26454 vss.n11020 vss.n11019 1118.26
R26455 vss.n11020 vss.n10999 1118.26
R26456 vss.n11034 vss.n10999 1118.26
R26457 vss.n11034 vss.n11000 1118.26
R26458 vss.n11026 vss.n11000 1118.26
R26459 vss.n11017 vss.n11006 1118.26
R26460 vss.n11021 vss.n11006 1118.26
R26461 vss.n11021 vss.n11008 1118.26
R26462 vss.n11008 vss.n11002 1118.26
R26463 vss.n11031 vss.n11002 1118.26
R26464 vss.n11031 vss.n11030 1118.26
R26465 vss.n10401 vss.n10400 1054.53
R26466 vss.n10400 vss.n10398 1054.53
R26467 vss.n2039 vss.n2035 1054.53
R26468 vss.n2040 vss.n2039 1054.53
R26469 vss.n2043 vss.n2036 1054.53
R26470 vss.n2043 vss.n2041 1054.53
R26471 vss.n12643 vss.n12634 1054.53
R26472 vss.n12634 vss.n12632 1054.53
R26473 vss.n12628 vss.n12624 1054.53
R26474 vss.n12629 vss.n12628 1054.53
R26475 vss.n12648 vss.n12625 1054.53
R26476 vss.n12648 vss.n12630 1054.53
R26477 vss.n11127 vss.n11118 1054.53
R26478 vss.n11118 vss.n11116 1054.53
R26479 vss.n11112 vss.n11108 1054.53
R26480 vss.n11113 vss.n11112 1054.53
R26481 vss.n11132 vss.n11109 1054.53
R26482 vss.n11132 vss.n11114 1054.53
R26483 vss.n10385 vss.n10377 1054.53
R26484 vss.n10386 vss.n10385 1054.53
R26485 vss.n12678 vss.n10388 1054.53
R26486 vss.n10388 vss.n10384 1054.53
R26487 vss.n12691 vss.n10378 1054.53
R26488 vss.n12691 vss.n12690 1054.53
R26489 vss.n11416 vss.n11408 1054.53
R26490 vss.n11417 vss.n11416 1054.53
R26491 vss.n11428 vss.n11419 1054.53
R26492 vss.n11419 vss.n11415 1054.53
R26493 vss.n11441 vss.n11409 1054.53
R26494 vss.n11441 vss.n11440 1054.53
R26495 vss.n11369 vss.n11361 1054.53
R26496 vss.n11370 vss.n11369 1054.53
R26497 vss.n11381 vss.n11372 1054.53
R26498 vss.n11372 vss.n11368 1054.53
R26499 vss.n11394 vss.n11362 1054.53
R26500 vss.n11394 vss.n11393 1054.53
R26501 vss.n10944 vss.n10936 1054.53
R26502 vss.n10945 vss.n10944 1054.53
R26503 vss.n10956 vss.n10947 1054.53
R26504 vss.n10947 vss.n10943 1054.53
R26505 vss.n10969 vss.n10937 1054.53
R26506 vss.n10969 vss.n10968 1054.53
R26507 vss.n10781 vss.n10773 1054.53
R26508 vss.n10782 vss.n10781 1054.53
R26509 vss.n10793 vss.n10784 1054.53
R26510 vss.n10784 vss.n10780 1054.53
R26511 vss.n10806 vss.n10774 1054.53
R26512 vss.n10806 vss.n10805 1054.53
R26513 vss.n10737 vss.n10729 1054.53
R26514 vss.n10738 vss.n10737 1054.53
R26515 vss.n10749 vss.n10740 1054.53
R26516 vss.n10740 vss.n10736 1054.53
R26517 vss.n10762 vss.n10730 1054.53
R26518 vss.n10762 vss.n10761 1054.53
R26519 vss.n11563 vss.n11555 1054.53
R26520 vss.n11564 vss.n11563 1054.53
R26521 vss.n11575 vss.n11566 1054.53
R26522 vss.n11566 vss.n11562 1054.53
R26523 vss.n11588 vss.n11556 1054.53
R26524 vss.n11588 vss.n11587 1054.53
R26525 vss.n10560 vss.n10552 1054.53
R26526 vss.n10561 vss.n10560 1054.53
R26527 vss.n10572 vss.n10563 1054.53
R26528 vss.n10563 vss.n10559 1054.53
R26529 vss.n10585 vss.n10553 1054.53
R26530 vss.n10585 vss.n10584 1054.53
R26531 vss.n10516 vss.n10508 1054.53
R26532 vss.n10517 vss.n10516 1054.53
R26533 vss.n10528 vss.n10519 1054.53
R26534 vss.n10519 vss.n10515 1054.53
R26535 vss.n10541 vss.n10509 1054.53
R26536 vss.n10541 vss.n10540 1054.53
R26537 vss.n11937 vss.n11929 1054.53
R26538 vss.n11938 vss.n11937 1054.53
R26539 vss.n11949 vss.n11940 1054.53
R26540 vss.n11940 vss.n11936 1054.53
R26541 vss.n11962 vss.n11930 1054.53
R26542 vss.n11962 vss.n11961 1054.53
R26543 vss.n11870 vss.n11867 1054.53
R26544 vss.n11870 vss.n11863 1054.53
R26545 vss.n11900 vss.n11896 1054.53
R26546 vss.n11900 vss.n11899 1054.53
R26547 vss.n12070 vss.n11895 1054.53
R26548 vss.n11895 vss.n11856 1054.53
R26549 vss.n12089 vss.n11857 1054.53
R26550 vss.n12090 vss.n12089 1054.53
R26551 vss.n12057 vss.n11904 1054.53
R26552 vss.n12057 vss.n11905 1054.53
R26553 vss.n11975 vss.n11914 1054.53
R26554 vss.n12052 vss.n11914 1054.53
R26555 vss.n11921 vss.n11920 1054.53
R26556 vss.n11920 vss.n11916 1054.53
R26557 vss.n12011 vss.n12010 1054.53
R26558 vss.n12010 vss.n11986 1054.53
R26559 vss.n12018 vss.n11985 1054.53
R26560 vss.n12029 vss.n11985 1054.53
R26561 vss.n12042 vss.n11981 1054.53
R26562 vss.n12042 vss.n11982 1054.53
R26563 vss.n12005 vss.n11992 1054.53
R26564 vss.n12005 vss.n11993 1054.53
R26565 vss.n10598 vss.n10594 1054.53
R26566 vss.n10599 vss.n10598 1054.53
R26567 vss.n10602 vss.n10595 1054.53
R26568 vss.n10602 vss.n10600 1054.53
R26569 vss.n10653 vss.n10652 1054.53
R26570 vss.n10652 vss.n10648 1054.53
R26571 vss.n10661 vss.n10649 1054.53
R26572 vss.n10663 vss.n10661 1054.53
R26573 vss.n12597 vss.n10607 1054.53
R26574 vss.n12597 vss.n10608 1054.53
R26575 vss.n10637 vss.n10632 1054.53
R26576 vss.n10637 vss.n10636 1054.53
R26577 vss.n10634 vss.n10629 1054.53
R26578 vss.n10634 vss.n10628 1054.53
R26579 vss.n11604 vss.n11602 1054.53
R26580 vss.n11605 vss.n11604 1054.53
R26581 vss.n10838 vss.n10837 1054.53
R26582 vss.n10837 vss.n10834 1054.53
R26583 vss.n10841 vss.n10839 1054.53
R26584 vss.n10841 vss.n10621 1054.53
R26585 vss.n11615 vss.n10622 1054.53
R26586 vss.n11616 vss.n11615 1054.53
R26587 vss.n10863 vss.n10825 1054.53
R26588 vss.n10825 vss.n10823 1054.53
R26589 vss.n10819 vss.n10815 1054.53
R26590 vss.n10820 vss.n10819 1054.53
R26591 vss.n10868 vss.n10816 1054.53
R26592 vss.n10868 vss.n10821 1054.53
R26593 vss.n11498 vss.n11497 1054.53
R26594 vss.n11497 vss.n10878 1054.53
R26595 vss.n11503 vss.n10877 1054.53
R26596 vss.n11514 vss.n10877 1054.53
R26597 vss.n11526 vss.n10873 1054.53
R26598 vss.n11526 vss.n10874 1054.53
R26599 vss.n11492 vss.n10883 1054.53
R26600 vss.n11492 vss.n10884 1054.53
R26601 vss.n10981 vss.n10893 1054.53
R26602 vss.n11487 vss.n10893 1054.53
R26603 vss.n10984 vss.n10983 1054.53
R26604 vss.n10983 vss.n10895 1054.53
R26605 vss.n10931 vss.n10930 1054.53
R26606 vss.n10930 vss.n10904 1054.53
R26607 vss.n11455 vss.n10903 1054.53
R26608 vss.n11466 vss.n10903 1054.53
R26609 vss.n11477 vss.n10899 1054.53
R26610 vss.n11477 vss.n10900 1054.53
R26611 vss.n10925 vss.n10912 1054.53
R26612 vss.n10925 vss.n10913 1054.53
R26613 vss.n10909 vss.n10336 1054.53
R26614 vss.n10909 vss.n10335 1054.53
R26615 vss.n12747 vss.n12745 1054.53
R26616 vss.n12748 vss.n12747 1054.53
R26617 vss.n10349 vss.n10345 1054.53
R26618 vss.n10349 vss.n10348 1054.53
R26619 vss.n12735 vss.n10344 1054.53
R26620 vss.n10344 vss.n10328 1054.53
R26621 vss.n12758 vss.n10329 1054.53
R26622 vss.n12759 vss.n12758 1054.53
R26623 vss.n12722 vss.n10353 1054.53
R26624 vss.n12722 vss.n10354 1054.53
R26625 vss.n12704 vss.n10363 1054.53
R26626 vss.n12717 vss.n10363 1054.53
R26627 vss.n10370 vss.n10369 1054.53
R26628 vss.n10369 vss.n10365 1054.53
R26629 vss.n13099 vss.n2089 1054.53
R26630 vss.n13099 vss.n2091 1054.53
R26631 vss.n2086 vss.n2084 1054.53
R26632 vss.n2086 vss.n2079 1054.53
R26633 vss.n2083 vss.n2082 1054.53
R26634 vss.n2082 vss.n2078 1054.53
R26635 vss.n10069 vss.n10060 1054.53
R26636 vss.n10070 vss.n10069 1054.53
R26637 vss.n10073 vss.n10072 1054.53
R26638 vss.n10073 vss.n10068 1054.53
R26639 vss.n10079 vss.n10076 1054.53
R26640 vss.n10079 vss.n10078 1054.53
R26641 vss.n12802 vss.n12796 1054.53
R26642 vss.n12802 vss.n12797 1054.53
R26643 vss.n12810 vss.n12788 1054.53
R26644 vss.n12819 vss.n12788 1054.53
R26645 vss.n12785 vss.n12778 1054.53
R26646 vss.n12785 vss.n12782 1054.53
R26647 vss.n12846 vss.n10307 1054.53
R26648 vss.n12852 vss.n10307 1054.53
R26649 vss.n11663 vss.n11657 1054.53
R26650 vss.n11672 vss.n11657 1054.53
R26651 vss.n11654 vss.n11647 1054.53
R26652 vss.n11654 vss.n11651 1054.53
R26653 vss.n11637 vss.n11636 1054.53
R26654 vss.n11636 vss.n11632 1054.53
R26655 vss.n12562 vss.n11701 1054.53
R26656 vss.n12563 vss.n12562 1054.53
R26657 vss.n11709 vss.n11708 1054.53
R26658 vss.n11709 vss.n11706 1054.53
R26659 vss.n12220 vss.n12214 1054.53
R26660 vss.n12220 vss.n12215 1054.53
R26661 vss.n12228 vss.n12206 1054.53
R26662 vss.n12237 vss.n12206 1054.53
R26663 vss.n12203 vss.n12196 1054.53
R26664 vss.n12203 vss.n12200 1054.53
R26665 vss.n12266 vss.n11784 1054.53
R26666 vss.n12272 vss.n11784 1054.53
R26667 vss.n12166 vss.n11788 1054.53
R26668 vss.n12167 vss.n12166 1054.53
R26669 vss.n11796 vss.n11795 1054.53
R26670 vss.n11796 vss.n11793 1054.53
R26671 vss.n12129 vss.n11824 1054.53
R26672 vss.n12135 vss.n11824 1054.53
R26673 vss.n13004 vss.n2250 1054.53
R26674 vss.n13004 vss.n2245 1054.53
R26675 vss.n2249 vss.n2248 1054.53
R26676 vss.n2248 vss.n2244 1054.53
R26677 vss.n2254 vss.n2252 1054.53
R26678 vss.n12999 vss.n2254 1054.53
R26679 vss.n2290 vss.n2278 1054.53
R26680 vss.n2290 vss.n2280 1054.53
R26681 vss.n2275 vss.n2273 1054.53
R26682 vss.n2275 vss.n2268 1054.53
R26683 vss.n2272 vss.n2271 1054.53
R26684 vss.n2271 vss.n2267 1054.53
R26685 vss.n13063 vss.n2136 1054.53
R26686 vss.n13063 vss.n2138 1054.53
R26687 vss.n2133 vss.n2131 1054.53
R26688 vss.n2133 vss.n2126 1054.53
R26689 vss.n2130 vss.n2129 1054.53
R26690 vss.n2129 vss.n2125 1054.53
R26691 vss.n14078 vss.n479 1054.53
R26692 vss.n14084 vss.n479 1054.53
R26693 vss.n490 vss.n486 1054.53
R26694 vss.n490 vss.n478 1054.53
R26695 vss.n446 vss.n445 1054.53
R26696 vss.n445 vss.n440 1054.53
R26697 vss.n447 vss.n443 1054.53
R26698 vss.n447 vss.n439 1054.53
R26699 vss.n453 vss.n450 1054.53
R26700 vss.n453 vss.n452 1054.53
R26701 vss.n628 vss.n623 1054.53
R26702 vss.n628 vss.n627 1054.53
R26703 vss.n625 vss.n620 1054.53
R26704 vss.n625 vss.n619 1054.53
R26705 vss.n650 vss.n648 1054.53
R26706 vss.n651 vss.n650 1054.53
R26707 vss.n2007 vss.n1998 1054.53
R26708 vss.n1998 vss.n1996 1054.53
R26709 vss.n1992 vss.n1988 1054.53
R26710 vss.n1993 vss.n1992 1054.53
R26711 vss.n2012 vss.n1989 1054.53
R26712 vss.n2012 vss.n1994 1054.53
R26713 vss.n1072 vss.n1063 1054.53
R26714 vss.n1063 vss.n1061 1054.53
R26715 vss.n1057 vss.n1053 1054.53
R26716 vss.n1058 vss.n1057 1054.53
R26717 vss.n1077 vss.n1054 1054.53
R26718 vss.n1077 vss.n1059 1054.53
R26719 vss.n1333 vss.n1324 1054.53
R26720 vss.n1324 vss.n1322 1054.53
R26721 vss.n1318 vss.n1314 1054.53
R26722 vss.n1319 vss.n1318 1054.53
R26723 vss.n1338 vss.n1315 1054.53
R26724 vss.n1338 vss.n1320 1054.53
R26725 vss.n1465 vss.n1456 1054.53
R26726 vss.n1456 vss.n1454 1054.53
R26727 vss.n1450 vss.n1446 1054.53
R26728 vss.n1451 vss.n1450 1054.53
R26729 vss.n1470 vss.n1447 1054.53
R26730 vss.n1470 vss.n1452 1054.53
R26731 vss.n1628 vss.n1619 1054.53
R26732 vss.n1619 vss.n1617 1054.53
R26733 vss.n1613 vss.n1609 1054.53
R26734 vss.n1614 vss.n1613 1054.53
R26735 vss.n1633 vss.n1610 1054.53
R26736 vss.n1633 vss.n1615 1054.53
R26737 vss.n1545 vss.n1536 1054.53
R26738 vss.n1536 vss.n1534 1054.53
R26739 vss.n1530 vss.n1526 1054.53
R26740 vss.n1531 vss.n1530 1054.53
R26741 vss.n1550 vss.n1527 1054.53
R26742 vss.n1550 vss.n1532 1054.53
R26743 vss.n895 vss.n894 1054.53
R26744 vss.n894 vss.n880 1054.53
R26745 vss.n899 vss.n881 1054.53
R26746 vss.n911 vss.n881 1054.53
R26747 vss.n888 vss.n887 1054.53
R26748 vss.n887 vss.n883 1054.53
R26749 vss.n851 vss.n850 1054.53
R26750 vss.n850 vss.n839 1054.53
R26751 vss.n855 vss.n841 1054.53
R26752 vss.n867 vss.n841 1054.53
R26753 vss.n848 vss.n847 1054.53
R26754 vss.n847 vss.n843 1054.53
R26755 vss.n825 vss.n824 1054.53
R26756 vss.n824 vss.n822 1054.53
R26757 vss.n602 vss.n598 1054.53
R26758 vss.n603 vss.n602 1054.53
R26759 vss.n606 vss.n599 1054.53
R26760 vss.n606 vss.n604 1054.53
R26761 vss.n13216 vss.n807 1054.53
R26762 vss.n807 vss.n805 1054.53
R26763 vss.n801 vss.n797 1054.53
R26764 vss.n802 vss.n801 1054.53
R26765 vss.n13221 vss.n798 1054.53
R26766 vss.n13221 vss.n803 1054.53
R26767 vss.n1675 vss.n1666 1054.53
R26768 vss.n1666 vss.n1664 1054.53
R26769 vss.n1660 vss.n1656 1054.53
R26770 vss.n1661 vss.n1660 1054.53
R26771 vss.n1680 vss.n1657 1054.53
R26772 vss.n1680 vss.n1662 1054.53
R26773 vss.n1380 vss.n1371 1054.53
R26774 vss.n1371 vss.n1369 1054.53
R26775 vss.n1365 vss.n1361 1054.53
R26776 vss.n1366 vss.n1365 1054.53
R26777 vss.n1385 vss.n1362 1054.53
R26778 vss.n1385 vss.n1367 1054.53
R26779 vss.n1181 vss.n1172 1054.53
R26780 vss.n1172 vss.n1170 1054.53
R26781 vss.n1166 vss.n1162 1054.53
R26782 vss.n1167 vss.n1166 1054.53
R26783 vss.n1186 vss.n1163 1054.53
R26784 vss.n1186 vss.n1168 1054.53
R26785 vss.n1117 vss.n1108 1054.53
R26786 vss.n1108 vss.n1106 1054.53
R26787 vss.n1102 vss.n1098 1054.53
R26788 vss.n1103 vss.n1102 1054.53
R26789 vss.n1122 vss.n1099 1054.53
R26790 vss.n1122 vss.n1104 1054.53
R26791 vss.n13195 vss.n13163 1054.53
R26792 vss.n13195 vss.n13166 1054.53
R26793 vss.n13169 vss.n13162 1054.53
R26794 vss.n13170 vss.n13169 1054.53
R26795 vss.n13181 vss.n13172 1054.53
R26796 vss.n13172 vss.n13168 1054.53
R26797 vss.n720 vss.n710 1054.53
R26798 vss.n721 vss.n720 1054.53
R26799 vss.n702 vss.n699 1054.53
R26800 vss.n702 vss.n695 1054.53
R26801 vss.n1929 vss.n1140 1054.53
R26802 vss.n1930 vss.n1929 1054.53
R26803 vss.n1156 vss.n1155 1054.53
R26804 vss.n1156 vss.n1151 1054.53
R26805 vss.n1858 vss.n1205 1054.53
R26806 vss.n1859 vss.n1858 1054.53
R26807 vss.n1221 vss.n1220 1054.53
R26808 vss.n1221 vss.n1216 1054.53
R26809 vss.n1240 vss.n1236 1054.53
R26810 vss.n1241 vss.n1240 1054.53
R26811 vss.n1274 vss.n1273 1054.53
R26812 vss.n1274 vss.n1269 1054.53
R26813 vss.n1754 vss.n1701 1054.53
R26814 vss.n1755 vss.n1754 1054.53
R26815 vss.n1717 vss.n1716 1054.53
R26816 vss.n1717 vss.n1712 1054.53
R26817 vss.n756 vss.n754 1054.53
R26818 vss.n756 vss.n749 1054.53
R26819 vss.n589 vss.n587 1054.53
R26820 vss.n589 vss.n582 1054.53
R26821 vss.n567 vss.n559 1054.53
R26822 vss.n568 vss.n567 1054.53
R26823 vss.n550 vss.n548 1054.53
R26824 vss.n550 vss.n543 1054.53
R26825 vss.n12 vss.n10 1054.53
R26826 vss.n12 vss.n5 1054.53
R26827 vss.n9 vss.n8 1054.53
R26828 vss.n8 vss.n4 1054.53
R26829 vss.n183 vss.n177 1054.53
R26830 vss.n183 vss.n178 1054.53
R26831 vss.n14716 vss.n14704 1054.53
R26832 vss.n14716 vss.n14706 1054.53
R26833 vss.n14701 vss.n14699 1054.53
R26834 vss.n14701 vss.n14694 1054.53
R26835 vss.n14698 vss.n14697 1054.53
R26836 vss.n14697 vss.n14693 1054.53
R26837 vss.n14593 vss.n14574 1054.53
R26838 vss.n14593 vss.n14569 1054.53
R26839 vss.n14573 vss.n14572 1054.53
R26840 vss.n14572 vss.n14568 1054.53
R26841 vss.n14578 vss.n14576 1054.53
R26842 vss.n14588 vss.n14578 1054.53
R26843 vss.n14521 vss.n14509 1054.53
R26844 vss.n14521 vss.n14511 1054.53
R26845 vss.n14506 vss.n14504 1054.53
R26846 vss.n14506 vss.n14499 1054.53
R26847 vss.n14503 vss.n14502 1054.53
R26848 vss.n14502 vss.n14498 1054.53
R26849 vss.n14398 vss.n14379 1054.53
R26850 vss.n14398 vss.n14374 1054.53
R26851 vss.n14378 vss.n14377 1054.53
R26852 vss.n14377 vss.n14373 1054.53
R26853 vss.n14383 vss.n14381 1054.53
R26854 vss.n14393 vss.n14383 1054.53
R26855 vss.n14326 vss.n14314 1054.53
R26856 vss.n14326 vss.n14316 1054.53
R26857 vss.n14311 vss.n14309 1054.53
R26858 vss.n14311 vss.n14304 1054.53
R26859 vss.n14308 vss.n14307 1054.53
R26860 vss.n14307 vss.n14303 1054.53
R26861 vss.n345 vss.n326 1054.53
R26862 vss.n345 vss.n321 1054.53
R26863 vss.n325 vss.n324 1054.53
R26864 vss.n324 vss.n320 1054.53
R26865 vss.n330 vss.n328 1054.53
R26866 vss.n340 vss.n330 1054.53
R26867 vss.n14207 vss.n14195 1054.53
R26868 vss.n14207 vss.n14197 1054.53
R26869 vss.n14192 vss.n14190 1054.53
R26870 vss.n14192 vss.n14185 1054.53
R26871 vss.n14189 vss.n14188 1054.53
R26872 vss.n14188 vss.n14184 1054.53
R26873 vss.n14124 vss.n14105 1054.53
R26874 vss.n14124 vss.n14100 1054.53
R26875 vss.n14104 vss.n14103 1054.53
R26876 vss.n14103 vss.n14099 1054.53
R26877 vss.n14109 vss.n14107 1054.53
R26878 vss.n14119 vss.n14109 1054.53
R26879 vss.n14233 vss.n423 1054.53
R26880 vss.n14233 vss.n418 1054.53
R26881 vss.n422 vss.n421 1054.53
R26882 vss.n421 vss.n417 1054.53
R26883 vss.n427 vss.n425 1054.53
R26884 vss.n14228 vss.n427 1054.53
R26885 vss.n14280 vss.n14268 1054.53
R26886 vss.n14280 vss.n14270 1054.53
R26887 vss.n14265 vss.n14263 1054.53
R26888 vss.n14265 vss.n14258 1054.53
R26889 vss.n14262 vss.n14261 1054.53
R26890 vss.n14261 vss.n14257 1054.53
R26891 vss.n14352 vss.n300 1054.53
R26892 vss.n14352 vss.n295 1054.53
R26893 vss.n299 vss.n298 1054.53
R26894 vss.n298 vss.n294 1054.53
R26895 vss.n304 vss.n302 1054.53
R26896 vss.n14347 vss.n304 1054.53
R26897 vss.n14475 vss.n14463 1054.53
R26898 vss.n14475 vss.n14465 1054.53
R26899 vss.n14460 vss.n14458 1054.53
R26900 vss.n14460 vss.n14453 1054.53
R26901 vss.n14457 vss.n14456 1054.53
R26902 vss.n14456 vss.n14452 1054.53
R26903 vss.n14547 vss.n241 1054.53
R26904 vss.n14547 vss.n236 1054.53
R26905 vss.n240 vss.n239 1054.53
R26906 vss.n239 vss.n235 1054.53
R26907 vss.n245 vss.n243 1054.53
R26908 vss.n14542 vss.n245 1054.53
R26909 vss.n14670 vss.n14658 1054.53
R26910 vss.n14670 vss.n14660 1054.53
R26911 vss.n14655 vss.n14653 1054.53
R26912 vss.n14655 vss.n14648 1054.53
R26913 vss.n14652 vss.n14651 1054.53
R26914 vss.n14651 vss.n14647 1054.53
R26915 vss.n14742 vss.n164 1054.53
R26916 vss.n14742 vss.n159 1054.53
R26917 vss.n163 vss.n162 1054.53
R26918 vss.n162 vss.n158 1054.53
R26919 vss.n168 vss.n166 1054.53
R26920 vss.n14737 vss.n168 1054.53
R26921 vss.n13576 vss.n13570 1054.53
R26922 vss.n13576 vss.n13571 1054.53
R26923 vss.n472 vss.n465 1054.53
R26924 vss.n472 vss.n469 1054.53
R26925 vss.n467 vss.n461 1054.53
R26926 vss.n468 vss.n467 1054.53
R26927 vss.n13595 vss.n13564 1054.53
R26928 vss.n13595 vss.n13584 1054.53
R26929 vss.n13561 vss.n13559 1054.53
R26930 vss.n13561 vss.n13554 1054.53
R26931 vss.n13558 vss.n13557 1054.53
R26932 vss.n13557 vss.n13553 1054.53
R26933 vss.n13625 vss.n13623 1054.53
R26934 vss.n13626 vss.n13625 1054.53
R26935 vss.n13635 vss.n13521 1054.53
R26936 vss.n13644 vss.n13521 1054.53
R26937 vss.n13518 vss.n13511 1054.53
R26938 vss.n13518 vss.n13515 1054.53
R26939 vss.n13679 vss.n13677 1054.53
R26940 vss.n13680 vss.n13679 1054.53
R26941 vss.n13690 vss.n13482 1054.53
R26942 vss.n13699 vss.n13482 1054.53
R26943 vss.n13479 vss.n13472 1054.53
R26944 vss.n13479 vss.n13476 1054.53
R26945 vss.n13730 vss.n13728 1054.53
R26946 vss.n13731 vss.n13730 1054.53
R26947 vss.n13740 vss.n13441 1054.53
R26948 vss.n13749 vss.n13441 1054.53
R26949 vss.n13438 vss.n13431 1054.53
R26950 vss.n13438 vss.n13435 1054.53
R26951 vss.n13784 vss.n13782 1054.53
R26952 vss.n13785 vss.n13784 1054.53
R26953 vss.n13795 vss.n13402 1054.53
R26954 vss.n13804 vss.n13402 1054.53
R26955 vss.n13399 vss.n13392 1054.53
R26956 vss.n13399 vss.n13396 1054.53
R26957 vss.n13835 vss.n13833 1054.53
R26958 vss.n13836 vss.n13835 1054.53
R26959 vss.n13845 vss.n13361 1054.53
R26960 vss.n13854 vss.n13361 1054.53
R26961 vss.n13358 vss.n13351 1054.53
R26962 vss.n13358 vss.n13355 1054.53
R26963 vss.n13889 vss.n13887 1054.53
R26964 vss.n13890 vss.n13889 1054.53
R26965 vss.n13900 vss.n13322 1054.53
R26966 vss.n13909 vss.n13322 1054.53
R26967 vss.n13316 vss.n13309 1054.53
R26968 vss.n13316 vss.n13313 1054.53
R26969 vss.n13311 vss.n13305 1054.53
R26970 vss.n13312 vss.n13311 1054.53
R26971 vss.n13337 vss.n13332 1054.53
R26972 vss.n13337 vss.n13331 1054.53
R26973 vss.n13340 vss.n13335 1054.53
R26974 vss.n13340 vss.n13339 1054.53
R26975 vss.n13353 vss.n13347 1054.53
R26976 vss.n13354 vss.n13353 1054.53
R26977 vss.n13378 vss.n13373 1054.53
R26978 vss.n13378 vss.n13372 1054.53
R26979 vss.n13381 vss.n13376 1054.53
R26980 vss.n13381 vss.n13380 1054.53
R26981 vss.n13394 vss.n13388 1054.53
R26982 vss.n13395 vss.n13394 1054.53
R26983 vss.n13417 vss.n13412 1054.53
R26984 vss.n13417 vss.n13411 1054.53
R26985 vss.n13420 vss.n13415 1054.53
R26986 vss.n13420 vss.n13419 1054.53
R26987 vss.n13433 vss.n13427 1054.53
R26988 vss.n13434 vss.n13433 1054.53
R26989 vss.n13458 vss.n13453 1054.53
R26990 vss.n13458 vss.n13452 1054.53
R26991 vss.n13461 vss.n13456 1054.53
R26992 vss.n13461 vss.n13460 1054.53
R26993 vss.n13474 vss.n13468 1054.53
R26994 vss.n13475 vss.n13474 1054.53
R26995 vss.n13497 vss.n13492 1054.53
R26996 vss.n13497 vss.n13491 1054.53
R26997 vss.n13500 vss.n13495 1054.53
R26998 vss.n13500 vss.n13499 1054.53
R26999 vss.n13513 vss.n13507 1054.53
R27000 vss.n13514 vss.n13513 1054.53
R27001 vss.n13538 vss.n13533 1054.53
R27002 vss.n13538 vss.n13532 1054.53
R27003 vss.n13541 vss.n13536 1054.53
R27004 vss.n13541 vss.n13540 1054.53
R27005 vss.n528 vss.n520 1054.53
R27006 vss.n529 vss.n528 1054.53
R27007 vss.n14007 vss.n531 1054.53
R27008 vss.n531 vss.n527 1054.53
R27009 vss.n14020 vss.n521 1054.53
R27010 vss.n14020 vss.n14019 1054.53
R27011 vss.n547 vss.n546 1054.53
R27012 vss.n546 vss.n542 1054.53
R27013 vss.n670 vss.n669 1054.53
R27014 vss.n669 vss.n665 1054.53
R27015 vss.n13972 vss.n570 1054.53
R27016 vss.n570 vss.n566 1054.53
R27017 vss.n13985 vss.n560 1054.53
R27018 vss.n13985 vss.n13984 1054.53
R27019 vss.n586 vss.n585 1054.53
R27020 vss.n585 vss.n581 1054.53
R27021 vss.n768 vss.n764 1054.53
R27022 vss.n769 vss.n768 1054.53
R27023 vss.n753 vss.n752 1054.53
R27024 vss.n752 vss.n748 1054.53
R27025 vss.n789 vss.n759 1054.53
R27026 vss.n789 vss.n788 1054.53
R27027 vss.n1723 vss.n1720 1054.53
R27028 vss.n1723 vss.n1722 1054.53
R27029 vss.n1713 vss.n1708 1054.53
R27030 vss.n1714 vss.n1713 1054.53
R27031 vss.n1784 vss.n1757 1054.53
R27032 vss.n1757 vss.n1753 1054.53
R27033 vss.n1797 vss.n1702 1054.53
R27034 vss.n1797 vss.n1796 1054.53
R27035 vss.n1770 vss.n1769 1054.53
R27036 vss.n1769 vss.n1767 1054.53
R27037 vss.n1270 vss.n1265 1054.53
R27038 vss.n1271 vss.n1270 1054.53
R27039 vss.n1829 vss.n1235 1054.53
R27040 vss.n1238 vss.n1235 1054.53
R27041 vss.n1249 vss.n1244 1054.53
R27042 vss.n1250 vss.n1249 1054.53
R27043 vss.n1227 vss.n1224 1054.53
R27044 vss.n1227 vss.n1226 1054.53
R27045 vss.n1217 vss.n1212 1054.53
R27046 vss.n1218 vss.n1217 1054.53
R27047 vss.n1888 vss.n1861 1054.53
R27048 vss.n1861 vss.n1857 1054.53
R27049 vss.n1901 vss.n1206 1054.53
R27050 vss.n1901 vss.n1900 1054.53
R27051 vss.n1874 vss.n1873 1054.53
R27052 vss.n1873 vss.n1871 1054.53
R27053 vss.n1152 vss.n1147 1054.53
R27054 vss.n1153 vss.n1152 1054.53
R27055 vss.n1959 vss.n1932 1054.53
R27056 vss.n1932 vss.n1928 1054.53
R27057 vss.n1972 vss.n1141 1054.53
R27058 vss.n1972 vss.n1971 1054.53
R27059 vss.n1945 vss.n1944 1054.53
R27060 vss.n1944 vss.n1942 1054.53
R27061 vss.n701 vss.n700 1054.53
R27062 vss.n700 vss.n696 1054.53
R27063 vss.n13271 vss.n723 1054.53
R27064 vss.n723 vss.n719 1054.53
R27065 vss.n13284 vss.n711 1054.53
R27066 vss.n13284 vss.n13283 1054.53
R27067 vss.n9614 vss.n9595 1054.53
R27068 vss.n9614 vss.n9590 1054.53
R27069 vss.n9594 vss.n9593 1054.53
R27070 vss.n9593 vss.n9589 1054.53
R27071 vss.n9599 vss.n9597 1054.53
R27072 vss.n9609 vss.n9599 1054.53
R27073 vss.n7522 vss.n7510 1054.53
R27074 vss.n7522 vss.n7512 1054.53
R27075 vss.n7507 vss.n7505 1054.53
R27076 vss.n7507 vss.n7500 1054.53
R27077 vss.n7504 vss.n7503 1054.53
R27078 vss.n7503 vss.n7499 1054.53
R27079 vss.n8934 vss.n8922 1054.53
R27080 vss.n8934 vss.n8924 1054.53
R27081 vss.n8919 vss.n8917 1054.53
R27082 vss.n8919 vss.n8912 1054.53
R27083 vss.n8916 vss.n8915 1054.53
R27084 vss.n8915 vss.n8911 1054.53
R27085 vss.n7573 vss.n7554 1054.53
R27086 vss.n7573 vss.n7549 1054.53
R27087 vss.n7553 vss.n7552 1054.53
R27088 vss.n7552 vss.n7548 1054.53
R27089 vss.n7558 vss.n7556 1054.53
R27090 vss.n7568 vss.n7558 1054.53
R27091 vss.n8815 vss.n8803 1054.53
R27092 vss.n8815 vss.n8805 1054.53
R27093 vss.n8800 vss.n8798 1054.53
R27094 vss.n8800 vss.n8793 1054.53
R27095 vss.n8797 vss.n8796 1054.53
R27096 vss.n8796 vss.n8792 1054.53
R27097 vss.n7716 vss.n7697 1054.53
R27098 vss.n7716 vss.n7692 1054.53
R27099 vss.n7696 vss.n7695 1054.53
R27100 vss.n7695 vss.n7691 1054.53
R27101 vss.n7701 vss.n7699 1054.53
R27102 vss.n7711 vss.n7701 1054.53
R27103 vss.n7796 vss.n7777 1054.53
R27104 vss.n7796 vss.n7772 1054.53
R27105 vss.n7776 vss.n7775 1054.53
R27106 vss.n7775 vss.n7771 1054.53
R27107 vss.n7781 vss.n7779 1054.53
R27108 vss.n7791 vss.n7781 1054.53
R27109 vss.n7937 vss.n7918 1054.53
R27110 vss.n7937 vss.n7913 1054.53
R27111 vss.n7917 vss.n7916 1054.53
R27112 vss.n7916 vss.n7912 1054.53
R27113 vss.n7922 vss.n7920 1054.53
R27114 vss.n7932 vss.n7922 1054.53
R27115 vss.n8205 vss.n8193 1054.53
R27116 vss.n8205 vss.n8195 1054.53
R27117 vss.n8190 vss.n8188 1054.53
R27118 vss.n8190 vss.n8183 1054.53
R27119 vss.n8187 vss.n8186 1054.53
R27120 vss.n8186 vss.n8182 1054.53
R27121 vss.n8231 vss.n8001 1054.53
R27122 vss.n8231 vss.n7996 1054.53
R27123 vss.n8000 vss.n7999 1054.53
R27124 vss.n7999 vss.n7995 1054.53
R27125 vss.n8005 vss.n8003 1054.53
R27126 vss.n8226 vss.n8005 1054.53
R27127 vss.n8993 vss.n7316 1054.53
R27128 vss.n8993 vss.n7318 1054.53
R27129 vss.n7313 vss.n7311 1054.53
R27130 vss.n7313 vss.n7306 1054.53
R27131 vss.n7310 vss.n7309 1054.53
R27132 vss.n7309 vss.n7305 1054.53
R27133 vss.n8722 vss.n7858 1054.53
R27134 vss.n8722 vss.n7853 1054.53
R27135 vss.n7857 vss.n7856 1054.53
R27136 vss.n7856 vss.n7852 1054.53
R27137 vss.n7862 vss.n7860 1054.53
R27138 vss.n8717 vss.n7862 1054.53
R27139 vss.n8769 vss.n8757 1054.53
R27140 vss.n8769 vss.n8759 1054.53
R27141 vss.n8754 vss.n8752 1054.53
R27142 vss.n8754 vss.n8747 1054.53
R27143 vss.n8751 vss.n8750 1054.53
R27144 vss.n8750 vss.n8746 1054.53
R27145 vss.n8841 vss.n7671 1054.53
R27146 vss.n8841 vss.n7666 1054.53
R27147 vss.n7670 vss.n7669 1054.53
R27148 vss.n7669 vss.n7665 1054.53
R27149 vss.n7675 vss.n7673 1054.53
R27150 vss.n8836 vss.n7675 1054.53
R27151 vss.n8888 vss.n8876 1054.53
R27152 vss.n8888 vss.n8878 1054.53
R27153 vss.n8873 vss.n8871 1054.53
R27154 vss.n8873 vss.n8866 1054.53
R27155 vss.n8870 vss.n8869 1054.53
R27156 vss.n8869 vss.n8865 1054.53
R27157 vss.n8960 vss.n7482 1054.53
R27158 vss.n8960 vss.n7477 1054.53
R27159 vss.n7481 vss.n7480 1054.53
R27160 vss.n7480 vss.n7476 1054.53
R27161 vss.n7486 vss.n7484 1054.53
R27162 vss.n8955 vss.n7486 1054.53
R27163 vss.n8067 vss.n8066 1054.53
R27164 vss.n8066 vss.n8062 1054.53
R27165 vss.n8068 vss.n8065 1054.53
R27166 vss.n8068 vss.n8061 1054.53
R27167 vss.n8074 vss.n8071 1054.53
R27168 vss.n8074 vss.n8073 1054.53
R27169 vss.n9343 vss.n9333 1054.53
R27170 vss.n9333 vss.n9331 1054.53
R27171 vss.n9327 vss.n9323 1054.53
R27172 vss.n9328 vss.n9327 1054.53
R27173 vss.n9348 vss.n9324 1054.53
R27174 vss.n9348 vss.n9329 1054.53
R27175 vss.n6347 vss.n6337 1054.53
R27176 vss.n6337 vss.n6335 1054.53
R27177 vss.n6331 vss.n6327 1054.53
R27178 vss.n6332 vss.n6331 1054.53
R27179 vss.n6352 vss.n6328 1054.53
R27180 vss.n6352 vss.n6333 1054.53
R27181 vss.n6425 vss.n6415 1054.53
R27182 vss.n6415 vss.n6413 1054.53
R27183 vss.n6409 vss.n6405 1054.53
R27184 vss.n6410 vss.n6409 1054.53
R27185 vss.n6430 vss.n6406 1054.53
R27186 vss.n6430 vss.n6411 1054.53
R27187 vss.n6961 vss.n6951 1054.53
R27188 vss.n6951 vss.n6949 1054.53
R27189 vss.n6945 vss.n6941 1054.53
R27190 vss.n6946 vss.n6945 1054.53
R27191 vss.n6966 vss.n6942 1054.53
R27192 vss.n6966 vss.n6947 1054.53
R27193 vss.n6652 vss.n6642 1054.53
R27194 vss.n6642 vss.n6640 1054.53
R27195 vss.n6636 vss.n6632 1054.53
R27196 vss.n6637 vss.n6636 1054.53
R27197 vss.n6657 vss.n6633 1054.53
R27198 vss.n6657 vss.n6638 1054.53
R27199 vss.n7150 vss.n7140 1054.53
R27200 vss.n7140 vss.n7138 1054.53
R27201 vss.n7134 vss.n7130 1054.53
R27202 vss.n7135 vss.n7134 1054.53
R27203 vss.n7155 vss.n7131 1054.53
R27204 vss.n7155 vss.n7136 1054.53
R27205 vss.n9414 vss.n9409 1054.53
R27206 vss.n9414 vss.n9413 1054.53
R27207 vss.n9411 vss.n9406 1054.53
R27208 vss.n9411 vss.n9405 1054.53
R27209 vss.n9436 vss.n9434 1054.53
R27210 vss.n9437 vss.n9436 1054.53
R27211 vss.n6031 vss.n6021 1054.53
R27212 vss.n6021 vss.n6019 1054.53
R27213 vss.n6015 vss.n6011 1054.53
R27214 vss.n6016 vss.n6015 1054.53
R27215 vss.n6036 vss.n6012 1054.53
R27216 vss.n6036 vss.n6017 1054.53
R27217 vss.n9458 vss.n9453 1054.53
R27218 vss.n9458 vss.n9457 1054.53
R27219 vss.n9472 vss.n9452 1054.53
R27220 vss.n9452 vss.n9450 1054.53
R27221 vss.n9478 vss.n9476 1054.53
R27222 vss.n9479 vss.n9478 1054.53
R27223 vss.n6158 vss.n6148 1054.53
R27224 vss.n6148 vss.n6146 1054.53
R27225 vss.n6142 vss.n6138 1054.53
R27226 vss.n6143 vss.n6142 1054.53
R27227 vss.n6163 vss.n6139 1054.53
R27228 vss.n6163 vss.n6144 1054.53
R27229 vss.n7201 vss.n7191 1054.53
R27230 vss.n7191 vss.n7189 1054.53
R27231 vss.n7185 vss.n7181 1054.53
R27232 vss.n7186 vss.n7185 1054.53
R27233 vss.n7206 vss.n7182 1054.53
R27234 vss.n7206 vss.n7187 1054.53
R27235 vss.n6696 vss.n6686 1054.53
R27236 vss.n6686 vss.n6684 1054.53
R27237 vss.n6680 vss.n6676 1054.53
R27238 vss.n6681 vss.n6680 1054.53
R27239 vss.n6701 vss.n6677 1054.53
R27240 vss.n6701 vss.n6682 1054.53
R27241 vss.n7010 vss.n7000 1054.53
R27242 vss.n7000 vss.n6998 1054.53
R27243 vss.n6994 vss.n6990 1054.53
R27244 vss.n6995 vss.n6994 1054.53
R27245 vss.n7015 vss.n6991 1054.53
R27246 vss.n7015 vss.n6996 1054.53
R27247 vss.n6470 vss.n6460 1054.53
R27248 vss.n6460 vss.n6458 1054.53
R27249 vss.n6454 vss.n6450 1054.53
R27250 vss.n6455 vss.n6454 1054.53
R27251 vss.n6475 vss.n6451 1054.53
R27252 vss.n6475 vss.n6456 1054.53
R27253 vss.n9173 vss.n9163 1054.53
R27254 vss.n9163 vss.n9161 1054.53
R27255 vss.n9157 vss.n9153 1054.53
R27256 vss.n9158 vss.n9157 1054.53
R27257 vss.n9178 vss.n9154 1054.53
R27258 vss.n9178 vss.n9159 1054.53
R27259 vss.n6199 vss.n6194 1054.53
R27260 vss.n6199 vss.n6198 1054.53
R27261 vss.n6196 vss.n6191 1054.53
R27262 vss.n6196 vss.n6190 1054.53
R27263 vss.n9374 vss.n9372 1054.53
R27264 vss.n9375 vss.n9374 1054.53
R27265 vss.n9110 vss.n9107 1054.53
R27266 vss.n9110 vss.n9103 1054.53
R27267 vss.n9057 vss.n6550 1054.53
R27268 vss.n9058 vss.n9057 1054.53
R27269 vss.n6540 vss.n6537 1054.53
R27270 vss.n6540 vss.n6533 1054.53
R27271 vss.n6522 vss.n6520 1054.53
R27272 vss.n6522 vss.n6515 1054.53
R27273 vss.n6501 vss.n6493 1054.53
R27274 vss.n6502 vss.n6501 1054.53
R27275 vss.n6862 vss.n6860 1054.53
R27276 vss.n6862 vss.n6855 1054.53
R27277 vss.n6839 vss.n6836 1054.53
R27278 vss.n6839 vss.n6832 1054.53
R27279 vss.n6811 vss.n6809 1054.53
R27280 vss.n6811 vss.n6804 1054.53
R27281 vss.n6790 vss.n6721 1054.53
R27282 vss.n6791 vss.n6790 1054.53
R27283 vss.n6737 vss.n6736 1054.53
R27284 vss.n6737 vss.n6732 1054.53
R27285 vss.n6593 vss.n6590 1054.53
R27286 vss.n6593 vss.n6586 1054.53
R27287 vss.n6129 vss.n6127 1054.53
R27288 vss.n6129 vss.n6122 1054.53
R27289 vss.n6107 vss.n6099 1054.53
R27290 vss.n6108 vss.n6107 1054.53
R27291 vss.n6090 vss.n6088 1054.53
R27292 vss.n6090 vss.n6083 1054.53
R27293 vss.n8029 vss.n8028 1054.53
R27294 vss.n8028 vss.n8024 1054.53
R27295 vss.n8023 vss.n8018 1054.53
R27296 vss.n8041 vss.n8023 1054.53
R27297 vss.n8020 vss.n8014 1054.53
R27298 vss.n8021 vss.n8020 1054.53
R27299 vss.n8131 vss.n8127 1054.53
R27300 vss.n8141 vss.n8131 1054.53
R27301 vss.n8144 vss.n8126 1054.53
R27302 vss.n8126 vss.n6000 1054.53
R27303 vss.n9655 vss.n5990 1054.53
R27304 vss.n9655 vss.n5992 1054.53
R27305 vss.n5987 vss.n5985 1054.53
R27306 vss.n5987 vss.n5980 1054.53
R27307 vss.n5984 vss.n5983 1054.53
R27308 vss.n5983 vss.n5979 1054.53
R27309 vss.n9646 vss.n5997 1054.53
R27310 vss.n9646 vss.n9645 1054.53
R27311 vss.n8111 vss.n8110 1054.53
R27312 vss.n8110 vss.n8106 1054.53
R27313 vss.n8112 vss.n8109 1054.53
R27314 vss.n8112 vss.n8105 1054.53
R27315 vss.n8118 vss.n8115 1054.53
R27316 vss.n8118 vss.n8117 1054.53
R27317 vss.n8541 vss.n8497 1054.53
R27318 vss.n8541 vss.n8498 1054.53
R27319 vss.n8518 vss.n8504 1054.53
R27320 vss.n8529 vss.n8504 1054.53
R27321 vss.n9024 vss.n7284 1054.53
R27322 vss.n9024 vss.n7286 1054.53
R27323 vss.n7281 vss.n7279 1054.53
R27324 vss.n7281 vss.n7274 1054.53
R27325 vss.n7278 vss.n7277 1054.53
R27326 vss.n7277 vss.n7273 1054.53
R27327 vss.n9015 vss.n7291 1054.53
R27328 vss.n9015 vss.n7292 1054.53
R27329 vss.n8269 vss.n8267 1054.53
R27330 vss.n8269 vss.n8262 1054.53
R27331 vss.n8266 vss.n8265 1054.53
R27332 vss.n8265 vss.n8260 1054.53
R27333 vss.n7889 vss.n7888 1054.53
R27334 vss.n7888 vss.n7884 1054.53
R27335 vss.n7890 vss.n7887 1054.53
R27336 vss.n7890 vss.n7883 1054.53
R27337 vss.n7896 vss.n7893 1054.53
R27338 vss.n7896 vss.n7895 1054.53
R27339 vss.n8308 vss.n8307 1054.53
R27340 vss.n8307 vss.n7876 1054.53
R27341 vss.n8309 vss.n8306 1054.53
R27342 vss.n8309 vss.n7875 1054.53
R27343 vss.n8315 vss.n8312 1054.53
R27344 vss.n8315 vss.n8314 1054.53
R27345 vss.n8342 vss.n8337 1054.53
R27346 vss.n8342 vss.n8332 1054.53
R27347 vss.n8336 vss.n8331 1054.53
R27348 vss.n8681 vss.n8331 1054.53
R27349 vss.n8686 vss.n8319 1054.53
R27350 vss.n8686 vss.n8320 1054.53
R27351 vss.n8671 vss.n8349 1054.53
R27352 vss.n8671 vss.n8350 1054.53
R27353 vss.n8359 vss.n8353 1054.53
R27354 vss.n8660 vss.n8353 1054.53
R27355 vss.n8360 vss.n8358 1054.53
R27356 vss.n8360 vss.n8354 1054.53
R27357 vss.n8392 vss.n8387 1054.53
R27358 vss.n8392 vss.n8382 1054.53
R27359 vss.n8386 vss.n8381 1054.53
R27360 vss.n8638 vss.n8381 1054.53
R27361 vss.n8643 vss.n8364 1054.53
R27362 vss.n8643 vss.n8365 1054.53
R27363 vss.n8628 vss.n8399 1054.53
R27364 vss.n8628 vss.n8400 1054.53
R27365 vss.n8412 vss.n8406 1054.53
R27366 vss.n8616 vss.n8406 1054.53
R27367 vss.n8413 vss.n8411 1054.53
R27368 vss.n8413 vss.n8407 1054.53
R27369 vss.n8440 vss.n8435 1054.53
R27370 vss.n8440 vss.n8430 1054.53
R27371 vss.n8434 vss.n8429 1054.53
R27372 vss.n8594 vss.n8429 1054.53
R27373 vss.n8599 vss.n8417 1054.53
R27374 vss.n8599 vss.n8418 1054.53
R27375 vss.n8584 vss.n8447 1054.53
R27376 vss.n8584 vss.n8448 1054.53
R27377 vss.n8457 vss.n8451 1054.53
R27378 vss.n8573 vss.n8451 1054.53
R27379 vss.n8458 vss.n8456 1054.53
R27380 vss.n8458 vss.n8452 1054.53
R27381 vss.n8490 vss.n8485 1054.53
R27382 vss.n8490 vss.n8480 1054.53
R27383 vss.n8484 vss.n8479 1054.53
R27384 vss.n8551 vss.n8479 1054.53
R27385 vss.n8556 vss.n8462 1054.53
R27386 vss.n8556 vss.n8463 1054.53
R27387 vss.n8513 vss.n8512 1054.53
R27388 vss.n8512 vss.n8505 1054.53
R27389 vss.n6068 vss.n6059 1054.53
R27390 vss.n6069 vss.n6068 1054.53
R27391 vss.n9556 vss.n6071 1054.53
R27392 vss.n6071 vss.n6067 1054.53
R27393 vss.n9569 vss.n6060 1054.53
R27394 vss.n9569 vss.n9568 1054.53
R27395 vss.n6087 vss.n6086 1054.53
R27396 vss.n6086 vss.n6082 1054.53
R27397 vss.n7258 vss.n7257 1054.53
R27398 vss.n7257 vss.n7253 1054.53
R27399 vss.n9521 vss.n6110 1054.53
R27400 vss.n6110 vss.n6106 1054.53
R27401 vss.n9534 vss.n6100 1054.53
R27402 vss.n9534 vss.n9533 1054.53
R27403 vss.n6126 vss.n6125 1054.53
R27404 vss.n6125 vss.n6121 1054.53
R27405 vss.n7239 vss.n7238 1054.53
R27406 vss.n7238 vss.n6580 1054.53
R27407 vss.n6761 vss.n6751 1054.53
R27408 vss.n6752 vss.n6751 1054.53
R27409 vss.n6592 vss.n6591 1054.53
R27410 vss.n6591 vss.n6587 1054.53
R27411 vss.n6743 vss.n6740 1054.53
R27412 vss.n6743 vss.n6742 1054.53
R27413 vss.n6733 vss.n6728 1054.53
R27414 vss.n6734 vss.n6733 1054.53
R27415 vss.n7066 vss.n6793 1054.53
R27416 vss.n6793 vss.n6789 1054.53
R27417 vss.n7079 vss.n6722 1054.53
R27418 vss.n7079 vss.n7078 1054.53
R27419 vss.n6808 vss.n6807 1054.53
R27420 vss.n6807 vss.n6803 1054.53
R27421 vss.n6816 vss.n6814 1054.53
R27422 vss.n6817 vss.n6816 1054.53
R27423 vss.n6845 vss.n6842 1054.53
R27424 vss.n6845 vss.n6844 1054.53
R27425 vss.n6838 vss.n6837 1054.53
R27426 vss.n6837 vss.n6833 1054.53
R27427 vss.n6859 vss.n6858 1054.53
R27428 vss.n6858 vss.n6854 1054.53
R27429 vss.n6867 vss.n6865 1054.53
R27430 vss.n6868 vss.n6867 1054.53
R27431 vss.n9229 vss.n6504 1054.53
R27432 vss.n6504 vss.n6500 1054.53
R27433 vss.n9242 vss.n6494 1054.53
R27434 vss.n9242 vss.n9241 1054.53
R27435 vss.n6519 vss.n6518 1054.53
R27436 vss.n6518 vss.n6514 1054.53
R27437 vss.n6527 vss.n6525 1054.53
R27438 vss.n6558 vss.n6527 1054.53
R27439 vss.n9079 vss.n9069 1054.53
R27440 vss.n9070 vss.n9069 1054.53
R27441 vss.n6539 vss.n6538 1054.53
R27442 vss.n6538 vss.n6534 1054.53
R27443 vss.n9087 vss.n9060 1054.53
R27444 vss.n9060 vss.n9056 1054.53
R27445 vss.n6554 vss.n6551 1054.53
R27446 vss.n9051 vss.n6554 1054.53
R27447 vss.n9116 vss.n9113 1054.53
R27448 vss.n9116 vss.n9115 1054.53
R27449 vss.n9109 vss.n9108 1054.53
R27450 vss.n9108 vss.n9104 1054.53
R27451 vss.n5964 vss.n5946 1054.53
R27452 vss.n5964 vss.n5941 1054.53
R27453 vss.n5945 vss.n5944 1054.53
R27454 vss.n5944 vss.n5940 1054.53
R27455 vss.n5950 vss.n5948 1054.53
R27456 vss.n5959 vss.n5950 1054.53
R27457 vss.n9882 vss.n2760 1054.53
R27458 vss.n9882 vss.n2762 1054.53
R27459 vss.n2757 vss.n2755 1054.53
R27460 vss.n2757 vss.n2750 1054.53
R27461 vss.n2754 vss.n2753 1054.53
R27462 vss.n2753 vss.n2749 1054.53
R27463 vss.n9714 vss.n9694 1054.53
R27464 vss.n9714 vss.n9689 1054.53
R27465 vss.n9693 vss.n9692 1054.53
R27466 vss.n9692 vss.n9688 1054.53
R27467 vss.n9698 vss.n9696 1054.53
R27468 vss.n9709 vss.n9698 1054.53
R27469 vss.n3295 vss.n3272 1054.53
R27470 vss.n3295 vss.n3267 1054.53
R27471 vss.n3271 vss.n3270 1054.53
R27472 vss.n3270 vss.n3266 1054.53
R27473 vss.n3276 vss.n3274 1054.53
R27474 vss.n3287 vss.n3276 1054.53
R27475 vss.n2585 vss.n2567 1054.53
R27476 vss.n2585 vss.n2562 1054.53
R27477 vss.n2566 vss.n2565 1054.53
R27478 vss.n2565 vss.n2561 1054.53
R27479 vss.n2571 vss.n2569 1054.53
R27480 vss.n2580 vss.n2571 1054.53
R27481 vss.n5912 vss.n5902 1054.53
R27482 vss.n5902 vss.n5900 1054.53
R27483 vss.n5896 vss.n5892 1054.53
R27484 vss.n5897 vss.n5896 1054.53
R27485 vss.n5917 vss.n5893 1054.53
R27486 vss.n5917 vss.n5898 1054.53
R27487 vss.n9775 vss.n9748 1054.53
R27488 vss.n9781 vss.n9748 1054.53
R27489 vss.n9757 vss.n9753 1054.53
R27490 vss.n9757 vss.n9747 1054.53
R27491 vss.n9759 vss.n9755 1054.53
R27492 vss.n9768 vss.n9759 1054.53
R27493 vss.n3215 vss.n3188 1054.53
R27494 vss.n3221 vss.n3188 1054.53
R27495 vss.n3197 vss.n3193 1054.53
R27496 vss.n3197 vss.n3187 1054.53
R27497 vss.n3199 vss.n3195 1054.53
R27498 vss.n3208 vss.n3199 1054.53
R27499 vss.n3017 vss.n3010 1054.53
R27500 vss.n3023 vss.n3010 1054.53
R27501 vss.n3007 vss.n3000 1054.53
R27502 vss.n3007 vss.n3004 1054.53
R27503 vss.n3002 vss.n2996 1054.53
R27504 vss.n3003 vss.n3002 1054.53
R27505 vss.n5245 vss.n5218 1054.53
R27506 vss.n5251 vss.n5218 1054.53
R27507 vss.n5227 vss.n5223 1054.53
R27508 vss.n5227 vss.n5217 1054.53
R27509 vss.n5229 vss.n5225 1054.53
R27510 vss.n5238 vss.n5229 1054.53
R27511 vss.n3058 vss.n3031 1054.53
R27512 vss.n3064 vss.n3031 1054.53
R27513 vss.n3040 vss.n3036 1054.53
R27514 vss.n3040 vss.n3030 1054.53
R27515 vss.n3042 vss.n3038 1054.53
R27516 vss.n3051 vss.n3042 1054.53
R27517 vss.n5115 vss.n5088 1054.53
R27518 vss.n5121 vss.n5088 1054.53
R27519 vss.n5097 vss.n5093 1054.53
R27520 vss.n5097 vss.n5087 1054.53
R27521 vss.n5099 vss.n5095 1054.53
R27522 vss.n5108 vss.n5099 1054.53
R27523 vss.n5304 vss.n5277 1054.53
R27524 vss.n5310 vss.n5277 1054.53
R27525 vss.n5286 vss.n5282 1054.53
R27526 vss.n5286 vss.n5276 1054.53
R27527 vss.n5288 vss.n5284 1054.53
R27528 vss.n5297 vss.n5288 1054.53
R27529 vss.n5032 vss.n5005 1054.53
R27530 vss.n5038 vss.n5005 1054.53
R27531 vss.n5014 vss.n5010 1054.53
R27532 vss.n5014 vss.n5004 1054.53
R27533 vss.n5016 vss.n5012 1054.53
R27534 vss.n5025 vss.n5016 1054.53
R27535 vss.n4913 vss.n4886 1054.53
R27536 vss.n4919 vss.n4886 1054.53
R27537 vss.n4895 vss.n4891 1054.53
R27538 vss.n4895 vss.n4885 1054.53
R27539 vss.n4897 vss.n4893 1054.53
R27540 vss.n4906 vss.n4897 1054.53
R27541 vss.n5394 vss.n5350 1054.53
R27542 vss.n5394 vss.n5351 1054.53
R27543 vss.n5371 vss.n5357 1054.53
R27544 vss.n5382 vss.n5357 1054.53
R27545 vss.n9916 vss.n2725 1054.53
R27546 vss.n9916 vss.n2727 1054.53
R27547 vss.n2722 vss.n2720 1054.53
R27548 vss.n2722 vss.n2715 1054.53
R27549 vss.n2719 vss.n2718 1054.53
R27550 vss.n2718 vss.n2714 1054.53
R27551 vss.n9907 vss.n2732 1054.53
R27552 vss.n9907 vss.n2733 1054.53
R27553 vss.n4653 vss.n4651 1054.53
R27554 vss.n4653 vss.n4646 1054.53
R27555 vss.n4650 vss.n4649 1054.53
R27556 vss.n4649 vss.n4644 1054.53
R27557 vss.n5618 vss.n4677 1054.53
R27558 vss.n5618 vss.n4679 1054.53
R27559 vss.n4674 vss.n4672 1054.53
R27560 vss.n4674 vss.n4636 1054.53
R27561 vss.n4671 vss.n4670 1054.53
R27562 vss.n4670 vss.n4635 1054.53
R27563 vss.n5609 vss.n4684 1054.53
R27564 vss.n5609 vss.n4685 1054.53
R27565 vss.n4694 vss.n4688 1054.53
R27566 vss.n5598 vss.n4688 1054.53
R27567 vss.n4695 vss.n4693 1054.53
R27568 vss.n4695 vss.n4689 1054.53
R27569 vss.n4720 vss.n4715 1054.53
R27570 vss.n4720 vss.n4710 1054.53
R27571 vss.n4714 vss.n4709 1054.53
R27572 vss.n5576 vss.n4709 1054.53
R27573 vss.n5581 vss.n4699 1054.53
R27574 vss.n5581 vss.n4700 1054.53
R27575 vss.n5566 vss.n4727 1054.53
R27576 vss.n5566 vss.n4728 1054.53
R27577 vss.n4737 vss.n4731 1054.53
R27578 vss.n5555 vss.n4731 1054.53
R27579 vss.n4738 vss.n4736 1054.53
R27580 vss.n4738 vss.n4732 1054.53
R27581 vss.n4763 vss.n4758 1054.53
R27582 vss.n4763 vss.n4753 1054.53
R27583 vss.n4757 vss.n4752 1054.53
R27584 vss.n5533 vss.n4752 1054.53
R27585 vss.n5538 vss.n4742 1054.53
R27586 vss.n5538 vss.n4743 1054.53
R27587 vss.n5523 vss.n4770 1054.53
R27588 vss.n5523 vss.n4771 1054.53
R27589 vss.n4780 vss.n4774 1054.53
R27590 vss.n5512 vss.n4774 1054.53
R27591 vss.n4781 vss.n4779 1054.53
R27592 vss.n4781 vss.n4775 1054.53
R27593 vss.n4806 vss.n4801 1054.53
R27594 vss.n4806 vss.n4796 1054.53
R27595 vss.n4800 vss.n4795 1054.53
R27596 vss.n5490 vss.n4795 1054.53
R27597 vss.n5495 vss.n4785 1054.53
R27598 vss.n5495 vss.n4786 1054.53
R27599 vss.n5480 vss.n4813 1054.53
R27600 vss.n5480 vss.n4814 1054.53
R27601 vss.n4823 vss.n4817 1054.53
R27602 vss.n5469 vss.n4817 1054.53
R27603 vss.n4824 vss.n4822 1054.53
R27604 vss.n4824 vss.n4818 1054.53
R27605 vss.n4849 vss.n4844 1054.53
R27606 vss.n4849 vss.n4839 1054.53
R27607 vss.n4843 vss.n4838 1054.53
R27608 vss.n5447 vss.n4838 1054.53
R27609 vss.n5452 vss.n4828 1054.53
R27610 vss.n5452 vss.n4829 1054.53
R27611 vss.n5437 vss.n4856 1054.53
R27612 vss.n5437 vss.n4857 1054.53
R27613 vss.n4866 vss.n4860 1054.53
R27614 vss.n5426 vss.n4860 1054.53
R27615 vss.n4867 vss.n4865 1054.53
R27616 vss.n4867 vss.n4861 1054.53
R27617 vss.n5343 vss.n5338 1054.53
R27618 vss.n5343 vss.n5333 1054.53
R27619 vss.n5337 vss.n5332 1054.53
R27620 vss.n5404 vss.n5332 1054.53
R27621 vss.n5409 vss.n4871 1054.53
R27622 vss.n5409 vss.n4872 1054.53
R27623 vss.n5366 vss.n5365 1054.53
R27624 vss.n5365 vss.n5358 1054.53
R27625 vss.n9834 vss.n2876 1054.53
R27626 vss.n9840 vss.n2876 1054.53
R27627 vss.n2885 vss.n2881 1054.53
R27628 vss.n2885 vss.n2875 1054.53
R27629 vss.n2887 vss.n2883 1054.53
R27630 vss.n9827 vss.n2887 1054.53
R27631 vss.n2960 vss.n2953 1054.53
R27632 vss.n2966 vss.n2953 1054.53
R27633 vss.n2950 vss.n2943 1054.53
R27634 vss.n2950 vss.n2947 1054.53
R27635 vss.n2945 vss.n2939 1054.53
R27636 vss.n2946 vss.n2945 1054.53
R27637 vss.n2913 vss.n2906 1054.53
R27638 vss.n2919 vss.n2906 1054.53
R27639 vss.n2903 vss.n2896 1054.53
R27640 vss.n2903 vss.n2900 1054.53
R27641 vss.n2898 vss.n2892 1054.53
R27642 vss.n2899 vss.n2898 1054.53
R27643 vss.n4954 vss.n4927 1054.53
R27644 vss.n4960 vss.n4927 1054.53
R27645 vss.n4936 vss.n4932 1054.53
R27646 vss.n4936 vss.n4926 1054.53
R27647 vss.n4938 vss.n4934 1054.53
R27648 vss.n4947 vss.n4938 1054.53
R27649 vss.n5156 vss.n5129 1054.53
R27650 vss.n5162 vss.n5129 1054.53
R27651 vss.n5138 vss.n5134 1054.53
R27652 vss.n5138 vss.n5128 1054.53
R27653 vss.n5140 vss.n5136 1054.53
R27654 vss.n5149 vss.n5140 1054.53
R27655 vss.n3137 vss.n3109 1054.53
R27656 vss.n3143 vss.n3109 1054.53
R27657 vss.n3118 vss.n3114 1054.53
R27658 vss.n3118 vss.n3108 1054.53
R27659 vss.n3120 vss.n3116 1054.53
R27660 vss.n3130 vss.n3120 1054.53
R27661 vss.n4472 vss.n4464 1054.53
R27662 vss.n4473 vss.n4472 1054.53
R27663 vss.n4485 vss.n4475 1054.53
R27664 vss.n4475 vss.n4471 1054.53
R27665 vss.n4498 vss.n4465 1054.53
R27666 vss.n4498 vss.n4497 1054.53
R27667 vss.n4380 vss.n4372 1054.53
R27668 vss.n4381 vss.n4380 1054.53
R27669 vss.n4393 vss.n4383 1054.53
R27670 vss.n4383 vss.n4379 1054.53
R27671 vss.n4406 vss.n4373 1054.53
R27672 vss.n4406 vss.n4405 1054.53
R27673 vss.n4332 vss.n4324 1054.53
R27674 vss.n4333 vss.n4332 1054.53
R27675 vss.n4345 vss.n4335 1054.53
R27676 vss.n4335 vss.n4331 1054.53
R27677 vss.n4358 vss.n4325 1054.53
R27678 vss.n4358 vss.n4357 1054.53
R27679 vss.n3732 vss.n3724 1054.53
R27680 vss.n3733 vss.n3732 1054.53
R27681 vss.n3745 vss.n3735 1054.53
R27682 vss.n3735 vss.n3731 1054.53
R27683 vss.n3758 vss.n3725 1054.53
R27684 vss.n3758 vss.n3757 1054.53
R27685 vss.n4034 vss.n4026 1054.53
R27686 vss.n4035 vss.n4034 1054.53
R27687 vss.n4047 vss.n4037 1054.53
R27688 vss.n4037 vss.n4033 1054.53
R27689 vss.n4060 vss.n4027 1054.53
R27690 vss.n4060 vss.n4059 1054.53
R27691 vss.n3687 vss.n3679 1054.53
R27692 vss.n3688 vss.n3687 1054.53
R27693 vss.n3700 vss.n3690 1054.53
R27694 vss.n3690 vss.n3686 1054.53
R27695 vss.n3713 vss.n3680 1054.53
R27696 vss.n3713 vss.n3712 1054.53
R27697 vss.n4088 vss.n4080 1054.53
R27698 vss.n4089 vss.n4088 1054.53
R27699 vss.n4101 vss.n4091 1054.53
R27700 vss.n4091 vss.n4087 1054.53
R27701 vss.n4114 vss.n4081 1054.53
R27702 vss.n4114 vss.n4113 1054.53
R27703 vss.n3512 vss.n3504 1054.53
R27704 vss.n3513 vss.n3512 1054.53
R27705 vss.n3525 vss.n3515 1054.53
R27706 vss.n3515 vss.n3511 1054.53
R27707 vss.n3538 vss.n3505 1054.53
R27708 vss.n3538 vss.n3537 1054.53
R27709 vss.n3467 vss.n3459 1054.53
R27710 vss.n3468 vss.n3467 1054.53
R27711 vss.n3480 vss.n3470 1054.53
R27712 vss.n3470 vss.n3466 1054.53
R27713 vss.n3493 vss.n3460 1054.53
R27714 vss.n3493 vss.n3492 1054.53
R27715 vss.n5755 vss.n5747 1054.53
R27716 vss.n5756 vss.n5755 1054.53
R27717 vss.n5768 vss.n5758 1054.53
R27718 vss.n5758 vss.n5754 1054.53
R27719 vss.n5781 vss.n5748 1054.53
R27720 vss.n5781 vss.n5780 1054.53
R27721 vss.n5704 vss.n5701 1054.53
R27722 vss.n5704 vss.n5697 1054.53
R27723 vss.n5651 vss.n3606 1054.53
R27724 vss.n5652 vss.n5651 1054.53
R27725 vss.n3596 vss.n3593 1054.53
R27726 vss.n3596 vss.n3589 1054.53
R27727 vss.n3576 vss.n3574 1054.53
R27728 vss.n3576 vss.n3569 1054.53
R27729 vss.n3555 vss.n3547 1054.53
R27730 vss.n3556 vss.n3555 1054.53
R27731 vss.n3905 vss.n3903 1054.53
R27732 vss.n3905 vss.n3898 1054.53
R27733 vss.n3882 vss.n3879 1054.53
R27734 vss.n3882 vss.n3875 1054.53
R27735 vss.n3853 vss.n3851 1054.53
R27736 vss.n3853 vss.n3846 1054.53
R27737 vss.n3832 vss.n3806 1054.53
R27738 vss.n3833 vss.n3832 1054.53
R27739 vss.n3797 vss.n3795 1054.53
R27740 vss.n3797 vss.n3790 1054.53
R27741 vss.n3776 vss.n3766 1054.53
R27742 vss.n3777 vss.n3776 1054.53
R27743 vss.n3643 vss.n3640 1054.53
R27744 vss.n3643 vss.n3636 1054.53
R27745 vss.n4562 vss.n4416 1054.53
R27746 vss.n4563 vss.n4562 1054.53
R27747 vss.n4433 vss.n4432 1054.53
R27748 vss.n4433 vss.n4428 1054.53
R27749 vss.n4452 vss.n4448 1054.53
R27750 vss.n4453 vss.n4452 1054.53
R27751 vss.n4533 vss.n4447 1054.53
R27752 vss.n4450 vss.n4447 1054.53
R27753 vss.n4512 vss.n4456 1054.53
R27754 vss.n4513 vss.n4512 1054.53
R27755 vss.n4439 vss.n4436 1054.53
R27756 vss.n4439 vss.n4438 1054.53
R27757 vss.n4429 vss.n4424 1054.53
R27758 vss.n4430 vss.n4429 1054.53
R27759 vss.n4592 vss.n4565 1054.53
R27760 vss.n4565 vss.n4561 1054.53
R27761 vss.n4605 vss.n4417 1054.53
R27762 vss.n4605 vss.n4604 1054.53
R27763 vss.n4578 vss.n4577 1054.53
R27764 vss.n4577 vss.n4575 1054.53
R27765 vss.n3642 vss.n3641 1054.53
R27766 vss.n3641 vss.n3637 1054.53
R27767 vss.n4189 vss.n3779 1054.53
R27768 vss.n3779 vss.n3775 1054.53
R27769 vss.n4202 vss.n3767 1054.53
R27770 vss.n4202 vss.n4201 1054.53
R27771 vss.n3794 vss.n3793 1054.53
R27772 vss.n3793 vss.n3789 1054.53
R27773 vss.n3817 vss.n3813 1054.53
R27774 vss.n3818 vss.n3817 1054.53
R27775 vss.n4154 vss.n3835 1054.53
R27776 vss.n3835 vss.n3831 1054.53
R27777 vss.n4167 vss.n3807 1054.53
R27778 vss.n4167 vss.n4166 1054.53
R27779 vss.n3850 vss.n3849 1054.53
R27780 vss.n3849 vss.n3845 1054.53
R27781 vss.n3859 vss.n3857 1054.53
R27782 vss.n3860 vss.n3859 1054.53
R27783 vss.n3888 vss.n3885 1054.53
R27784 vss.n3888 vss.n3887 1054.53
R27785 vss.n3881 vss.n3880 1054.53
R27786 vss.n3880 vss.n3876 1054.53
R27787 vss.n3902 vss.n3901 1054.53
R27788 vss.n3901 vss.n3897 1054.53
R27789 vss.n3910 vss.n3908 1054.53
R27790 vss.n3911 vss.n3910 1054.53
R27791 vss.n5821 vss.n3558 1054.53
R27792 vss.n3558 vss.n3554 1054.53
R27793 vss.n5834 vss.n3548 1054.53
R27794 vss.n5834 vss.n5833 1054.53
R27795 vss.n3573 vss.n3572 1054.53
R27796 vss.n3572 vss.n3568 1054.53
R27797 vss.n3583 vss.n3581 1054.53
R27798 vss.n3614 vss.n3583 1054.53
R27799 vss.n5673 vss.n5663 1054.53
R27800 vss.n5664 vss.n5663 1054.53
R27801 vss.n3595 vss.n3594 1054.53
R27802 vss.n3594 vss.n3590 1054.53
R27803 vss.n5681 vss.n5654 1054.53
R27804 vss.n5654 vss.n5650 1054.53
R27805 vss.n3610 vss.n3607 1054.53
R27806 vss.n5645 vss.n3610 1054.53
R27807 vss.n5710 vss.n5707 1054.53
R27808 vss.n5710 vss.n5709 1054.53
R27809 vss.n5703 vss.n5702 1054.53
R27810 vss.n5702 vss.n5698 1054.53
R27811 vss.n9959 vss.n2634 1054.53
R27812 vss.n9960 vss.n9959 1054.53
R27813 vss.n9972 vss.n9962 1054.53
R27814 vss.n9962 vss.n9958 1054.53
R27815 vss.n9985 vss.n2635 1054.53
R27816 vss.n9985 vss.n9984 1054.53
R27817 vss.n2652 vss.n2649 1054.53
R27818 vss.n2652 vss.n2645 1054.53
R27819 vss.n2658 vss.n2655 1054.53
R27820 vss.n2658 vss.n2657 1054.53
R27821 vss.n2651 vss.n2650 1054.53
R27822 vss.n2650 vss.n2646 1054.53
R27823 vss.n3392 vss.n3384 1054.53
R27824 vss.n3393 vss.n3392 1054.53
R27825 vss.n3405 vss.n3395 1054.53
R27826 vss.n3395 vss.n3391 1054.53
R27827 vss.n3418 vss.n3385 1054.53
R27828 vss.n3418 vss.n3417 1054.53
R27829 vss.n3989 vss.n3981 1054.53
R27830 vss.n3990 vss.n3989 1054.53
R27831 vss.n4002 vss.n3992 1054.53
R27832 vss.n3992 vss.n3988 1054.53
R27833 vss.n4015 vss.n3982 1054.53
R27834 vss.n4015 vss.n4014 1054.53
R27835 vss.n4256 vss.n4248 1054.53
R27836 vss.n4257 vss.n4256 1054.53
R27837 vss.n4269 vss.n4259 1054.53
R27838 vss.n4259 vss.n4255 1054.53
R27839 vss.n4282 vss.n4249 1054.53
R27840 vss.n4282 vss.n4281 1054.53
R27841 vss.n492 vss.n488 1054.53
R27842 vss.n14071 vss.n492 1054.53
R27843 vss.n10133 vss.n10106 1054.53
R27844 vss.n10139 vss.n10106 1054.53
R27845 vss.n10115 vss.n10111 1054.53
R27846 vss.n10115 vss.n10105 1054.53
R27847 vss.n10117 vss.n10113 1054.53
R27848 vss.n10126 vss.n10117 1054.53
R27849 vss.n12891 vss.n12864 1054.53
R27850 vss.n12897 vss.n12864 1054.53
R27851 vss.n12873 vss.n12869 1054.53
R27852 vss.n12873 vss.n12863 1054.53
R27853 vss.n12875 vss.n12871 1054.53
R27854 vss.n12884 vss.n12875 1054.53
R27855 vss.n10174 vss.n10147 1054.53
R27856 vss.n10180 vss.n10147 1054.53
R27857 vss.n10156 vss.n10152 1054.53
R27858 vss.n10156 vss.n10146 1054.53
R27859 vss.n10158 vss.n10154 1054.53
R27860 vss.n10167 vss.n10158 1054.53
R27861 vss.n12440 vss.n12413 1054.53
R27862 vss.n12446 vss.n12413 1054.53
R27863 vss.n12422 vss.n12418 1054.53
R27864 vss.n12422 vss.n12412 1054.53
R27865 vss.n12424 vss.n12420 1054.53
R27866 vss.n12433 vss.n12424 1054.53
R27867 vss.n11769 vss.n11742 1054.53
R27868 vss.n11775 vss.n11742 1054.53
R27869 vss.n11751 vss.n11747 1054.53
R27870 vss.n11751 vss.n11741 1054.53
R27871 vss.n11753 vss.n11749 1054.53
R27872 vss.n11762 vss.n11753 1054.53
R27873 vss.n12485 vss.n12458 1054.53
R27874 vss.n12491 vss.n12458 1054.53
R27875 vss.n12467 vss.n12463 1054.53
R27876 vss.n12467 vss.n12457 1054.53
R27877 vss.n12469 vss.n12465 1054.53
R27878 vss.n12478 vss.n12469 1054.53
R27879 vss.n2330 vss.n2323 1054.53
R27880 vss.n2336 vss.n2323 1054.53
R27881 vss.n2320 vss.n2313 1054.53
R27882 vss.n2320 vss.n2317 1054.53
R27883 vss.n2315 vss.n2309 1054.53
R27884 vss.n2316 vss.n2315 1054.53
R27885 vss.n12310 vss.n12283 1054.53
R27886 vss.n12316 vss.n12283 1054.53
R27887 vss.n12292 vss.n12288 1054.53
R27888 vss.n12292 vss.n12282 1054.53
R27889 vss.n12294 vss.n12290 1054.53
R27890 vss.n12303 vss.n12294 1054.53
R27891 vss.n12355 vss.n12328 1054.53
R27892 vss.n12361 vss.n12328 1054.53
R27893 vss.n12337 vss.n12333 1054.53
R27894 vss.n12337 vss.n12327 1054.53
R27895 vss.n12339 vss.n12335 1054.53
R27896 vss.n12348 vss.n12339 1054.53
R27897 vss.n10251 vss.n10224 1054.53
R27898 vss.n10257 vss.n10224 1054.53
R27899 vss.n10233 vss.n10229 1054.53
R27900 vss.n10233 vss.n10223 1054.53
R27901 vss.n10235 vss.n10231 1054.53
R27902 vss.n10244 vss.n10235 1054.53
R27903 vss.n2431 vss.n2404 1054.53
R27904 vss.n2437 vss.n2404 1054.53
R27905 vss.n2413 vss.n2409 1054.53
R27906 vss.n2413 vss.n2403 1054.53
R27907 vss.n2415 vss.n2411 1054.53
R27908 vss.n2424 vss.n2415 1054.53
R27909 vss.n2390 vss.n2383 1054.53
R27910 vss.n2396 vss.n2383 1054.53
R27911 vss.n2380 vss.n2373 1054.53
R27912 vss.n2380 vss.n2377 1054.53
R27913 vss.n2375 vss.n2369 1054.53
R27914 vss.n2376 vss.n2375 1054.53
R27915 vss.n10052 vss.n10026 1054.53
R27916 vss.n10052 vss.n10021 1054.53
R27917 vss.n10025 vss.n10024 1054.53
R27918 vss.n10024 vss.n10020 1054.53
R27919 vss.n10030 vss.n10028 1054.53
R27920 vss.n10047 vss.n10030 1054.53
R27921 vss.n2112 vss.n2107 1054.53
R27922 vss.n2112 vss.n2102 1054.53
R27923 vss.n2106 vss.n2101 1054.53
R27924 vss.n13085 vss.n2101 1054.53
R27925 vss.n13090 vss.n2096 1054.53
R27926 vss.n13090 vss.n2097 1054.53
R27927 vss.n2511 vss.n2483 1054.53
R27928 vss.n2517 vss.n2483 1054.53
R27929 vss.n2492 vss.n2488 1054.53
R27930 vss.n2492 vss.n2482 1054.53
R27931 vss.n2494 vss.n2490 1054.53
R27932 vss.n2504 vss.n2494 1054.53
R27933 vss.n12113 vss.n11829 1054.53
R27934 vss.n12114 vss.n12113 1054.53
R27935 vss.n11840 vss.n11839 1054.53
R27936 vss.n11840 vss.n11837 1054.53
R27937 vss.n11846 vss.n11843 1054.53
R27938 vss.n11846 vss.n11845 1054.53
R27939 vss.n11821 vss.n11814 1054.53
R27940 vss.n11821 vss.n11818 1054.53
R27941 vss.n11816 vss.n11810 1054.53
R27942 vss.n11817 vss.n11816 1054.53
R27943 vss.n11802 vss.n11799 1054.53
R27944 vss.n11802 vss.n11801 1054.53
R27945 vss.n12184 vss.n12180 1054.53
R27946 vss.n12184 vss.n11783 1054.53
R27947 vss.n12258 vss.n12182 1054.53
R27948 vss.n12259 vss.n12258 1054.53
R27949 vss.n12198 vss.n12192 1054.53
R27950 vss.n12199 vss.n12198 1054.53
R27951 vss.n11733 vss.n11726 1054.53
R27952 vss.n11733 vss.n11730 1054.53
R27953 vss.n11728 vss.n11722 1054.53
R27954 vss.n11729 vss.n11728 1054.53
R27955 vss.n11715 vss.n11712 1054.53
R27956 vss.n11715 vss.n11714 1054.53
R27957 vss.n11693 vss.n11630 1054.53
R27958 vss.n12579 vss.n11630 1054.53
R27959 vss.n11689 vss.n11688 1054.53
R27960 vss.n11688 vss.n11629 1054.53
R27961 vss.n11649 vss.n11643 1054.53
R27962 vss.n11650 vss.n11649 1054.53
R27963 vss.n10316 vss.n10312 1054.53
R27964 vss.n10316 vss.n10306 1054.53
R27965 vss.n12838 vss.n10314 1054.53
R27966 vss.n12839 vss.n12838 1054.53
R27967 vss.n12780 vss.n12774 1054.53
R27968 vss.n12781 vss.n12780 1054.53
R27969 vss.n10098 vss.n10091 1054.53
R27970 vss.n10098 vss.n10095 1054.53
R27971 vss.n10093 vss.n10087 1054.53
R27972 vss.n10094 vss.n10093 1054.53
R27973 vss.n11876 vss.n11873 1054.53
R27974 vss.n11876 vss.n11875 1054.53
R27975 vss.n11869 vss.n11868 1054.53
R27976 vss.n11868 vss.n11864 1054.53
R27977 vss.n10472 vss.n10464 1054.53
R27978 vss.n10473 vss.n10472 1054.53
R27979 vss.n10484 vss.n10475 1054.53
R27980 vss.n10475 vss.n10471 1054.53
R27981 vss.n10497 vss.n10465 1054.53
R27982 vss.n10497 vss.n10496 1054.53
R27983 vss.n10693 vss.n10685 1054.53
R27984 vss.n10694 vss.n10693 1054.53
R27985 vss.n10705 vss.n10696 1054.53
R27986 vss.n10696 vss.n10692 1054.53
R27987 vss.n10718 vss.n10686 1054.53
R27988 vss.n10718 vss.n10717 1054.53
R27989 vss.n11007 vss.n10999 1054.53
R27990 vss.n11008 vss.n11007 1054.53
R27991 vss.n11019 vss.n11010 1054.53
R27992 vss.n11010 vss.n11006 1054.53
R27993 vss.n11032 vss.n11000 1054.53
R27994 vss.n11032 vss.n11031 1054.53
R27995 vss.n13114 vss.n13113 854.47
R27996 vss.n5643 vss.n3611 814.227
R27997 vss.n9049 vss.n6555 814.227
R27998 vss.n8122 vss.n5973 814.227
R27999 vss.n13922 vss.n13921 814.227
R28000 vss.n12099 vss.n12098 814.227
R28001 vss.n11076 vss.n10433 759.029
R28002 vss.n11091 vss.n11083 759.029
R28003 vss.n11092 vss.n11091 759.029
R28004 vss.n11092 vss.n11089 759.029
R28005 vss.n11076 vss.n10432 759.029
R28006 vss.n11081 vss.n10432 759.029
R28007 vss.n11081 vss.n10431 759.029
R28008 vss.n11078 vss.n10431 759.029
R28009 vss.n11096 vss.n11089 759.029
R28010 vss.n11097 vss.n11096 759.029
R28011 vss.n11098 vss.n11097 759.029
R28012 vss.n11078 vss.n10430 759.029
R28013 vss.n11072 vss.n10436 759.029
R28014 vss.n11161 vss.n11158 759.029
R28015 vss.n11167 vss.n11161 759.029
R28016 vss.n11167 vss.n11166 759.029
R28017 vss.n11072 vss.n10435 759.029
R28018 vss.n11156 vss.n10435 759.029
R28019 vss.n11156 vss.n10434 759.029
R28020 vss.n11074 vss.n10434 759.029
R28021 vss.n11166 vss.n11165 759.029
R28022 vss.n11165 vss.n11162 759.029
R28023 vss.n11162 vss.n11047 759.029
R28024 vss.n11074 vss.n10429 759.029
R28025 vss.n11068 vss.n10439 759.029
R28026 vss.n11186 vss.n11178 759.029
R28027 vss.n11187 vss.n11186 759.029
R28028 vss.n11187 vss.n11184 759.029
R28029 vss.n11068 vss.n10438 759.029
R28030 vss.n11176 vss.n10438 759.029
R28031 vss.n11176 vss.n10437 759.029
R28032 vss.n11070 vss.n10437 759.029
R28033 vss.n11191 vss.n11184 759.029
R28034 vss.n11192 vss.n11191 759.029
R28035 vss.n11193 vss.n11192 759.029
R28036 vss.n11070 vss.n10428 759.029
R28037 vss.n11064 vss.n10442 759.029
R28038 vss.n11217 vss.n11209 759.029
R28039 vss.n11218 vss.n11217 759.029
R28040 vss.n11218 vss.n11215 759.029
R28041 vss.n11064 vss.n10441 759.029
R28042 vss.n11207 vss.n10441 759.029
R28043 vss.n11207 vss.n10440 759.029
R28044 vss.n11066 vss.n10440 759.029
R28045 vss.n11222 vss.n11215 759.029
R28046 vss.n11223 vss.n11222 759.029
R28047 vss.n11224 vss.n11223 759.029
R28048 vss.n11066 vss.n10427 759.029
R28049 vss.n11060 vss.n10445 759.029
R28050 vss.n11243 vss.n11240 759.029
R28051 vss.n11258 vss.n11243 759.029
R28052 vss.n11258 vss.n11257 759.029
R28053 vss.n11060 vss.n10444 759.029
R28054 vss.n11238 vss.n10444 759.029
R28055 vss.n11238 vss.n10443 759.029
R28056 vss.n11062 vss.n10443 759.029
R28057 vss.n11257 vss.n11256 759.029
R28058 vss.n11256 vss.n11244 759.029
R28059 vss.n11252 vss.n11244 759.029
R28060 vss.n11062 vss.n10426 759.029
R28061 vss.n11056 vss.n10448 759.029
R28062 vss.n11278 vss.n11270 759.029
R28063 vss.n11279 vss.n11278 759.029
R28064 vss.n11279 vss.n11276 759.029
R28065 vss.n11056 vss.n10447 759.029
R28066 vss.n11268 vss.n10447 759.029
R28067 vss.n11268 vss.n10446 759.029
R28068 vss.n11058 vss.n10446 759.029
R28069 vss.n11283 vss.n11276 759.029
R28070 vss.n11284 vss.n11283 759.029
R28071 vss.n11285 vss.n11284 759.029
R28072 vss.n11058 vss.n10425 759.029
R28073 vss.n11052 vss.n10451 759.029
R28074 vss.n11304 vss.n11301 759.029
R28075 vss.n11319 vss.n11304 759.029
R28076 vss.n11319 vss.n11318 759.029
R28077 vss.n11052 vss.n10450 759.029
R28078 vss.n11299 vss.n10450 759.029
R28079 vss.n11299 vss.n10449 759.029
R28080 vss.n11054 vss.n10449 759.029
R28081 vss.n11318 vss.n11317 759.029
R28082 vss.n11317 vss.n11305 759.029
R28083 vss.n11313 vss.n11305 759.029
R28084 vss.n11054 vss.n10424 759.029
R28085 vss.n3330 vss.n2603 759.029
R28086 vss.n3335 vss.n3325 759.029
R28087 vss.n3325 vss.n3311 759.029
R28088 vss.n5884 vss.n3311 759.029
R28089 vss.n3330 vss.n2602 759.029
R28090 vss.n5885 vss.n2602 759.029
R28091 vss.n5885 vss.n2601 759.029
R28092 vss.n3316 vss.n2601 759.029
R28093 vss.n5884 vss.n5883 759.029
R28094 vss.n5883 vss.n3312 759.029
R28095 vss.n3323 vss.n3312 759.029
R28096 vss.n3316 vss.n2599 759.029
R28097 vss.n4310 vss.n2606 759.029
R28098 vss.n4309 vss.n3339 759.029
R28099 vss.n4309 vss.n3338 759.029
R28100 vss.n4316 vss.n3338 759.029
R28101 vss.n4310 vss.n2605 759.029
R28102 vss.n4317 vss.n2605 759.029
R28103 vss.n4317 vss.n2604 759.029
R28104 vss.n4299 vss.n2604 759.029
R28105 vss.n4316 vss.n3337 759.029
R28106 vss.n4298 vss.n3337 759.029
R28107 vss.n4298 vss.n3336 759.029
R28108 vss.n4299 vss.n2598 759.029
R28109 vss.n4234 vss.n2609 759.029
R28110 vss.n4233 vss.n3343 759.029
R28111 vss.n4233 vss.n3342 759.029
R28112 vss.n4240 vss.n3342 759.029
R28113 vss.n4234 vss.n2608 759.029
R28114 vss.n4241 vss.n2608 759.029
R28115 vss.n4241 vss.n2607 759.029
R28116 vss.n4223 vss.n2607 759.029
R28117 vss.n4240 vss.n3341 759.029
R28118 vss.n4222 vss.n3341 759.029
R28119 vss.n4222 vss.n3340 759.029
R28120 vss.n4223 vss.n2597 759.029
R28121 vss.n3665 vss.n2612 759.029
R28122 vss.n3664 vss.n3347 759.029
R28123 vss.n3664 vss.n3346 759.029
R28124 vss.n3671 vss.n3346 759.029
R28125 vss.n3665 vss.n2611 759.029
R28126 vss.n3672 vss.n2611 759.029
R28127 vss.n3672 vss.n2610 759.029
R28128 vss.n3654 vss.n2610 759.029
R28129 vss.n3671 vss.n3345 759.029
R28130 vss.n3653 vss.n3345 759.029
R28131 vss.n3653 vss.n3344 759.029
R28132 vss.n3654 vss.n2596 759.029
R28133 vss.n3967 vss.n2615 759.029
R28134 vss.n3966 vss.n3351 759.029
R28135 vss.n3966 vss.n3350 759.029
R28136 vss.n3973 vss.n3350 759.029
R28137 vss.n3967 vss.n2614 759.029
R28138 vss.n3974 vss.n2614 759.029
R28139 vss.n3974 vss.n2613 759.029
R28140 vss.n3956 vss.n2613 759.029
R28141 vss.n3973 vss.n3349 759.029
R28142 vss.n3955 vss.n3349 759.029
R28143 vss.n3955 vss.n3348 759.029
R28144 vss.n3956 vss.n2595 759.029
R28145 vss.n3445 vss.n2618 759.029
R28146 vss.n3444 vss.n3355 759.029
R28147 vss.n3444 vss.n3354 759.029
R28148 vss.n3451 vss.n3354 759.029
R28149 vss.n3445 vss.n2617 759.029
R28150 vss.n3452 vss.n2617 759.029
R28151 vss.n3452 vss.n2616 759.029
R28152 vss.n3434 vss.n2616 759.029
R28153 vss.n3451 vss.n3353 759.029
R28154 vss.n3433 vss.n3353 759.029
R28155 vss.n3433 vss.n3352 759.029
R28156 vss.n3434 vss.n2594 759.029
R28157 vss.n5852 vss.n2621 759.029
R28158 vss.n5857 vss.n3360 759.029
R28159 vss.n3360 vss.n3358 759.029
R28160 vss.n3377 vss.n3358 759.029
R28161 vss.n5852 vss.n2620 759.029
R28162 vss.n3378 vss.n2620 759.029
R28163 vss.n3378 vss.n2619 759.029
R28164 vss.n3371 vss.n2619 759.029
R28165 vss.n3377 vss.n3357 759.029
R28166 vss.n3370 vss.n3357 759.029
R28167 vss.n3370 vss.n3356 759.029
R28168 vss.n3371 vss.n2593 759.029
R28169 vss.n9998 vss.n2625 759.029
R28170 vss.n5881 vss.n5865 759.029
R28171 vss.n5865 vss.n5863 759.029
R28172 vss.n5863 vss.n5862 759.029
R28173 vss.n2625 vss.n2623 759.029
R28174 vss.n5860 vss.n2623 759.029
R28175 vss.n5860 vss.n2622 759.029
R28176 vss.n5872 vss.n2622 759.029
R28177 vss.n5862 vss.n5859 759.029
R28178 vss.n5871 vss.n5859 759.029
R28179 vss.n5871 vss.n5858 759.029
R28180 vss.n5872 vss.n2592 759.029
R28181 vss.n2235 vss.n2234 759.029
R28182 vss.n2228 vss.n2210 759.029
R28183 vss.n2229 vss.n2228 759.029
R28184 vss.n2230 vss.n2229 759.029
R28185 vss.n2217 vss.n2216 759.029
R28186 vss.n2216 vss.n2207 759.029
R28187 vss.n2236 vss.n2207 759.029
R28188 vss.n2236 vss.n2235 759.029
R28189 vss.n2218 vss.n2217 759.029
R28190 vss.n2223 vss.n2222 759.029
R28191 vss.n2224 vss.n2223 759.029
R28192 vss.n2224 vss.n2210 759.029
R28193 vss.n12398 vss.n12397 759.029
R28194 vss.n12391 vss.n12373 759.029
R28195 vss.n12392 vss.n12391 759.029
R28196 vss.n12393 vss.n12392 759.029
R28197 vss.n12380 vss.n12379 759.029
R28198 vss.n12379 vss.n12370 759.029
R28199 vss.n12399 vss.n12370 759.029
R28200 vss.n12399 vss.n12398 759.029
R28201 vss.n12381 vss.n12380 759.029
R28202 vss.n12386 vss.n12385 759.029
R28203 vss.n12387 vss.n12386 759.029
R28204 vss.n12387 vss.n12373 759.029
R28205 vss.n12527 vss.n12526 759.029
R28206 vss.n12520 vss.n12502 759.029
R28207 vss.n12521 vss.n12520 759.029
R28208 vss.n12522 vss.n12521 759.029
R28209 vss.n12509 vss.n12508 759.029
R28210 vss.n12508 vss.n12499 759.029
R28211 vss.n12528 vss.n12499 759.029
R28212 vss.n12528 vss.n12527 759.029
R28213 vss.n12510 vss.n12509 759.029
R28214 vss.n12515 vss.n12514 759.029
R28215 vss.n12516 vss.n12515 759.029
R28216 vss.n12516 vss.n12502 759.029
R28217 vss.n10294 vss.n10293 759.029
R28218 vss.n10287 vss.n10269 759.029
R28219 vss.n10288 vss.n10287 759.029
R28220 vss.n10289 vss.n10288 759.029
R28221 vss.n10276 vss.n10275 759.029
R28222 vss.n10275 vss.n10266 759.029
R28223 vss.n10295 vss.n10266 759.029
R28224 vss.n10295 vss.n10294 759.029
R28225 vss.n10277 vss.n10276 759.029
R28226 vss.n10282 vss.n10281 759.029
R28227 vss.n10283 vss.n10282 759.029
R28228 vss.n10283 vss.n10269 759.029
R28229 vss.n10216 vss.n10215 759.029
R28230 vss.n10209 vss.n10191 759.029
R28231 vss.n10210 vss.n10209 759.029
R28232 vss.n10211 vss.n10210 759.029
R28233 vss.n10198 vss.n10197 759.029
R28234 vss.n10197 vss.n10188 759.029
R28235 vss.n10217 vss.n10188 759.029
R28236 vss.n10217 vss.n10216 759.029
R28237 vss.n10199 vss.n10198 759.029
R28238 vss.n10204 vss.n10203 759.029
R28239 vss.n10205 vss.n10204 759.029
R28240 vss.n10205 vss.n10191 759.029
R28241 vss.n2474 vss.n2473 759.029
R28242 vss.n2467 vss.n2449 759.029
R28243 vss.n2468 vss.n2467 759.029
R28244 vss.n2469 vss.n2468 759.029
R28245 vss.n2456 vss.n2455 759.029
R28246 vss.n2455 vss.n2446 759.029
R28247 vss.n2475 vss.n2446 759.029
R28248 vss.n2475 vss.n2474 759.029
R28249 vss.n2457 vss.n2456 759.029
R28250 vss.n2462 vss.n2461 759.029
R28251 vss.n2463 vss.n2462 759.029
R28252 vss.n2463 vss.n2449 759.029
R28253 vss.n2553 vss.n2552 759.029
R28254 vss.n2546 vss.n2528 759.029
R28255 vss.n2547 vss.n2546 759.029
R28256 vss.n2548 vss.n2547 759.029
R28257 vss.n2535 vss.n2534 759.029
R28258 vss.n2534 vss.n2525 759.029
R28259 vss.n2554 vss.n2525 759.029
R28260 vss.n2554 vss.n2553 759.029
R28261 vss.n2536 vss.n2535 759.029
R28262 vss.n2541 vss.n2540 759.029
R28263 vss.n2542 vss.n2541 759.029
R28264 vss.n2542 vss.n2528 759.029
R28265 vss.n7413 vss.n7403 759.029
R28266 vss.n7426 vss.n7416 759.029
R28267 vss.n7431 vss.n7426 759.029
R28268 vss.n7431 vss.n7430 759.029
R28269 vss.n7407 vss.n7405 759.029
R28270 vss.n7414 vss.n7405 759.029
R28271 vss.n7414 vss.n7404 759.029
R28272 vss.n7413 vss.n7404 759.029
R28273 vss.n8984 vss.n7407 759.029
R28274 vss.n7421 vss.n7419 759.029
R28275 vss.n7422 vss.n7421 759.029
R28276 vss.n7422 vss.n7416 759.029
R28277 vss.n7439 vss.n7399 759.029
R28278 vss.n7460 vss.n7440 759.029
R28279 vss.n7465 vss.n7460 759.029
R28280 vss.n7465 vss.n7464 759.029
R28281 vss.n7446 vss.n7401 759.029
R28282 vss.n7441 vss.n7401 759.029
R28283 vss.n7441 vss.n7400 759.029
R28284 vss.n7439 vss.n7400 759.029
R28285 vss.n7446 vss.n7402 759.029
R28286 vss.n7455 vss.n7445 759.029
R28287 vss.n7456 vss.n7455 759.029
R28288 vss.n7456 vss.n7440 759.029
R28289 vss.n7593 vss.n7395 759.029
R28290 vss.n7614 vss.n7594 759.029
R28291 vss.n7619 vss.n7614 759.029
R28292 vss.n7619 vss.n7618 759.029
R28293 vss.n7600 vss.n7397 759.029
R28294 vss.n7595 vss.n7397 759.029
R28295 vss.n7595 vss.n7396 759.029
R28296 vss.n7593 vss.n7396 759.029
R28297 vss.n7600 vss.n7398 759.029
R28298 vss.n7609 vss.n7599 759.029
R28299 vss.n7610 vss.n7609 759.029
R28300 vss.n7610 vss.n7594 759.029
R28301 vss.n7628 vss.n7391 759.029
R28302 vss.n7649 vss.n7629 759.029
R28303 vss.n7654 vss.n7649 759.029
R28304 vss.n7654 vss.n7653 759.029
R28305 vss.n7635 vss.n7393 759.029
R28306 vss.n7630 vss.n7393 759.029
R28307 vss.n7630 vss.n7392 759.029
R28308 vss.n7628 vss.n7392 759.029
R28309 vss.n7635 vss.n7394 759.029
R28310 vss.n7644 vss.n7634 759.029
R28311 vss.n7645 vss.n7644 759.029
R28312 vss.n7645 vss.n7629 759.029
R28313 vss.n7736 vss.n7387 759.029
R28314 vss.n7757 vss.n7737 759.029
R28315 vss.n7762 vss.n7757 759.029
R28316 vss.n7762 vss.n7761 759.029
R28317 vss.n7743 vss.n7389 759.029
R28318 vss.n7738 vss.n7389 759.029
R28319 vss.n7738 vss.n7388 759.029
R28320 vss.n7736 vss.n7388 759.029
R28321 vss.n7743 vss.n7390 759.029
R28322 vss.n7752 vss.n7742 759.029
R28323 vss.n7753 vss.n7752 759.029
R28324 vss.n7753 vss.n7737 759.029
R28325 vss.n7815 vss.n7383 759.029
R28326 vss.n7836 vss.n7816 759.029
R28327 vss.n7841 vss.n7836 759.029
R28328 vss.n7841 vss.n7840 759.029
R28329 vss.n7822 vss.n7385 759.029
R28330 vss.n7817 vss.n7385 759.029
R28331 vss.n7817 vss.n7384 759.029
R28332 vss.n7815 vss.n7384 759.029
R28333 vss.n7822 vss.n7386 759.029
R28334 vss.n7831 vss.n7821 759.029
R28335 vss.n7832 vss.n7831 759.029
R28336 vss.n7832 vss.n7816 759.029
R28337 vss.n7957 vss.n7379 759.029
R28338 vss.n7978 vss.n7958 759.029
R28339 vss.n7983 vss.n7978 759.029
R28340 vss.n7983 vss.n7982 759.029
R28341 vss.n7964 vss.n7381 759.029
R28342 vss.n7959 vss.n7381 759.029
R28343 vss.n7959 vss.n7380 759.029
R28344 vss.n7957 vss.n7380 759.029
R28345 vss.n7964 vss.n7382 759.029
R28346 vss.n7973 vss.n7963 759.029
R28347 vss.n7974 vss.n7973 759.029
R28348 vss.n7974 vss.n7958 759.029
R28349 vss.n7370 vss.n7348 759.029
R28350 vss.n7360 vss.n7359 759.029
R28351 vss.n7360 vss.n7349 759.029
R28352 vss.n7365 vss.n7349 759.029
R28353 vss.n7342 vss.n7340 759.029
R28354 vss.n7347 vss.n7340 759.029
R28355 vss.n7371 vss.n7347 759.029
R28356 vss.n7371 vss.n7370 759.029
R28357 vss.n7378 vss.n7342 759.029
R28358 vss.n7354 vss.n7353 759.029
R28359 vss.n7358 vss.n7353 759.029
R28360 vss.n7359 vss.n7358 759.029
R28361 vss.n14045 vss.n500 759.029
R28362 vss.n14050 vss.n510 759.029
R28363 vss.n14050 vss.n514 759.029
R28364 vss.n514 vss.n513 759.029
R28365 vss.n504 vss.n502 759.029
R28366 vss.n14036 vss.n502 759.029
R28367 vss.n14036 vss.n501 759.029
R28368 vss.n14045 vss.n501 759.029
R28369 vss.n14053 vss.n509 759.029
R28370 vss.n14053 vss.n14052 759.029
R28371 vss.n14052 vss.n510 759.029
R28372 vss.n14058 vss.n504 759.029
R28373 vss.n968 vss.n935 759.029
R28374 vss.n942 vss.n941 759.029
R28375 vss.n946 vss.n941 759.029
R28376 vss.n960 vss.n946 759.029
R28377 vss.n935 vss.n933 759.029
R28378 vss.n961 vss.n933 759.029
R28379 vss.n961 vss.n932 759.029
R28380 vss.n954 vss.n932 759.029
R28381 vss.n960 vss.n959 759.029
R28382 vss.n959 vss.n947 759.029
R28383 vss.n949 vss.n947 759.029
R28384 vss.n954 vss.n931 759.029
R28385 vss.n1499 vss.n971 759.029
R28386 vss.n1494 vss.n1492 759.029
R28387 vss.n1504 vss.n1492 759.029
R28388 vss.n1518 vss.n1504 759.029
R28389 vss.n1499 vss.n970 759.029
R28390 vss.n1519 vss.n970 759.029
R28391 vss.n1519 vss.n969 759.029
R28392 vss.n1512 vss.n969 759.029
R28393 vss.n1518 vss.n1517 759.029
R28394 vss.n1517 vss.n1505 759.029
R28395 vss.n1507 vss.n1505 759.029
R28396 vss.n1512 vss.n930 759.029
R28397 vss.n1582 vss.n974 759.029
R28398 vss.n1577 vss.n1575 759.029
R28399 vss.n1587 vss.n1575 759.029
R28400 vss.n1601 vss.n1587 759.029
R28401 vss.n1582 vss.n973 759.029
R28402 vss.n1602 vss.n973 759.029
R28403 vss.n1602 vss.n972 759.029
R28404 vss.n1595 vss.n972 759.029
R28405 vss.n1601 vss.n1600 759.029
R28406 vss.n1600 vss.n1588 759.029
R28407 vss.n1590 vss.n1588 759.029
R28408 vss.n1595 vss.n929 759.029
R28409 vss.n1419 vss.n977 759.029
R28410 vss.n1414 vss.n1412 759.029
R28411 vss.n1424 vss.n1412 759.029
R28412 vss.n1438 vss.n1424 759.029
R28413 vss.n1419 vss.n976 759.029
R28414 vss.n1439 vss.n976 759.029
R28415 vss.n1439 vss.n975 759.029
R28416 vss.n1432 vss.n975 759.029
R28417 vss.n1438 vss.n1437 759.029
R28418 vss.n1437 vss.n1425 759.029
R28419 vss.n1427 vss.n1425 759.029
R28420 vss.n1432 vss.n928 759.029
R28421 vss.n1287 vss.n980 759.029
R28422 vss.n1282 vss.n1280 759.029
R28423 vss.n1292 vss.n1280 759.029
R28424 vss.n1306 vss.n1292 759.029
R28425 vss.n1287 vss.n979 759.029
R28426 vss.n1307 vss.n979 759.029
R28427 vss.n1307 vss.n978 759.029
R28428 vss.n1300 vss.n978 759.029
R28429 vss.n1306 vss.n1305 759.029
R28430 vss.n1305 vss.n1293 759.029
R28431 vss.n1295 vss.n1293 759.029
R28432 vss.n1300 vss.n927 759.029
R28433 vss.n1026 vss.n983 759.029
R28434 vss.n1021 vss.n1019 759.029
R28435 vss.n1031 vss.n1019 759.029
R28436 vss.n1045 vss.n1031 759.029
R28437 vss.n1026 vss.n982 759.029
R28438 vss.n1046 vss.n982 759.029
R28439 vss.n1046 vss.n981 759.029
R28440 vss.n1039 vss.n981 759.029
R28441 vss.n1045 vss.n1044 759.029
R28442 vss.n1044 vss.n1032 759.029
R28443 vss.n1034 vss.n1032 759.029
R28444 vss.n1039 vss.n926 759.029
R28445 vss.n13208 vss.n987 759.029
R28446 vss.n994 vss.n993 759.029
R28447 vss.n998 vss.n993 759.029
R28448 vss.n1012 vss.n998 759.029
R28449 vss.n987 vss.n985 759.029
R28450 vss.n1013 vss.n985 759.029
R28451 vss.n1013 vss.n984 759.029
R28452 vss.n1006 vss.n984 759.029
R28453 vss.n1012 vss.n1011 759.029
R28454 vss.n1011 vss.n999 759.029
R28455 vss.n1001 vss.n999 759.029
R28456 vss.n1006 vss.n925 759.029
R28457 vss.n405 vss.n64 759.029
R28458 vss.n384 vss.n72 759.029
R28459 vss.n406 vss.n72 759.029
R28460 vss.n406 vss.n71 759.029
R28461 vss.n387 vss.n62 759.029
R28462 vss.n383 vss.n62 759.029
R28463 vss.n383 vss.n63 759.029
R28464 vss.n405 vss.n63 759.029
R28465 vss.n387 vss.n61 759.029
R28466 vss.n388 vss.n74 759.029
R28467 vss.n388 vss.n73 759.029
R28468 vss.n384 vss.n73 759.029
R28469 vss.n282 vss.n57 759.029
R28470 vss.n261 vss.n78 759.029
R28471 vss.n283 vss.n78 759.029
R28472 vss.n283 vss.n77 759.029
R28473 vss.n264 vss.n55 759.029
R28474 vss.n260 vss.n55 759.029
R28475 vss.n260 vss.n56 759.029
R28476 vss.n282 vss.n56 759.029
R28477 vss.n264 vss.n54 759.029
R28478 vss.n265 vss.n80 759.029
R28479 vss.n265 vss.n79 759.029
R28480 vss.n261 vss.n79 759.029
R28481 vss.n14439 vss.n53 759.029
R28482 vss.n14418 vss.n82 759.029
R28483 vss.n14440 vss.n82 759.029
R28484 vss.n14440 vss.n81 759.029
R28485 vss.n14421 vss.n51 759.029
R28486 vss.n14417 vss.n51 759.029
R28487 vss.n14417 vss.n52 759.029
R28488 vss.n14439 vss.n52 759.029
R28489 vss.n14421 vss.n50 759.029
R28490 vss.n14422 vss.n84 759.029
R28491 vss.n14422 vss.n83 759.029
R28492 vss.n14418 vss.n83 759.029
R28493 vss.n223 vss.n49 759.029
R28494 vss.n202 vss.n86 759.029
R28495 vss.n224 vss.n86 759.029
R28496 vss.n224 vss.n85 759.029
R28497 vss.n205 vss.n47 759.029
R28498 vss.n201 vss.n47 759.029
R28499 vss.n201 vss.n48 759.029
R28500 vss.n223 vss.n48 759.029
R28501 vss.n205 vss.n46 759.029
R28502 vss.n206 vss.n88 759.029
R28503 vss.n206 vss.n87 759.029
R28504 vss.n202 vss.n87 759.029
R28505 vss.n14634 vss.n45 759.029
R28506 vss.n14613 vss.n90 759.029
R28507 vss.n14635 vss.n90 759.029
R28508 vss.n14635 vss.n89 759.029
R28509 vss.n14616 vss.n43 759.029
R28510 vss.n14612 vss.n43 759.029
R28511 vss.n14612 vss.n44 759.029
R28512 vss.n14634 vss.n44 759.029
R28513 vss.n14616 vss.n42 759.029
R28514 vss.n14617 vss.n92 759.029
R28515 vss.n14617 vss.n91 759.029
R28516 vss.n14613 vss.n91 759.029
R28517 vss.n146 vss.n41 759.029
R28518 vss.n125 vss.n94 759.029
R28519 vss.n147 vss.n94 759.029
R28520 vss.n147 vss.n93 759.029
R28521 vss.n128 vss.n39 759.029
R28522 vss.n124 vss.n39 759.029
R28523 vss.n124 vss.n40 759.029
R28524 vss.n146 vss.n40 759.029
R28525 vss.n128 vss.n38 759.029
R28526 vss.n129 vss.n96 759.029
R28527 vss.n129 vss.n95 759.029
R28528 vss.n125 vss.n95 759.029
R28529 vss.n116 vss.n37 759.029
R28530 vss.n106 vss.n98 759.029
R28531 vss.n117 vss.n98 759.029
R28532 vss.n117 vss.n97 759.029
R28533 vss.n14766 vss.n35 759.029
R28534 vss.n105 vss.n35 759.029
R28535 vss.n105 vss.n36 759.029
R28536 vss.n116 vss.n36 759.029
R28537 vss.n14766 vss.n34 759.029
R28538 vss.n14771 vss.n101 759.029
R28539 vss.n101 vss.n99 759.029
R28540 vss.n106 vss.n99 759.029
R28541 vss.n14781 vss.n65 759.029
R28542 vss.n14773 vss.n70 759.029
R28543 vss.n14774 vss.n14773 759.029
R28544 vss.n14774 vss.n67 759.029
R28545 vss.n365 vss.n59 759.029
R28546 vss.n362 vss.n59 759.029
R28547 vss.n362 vss.n60 759.029
R28548 vss.n65 vss.n60 759.029
R28549 vss.n366 vss.n76 759.029
R28550 vss.n366 vss.n75 759.029
R28551 vss.n75 vss.n70 759.029
R28552 vss.n365 vss.n58 759.029
R28553 vss.n9858 vss.n9857 759.029
R28554 vss.n9866 vss.n9865 759.029
R28555 vss.n9865 vss.n2831 759.029
R28556 vss.n2832 vss.n2831 759.029
R28557 vss.n9855 vss.n9850 759.029
R28558 vss.n9856 vss.n9855 759.029
R28559 vss.n9859 vss.n9856 759.029
R28560 vss.n9859 vss.n9858 759.029
R28561 vss.n9850 vss.n2825 759.029
R28562 vss.n2830 vss.n2826 759.029
R28563 vss.n9867 vss.n2830 759.029
R28564 vss.n9867 vss.n9866 759.029
R28565 vss.n2866 vss.n2865 759.029
R28566 vss.n2859 vss.n2841 759.029
R28567 vss.n2860 vss.n2859 759.029
R28568 vss.n2861 vss.n2860 759.029
R28569 vss.n2848 vss.n2847 759.029
R28570 vss.n2847 vss.n2838 759.029
R28571 vss.n2867 vss.n2838 759.029
R28572 vss.n2867 vss.n2866 759.029
R28573 vss.n2849 vss.n2848 759.029
R28574 vss.n2854 vss.n2853 759.029
R28575 vss.n2855 vss.n2854 759.029
R28576 vss.n2855 vss.n2841 759.029
R28577 vss.n4997 vss.n4996 759.029
R28578 vss.n4990 vss.n4972 759.029
R28579 vss.n4991 vss.n4990 759.029
R28580 vss.n4992 vss.n4991 759.029
R28581 vss.n4979 vss.n4978 759.029
R28582 vss.n4978 vss.n4969 759.029
R28583 vss.n4998 vss.n4969 759.029
R28584 vss.n4998 vss.n4997 759.029
R28585 vss.n4980 vss.n4979 759.029
R28586 vss.n4985 vss.n4984 759.029
R28587 vss.n4986 vss.n4985 759.029
R28588 vss.n4986 vss.n4972 759.029
R28589 vss.n5074 vss.n5073 759.029
R28590 vss.n5067 vss.n5049 759.029
R28591 vss.n5068 vss.n5067 759.029
R28592 vss.n5069 vss.n5068 759.029
R28593 vss.n5056 vss.n5055 759.029
R28594 vss.n5055 vss.n5046 759.029
R28595 vss.n5075 vss.n5046 759.029
R28596 vss.n5075 vss.n5074 759.029
R28597 vss.n5057 vss.n5056 759.029
R28598 vss.n5062 vss.n5061 759.029
R28599 vss.n5063 vss.n5062 759.029
R28600 vss.n5063 vss.n5049 759.029
R28601 vss.n5199 vss.n5198 759.029
R28602 vss.n5192 vss.n5174 759.029
R28603 vss.n5193 vss.n5192 759.029
R28604 vss.n5194 vss.n5193 759.029
R28605 vss.n5181 vss.n5180 759.029
R28606 vss.n5180 vss.n5171 759.029
R28607 vss.n5200 vss.n5171 759.029
R28608 vss.n5200 vss.n5199 759.029
R28609 vss.n5182 vss.n5181 759.029
R28610 vss.n5187 vss.n5186 759.029
R28611 vss.n5188 vss.n5187 759.029
R28612 vss.n5188 vss.n5174 759.029
R28613 vss.n3100 vss.n3099 759.029
R28614 vss.n3093 vss.n3075 759.029
R28615 vss.n3094 vss.n3093 759.029
R28616 vss.n3095 vss.n3094 759.029
R28617 vss.n3082 vss.n3081 759.029
R28618 vss.n3081 vss.n3072 759.029
R28619 vss.n3101 vss.n3072 759.029
R28620 vss.n3101 vss.n3100 759.029
R28621 vss.n3083 vss.n3082 759.029
R28622 vss.n3088 vss.n3087 759.029
R28623 vss.n3089 vss.n3088 759.029
R28624 vss.n3089 vss.n3075 759.029
R28625 vss.n3180 vss.n3179 759.029
R28626 vss.n3173 vss.n3155 759.029
R28627 vss.n3174 vss.n3173 759.029
R28628 vss.n3175 vss.n3174 759.029
R28629 vss.n3162 vss.n3161 759.029
R28630 vss.n3161 vss.n3152 759.029
R28631 vss.n3181 vss.n3152 759.029
R28632 vss.n3181 vss.n3180 759.029
R28633 vss.n3163 vss.n3162 759.029
R28634 vss.n3168 vss.n3167 759.029
R28635 vss.n3169 vss.n3168 759.029
R28636 vss.n3169 vss.n3155 759.029
R28637 vss.n3257 vss.n3256 759.029
R28638 vss.n3250 vss.n3232 759.029
R28639 vss.n3251 vss.n3250 759.029
R28640 vss.n3252 vss.n3251 759.029
R28641 vss.n3239 vss.n3238 759.029
R28642 vss.n3238 vss.n3229 759.029
R28643 vss.n3258 vss.n3229 759.029
R28644 vss.n3258 vss.n3257 759.029
R28645 vss.n3240 vss.n3239 759.029
R28646 vss.n3245 vss.n3244 759.029
R28647 vss.n3246 vss.n3245 759.029
R28648 vss.n3246 vss.n3232 759.029
R28649 vss.n6229 vss.n6226 759.029
R28650 vss.n6235 vss.n6225 759.029
R28651 vss.n6240 vss.n6235 759.029
R28652 vss.n6241 vss.n6240 759.029
R28653 vss.n6252 vss.n6229 759.029
R28654 vss.n6252 vss.n6251 759.029
R28655 vss.n6251 vss.n6250 759.029
R28656 vss.n6250 vss.n6230 759.029
R28657 vss.n6242 vss.n6241 759.029
R28658 vss.n6243 vss.n6242 759.029
R28659 vss.n6244 vss.n6243 759.029
R28660 vss.n6231 vss.n6230 759.029
R28661 vss.n6267 vss.n6263 759.029
R28662 vss.n6273 vss.n6262 759.029
R28663 vss.n6278 vss.n6273 759.029
R28664 vss.n6279 vss.n6278 759.029
R28665 vss.n6290 vss.n6267 759.029
R28666 vss.n6290 vss.n6289 759.029
R28667 vss.n6289 vss.n6288 759.029
R28668 vss.n6288 vss.n6268 759.029
R28669 vss.n6280 vss.n6279 759.029
R28670 vss.n6281 vss.n6280 759.029
R28671 vss.n6282 vss.n6281 759.029
R28672 vss.n6269 vss.n6268 759.029
R28673 vss.n7109 vss.n7108 759.029
R28674 vss.n7102 vss.n7098 759.029
R28675 vss.n7122 vss.n7098 759.029
R28676 vss.n7122 vss.n7121 759.029
R28677 vss.n7110 vss.n7109 759.029
R28678 vss.n7111 vss.n7110 759.029
R28679 vss.n7112 vss.n7111 759.029
R28680 vss.n7113 vss.n7112 759.029
R28681 vss.n7121 vss.n7120 759.029
R28682 vss.n7120 vss.n7119 759.029
R28683 vss.n7119 vss.n7118 759.029
R28684 vss.n7114 vss.n7113 759.029
R28685 vss.n6611 vss.n6610 759.029
R28686 vss.n6604 vss.n6600 759.029
R28687 vss.n6624 vss.n6600 759.029
R28688 vss.n6624 vss.n6623 759.029
R28689 vss.n6612 vss.n6611 759.029
R28690 vss.n6613 vss.n6612 759.029
R28691 vss.n6614 vss.n6613 759.029
R28692 vss.n6615 vss.n6614 759.029
R28693 vss.n6623 vss.n6622 759.029
R28694 vss.n6622 vss.n6621 759.029
R28695 vss.n6621 vss.n6620 759.029
R28696 vss.n6616 vss.n6615 759.029
R28697 vss.n6920 vss.n6919 759.029
R28698 vss.n6913 vss.n6909 759.029
R28699 vss.n6933 vss.n6909 759.029
R28700 vss.n6933 vss.n6932 759.029
R28701 vss.n6921 vss.n6920 759.029
R28702 vss.n6922 vss.n6921 759.029
R28703 vss.n6923 vss.n6922 759.029
R28704 vss.n6924 vss.n6923 759.029
R28705 vss.n6932 vss.n6931 759.029
R28706 vss.n6931 vss.n6930 759.029
R28707 vss.n6930 vss.n6929 759.029
R28708 vss.n6925 vss.n6924 759.029
R28709 vss.n6384 vss.n6383 759.029
R28710 vss.n6377 vss.n6373 759.029
R28711 vss.n6397 vss.n6373 759.029
R28712 vss.n6397 vss.n6396 759.029
R28713 vss.n6385 vss.n6384 759.029
R28714 vss.n6386 vss.n6385 759.029
R28715 vss.n6387 vss.n6386 759.029
R28716 vss.n6388 vss.n6387 759.029
R28717 vss.n6396 vss.n6395 759.029
R28718 vss.n6395 vss.n6394 759.029
R28719 vss.n6394 vss.n6393 759.029
R28720 vss.n6389 vss.n6388 759.029
R28721 vss.n9258 vss.n6321 759.029
R28722 vss.n9264 vss.n6320 759.029
R28723 vss.n9269 vss.n9264 759.029
R28724 vss.n9270 vss.n9269 759.029
R28725 vss.n9281 vss.n9258 759.029
R28726 vss.n9281 vss.n9280 759.029
R28727 vss.n9280 vss.n9279 759.029
R28728 vss.n9279 vss.n9259 759.029
R28729 vss.n9271 vss.n9270 759.029
R28730 vss.n9272 vss.n9271 759.029
R28731 vss.n9273 vss.n9272 759.029
R28732 vss.n9260 vss.n9259 759.029
R28733 vss.n9306 vss.n9305 759.029
R28734 vss.n9308 vss.n9303 759.029
R28735 vss.n9309 vss.n9308 759.029
R28736 vss.n9309 vss.n6217 759.029
R28737 vss.n9305 vss.n9304 759.029
R28738 vss.n9304 vss.n6218 759.029
R28739 vss.n9289 vss.n6218 759.029
R28740 vss.n9290 vss.n9289 759.029
R28741 vss.n9291 vss.n6217 759.029
R28742 vss.n9291 vss.n9288 759.029
R28743 vss.n9295 vss.n9288 759.029
R28744 vss.n9294 vss.n9290 759.029
R28745 vss.n13047 vss.n2201 759.029
R28746 vss.n13034 vss.n2203 759.029
R28747 vss.n13052 vss.n2203 759.029
R28748 vss.n13052 vss.n13051 759.029
R28749 vss.n13042 vss.n13024 759.029
R28750 vss.n13043 vss.n13042 759.029
R28751 vss.n13044 vss.n13043 759.029
R28752 vss.n13044 vss.n2201 759.029
R28753 vss.n13033 vss.n13032 759.029
R28754 vss.n13035 vss.n13033 759.029
R28755 vss.n13035 vss.n13034 759.029
R28756 vss.n13028 vss.n13024 759.029
R28757 vss.n11343 vss.n11329 759.029
R28758 vss.n11050 vss.n10453 759.029
R28759 vss.n11349 vss.n10453 759.029
R28760 vss.n11349 vss.n10452 759.029
R28761 vss.n11337 vss.n11332 759.029
R28762 vss.n11338 vss.n11337 759.029
R28763 vss.n11339 vss.n11338 759.029
R28764 vss.n11339 vss.n11329 759.029
R28765 vss.n12670 vss.n10456 759.029
R28766 vss.n10456 vss.n10454 759.029
R28767 vss.n11050 vss.n10454 759.029
R28768 vss.n11333 vss.n11332 759.029
R28769 vss.n8174 vss.n8173 727.362
R28770 vss.t244 vss.n9604 704.146
R28771 vss.t244 vss.n9598 704.146
R28772 vss.t1139 vss.n9598 704.146
R28773 vss.t1139 vss.n9591 704.146
R28774 vss.t1140 vss.n9591 704.146
R28775 vss.t1140 vss.n9592 704.146
R28776 vss.t1016 vss.n9592 704.146
R28777 vss.t1016 vss.n495 704.146
R28778 vss.n9668 vss.t1121 704.146
R28779 vss.n5981 vss.t1121 704.146
R28780 vss.t735 vss.n5981 704.146
R28781 vss.t735 vss.n5982 704.146
R28782 vss.t736 vss.n5982 704.146
R28783 vss.t736 vss.n9656 704.146
R28784 vss.n9656 vss.t41 704.146
R28785 vss.n9649 vss.t41 704.146
R28786 vss.t1271 vss.n2784 704.146
R28787 vss.t1271 vss.n5949 704.146
R28788 vss.t563 vss.n5949 704.146
R28789 vss.t563 vss.n5942 704.146
R28790 vss.t564 vss.n5942 704.146
R28791 vss.t564 vss.n5943 704.146
R28792 vss.t1214 vss.n5943 704.146
R28793 vss.t1214 vss.n9673 704.146
R28794 vss.t1180 vss.n2160 704.146
R28795 vss.t1180 vss.n2570 704.146
R28796 vss.t1200 vss.n2570 704.146
R28797 vss.t1200 vss.n2563 704.146
R28798 vss.t1201 vss.n2563 704.146
R28799 vss.t1201 vss.n2564 704.146
R28800 vss.t1014 vss.n2564 704.146
R28801 vss.t1014 vss.n10001 704.146
R28802 vss.t1398 vss.n9704 704.146
R28803 vss.t1398 vss.n9697 704.146
R28804 vss.t1444 vss.n9697 704.146
R28805 vss.t1444 vss.n9690 704.146
R28806 vss.t1445 vss.n9690 704.146
R28807 vss.t1445 vss.n9691 704.146
R28808 vss.t39 vss.n9691 704.146
R28809 vss.t39 vss.n9720 704.146
R28810 vss.t734 vss.n14063 704.146
R28811 vss.t734 vss.n489 704.146
R28812 vss.t920 vss.n489 704.146
R28813 vss.t920 vss.n491 704.146
R28814 vss.n491 vss.t921 704.146
R28815 vss.n480 vss.t921 704.146
R28816 vss.t35 vss.n480 704.146
R28817 vss.n482 vss.t35 704.146
R28818 vss.n13112 vss.t776 704.146
R28819 vss.n2080 vss.t776 704.146
R28820 vss.t1181 vss.n2080 704.146
R28821 vss.t1181 vss.n2081 704.146
R28822 vss.t1182 vss.n2081 704.146
R28823 vss.t1182 vss.n13100 704.146
R28824 vss.n13100 vss.t37 704.146
R28825 vss.n13093 vss.t37 704.146
R28826 vss.t176 vss.n12060 691.532
R28827 vss.t176 vss.n11897 691.532
R28828 vss.t126 vss.n11897 691.532
R28829 vss.t126 vss.n11898 691.532
R28830 vss.n11898 vss.t128 691.532
R28831 vss.n12088 vss.t128 691.532
R28832 vss.n10670 vss.t444 691.532
R28833 vss.n10651 vss.t444 691.532
R28834 vss.n10651 vss.t869 691.532
R28835 vss.n10660 vss.t869 691.532
R28836 vss.n10660 vss.t871 691.532
R28837 vss.n12598 vss.t871 691.532
R28838 vss.t861 vss.n11495 691.532
R28839 vss.t861 vss.n11496 691.532
R28840 vss.n11496 vss.t376 691.532
R28841 vss.t376 vss.n10879 691.532
R28842 vss.n10879 vss.t378 691.532
R28843 vss.n11527 vss.t378 691.532
R28844 vss.t655 vss.n12725 691.532
R28845 vss.t655 vss.n10346 691.532
R28846 vss.t1216 vss.n10346 691.532
R28847 vss.t1216 vss.n10347 691.532
R28848 vss.n10347 vss.t1218 691.532
R28849 vss.n12757 vss.t1218 691.532
R28850 vss.t681 vss.n13336 691.532
R28851 vss.t681 vss.n13338 691.532
R28852 vss.n13338 vss.t679 691.532
R28853 vss.n13888 vss.t679 691.532
R28854 vss.n13888 vss.t820 691.532
R28855 vss.n13897 vss.t820 691.532
R28856 vss.t307 vss.n13416 691.532
R28857 vss.t307 vss.n13418 691.532
R28858 vss.n13418 vss.t308 691.532
R28859 vss.n13783 vss.t308 691.532
R28860 vss.n13783 vss.t795 691.532
R28861 vss.n13792 vss.t795 691.532
R28862 vss.t271 vss.n13496 691.532
R28863 vss.t271 vss.n13498 691.532
R28864 vss.n13498 vss.t269 691.532
R28865 vss.n13678 vss.t269 691.532
R28866 vss.n13678 vss.t826 691.532
R28867 vss.n13687 vss.t826 691.532
R28868 vss.t1272 vss.n457 691.532
R28869 vss.t1272 vss.n466 691.532
R28870 vss.t1273 vss.n466 691.532
R28871 vss.n13575 vss.t1273 691.532
R28872 vss.n13575 vss.t816 691.532
R28873 vss.n13582 vss.t816 691.532
R28874 vss.n14001 vss.t653 691.532
R28875 vss.n544 vss.t653 691.532
R28876 vss.t673 vss.n544 691.532
R28877 vss.t673 vss.n545 691.532
R28878 vss.t675 vss.n545 691.532
R28879 vss.t675 vss.n668 691.532
R28880 vss.t657 vss.n1728 691.532
R28881 vss.t657 vss.n1721 691.532
R28882 vss.t908 vss.n1721 691.532
R28883 vss.t908 vss.n1715 691.532
R28884 vss.t907 vss.n1715 691.532
R28885 vss.t907 vss.n1706 691.532
R28886 vss.t174 vss.n1832 691.532
R28887 vss.t174 vss.n1225 691.532
R28888 vss.t1455 vss.n1225 691.532
R28889 vss.t1455 vss.n1219 691.532
R28890 vss.t1457 vss.n1219 691.532
R28891 vss.t1457 vss.n1210 691.532
R28892 vss.n1953 vss.t824 691.532
R28893 vss.n1943 vss.t824 691.532
R28894 vss.t114 vss.n1943 691.532
R28895 vss.t114 vss.n697 691.532
R28896 vss.t116 vss.n697 691.532
R28897 vss.t116 vss.n698 691.532
R28898 vss.t811 vss.n7894 691.532
R28899 vss.t811 vss.n7885 691.532
R28900 vss.t809 vss.n7885 691.532
R28901 vss.t809 vss.n7886 691.532
R28902 vss.n7886 vss.t65 691.532
R28903 vss.n8303 vss.t65 691.532
R28904 vss.n8644 vss.t608 691.532
R28905 vss.n8384 vss.t608 691.532
R28906 vss.t606 vss.n8384 691.532
R28907 vss.t606 vss.n8385 691.532
R28908 vss.t865 vss.n8385 691.532
R28909 vss.t865 vss.n8631 691.532
R28910 vss.n8557 vss.t794 691.532
R28911 vss.n8482 vss.t794 691.532
R28912 vss.t792 vss.n8482 691.532
R28913 vss.t792 vss.n8483 691.532
R28914 vss.t178 vss.n8483 691.532
R28915 vss.t178 vss.n8544 691.532
R28916 vss.n9550 vss.t822 691.532
R28917 vss.n6084 vss.t822 691.532
R28918 vss.t903 vss.n6084 691.532
R28919 vss.t903 vss.n6085 691.532
R28920 vss.t905 vss.n6085 691.532
R28921 vss.t905 vss.n7256 691.532
R28922 vss.t446 vss.n6764 691.532
R28923 vss.t446 vss.n6741 691.532
R28924 vss.t246 vss.n6741 691.532
R28925 vss.t246 vss.n6735 691.532
R28926 vss.t245 vss.n6735 691.532
R28927 vss.t245 vss.n6726 691.532
R28928 vss.n6892 vss.t797 691.532
R28929 vss.n6856 vss.t797 691.532
R28930 vss.t140 vss.n6856 691.532
R28931 vss.t140 vss.n6857 691.532
R28932 vss.t139 vss.n6857 691.532
R28933 vss.t139 vss.n6880 691.532
R28934 vss.t859 vss.n9082 691.532
R28935 vss.t859 vss.n9059 691.532
R28936 vss.t460 vss.n9059 691.532
R28937 vss.t460 vss.n6552 691.532
R28938 vss.t459 vss.n6552 691.532
R28939 vss.t459 vss.n9141 691.532
R28940 vss.t777 vss.n2716 691.532
R28941 vss.t777 vss.n2717 691.532
R28942 vss.t778 vss.n2717 691.532
R28943 vss.t778 vss.n9917 691.532
R28944 vss.n9917 vss.t69 691.532
R28945 vss.n9910 vss.t69 691.532
R28946 vss.n5582 vss.t1232 691.532
R28947 vss.n4712 vss.t1232 691.532
R28948 vss.t1233 vss.n4712 691.532
R28949 vss.t1233 vss.n4713 691.532
R28950 vss.t67 vss.n4713 691.532
R28951 vss.t67 vss.n5569 691.532
R28952 vss.n5496 vss.t1539 691.532
R28953 vss.n4798 vss.t1539 691.532
R28954 vss.t1537 vss.n4798 691.532
R28955 vss.t1537 vss.n4799 691.532
R28956 vss.t818 vss.n4799 691.532
R28957 vss.t818 vss.n5483 691.532
R28958 vss.n5410 vss.t191 691.532
R28959 vss.n5335 vss.t191 691.532
R28960 vss.t192 vss.n5335 691.532
R28961 vss.t192 vss.n5336 691.532
R28962 vss.t180 vss.n5336 691.532
R28963 vss.t180 vss.n5397 691.532
R28964 vss.t442 vss.n4536 691.532
R28965 vss.t442 vss.n4437 691.532
R28966 vss.t456 vss.n4437 691.532
R28967 vss.t456 vss.n4431 691.532
R28968 vss.t458 vss.n4431 691.532
R28969 vss.t458 vss.n4421 691.532
R28970 vss.n4183 vss.t867 691.532
R28971 vss.n3791 vss.t867 691.532
R28972 vss.t373 vss.n3791 691.532
R28973 vss.t373 vss.n3792 691.532
R28974 vss.t375 vss.n3792 691.532
R28975 vss.t375 vss.n3811 691.532
R28976 vss.n3935 vss.t448 691.532
R28977 vss.n3899 vss.t448 691.532
R28978 vss.t117 vss.n3899 691.532
R28979 vss.t117 vss.n3900 691.532
R28980 vss.t119 vss.n3900 691.532
R28981 vss.t119 vss.n3923 691.532
R28982 vss.t63 vss.n5676 691.532
R28983 vss.t63 vss.n5653 691.532
R28984 vss.t1513 vss.n5653 691.532
R28985 vss.t1513 vss.n3608 691.532
R28986 vss.t1515 vss.n3608 691.532
R28987 vss.t1515 vss.n5735 691.532
R28988 vss.t1058 vss.n8116 691.532
R28989 vss.t1058 vss.n8107 691.532
R28990 vss.t1059 vss.n8107 691.532
R28991 vss.t1059 vss.n8108 691.532
R28992 vss.n8108 vss.t863 691.532
R28993 vss.n8173 vss.t863 691.532
R28994 vss.t342 vss.n11806 691.532
R28995 vss.t342 vss.n11815 691.532
R28996 vss.t340 vss.n11815 691.532
R28997 vss.n11825 vss.t340 691.532
R28998 vss.t799 vss.n11825 691.532
R28999 vss.n12123 vss.t799 691.532
R29000 vss.t145 vss.n11719 691.532
R29001 vss.t145 vss.n11727 691.532
R29002 vss.t143 vss.n11727 691.532
R29003 vss.n12219 vss.t143 691.532
R29004 vss.n12219 vss.t71 691.532
R29005 vss.n12226 vss.t71 691.532
R29006 vss.t284 vss.n10315 691.532
R29007 vss.t284 vss.n10317 691.532
R29008 vss.n10317 vss.t282 691.532
R29009 vss.n10308 vss.t282 691.532
R29010 vss.t801 vss.n10308 691.532
R29011 vss.n11661 vss.t801 691.532
R29012 vss.t1520 vss.n10029 691.532
R29013 vss.t1520 vss.n10022 691.532
R29014 vss.t1518 vss.n10022 691.532
R29015 vss.t1518 vss.n10023 691.532
R29016 vss.t857 vss.n10023 691.532
R29017 vss.t857 vss.n12943 691.532
R29018 vss.n8986 vss.n498 676.971
R29019 vss.t1374 vss.n10410 669.716
R29020 vss.t1374 vss.n12633 669.716
R29021 vss.t121 vss.n12633 669.716
R29022 vss.t121 vss.n12626 669.716
R29023 vss.t123 vss.n12626 669.716
R29024 vss.t123 vss.n12627 669.716
R29025 vss.t971 vss.n12627 669.716
R29026 vss.t971 vss.n2049 669.716
R29027 vss.t574 vss.n12673 669.716
R29028 vss.t574 vss.n10387 669.716
R29029 vss.t1095 vss.n10387 669.716
R29030 vss.t1095 vss.n10379 669.716
R29031 vss.t1094 vss.n10379 669.716
R29032 vss.t1094 vss.n12692 669.716
R29033 vss.n12692 vss.t1063 669.716
R29034 vss.t1063 vss.n2068 669.716
R29035 vss.t207 vss.n10411 669.716
R29036 vss.t207 vss.n11418 669.716
R29037 vss.t102 vss.n11418 669.716
R29038 vss.t102 vss.n11410 669.716
R29039 vss.t101 vss.n11410 669.716
R29040 vss.t101 vss.n11442 669.716
R29041 vss.n11442 vss.t1048 669.716
R29042 vss.t1048 vss.n2065 669.716
R29043 vss.t19 vss.n10412 669.716
R29044 vss.t19 vss.n11371 669.716
R29045 vss.t420 vss.n11371 669.716
R29046 vss.t420 vss.n11363 669.716
R29047 vss.t422 vss.n11363 669.716
R29048 vss.t422 vss.n11395 669.716
R29049 vss.n11395 vss.t1463 669.716
R29050 vss.t1463 vss.n2067 669.716
R29051 vss.t1368 vss.n10413 669.716
R29052 vss.t1368 vss.n10946 669.716
R29053 vss.t813 vss.n10946 669.716
R29054 vss.t813 vss.n10938 669.716
R29055 vss.t815 vss.n10938 669.716
R29056 vss.t815 vss.n10970 669.716
R29057 vss.n10970 vss.t1311 669.716
R29058 vss.t1311 vss.n2062 669.716
R29059 vss.t21 vss.n10414 669.716
R29060 vss.t21 vss.n10783 669.716
R29061 vss.t168 vss.n10783 669.716
R29062 vss.t168 vss.n10775 669.716
R29063 vss.t170 vss.n10775 669.716
R29064 vss.t170 vss.n10807 669.716
R29065 vss.n10807 vss.t276 669.716
R29066 vss.t276 vss.n2059 669.716
R29067 vss.t576 vss.n10415 669.716
R29068 vss.t576 vss.n10739 669.716
R29069 vss.t319 vss.n10739 669.716
R29070 vss.t319 vss.n10731 669.716
R29071 vss.t321 vss.n10731 669.716
R29072 vss.t321 vss.n10763 669.716
R29073 vss.n10763 vss.t81 669.716
R29074 vss.t81 vss.n2061 669.716
R29075 vss.t1364 vss.n10416 669.716
R29076 vss.t1364 vss.n11565 669.716
R29077 vss.t663 vss.n11565 669.716
R29078 vss.t663 vss.n11557 669.716
R29079 vss.t665 vss.n11557 669.716
R29080 vss.t665 vss.n11589 669.716
R29081 vss.n11589 vss.t120 669.716
R29082 vss.t120 vss.n2056 669.716
R29083 vss.t201 vss.n10417 669.716
R29084 vss.t201 vss.n10562 669.716
R29085 vss.t1143 vss.n10562 669.716
R29086 vss.t1143 vss.n10554 669.716
R29087 vss.t1142 vss.n10554 669.716
R29088 vss.t1142 vss.n10586 669.716
R29089 vss.n10586 vss.t1145 669.716
R29090 vss.t1145 vss.n2053 669.716
R29091 vss.t11 vss.n10418 669.716
R29092 vss.t11 vss.n10518 669.716
R29093 vss.t1388 vss.n10518 669.716
R29094 vss.t1388 vss.n10510 669.716
R29095 vss.t1390 vss.n10510 669.716
R29096 vss.t1390 vss.n10542 669.716
R29097 vss.n10542 vss.t104 669.716
R29098 vss.t104 vss.n2055 669.716
R29099 vss.t1481 vss.n10419 669.716
R29100 vss.t1481 vss.n11939 669.716
R29101 vss.t1068 vss.n11939 669.716
R29102 vss.t1068 vss.n11931 669.716
R29103 vss.t1070 vss.n11931 669.716
R29104 vss.t1070 vss.n11963 669.716
R29105 vss.n11963 vss.t113 669.716
R29106 vss.t113 vss.n2050 669.716
R29107 vss.t1471 vss.n12008 669.716
R29108 vss.t1471 vss.n12009 669.716
R29109 vss.n12009 vss.t700 669.716
R29110 vss.t700 vss.n11987 669.716
R29111 vss.n11987 vss.t702 669.716
R29112 vss.n12043 vss.t702 669.716
R29113 vss.n12006 vss.t237 669.716
R29114 vss.t237 vss.n10596 669.716
R29115 vss.t239 vss.n10596 669.716
R29116 vss.t239 vss.n10597 669.716
R29117 vss.t1161 vss.n10597 669.716
R29118 vss.n12600 vss.t1161 669.716
R29119 vss.n10857 vss.t1393 669.716
R29120 vss.n10835 vss.t1393 669.716
R29121 vss.t683 vss.n10835 669.716
R29122 vss.t683 vss.n10836 669.716
R29123 vss.n10836 vss.t682 669.716
R29124 vss.n11614 vss.t682 669.716
R29125 vss.t401 vss.n10824 669.716
R29126 vss.t401 vss.n10817 669.716
R29127 vss.t400 vss.n10817 669.716
R29128 vss.t400 vss.n10818 669.716
R29129 vss.t403 vss.n10818 669.716
R29130 vss.n11529 vss.t403 669.716
R29131 vss.t593 vss.n10928 669.716
R29132 vss.t593 vss.n10929 669.716
R29133 vss.n10929 vss.t1099 669.716
R29134 vss.t1099 vss.n10905 669.716
R29135 vss.n10905 vss.t1098 669.716
R29136 vss.n11478 vss.t1098 669.716
R29137 vss.n10926 vss.t976 669.716
R29138 vss.t976 vss.n10910 669.716
R29139 vss.n10910 vss.t978 669.716
R29140 vss.n12746 vss.t978 669.716
R29141 vss.n12746 vss.t317 669.716
R29142 vss.n12755 vss.t317 669.716
R29143 vss.n2303 vss.t1241 669.716
R29144 vss.n2269 vss.t1241 669.716
R29145 vss.t187 vss.n2269 669.716
R29146 vss.t187 vss.n2270 669.716
R29147 vss.t185 vss.n2270 669.716
R29148 vss.t185 vss.n2291 669.716
R29149 vss.n2291 vss.t1511 669.716
R29150 vss.t1511 vss.n2143 669.716
R29151 vss.t926 vss.n12994 669.716
R29152 vss.t926 vss.n2253 669.716
R29153 vss.t644 vss.n2253 669.716
R29154 vss.t644 vss.n2246 669.716
R29155 vss.t642 vss.n2246 669.716
R29156 vss.t642 vss.n2247 669.716
R29157 vss.t500 vss.n2247 669.716
R29158 vss.t500 vss.n2144 669.716
R29159 vss.n13872 vss.t1454 669.716
R29160 vss.t1454 vss.n13345 669.716
R29161 vss.t806 vss.n13345 669.716
R29162 vss.t806 vss.n13352 669.716
R29163 vss.t807 vss.n13352 669.716
R29164 vss.n13364 vss.t807 669.716
R29165 vss.t1415 vss.n13377 669.716
R29166 vss.t1415 vss.n13379 669.716
R29167 vss.n13379 vss.t1413 669.716
R29168 vss.n13834 vss.t1413 669.716
R29169 vss.n13834 vss.t111 669.716
R29170 vss.n13843 vss.t111 669.716
R29171 vss.n13767 vss.t1470 669.716
R29172 vss.t1470 vss.n13425 669.716
R29173 vss.t1416 vss.n13425 669.716
R29174 vss.t1416 vss.n13432 669.716
R29175 vss.t1417 vss.n13432 669.716
R29176 vss.n13444 vss.t1417 669.716
R29177 vss.t1432 vss.n13457 669.716
R29178 vss.t1432 vss.n13459 669.716
R29179 vss.n13459 vss.t1433 669.716
R29180 vss.n13729 vss.t1433 669.716
R29181 vss.n13729 vss.t1391 669.716
R29182 vss.n13738 vss.t1391 669.716
R29183 vss.n13662 vss.t261 669.716
R29184 vss.t261 vss.n13505 669.716
R29185 vss.t630 vss.n13505 669.716
R29186 vss.t630 vss.n13512 669.716
R29187 vss.t631 vss.n13512 669.716
R29188 vss.n13524 vss.t631 669.716
R29189 vss.t1383 vss.n13537 669.716
R29190 vss.t1383 vss.n13539 669.716
R29191 vss.n13539 vss.t1384 669.716
R29192 vss.n13624 vss.t1384 669.716
R29193 vss.n13624 vss.t107 669.716
R29194 vss.n13633 vss.t107 669.716
R29195 vss.t1192 vss.n14732 669.716
R29196 vss.t1192 vss.n167 669.716
R29197 vss.t1111 vss.n167 669.716
R29198 vss.t1111 vss.n160 669.716
R29199 vss.t1112 vss.n160 669.716
R29200 vss.t1112 vss.n161 669.716
R29201 vss.t613 vss.n161 669.716
R29202 vss.t613 vss.n19 669.716
R29203 vss.n14683 vss.t430 669.716
R29204 vss.n14649 vss.t430 669.716
R29205 vss.t1052 vss.n14649 669.716
R29206 vss.t1052 vss.n14650 669.716
R29207 vss.t1050 vss.n14650 669.716
R29208 vss.t1050 vss.n14671 669.716
R29209 vss.n14671 vss.t1497 669.716
R29210 vss.t1497 vss.n20 669.716
R29211 vss.t1168 vss.n14537 669.716
R29212 vss.t1168 vss.n244 669.716
R29213 vss.t364 vss.n244 669.716
R29214 vss.t364 vss.n237 669.716
R29215 vss.t362 vss.n237 669.716
R29216 vss.t362 vss.n238 669.716
R29217 vss.t1324 vss.n238 669.716
R29218 vss.t1324 vss.n21 669.716
R29219 vss.n14488 vss.t1285 669.716
R29220 vss.n14454 vss.t1285 669.716
R29221 vss.t833 vss.n14454 669.716
R29222 vss.t833 vss.n14455 669.716
R29223 vss.t834 vss.n14455 669.716
R29224 vss.t834 vss.n14476 669.716
R29225 vss.n14476 vss.t381 669.716
R29226 vss.t381 vss.n22 669.716
R29227 vss.t1049 vss.n14342 669.716
R29228 vss.t1049 vss.n303 669.716
R29229 vss.t1101 vss.n303 669.716
R29230 vss.t1101 vss.n296 669.716
R29231 vss.t1102 vss.n296 669.716
R29232 vss.t1102 vss.n297 669.716
R29233 vss.t1350 vss.n297 669.716
R29234 vss.t1350 vss.n23 669.716
R29235 vss.n14293 vss.t300 669.716
R29236 vss.n14259 vss.t300 669.716
R29237 vss.t158 vss.n14259 669.716
R29238 vss.t158 vss.n14260 669.716
R29239 vss.t156 vss.n14260 669.716
R29240 vss.t156 vss.n14281 669.716
R29241 vss.n14281 vss.t502 669.716
R29242 vss.t502 vss.n24 669.716
R29243 vss.t429 vss.n14223 669.716
R29244 vss.t429 vss.n426 669.716
R29245 vss.t1188 vss.n426 669.716
R29246 vss.t1188 vss.n419 669.716
R29247 vss.t1189 vss.n419 669.716
R29248 vss.t1189 vss.n420 669.716
R29249 vss.t1332 vss.n420 669.716
R29250 vss.t1332 vss.n25 669.716
R29251 vss.n14220 vss.t1524 669.716
R29252 vss.n14186 vss.t1524 669.716
R29253 vss.t1521 vss.n14186 669.716
R29254 vss.t1521 vss.n14187 669.716
R29255 vss.t1522 vss.n14187 669.716
R29256 vss.t1522 vss.n14208 669.716
R29257 vss.n14208 vss.t1316 669.716
R29258 vss.t1316 vss.n27 669.716
R29259 vss.t88 vss.n335 669.716
R29260 vss.t88 vss.n329 669.716
R29261 vss.t1403 vss.n329 669.716
R29262 vss.t1403 vss.n322 669.716
R29263 vss.t1404 vss.n322 669.716
R29264 vss.t1404 vss.n323 669.716
R29265 vss.t1352 vss.n323 669.716
R29266 vss.t1352 vss.n28 669.716
R29267 vss.n14339 vss.t368 669.716
R29268 vss.n14305 vss.t368 669.716
R29269 vss.t753 vss.n14305 669.716
R29270 vss.t753 vss.n14306 669.716
R29271 vss.t754 vss.n14306 669.716
R29272 vss.t754 vss.n14327 669.716
R29273 vss.n14327 vss.t1477 669.716
R29274 vss.t1477 vss.n29 669.716
R29275 vss.t1312 vss.n14388 669.716
R29276 vss.t1312 vss.n14382 669.716
R29277 vss.t1207 vss.n14382 669.716
R29278 vss.t1207 vss.n14375 669.716
R29279 vss.t1208 vss.n14375 669.716
R29280 vss.t1208 vss.n14376 669.716
R29281 vss.t466 vss.n14376 669.716
R29282 vss.t466 vss.n30 669.716
R29283 vss.n14534 vss.t1053 669.716
R29284 vss.n14500 vss.t1053 669.716
R29285 vss.t265 vss.n14500 669.716
R29286 vss.t265 vss.n14501 669.716
R29287 vss.t266 vss.n14501 669.716
R29288 vss.t266 vss.n14522 669.716
R29289 vss.n14522 vss.t1077 669.716
R29290 vss.t1077 vss.n31 669.716
R29291 vss.t984 vss.n14583 669.716
R29292 vss.t984 vss.n14577 669.716
R29293 vss.t73 vss.n14577 669.716
R29294 vss.t73 vss.n14570 669.716
R29295 vss.t74 vss.n14570 669.716
R29296 vss.t74 vss.n14571 669.716
R29297 vss.t1336 vss.n14571 669.716
R29298 vss.t1336 vss.n32 669.716
R29299 vss.n14729 vss.t562 669.716
R29300 vss.n14695 vss.t562 669.716
R29301 vss.t345 vss.n14695 669.716
R29302 vss.t345 vss.n14696 669.716
R29303 vss.t346 vss.n14696 669.716
R29304 vss.t346 vss.n14717 669.716
R29305 vss.n14717 vss.t474 669.716
R29306 vss.t474 vss.n33 669.716
R29307 vss.n189 vss.t853 669.716
R29308 vss.n182 vss.t853 669.716
R29309 vss.n182 vss.t1108 669.716
R29310 vss.t1108 vss.n6 669.716
R29311 vss.t1109 vss.n6 669.716
R29312 vss.t1109 vss.n7 669.716
R29313 vss.t1081 vss.n7 669.716
R29314 vss.t1081 vss.n14784 669.716
R29315 vss.t301 vss.n569 669.716
R29316 vss.t301 vss.n561 669.716
R29317 vss.t303 vss.n561 669.716
R29318 vss.t303 vss.n13986 669.716
R29319 vss.n13986 vss.t553 669.716
R29320 vss.n666 vss.t553 669.716
R29321 vss.n13966 vss.t109 669.716
R29322 vss.n583 vss.t109 669.716
R29323 vss.t767 vss.n583 669.716
R29324 vss.t767 vss.n584 669.716
R29325 vss.t769 vss.n584 669.716
R29326 vss.t769 vss.n762 669.716
R29327 vss.t289 vss.n1756 669.716
R29328 vss.t289 vss.n1703 669.716
R29329 vss.t291 vss.n1703 669.716
R29330 vss.t291 vss.n1798 669.716
R29331 vss.n1798 vss.t982 669.716
R29332 vss.n1750 vss.t982 669.716
R29333 vss.n1778 vss.t1159 669.716
R29334 vss.n1768 vss.t1159 669.716
R29335 vss.t417 vss.n1768 669.716
R29336 vss.t417 vss.n1272 669.716
R29337 vss.t419 vss.n1272 669.716
R29338 vss.t419 vss.n1263 669.716
R29339 vss.t1276 vss.n1860 669.716
R29340 vss.t1276 vss.n1207 669.716
R29341 vss.t1278 vss.n1207 669.716
R29342 vss.t1278 vss.n1902 669.716
R29343 vss.n1902 vss.t669 669.716
R29344 vss.n1854 vss.t669 669.716
R29345 vss.n1882 vss.t599 669.716
R29346 vss.n1872 vss.t599 669.716
R29347 vss.t150 vss.n1872 669.716
R29348 vss.t150 vss.n1154 669.716
R29349 vss.t152 vss.n1154 669.716
R29350 vss.t152 vss.n1145 669.716
R29351 vss.t578 vss.n813 669.716
R29352 vss.t578 vss.n1107 669.716
R29353 vss.t323 vss.n1107 669.716
R29354 vss.t323 vss.n1100 669.716
R29355 vss.t325 vss.n1100 669.716
R29356 vss.t325 vss.n1101 669.716
R29357 vss.t1299 vss.n1101 669.716
R29358 vss.t1299 vss.n730 669.716
R29359 vss.t13 vss.n814 669.716
R29360 vss.t13 vss.n1171 669.716
R29361 vss.t542 vss.n1171 669.716
R29362 vss.t542 vss.n1164 669.716
R29363 vss.t544 vss.n1164 669.716
R29364 vss.t544 vss.n1165 669.716
R29365 vss.t1146 vss.n1165 669.716
R29366 vss.t1146 vss.n733 669.716
R29367 vss.t615 vss.n815 669.716
R29368 vss.t615 vss.n1370 669.716
R29369 vss.t1407 vss.n1370 669.716
R29370 vss.t1407 vss.n1363 669.716
R29371 vss.t1406 vss.n1363 669.716
R29372 vss.t1406 vss.n1364 669.716
R29373 vss.t549 vss.n1364 669.716
R29374 vss.t549 vss.n736 669.716
R29375 vss.t1360 vss.n816 669.716
R29376 vss.t1360 vss.n1665 669.716
R29377 vss.t1531 vss.n1665 669.716
R29378 vss.t1531 vss.n1658 669.716
R29379 vss.t1533 vss.n1658 669.716
R29380 vss.t1533 vss.n1659 669.716
R29381 vss.t1270 vss.n1659 669.716
R29382 vss.t1270 vss.n739 669.716
R29383 vss.t506 vss.n13211 669.716
R29384 vss.t506 vss.n806 669.716
R29385 vss.t1174 vss.n806 669.716
R29386 vss.t1174 vss.n799 669.716
R29387 vss.t1176 vss.n799 669.716
R29388 vss.t1176 vss.n800 669.716
R29389 vss.t1177 vss.n800 669.716
R29390 vss.t1177 vss.n742 669.716
R29391 vss.n833 vss.t17 669.716
R29392 vss.n823 vss.t17 669.716
R29393 vss.t358 vss.n823 669.716
R29394 vss.t358 vss.n600 669.716
R29395 vss.t360 vss.n600 669.716
R29396 vss.t360 vss.n601 669.716
R29397 vss.t222 vss.n601 669.716
R29398 vss.n13943 vss.t222 669.716
R29399 vss.n874 vss.t395 669.716
R29400 vss.n849 vss.t395 669.716
R29401 vss.n849 vss.t762 669.716
R29402 vss.n842 vss.t762 669.716
R29403 vss.t761 vss.n842 669.716
R29404 vss.n846 vss.t761 669.716
R29405 vss.n846 vss.t552 669.716
R29406 vss.t552 vss.n613 669.716
R29407 vss.n918 vss.t504 669.716
R29408 vss.n893 vss.t504 669.716
R29409 vss.n893 vss.t935 669.716
R29410 vss.n882 vss.t935 669.716
R29411 vss.t937 vss.n882 669.716
R29412 vss.n886 vss.t937 669.716
R29413 vss.n886 vss.t344 669.716
R29414 vss.t344 vss.n612 669.716
R29415 vss.t397 vss.n919 669.716
R29416 vss.t397 vss.n1535 669.716
R29417 vss.t1429 vss.n1535 669.716
R29418 vss.t1429 vss.n1528 669.716
R29419 vss.t1431 vss.n1528 669.716
R29420 vss.t1431 vss.n1529 669.716
R29421 vss.t983 vss.n1529 669.716
R29422 vss.n1555 vss.t983 669.716
R29423 vss.t621 vss.n920 669.716
R29424 vss.t621 vss.n1618 669.716
R29425 vss.t583 vss.n1618 669.716
R29426 vss.t583 vss.n1611 669.716
R29427 vss.t582 vss.n1611 669.716
R29428 vss.t582 vss.n1612 669.716
R29429 vss.t166 vss.n1612 669.716
R29430 vss.t166 vss.n741 669.716
R29431 vss.t498 vss.n921 669.716
R29432 vss.t498 vss.n1455 669.716
R29433 vss.t171 vss.n1455 669.716
R29434 vss.t171 vss.n1448 669.716
R29435 vss.t173 vss.n1448 669.716
R29436 vss.t173 vss.n1449 669.716
R29437 vss.t1266 vss.n1449 669.716
R29438 vss.t1266 vss.n738 669.716
R29439 vss.t1083 vss.n922 669.716
R29440 vss.t1083 vss.n1323 669.716
R29441 vss.t764 vss.n1323 669.716
R29442 vss.t764 vss.n1316 669.716
R29443 vss.t766 vss.n1316 669.716
R29444 vss.t766 vss.n1317 669.716
R29445 vss.t541 vss.n1317 669.716
R29446 vss.t541 vss.n735 669.716
R29447 vss.t1372 vss.n923 669.716
R29448 vss.t1372 vss.n1062 669.716
R29449 vss.t923 vss.n1062 669.716
R29450 vss.t923 vss.n1055 669.716
R29451 vss.t925 vss.n1055 669.716
R29452 vss.t925 vss.n1056 669.716
R29453 vss.t1007 vss.n1056 669.716
R29454 vss.t1007 vss.n732 669.716
R29455 vss.t1320 vss.n924 669.716
R29456 vss.t1320 vss.n1997 669.716
R29457 vss.t521 vss.n1997 669.716
R29458 vss.t521 vss.n1990 669.716
R29459 vss.t523 vss.n1990 669.716
R29460 vss.t523 vss.n1991 669.716
R29461 vss.t1210 vss.n1991 669.716
R29462 vss.t1210 vss.n729 669.716
R29463 vss.t719 vss.n7275 669.716
R29464 vss.t719 vss.n7276 669.716
R29465 vss.t720 vss.n7276 669.716
R29466 vss.t720 vss.n9025 669.716
R29467 vss.n9025 vss.t585 669.716
R29468 vss.n9018 vss.t585 669.716
R29469 vss.n8282 vss.t703 669.716
R29470 vss.n8263 vss.t703 669.716
R29471 vss.t772 vss.n8263 669.716
R29472 vss.t772 vss.n8264 669.716
R29473 vss.n8264 vss.t773 669.716
R29474 vss.n9016 vss.t773 669.716
R29475 vss.n8687 vss.t1227 669.716
R29476 vss.n8334 vss.t1227 669.716
R29477 vss.t1228 vss.n8334 669.716
R29478 vss.t1228 vss.n8335 669.716
R29479 vss.t1153 vss.n8335 669.716
R29480 vss.t1153 vss.n8674 669.716
R29481 vss.t1088 vss.n8646 669.716
R29482 vss.t1088 vss.n8356 669.716
R29483 vss.t666 vss.n8356 669.716
R29484 vss.t666 vss.n8357 669.716
R29485 vss.n8357 vss.t667 669.716
R29486 vss.n8672 vss.t667 669.716
R29487 vss.n8600 vss.t100 669.716
R29488 vss.n8432 vss.t100 669.716
R29489 vss.t98 vss.n8432 669.716
R29490 vss.t98 vss.n8433 669.716
R29491 vss.t595 vss.n8433 669.716
R29492 vss.t595 vss.n8587 669.716
R29493 vss.t686 vss.n8559 669.716
R29494 vss.t686 vss.n8454 669.716
R29495 vss.t943 vss.n8454 669.716
R29496 vss.t943 vss.n8455 669.716
R29497 vss.n8455 vss.t944 669.716
R29498 vss.n8585 vss.t944 669.716
R29499 vss.t258 vss.n6109 669.716
R29500 vss.t258 vss.n6101 669.716
R29501 vss.t260 vss.n6101 669.716
R29502 vss.t260 vss.n9535 669.716
R29503 vss.n9535 vss.t892 669.716
R29504 vss.n7254 vss.t892 669.716
R29505 vss.n9515 vss.t105 669.716
R29506 vss.n6123 vss.t105 669.716
R29507 vss.t453 vss.n6123 669.716
R29508 vss.t453 vss.n6124 669.716
R29509 vss.t452 vss.n6124 669.716
R29510 vss.t452 vss.n7237 669.716
R29511 vss.t327 vss.n6792 669.716
R29512 vss.t327 vss.n6723 669.716
R29513 vss.t326 vss.n6723 669.716
R29514 vss.t326 vss.n7080 669.716
R29515 vss.n7080 vss.t646 669.716
R29516 vss.n6786 vss.t646 669.716
R29517 vss.n7060 vss.t1157 669.716
R29518 vss.n6805 vss.t1157 669.716
R29519 vss.t555 vss.n6805 669.716
R29520 vss.t555 vss.n6806 669.716
R29521 vss.t554 vss.n6806 669.716
R29522 vss.t554 vss.n7046 669.716
R29523 vss.t255 vss.n6503 669.716
R29524 vss.t255 vss.n6495 669.716
R29525 vss.t254 vss.n6495 669.716
R29526 vss.t254 vss.n9243 669.716
R29527 vss.n9243 vss.t1458 669.716
R29528 vss.n6878 vss.t1458 669.716
R29529 vss.n9223 vss.t589 669.716
R29530 vss.n6516 vss.t589 669.716
R29531 vss.t1410 vss.n6516 669.716
R29532 vss.t1410 vss.n6517 669.716
R29533 vss.t1409 vss.n6517 669.716
R29534 vss.t1409 vss.n9209 669.716
R29535 vss.t472 vss.n9168 669.716
R29536 vss.t472 vss.n9162 669.716
R29537 vss.t897 vss.n9162 669.716
R29538 vss.t897 vss.n9155 669.716
R29539 vss.t896 vss.n9155 669.716
R29540 vss.t896 vss.n9156 669.716
R29541 vss.t899 vss.n9156 669.716
R29542 vss.t899 vss.n6182 669.716
R29543 vss.t1334 vss.n6465 669.716
R29544 vss.t1334 vss.n6459 669.716
R29545 vss.t1465 vss.n6459 669.716
R29546 vss.t1465 vss.n6452 669.716
R29547 vss.t1464 vss.n6452 669.716
R29548 vss.t1464 vss.n6453 669.716
R29549 vss.t771 vss.n6453 669.716
R29550 vss.t771 vss.n6179 669.716
R29551 vss.t1314 vss.n7005 669.716
R29552 vss.t1314 vss.n6999 669.716
R29553 vss.t333 vss.n6999 669.716
R29554 vss.t333 vss.n6992 669.716
R29555 vss.t332 vss.n6992 669.716
R29556 vss.t332 vss.n6993 669.716
R29557 vss.t87 vss.n6993 669.716
R29558 vss.t87 vss.n6176 669.716
R29559 vss.t1370 vss.n6691 669.716
R29560 vss.t1370 vss.n6685 669.716
R29561 vss.t985 vss.n6685 669.716
R29562 vss.t985 vss.n6678 669.716
R29563 vss.t987 vss.n6678 669.716
R29564 vss.t987 vss.n6679 669.716
R29565 vss.t1008 vss.n6679 669.716
R29566 vss.t1008 vss.n6173 669.716
R29567 vss.t213 vss.n7196 669.716
R29568 vss.t213 vss.n7190 669.716
R29569 vss.t85 vss.n7190 669.716
R29570 vss.t85 vss.n7183 669.716
R29571 vss.t84 vss.n7183 669.716
R29572 vss.t84 vss.n7184 669.716
R29573 vss.t314 vss.n7184 669.716
R29574 vss.t314 vss.n6170 669.716
R29575 vss.t1340 vss.n6153 669.716
R29576 vss.t1340 vss.n6147 669.716
R29577 vss.t1293 vss.n6147 669.716
R29578 vss.t1293 vss.n6140 669.716
R29579 vss.t1292 vss.n6140 669.716
R29580 vss.t1292 vss.n6141 669.716
R29581 vss.t1104 vss.n6141 669.716
R29582 vss.n9492 vss.t1104 669.716
R29583 vss.t510 vss.n9462 669.716
R29584 vss.t510 vss.n9455 669.716
R29585 vss.t230 vss.n9455 669.716
R29586 vss.t230 vss.n9456 669.716
R29587 vss.n9456 vss.t229 669.716
R29588 vss.n9477 vss.t229 669.716
R29589 vss.n9477 vss.t1254 669.716
R29590 vss.n9486 vss.t1254 669.716
R29591 vss.t211 vss.n6026 669.716
R29592 vss.t211 vss.n6020 669.716
R29593 vss.t731 vss.n6020 669.716
R29594 vss.t731 vss.n6013 669.716
R29595 vss.t733 vss.n6013 669.716
R29596 vss.t733 vss.n6014 669.716
R29597 vss.t1114 vss.n6014 669.716
R29598 vss.n6041 vss.t1114 669.716
R29599 vss.t1487 vss.n9418 669.716
R29600 vss.t1487 vss.n9410 669.716
R29601 vss.t941 vss.n9410 669.716
R29602 vss.t941 vss.n9412 669.716
R29603 vss.n9412 vss.t940 669.716
R29604 vss.n9435 vss.t940 669.716
R29605 vss.n9435 vss.t153 669.716
R29606 vss.n9444 vss.t153 669.716
R29607 vss.t1501 vss.n7145 669.716
R29608 vss.t1501 vss.n7139 669.716
R29609 vss.t1281 vss.n7139 669.716
R29610 vss.t1281 vss.n7132 669.716
R29611 vss.t1280 vss.n7132 669.716
R29612 vss.t1280 vss.n7133 669.716
R29613 vss.t1283 vss.n7133 669.716
R29614 vss.t1283 vss.n6168 669.716
R29615 vss.t1330 vss.n6647 669.716
R29616 vss.t1330 vss.n6641 669.716
R29617 vss.t1118 vss.n6641 669.716
R29618 vss.t1118 vss.n6634 669.716
R29619 vss.t1117 vss.n6634 669.716
R29620 vss.t1117 vss.n6635 669.716
R29621 vss.t1120 vss.n6635 669.716
R29622 vss.t1120 vss.n6171 669.716
R29623 vss.t482 vss.n6956 669.716
R29624 vss.t482 vss.n6950 669.716
R29625 vss.t547 vss.n6950 669.716
R29626 vss.t547 vss.n6943 669.716
R29627 vss.t546 vss.n6943 669.716
R29628 vss.t546 vss.n6944 669.716
R29629 vss.t550 vss.n6944 669.716
R29630 vss.t550 vss.n6174 669.716
R29631 vss.t1491 vss.n6420 669.716
R29632 vss.t1491 vss.n6414 669.716
R29633 vss.t900 vss.n6414 669.716
R29634 vss.t900 vss.n6407 669.716
R29635 vss.t902 vss.n6407 669.716
R29636 vss.t902 vss.n6408 669.716
R29637 vss.t1313 vss.n6408 669.716
R29638 vss.t1313 vss.n6177 669.716
R29639 vss.t1356 vss.n6342 669.716
R29640 vss.t1356 vss.n6336 669.716
R29641 vss.t189 vss.n6336 669.716
R29642 vss.t189 vss.n6329 669.716
R29643 vss.t188 vss.n6329 669.716
R29644 vss.t188 vss.n6330 669.716
R29645 vss.t1009 vss.n6330 669.716
R29646 vss.t1009 vss.n6180 669.716
R29647 vss.t609 vss.n9338 669.716
R29648 vss.t609 vss.n9332 669.716
R29649 vss.t535 vss.n9332 669.716
R29650 vss.t535 vss.n9325 669.716
R29651 vss.t534 vss.n9325 669.716
R29652 vss.t534 vss.n9326 669.716
R29653 vss.t1055 vss.n9326 669.716
R29654 vss.t1055 vss.n6183 669.716
R29655 vss.t641 vss.n2740 669.716
R29656 vss.t641 vss.n9756 669.716
R29657 vss.t712 vss.n9756 669.716
R29658 vss.t712 vss.n9758 669.716
R29659 vss.n9758 vss.t713 669.716
R29660 vss.n9749 vss.t713 669.716
R29661 vss.t476 vss.n9749 669.716
R29662 vss.t476 vss.n2768 669.716
R29663 vss.t451 vss.n2741 669.716
R29664 vss.t451 vss.n3196 669.716
R29665 vss.t494 vss.n3196 669.716
R29666 vss.t494 vss.n3198 669.716
R29667 vss.n3198 vss.t492 669.716
R29668 vss.n3189 vss.t492 669.716
R29669 vss.t1358 vss.n3189 669.716
R29670 vss.t1358 vss.n2769 669.716
R29671 vss.n9802 vss.t1056 669.716
R29672 vss.t1056 vss.n2994 669.716
R29673 vss.t968 vss.n2994 669.716
R29674 vss.t968 vss.n3001 669.716
R29675 vss.t969 vss.n3001 669.716
R29676 vss.n3011 vss.t969 669.716
R29677 vss.t625 vss.n3011 669.716
R29678 vss.t625 vss.n2770 669.716
R29679 vss.t399 vss.n2990 669.716
R29680 vss.t399 vss.n5226 669.716
R29681 vss.t1185 vss.n5226 669.716
R29682 vss.t1185 vss.n5228 669.716
R29683 vss.n5228 vss.t1186 669.716
R29684 vss.n5219 vss.t1186 669.716
R29685 vss.t480 vss.n5219 669.716
R29686 vss.t480 vss.n2771 669.716
R29687 vss.t517 vss.n2991 669.716
R29688 vss.t517 vss.n3039 669.716
R29689 vss.t198 vss.n3039 669.716
R29690 vss.t198 vss.n3041 669.716
R29691 vss.n3041 vss.t199 669.716
R29692 vss.n3032 vss.t199 669.716
R29693 vss.t1366 vss.n3032 669.716
R29694 vss.t1366 vss.n2772 669.716
R29695 vss.t441 vss.n2987 669.716
R29696 vss.t441 vss.n5096 669.716
R29697 vss.t0 vss.n5096 669.716
R29698 vss.t0 vss.n5098 669.716
R29699 vss.n5098 vss.t1 669.716
R29700 vss.n5089 vss.t1 669.716
R29701 vss.t1485 vss.n5089 669.716
R29702 vss.t1485 vss.n2773 669.716
R29703 vss.t707 vss.n2984 669.716
R29704 vss.t707 vss.n5285 669.716
R29705 vss.t704 vss.n5285 669.716
R29706 vss.t704 vss.n5287 669.716
R29707 vss.n5287 vss.t705 669.716
R29708 vss.n5278 vss.t705 669.716
R29709 vss.t1348 vss.n5278 669.716
R29710 vss.t1348 vss.n2774 669.716
R29711 vss.t637 vss.n2985 669.716
R29712 vss.t637 vss.n5013 669.716
R29713 vss.t1162 vss.n5013 669.716
R29714 vss.t1162 vss.n5015 669.716
R29715 vss.n5015 vss.t1163 669.716
R29716 vss.n5006 vss.t1163 669.716
R29717 vss.t1380 vss.n5006 669.716
R29718 vss.t1380 vss.n2775 669.716
R29719 vss.t436 vss.n2981 669.716
R29720 vss.t436 vss.n4894 669.716
R29721 vss.t603 vss.n4894 669.716
R29722 vss.t603 vss.n4896 669.716
R29723 vss.n4896 vss.t604 669.716
R29724 vss.n4887 vss.t604 669.716
R29725 vss.t1085 vss.n4887 669.716
R29726 vss.t1085 vss.n2776 669.716
R29727 vss.t749 vss.n4668 669.716
R29728 vss.t749 vss.n4669 669.716
R29729 vss.t750 vss.n4669 669.716
R29730 vss.t750 vss.n5619 669.716
R29731 vss.n5619 vss.t587 669.716
R29732 vss.n5612 vss.t587 669.716
R29733 vss.t253 vss.n5584 669.716
R29734 vss.t253 vss.n4691 669.716
R29735 vss.t1419 vss.n4691 669.716
R29736 vss.t1419 vss.n4692 669.716
R29737 vss.n4692 vss.t1420 669.716
R29738 vss.n5610 vss.t1420 669.716
R29739 vss.n5539 vss.t803 669.716
R29740 vss.n4755 vss.t803 669.716
R29741 vss.t804 vss.n4755 669.716
R29742 vss.t804 vss.n4756 669.716
R29743 vss.t1155 vss.n4756 669.716
R29744 vss.t1155 vss.n5526 669.716
R29745 vss.t1286 vss.n5498 669.716
R29746 vss.t1286 vss.n4777 669.716
R29747 vss.t1220 vss.n4777 669.716
R29748 vss.t1220 vss.n4778 669.716
R29749 vss.n4778 vss.t1221 669.716
R29750 vss.n5524 vss.t1221 669.716
R29751 vss.n5453 vss.t1525 669.716
R29752 vss.n4841 vss.t1525 669.716
R29753 vss.t1526 vss.n4841 669.716
R29754 vss.t1526 vss.n4842 669.716
R29755 vss.t601 vss.n4842 669.716
R29756 vss.t601 vss.n5440 669.716
R29757 vss.t934 vss.n5412 669.716
R29758 vss.t934 vss.n4863 669.716
R29759 vss.t1242 vss.n4863 669.716
R29760 vss.t1242 vss.n4864 669.716
R29761 vss.n4864 vss.t1243 669.716
R29762 vss.n5438 vss.t1243 669.716
R29763 vss.t154 vss.n9819 669.716
R29764 vss.t154 vss.n2884 669.716
R29765 vss.t410 vss.n2884 669.716
R29766 vss.t410 vss.n2886 669.716
R29767 vss.n2886 vss.t408 669.716
R29768 vss.n2877 vss.t408 669.716
R29769 vss.t15 vss.n2877 669.716
R29770 vss.t15 vss.n2777 669.716
R29771 vss.n2979 vss.t491 669.716
R29772 vss.t491 vss.n2937 669.716
R29773 vss.t1425 vss.n2937 669.716
R29774 vss.t1425 vss.n2944 669.716
R29775 vss.t1423 vss.n2944 669.716
R29776 vss.n2954 vss.t1423 669.716
R29777 vss.t1318 vss.n2954 669.716
R29778 vss.t1318 vss.n2778 669.716
R29779 vss.n2933 vss.t335 669.716
R29780 vss.t335 vss.n2890 669.716
R29781 vss.t789 vss.n2890 669.716
R29782 vss.t789 vss.n2897 669.716
R29783 vss.t790 vss.n2897 669.716
R29784 vss.n2907 vss.t790 669.716
R29785 vss.t470 vss.n2907 669.716
R29786 vss.t470 vss.n2779 669.716
R29787 vss.t832 vss.n2982 669.716
R29788 vss.t832 vss.n4935 669.716
R29789 vss.t1237 vss.n4935 669.716
R29790 vss.t1237 vss.n4937 669.716
R29791 vss.n4937 vss.t1235 669.716
R29792 vss.n4928 vss.t1235 669.716
R29793 vss.t1509 vss.n4928 669.716
R29794 vss.t1509 vss.n2780 669.716
R29795 vss.t146 vss.n2988 669.716
R29796 vss.t146 vss.n5137 669.716
R29797 vss.t1307 vss.n5137 669.716
R29798 vss.t1307 vss.n5139 669.716
R29799 vss.n5139 vss.t1308 669.716
R29800 vss.n5130 vss.t1308 669.716
R29801 vss.t508 vss.n5130 669.716
R29802 vss.t508 vss.n2781 669.716
R29803 vss.t240 vss.n3122 669.716
R29804 vss.t240 vss.n3117 669.716
R29805 vss.t710 vss.n3117 669.716
R29806 vss.t710 vss.n3119 669.716
R29807 vss.n3119 vss.t708 669.716
R29808 vss.n3110 vss.t708 669.716
R29809 vss.t1342 vss.n3110 669.716
R29810 vss.t1342 vss.n2782 669.716
R29811 vss.t580 vss.n4480 669.716
R29812 vss.t580 vss.n4474 669.716
R29813 vss.t159 vss.n4474 669.716
R29814 vss.t159 vss.n4466 669.716
R29815 vss.t161 vss.n4466 669.716
R29816 vss.t161 vss.n4499 669.716
R29817 vss.n4499 vss.t1206 669.716
R29818 vss.t1206 vss.n2703 669.716
R29819 vss.t568 vss.n4388 669.716
R29820 vss.t568 vss.n4382 669.716
R29821 vss.t488 vss.n4382 669.716
R29822 vss.t488 vss.n4374 669.716
R29823 vss.t490 vss.n4374 669.716
R29824 vss.t490 vss.n4407 669.716
R29825 vss.n4407 vss.t1062 669.716
R29826 vss.t1062 vss.n2700 669.716
R29827 vss.t1503 vss.n4340 669.716
R29828 vss.t1503 vss.n4334 669.716
R29829 vss.t1259 vss.n4334 669.716
R29830 vss.t1259 vss.n4326 669.716
R29831 vss.t1261 vss.n4326 669.716
R29832 vss.t1261 vss.n4359 669.716
R29833 vss.n4359 vss.t975 669.716
R29834 vss.t975 vss.n2702 669.716
R29835 vss.t1071 vss.n3740 669.716
R29836 vss.t1071 vss.n3734 669.716
R29837 vss.t1255 vss.n3734 669.716
R29838 vss.t1255 vss.n3726 669.716
R29839 vss.t1257 vss.n3726 669.716
R29840 vss.t1257 vss.n3759 669.716
R29841 vss.n3759 vss.t1116 669.716
R29842 vss.t1116 vss.n2697 669.716
R29843 vss.t623 vss.n4042 669.716
R29844 vss.t623 vss.n4036 669.716
R29845 vss.t1126 vss.n4036 669.716
R29846 vss.t1126 vss.n4028 669.716
R29847 vss.t1125 vss.n4028 669.716
R29848 vss.t1125 vss.n4061 669.716
R29849 vss.n4061 vss.t316 669.716
R29850 vss.t316 vss.n2694 669.716
R29851 vss.t1493 vss.n3695 669.716
R29852 vss.t1493 vss.n3689 669.716
R29853 vss.t1441 vss.n3689 669.716
R29854 vss.t1441 vss.n3681 669.716
R29855 vss.t1440 vss.n3681 669.716
R29856 vss.t1440 vss.n3714 669.716
R29857 vss.n3714 vss.t1443 669.716
R29858 vss.t1443 vss.n2696 669.716
R29859 vss.t1483 vss.n4096 669.716
R29860 vss.t1483 vss.n4090 669.716
R29861 vss.t352 vss.n4090 669.716
R29862 vss.t352 vss.n4082 669.716
R29863 vss.t354 vss.n4082 669.716
R29864 vss.t354 vss.n4115 669.716
R29865 vss.n4115 vss.t197 669.716
R29866 vss.t197 vss.n2691 669.716
R29867 vss.t566 vss.n3520 669.716
R29868 vss.t566 vss.n3514 669.716
R29869 vss.t727 vss.n3514 669.716
R29870 vss.t727 vss.n3506 669.716
R29871 vss.t729 vss.n3506 669.716
R29872 vss.t729 vss.n3539 669.716
R29873 vss.n3539 vss.t551 669.716
R29874 vss.t551 vss.n2688 669.716
R29875 vss.t617 vss.n3475 669.716
R29876 vss.t617 vss.n3469 669.716
R29877 vss.t1212 vss.n3469 669.716
R29878 vss.t1212 vss.n3461 669.716
R29879 vss.t1211 vss.n3461 669.716
R29880 vss.t1211 vss.n3494 669.716
R29881 vss.n3494 vss.t124 669.716
R29882 vss.t124 vss.n2690 669.716
R29883 vss.t379 vss.n5763 669.716
R29884 vss.t379 vss.n5757 669.716
R29885 vss.t746 vss.n5757 669.716
R29886 vss.t746 vss.n5749 669.716
R29887 vss.t748 vss.n5749 669.716
R29888 vss.t748 vss.n5782 669.716
R29889 vss.n5782 vss.t78 669.716
R29890 vss.t78 vss.n2685 669.716
R29891 vss.t695 vss.n4564 669.716
R29892 vss.t695 vss.n4418 669.716
R29893 vss.t697 vss.n4418 669.716
R29894 vss.t697 vss.n4606 669.716
R29895 vss.n4606 vss.t698 669.716
R29896 vss.n4558 vss.t698 669.716
R29897 vss.n4586 vss.t597 669.716
R29898 vss.n4576 vss.t597 669.716
R29899 vss.t1267 vss.n4576 669.716
R29900 vss.t1267 vss.n3638 669.716
R29901 vss.t1269 vss.n3638 669.716
R29902 vss.t1269 vss.n3639 669.716
R29903 vss.t525 vss.n3834 669.716
R29904 vss.t525 vss.n3808 669.716
R29905 vss.t524 vss.n3808 669.716
R29906 vss.t524 vss.n4168 669.716
R29907 vss.n4168 vss.t1193 669.716
R29908 vss.n3828 vss.t1193 669.716
R29909 vss.n4148 vss.t1151 669.716
R29910 vss.n3847 vss.t1151 669.716
R29911 vss.t426 vss.n3847 669.716
R29912 vss.t426 vss.n3848 669.716
R29913 vss.t428 vss.n3848 669.716
R29914 vss.t428 vss.n4136 669.716
R29915 vss.t329 vss.n3557 669.716
R29916 vss.t329 vss.n3549 669.716
R29917 vss.t331 vss.n3549 669.716
R29918 vss.t331 vss.n5835 669.716
R29919 vss.n5835 vss.t1306 669.716
R29920 vss.n3921 vss.t1306 669.716
R29921 vss.n5815 vss.t1475 669.716
R29922 vss.n3570 vss.t1475 669.716
R29923 vss.t738 vss.n3570 669.716
R29924 vss.t738 vss.n3571 669.716
R29925 vss.t740 vss.n3571 669.716
R29926 vss.t740 vss.n5803 669.716
R29927 vss.t1075 vss.n2662 669.716
R29928 vss.t1075 vss.n2656 669.716
R29929 vss.t405 vss.n2656 669.716
R29930 vss.t405 vss.n2647 669.716
R29931 vss.t407 vss.n2647 669.716
R29932 vss.t407 vss.n2648 669.716
R29933 vss.n2648 vss.t450 669.716
R29934 vss.n2684 vss.t450 669.716
R29935 vss.t3 vss.n3400 669.716
R29936 vss.t3 vss.n3394 669.716
R29937 vss.t647 vss.n3394 669.716
R29938 vss.t647 vss.n3386 669.716
R29939 vss.t649 vss.n3386 669.716
R29940 vss.t649 vss.n3419 669.716
R29941 vss.n3419 vss.t495 669.716
R29942 vss.t495 vss.n2687 669.716
R29943 vss.t391 vss.n3997 669.716
R29944 vss.t391 vss.n3991 669.716
R29945 vss.t431 vss.n3991 669.716
R29946 vss.t431 vss.n3983 669.716
R29947 vss.t433 vss.n3983 669.716
R29948 vss.t433 vss.n4016 669.716
R29949 vss.n4016 vss.t840 669.716
R29950 vss.t840 vss.n2693 669.716
R29951 vss.t486 vss.n4264 669.716
R29952 vss.t486 vss.n4258 669.716
R29953 vss.t1452 vss.n4258 669.716
R29954 vss.t1452 vss.n4250 669.716
R29955 vss.t1451 vss.n4250 669.716
R29956 vss.t1451 vss.n4283 669.716
R29957 vss.n4283 vss.t1253 669.716
R29958 vss.t1253 vss.n2699 669.716
R29959 vss.t478 vss.n5907 669.716
R29960 vss.t478 vss.n5901 669.716
R29961 vss.t1064 vss.n5901 669.716
R29962 vss.t1064 vss.n5894 669.716
R29963 vss.t1066 vss.n5894 669.716
R29964 vss.t1066 vss.n5895 669.716
R29965 vss.t236 vss.n5895 669.716
R29966 vss.t236 vss.n2705 669.716
R29967 vss.t1173 vss.n8950 669.716
R29968 vss.t1173 vss.n7485 669.716
R29969 vss.t264 vss.n7485 669.716
R29970 vss.t264 vss.n7478 669.716
R29971 vss.t262 vss.n7478 669.716
R29972 vss.t262 vss.n7479 669.716
R29973 vss.t1505 vss.n7479 669.716
R29974 vss.t1505 vss.n7325 669.716
R29975 vss.n8901 vss.t1517 669.716
R29976 vss.n8867 vss.t1517 669.716
R29977 vss.t194 vss.n8867 669.716
R29978 vss.t194 vss.n8868 669.716
R29979 vss.t195 vss.n8868 669.716
R29980 vss.t195 vss.n8889 669.716
R29981 vss.n8889 vss.t572 669.716
R29982 vss.t572 vss.n7326 669.716
R29983 vss.t786 vss.n8831 669.716
R29984 vss.t786 vss.n7674 669.716
R29985 vss.t783 vss.n7674 669.716
R29986 vss.t783 vss.n7667 669.716
R29987 vss.t784 vss.n7667 669.716
R29988 vss.t784 vss.n7668 669.716
R29989 vss.t1073 vss.n7668 669.716
R29990 vss.t1073 vss.n7327 669.716
R29991 vss.n8782 vss.t1134 669.716
R29992 vss.n8748 vss.t1134 669.716
R29993 vss.t1534 vss.n8748 669.716
R29994 vss.t1534 vss.n8749 669.716
R29995 vss.t1535 vss.n8749 669.716
R29996 vss.t1535 vss.n8770 669.716
R29997 vss.n8770 vss.t1376 669.716
R29998 vss.t1376 vss.n7328 669.716
R29999 vss.t1298 vss.n8712 669.716
R30000 vss.t1298 vss.n7861 669.716
R30001 vss.t1295 vss.n7861 669.716
R30002 vss.t1295 vss.n7854 669.716
R30003 vss.t1296 vss.n7854 669.716
R30004 vss.t1296 vss.n7855 669.716
R30005 vss.t611 vss.n7855 669.716
R30006 vss.t611 vss.n7329 669.716
R30007 vss.n9006 vss.t561 669.716
R30008 vss.n7307 vss.t561 669.716
R30009 vss.t411 vss.n7307 669.716
R30010 vss.t411 vss.n7308 669.716
R30011 vss.t412 vss.n7308 669.716
R30012 vss.t412 vss.n8994 669.716
R30013 vss.n8994 vss.t383 669.716
R30014 vss.n8987 vss.t383 669.716
R30015 vss.t440 vss.n8221 669.716
R30016 vss.t440 vss.n8004 669.716
R30017 vss.t558 vss.n8004 669.716
R30018 vss.t558 vss.n7997 669.716
R30019 vss.t559 vss.n7997 669.716
R30020 vss.t559 vss.n7998 669.716
R30021 vss.t1507 vss.n7998 669.716
R30022 vss.t1507 vss.n7330 669.716
R30023 vss.n8218 vss.t756 669.716
R30024 vss.n8184 vss.t756 669.716
R30025 vss.t370 vss.n8184 669.716
R30026 vss.t370 vss.n8185 669.716
R30027 vss.t371 vss.n8185 669.716
R30028 vss.t371 vss.n8206 669.716
R30029 vss.n8206 vss.t1346 669.716
R30030 vss.t1346 vss.n7331 669.716
R30031 vss.t241 vss.n7927 669.716
R30032 vss.t241 vss.n7921 669.716
R30033 vss.t650 vss.n7921 669.716
R30034 vss.t650 vss.n7914 669.716
R30035 vss.t651 vss.n7914 669.716
R30036 vss.t651 vss.n7915 669.716
R30037 vss.t484 vss.n7915 669.716
R30038 vss.t484 vss.n7333 669.716
R30039 vss.t165 vss.n7786 669.716
R30040 vss.t165 vss.n7780 669.716
R30041 vss.t162 vss.n7780 669.716
R30042 vss.t162 vss.n7773 669.716
R30043 vss.t163 vss.n7773 669.716
R30044 vss.t163 vss.n7774 669.716
R30045 vss.t496 vss.n7774 669.716
R30046 vss.t496 vss.n7334 669.716
R30047 vss.t425 vss.n7706 669.716
R30048 vss.t425 vss.n7700 669.716
R30049 vss.t225 vss.n7700 669.716
R30050 vss.t225 vss.n7693 669.716
R30051 vss.t223 vss.n7693 669.716
R30052 vss.t223 vss.n7694 669.716
R30053 vss.t5 vss.n7694 669.716
R30054 vss.t5 vss.n7335 669.716
R30055 vss.n8828 vss.t1013 669.716
R30056 vss.n8794 vss.t1013 669.716
R30057 vss.t1010 vss.n8794 669.716
R30058 vss.t1010 vss.n8795 669.716
R30059 vss.t1011 vss.n8795 669.716
R30060 vss.t1011 vss.n8816 669.716
R30061 vss.n8816 vss.t205 669.716
R30062 vss.t205 vss.n7336 669.716
R30063 vss.t1133 vss.n7563 669.716
R30064 vss.t1133 vss.n7557 669.716
R30065 vss.t838 vss.n7557 669.716
R30066 vss.t838 vss.n7550 669.716
R30067 vss.t836 vss.n7550 669.716
R30068 vss.t836 vss.n7551 669.716
R30069 vss.t633 vss.n7551 669.716
R30070 vss.t633 vss.n7337 669.716
R30071 vss.n8947 vss.t361 669.716
R30072 vss.n8913 vss.t361 669.716
R30073 vss.t312 vss.n8913 669.716
R30074 vss.t312 vss.n8914 669.716
R30075 vss.t310 vss.n8914 669.716
R30076 vss.t310 vss.n8935 669.716
R30077 vss.n8935 vss.t9 669.716
R30078 vss.t9 vss.n7338 669.716
R30079 vss.n7535 vss.t662 669.716
R30080 vss.n7501 vss.t662 669.716
R30081 vss.t1467 vss.n7501 669.716
R30082 vss.t1467 vss.n7502 669.716
R30083 vss.t1468 vss.n7502 669.716
R30084 vss.t1468 vss.n7523 669.716
R30085 vss.n7523 vss.t215 669.716
R30086 vss.t215 vss.n7339 669.716
R30087 vss.t23 vss.n512 669.716
R30088 vss.t23 vss.n624 669.716
R30089 vss.t136 vss.n624 669.716
R30090 vss.t136 vss.n626 669.716
R30091 vss.n626 vss.t138 669.716
R30092 vss.n649 vss.t138 669.716
R30093 vss.n649 vss.t132 669.716
R30094 vss.n658 vss.t132 669.716
R30095 vss.t828 vss.n2363 669.716
R30096 vss.t828 vss.n10114 669.716
R30097 vss.t1305 vss.n10114 669.716
R30098 vss.t1305 vss.n10116 669.716
R30099 vss.n10116 vss.t1303 669.716
R30100 vss.n10107 vss.t1303 669.716
R30101 vss.t468 vss.n10107 669.716
R30102 vss.t468 vss.n2146 669.716
R30103 vss.t252 vss.n2360 669.716
R30104 vss.t252 vss.n12872 669.716
R30105 vss.t288 vss.n12872 669.716
R30106 vss.t288 vss.n12874 669.716
R30107 vss.n12874 vss.t286 669.716
R30108 vss.n12865 vss.t286 669.716
R30109 vss.t1479 vss.n12865 669.716
R30110 vss.t1479 vss.n2147 669.716
R30111 vss.t1230 vss.n2361 669.716
R30112 vss.t1230 vss.n10155 669.716
R30113 vss.t299 vss.n10155 669.716
R30114 vss.t299 vss.n10157 669.716
R30115 vss.n10157 vss.t297 669.716
R30116 vss.n10148 vss.t297 669.716
R30117 vss.t385 vss.n10148 669.716
R30118 vss.t385 vss.n2148 669.716
R30119 vss.t1450 vss.n2357 669.716
R30120 vss.t1450 vss.n12421 669.716
R30121 vss.t464 vss.n12421 669.716
R30122 vss.t464 vss.n12423 669.716
R30123 vss.n12423 vss.t462 669.716
R30124 vss.n12414 vss.t462 669.716
R30125 vss.t7 vss.n12414 669.716
R30126 vss.t7 vss.n2149 669.716
R30127 vss.t627 vss.n2354 669.716
R30128 vss.t627 vss.n11750 669.716
R30129 vss.t228 vss.n11750 669.716
R30130 vss.t228 vss.n11752 669.716
R30131 vss.n11752 vss.t226 669.716
R30132 vss.n11743 vss.t226 669.716
R30133 vss.t209 vss.n11743 669.716
R30134 vss.t209 vss.n2150 669.716
R30135 vss.t369 vss.n2355 669.716
R30136 vss.t369 vss.n12466 669.716
R30137 vss.t221 vss.n12466 669.716
R30138 vss.t221 vss.n12468 669.716
R30139 vss.n12468 vss.t219 669.716
R30140 vss.n12459 vss.t219 669.716
R30141 vss.t1499 vss.n12459 669.716
R30142 vss.t1499 vss.n2151 669.716
R30143 vss.n2349 vss.t1287 669.716
R30144 vss.t1287 vss.n2307 669.716
R30145 vss.t981 vss.n2307 669.716
R30146 vss.t981 vss.n2314 669.716
R30147 vss.t979 vss.n2314 669.716
R30148 vss.n2324 vss.t979 669.716
R30149 vss.t1362 vss.n2324 669.716
R30150 vss.t1362 vss.n2152 669.716
R30151 vss.t404 vss.n2351 669.716
R30152 vss.t404 vss.n12291 669.716
R30153 vss.t1171 vss.n12291 669.716
R30154 vss.t1171 vss.n12293 669.716
R30155 vss.n12293 vss.t1169 669.716
R30156 vss.n12284 vss.t1169 669.716
R30157 vss.t1338 vss.n12284 669.716
R30158 vss.t1338 vss.n2153 669.716
R30159 vss.t243 vss.n2352 669.716
R30160 vss.t243 vss.n12336 669.716
R30161 vss.t933 vss.n12336 669.716
R30162 vss.t933 vss.n12338 669.716
R30163 vss.n12338 vss.t931 669.716
R30164 vss.n12329 vss.t931 669.716
R30165 vss.t1326 vss.n12329 669.716
R30166 vss.t1326 vss.n2154 669.716
R30167 vss.t1399 vss.n2358 669.716
R30168 vss.t1399 vss.n10232 669.716
R30169 vss.t439 vss.n10232 669.716
R30170 vss.t439 vss.n10234 669.716
R30171 vss.n10234 vss.t437 669.716
R30172 vss.n10225 vss.t437 669.716
R30173 vss.t1354 vss.n10225 669.716
R30174 vss.t1354 vss.n2155 669.716
R30175 vss.t1422 vss.n2364 669.716
R30176 vss.t1422 vss.n2412 669.716
R30177 vss.t135 vss.n2412 669.716
R30178 vss.t135 vss.n2414 669.716
R30179 vss.n2414 vss.t133 669.716
R30180 vss.n2405 vss.t133 669.716
R30181 vss.t389 vss.n2405 669.716
R30182 vss.t389 vss.n2156 669.716
R30183 vss.n12974 vss.t1150 669.716
R30184 vss.t1150 vss.n2367 669.716
R30185 vss.t1165 vss.n2367 669.716
R30186 vss.t1165 vss.n2374 669.716
R30187 vss.t1166 vss.n2374 669.716
R30188 vss.n2384 vss.t1166 669.716
R30189 vss.t203 vss.n2384 669.716
R30190 vss.t203 vss.n2157 669.716
R30191 vss.t723 vss.n2496 669.716
R30192 vss.t723 vss.n2491 669.716
R30193 vss.t61 vss.n2491 669.716
R30194 vss.t61 vss.n2493 669.716
R30195 vss.n2493 vss.t59 669.716
R30196 vss.n2484 vss.t59 669.716
R30197 vss.t570 vss.n2484 669.716
R30198 vss.t570 vss.n2158 669.716
R30199 vss.t745 vss.n12153 669.716
R30200 vss.t745 vss.n11800 669.716
R30201 vss.t1124 vss.n11800 669.716
R30202 vss.t1124 vss.n11794 669.716
R30203 vss.t1122 vss.n11794 669.716
R30204 vss.t1122 vss.n11786 669.716
R30205 vss.t416 vss.n12183 669.716
R30206 vss.t416 vss.n12185 669.716
R30207 vss.n12185 vss.t414 669.716
R30208 vss.n11785 vss.t414 669.716
R30209 vss.t591 vss.n11785 669.716
R30210 vss.n12176 vss.t591 669.716
R30211 vss.t1249 vss.n12549 669.716
R30212 vss.t1249 vss.n11713 669.716
R30213 vss.t1402 vss.n11713 669.716
R30214 vss.t1402 vss.n11707 669.716
R30215 vss.t1400 vss.n11707 669.716
R30216 vss.t1400 vss.n11699 669.716
R30217 vss.n11687 vss.t638 669.716
R30218 vss.n11631 vss.t638 669.716
R30219 vss.t639 vss.n11631 669.716
R30220 vss.n11635 vss.t639 669.716
R30221 vss.n11635 vss.t1395 669.716
R30222 vss.n12572 vss.t1395 669.716
R30223 vss.n12830 vss.t1310 669.716
R30224 vss.t1310 vss.n12772 669.716
R30225 vss.t1240 vss.n12772 669.716
R30226 vss.t1240 vss.n12779 669.716
R30227 vss.t1238 vss.n12779 669.716
R30228 vss.n12791 vss.t1238 669.716
R30229 vss.t1447 vss.n10083 669.716
R30230 vss.t1447 vss.n10092 669.716
R30231 vss.t1448 vss.n10092 669.716
R30232 vss.n12801 vss.t1448 669.716
R30233 vss.n12801 vss.t1473 669.716
R30234 vss.n12808 vss.t1473 669.716
R30235 vss.t387 vss.n10420 669.716
R30236 vss.t387 vss.n10474 669.716
R30237 vss.t758 vss.n10474 669.716
R30238 vss.t758 vss.n10466 669.716
R30239 vss.t760 vss.n10466 669.716
R30240 vss.t760 vss.n10498 669.716
R30241 vss.n10498 vss.t775 669.716
R30242 vss.t775 vss.n2052 669.716
R30243 vss.t1489 vss.n10421 669.716
R30244 vss.t1489 vss.n10695 669.716
R30245 vss.t1129 vss.n10695 669.716
R30246 vss.t1129 vss.n10687 669.716
R30247 vss.t1131 vss.n10687 669.716
R30248 vss.t1131 vss.n10719 669.716
R30249 vss.n10719 vss.t167 669.716
R30250 vss.t167 vss.n2058 669.716
R30251 vss.t1328 vss.n10422 669.716
R30252 vss.t1328 vss.n11009 669.716
R30253 vss.t927 vss.n11009 669.716
R30254 vss.t927 vss.n11001 669.716
R30255 vss.t929 vss.n11001 669.716
R30256 vss.t929 vss.n11033 669.716
R30257 vss.n11033 vss.t930 669.716
R30258 vss.t930 vss.n2064 669.716
R30259 vss.t1378 vss.n10423 669.716
R30260 vss.t1378 vss.n11117 669.716
R30261 vss.t355 vss.n11117 669.716
R30262 vss.t355 vss.n11110 669.716
R30263 vss.t357 vss.n11110 669.716
R30264 vss.t357 vss.n11111 669.716
R30265 vss.t911 vss.n11111 669.716
R30266 vss.t911 vss.n2070 669.716
R30267 vss.n12058 vss.t305 649.236
R30268 vss.n11915 vss.t305 649.236
R30269 vss.t304 vss.n11915 649.236
R30270 vss.n11919 vss.t304 649.236
R30271 vss.n11919 vss.t939 649.236
R30272 vss.n12045 vss.t939 649.236
R30273 vss.t1245 vss.n10633 649.236
R30274 vss.t1245 vss.n10635 649.236
R30275 vss.n10635 vss.t1247 649.236
R30276 vss.n11603 vss.t1247 649.236
R30277 vss.n11603 vss.t1248 649.236
R30278 vss.n11612 vss.t1248 649.236
R30279 vss.n11493 vss.t693 649.236
R30280 vss.n10894 vss.t693 649.236
R30281 vss.t692 vss.n10894 649.236
R30282 vss.n10982 vss.t692 649.236
R30283 vss.n10982 vss.t711 649.236
R30284 vss.n11480 vss.t711 649.236
R30285 vss.n12723 vss.t1250 649.236
R30286 vss.n10364 vss.t1250 649.236
R30287 vss.t1252 vss.n10364 649.236
R30288 vss.n10368 vss.t1252 649.236
R30289 vss.n10368 vss.t1172 649.236
R30290 vss.n12710 vss.t1172 649.236
R30291 vss.n13920 vss.t434 649.236
R30292 vss.t434 vss.n13303 649.236
R30293 vss.t249 vss.n13303 649.236
R30294 vss.t249 vss.n13310 649.236
R30295 vss.t250 vss.n13310 649.236
R30296 vss.n13325 vss.t250 649.236
R30297 vss.n13818 vss.t730 649.236
R30298 vss.t730 vss.n13386 649.236
R30299 vss.t715 vss.n13386 649.236
R30300 vss.t715 vss.n13393 649.236
R30301 vss.t716 vss.n13393 649.236
R30302 vss.n13405 vss.t716 649.236
R30303 vss.n13713 vss.t1386 649.236
R30304 vss.t1386 vss.n13466 649.236
R30305 vss.t1288 vss.n13466 649.236
R30306 vss.t1288 vss.n13473 649.236
R30307 vss.t1289 vss.n13473 649.236
R30308 vss.n13485 vss.t1289 649.236
R30309 vss.n13608 vss.t770 649.236
R30310 vss.n13555 vss.t770 649.236
R30311 vss.t1264 vss.n13555 649.236
R30312 vss.t1264 vss.n13556 649.236
R30313 vss.t1262 vss.n13556 649.236
R30314 vss.t1262 vss.n13596 649.236
R30315 vss.t294 vss.n530 649.236
R30316 vss.t294 vss.n522 649.236
R30317 vss.t296 vss.n522 649.236
R30318 vss.t296 vss.n14021 649.236
R30319 vss.n14021 vss.t512 649.236
R30320 vss.n659 vss.t512 649.236
R30321 vss.t527 vss.n750 649.236
R30322 vss.t527 vss.n751 649.236
R30323 vss.t529 vss.n751 649.236
R30324 vss.t529 vss.n790 649.236
R30325 vss.n790 vss.t125 649.236
R30326 vss.n779 vss.t125 649.236
R30327 vss.t279 vss.n1231 649.236
R30328 vss.t279 vss.n1827 649.236
R30329 vss.n1827 vss.t278 649.236
R30330 vss.t278 vss.n1243 649.236
R30331 vss.t281 vss.n1243 649.236
R30332 vss.t281 vss.n1821 649.236
R30333 vss.t365 vss.n1931 649.236
R30334 vss.t365 vss.n1142 649.236
R30335 vss.t367 vss.n1142 649.236
R30336 vss.t367 vss.n1973 649.236
R30337 vss.n1973 vss.t62 649.236
R30338 vss.n1925 vss.t62 649.236
R30339 vss.t80 vss.n8689 649.236
R30340 vss.t80 vss.n8313 649.236
R30341 vss.t97 vss.n8313 649.236
R30342 vss.t97 vss.n7877 649.236
R30343 vss.t95 vss.n7877 649.236
R30344 vss.t95 vss.n8305 649.236
R30345 vss.t82 vss.n8602 649.236
R30346 vss.t82 vss.n8409 649.236
R30347 vss.t147 vss.n8409 649.236
R30348 vss.t147 vss.n8410 649.236
R30349 vss.n8410 vss.t148 649.236
R30350 vss.n8629 vss.t148 649.236
R30351 vss.t292 vss.n8510 649.236
R30352 vss.t292 vss.n8511 649.236
R30353 vss.n8511 vss.t1105 649.236
R30354 vss.t1105 vss.n8506 649.236
R30355 vss.n8506 vss.t1106 649.236
R30356 vss.n8542 vss.t1106 649.236
R30357 vss.t1300 vss.n6070 649.236
R30358 vss.t1300 vss.n6061 649.236
R30359 vss.t1302 vss.n6061 649.236
R30360 vss.t1302 vss.n9570 649.236
R30361 vss.n9570 vss.t1291 649.236
R30362 vss.n6064 vss.t1291 649.236
R30363 vss.t532 vss.n6747 649.236
R30364 vss.t532 vss.n6588 649.236
R30365 vss.t531 vss.n6588 649.236
R30366 vss.t531 vss.n6589 649.236
R30367 vss.n6589 vss.t1516 649.236
R30368 vss.n7235 vss.t1516 649.236
R30369 vss.t670 vss.n6843 649.236
R30370 vss.t670 vss.n6834 649.236
R30371 vss.t672 vss.n6834 649.236
R30372 vss.t672 vss.n6835 649.236
R30373 vss.n6835 vss.t33 649.236
R30374 vss.n7044 vss.t33 649.236
R30375 vss.t1204 vss.n9065 649.236
R30376 vss.t1204 vss.n6535 649.236
R30377 vss.t1203 vss.n6535 649.236
R30378 vss.t1203 vss.n6536 649.236
R30379 vss.n6536 vss.t1138 649.236
R30380 vss.n9207 vss.t1138 649.236
R30381 vss.n4666 vss.t31 649.236
R30382 vss.n4647 vss.t31 649.236
R30383 vss.t30 vss.n4647 649.236
R30384 vss.t30 vss.n4648 649.236
R30385 vss.n4648 vss.t28 649.236
R30386 vss.n9908 vss.t28 649.236
R30387 vss.t313 vss.n5541 649.236
R30388 vss.t313 vss.n4734 649.236
R30389 vss.t661 vss.n4734 649.236
R30390 vss.t661 vss.n4735 649.236
R30391 vss.n4735 vss.t659 649.236
R30392 vss.n5567 vss.t659 649.236
R30393 vss.t34 vss.n5455 649.236
R30394 vss.t34 vss.n4820 649.236
R30395 vss.t336 vss.n4820 649.236
R30396 vss.t336 vss.n4821 649.236
R30397 vss.n4821 vss.t337 649.236
R30398 vss.n5481 vss.t337 649.236
R30399 vss.t744 vss.n5363 649.236
R30400 vss.t744 vss.n5364 649.236
R30401 vss.n5364 vss.t741 649.236
R30402 vss.t741 vss.n5359 649.236
R30403 vss.n5359 vss.t742 649.236
R30404 vss.n5395 vss.t742 649.236
R30405 vss.t724 vss.n4443 649.236
R30406 vss.t724 vss.n4531 649.236
R30407 vss.n4531 vss.t726 649.236
R30408 vss.t726 vss.n4455 649.236
R30409 vss.t1178 vss.n4455 649.236
R30410 vss.t1178 vss.n2707 649.236
R30411 vss.t234 vss.n3778 649.236
R30412 vss.t234 vss.n3768 649.236
R30413 vss.t233 vss.n3768 649.236
R30414 vss.t233 vss.n4203 649.236
R30415 vss.n4203 vss.t89 649.236
R30416 vss.n3772 vss.t89 649.236
R30417 vss.t1194 vss.n3886 649.236
R30418 vss.t1194 vss.n3877 649.236
R30419 vss.t1196 vss.n3877 649.236
R30420 vss.t1196 vss.n3878 649.236
R30421 vss.n3878 vss.t1428 649.236
R30422 vss.n4134 vss.t1428 649.236
R30423 vss.t1136 vss.n5659 649.236
R30424 vss.t1136 vss.n3591 649.236
R30425 vss.t1135 vss.n3591 649.236
R30426 vss.t1135 vss.n3592 649.236
R30427 vss.n3592 vss.t906 649.236
R30428 vss.n5801 vss.t906 649.236
R30429 vss.t537 vss.n8079 649.236
R30430 vss.t537 vss.n8072 649.236
R30431 vss.t182 vss.n8072 649.236
R30432 vss.t182 vss.n8063 649.236
R30433 vss.t183 vss.n8063 649.236
R30434 vss.t183 vss.n8064 649.236
R30435 vss.t435 vss.n12100 649.236
R30436 vss.t435 vss.n11844 649.236
R30437 vss.t540 vss.n11844 649.236
R30438 vss.t540 vss.n11838 649.236
R30439 vss.t538 vss.n11838 649.236
R30440 vss.t538 vss.n11826 649.236
R30441 vss.n12250 vss.t455 649.236
R30442 vss.t455 vss.n12190 649.236
R30443 vss.t93 vss.n12190 649.236
R30444 vss.t93 vss.n12197 649.236
R30445 vss.t91 vss.n12197 649.236
R30446 vss.n12209 vss.t91 649.236
R30447 vss.n11685 vss.t1184 649.236
R30448 vss.t1184 vss.n11641 649.236
R30449 vss.t831 vss.n11641 649.236
R30450 vss.t831 vss.n11648 649.236
R30451 vss.t829 vss.n11648 649.236
R30452 vss.n11660 vss.t829 649.236
R30453 vss.t1231 vss.n12922 649.236
R30454 vss.t1231 vss.n10077 649.236
R30455 vss.t275 vss.n10077 649.236
R30456 vss.t275 vss.n10071 649.236
R30457 vss.t273 vss.n10071 649.236
R30458 vss.t273 vss.n10058 649.236
R30459 vss.n8064 vss.t960 589.682
R30460 vss.n8219 vss.n8051 562.532
R30461 vss.n8219 vss.n8174 537.46
R30462 vss.n10409 vss.t1344 501.3
R30463 vss.n10399 vss.t1344 501.3
R30464 vss.t1460 vss.n10399 501.3
R30465 vss.t1460 vss.n2037 501.3
R30466 vss.t1462 vss.n2037 501.3
R30467 vss.t1462 vss.n2038 501.3
R30468 vss.t1439 vss.n2038 501.3
R30469 vss.n13138 vss.t1439 501.3
R30470 vss.t1495 vss.n812 501.3
R30471 vss.t1495 vss.n13171 501.3
R30472 vss.t348 vss.n13171 501.3
R30473 vss.t348 vss.n13164 501.3
R30474 vss.t350 vss.n13164 501.3
R30475 vss.t350 vss.n13196 501.3
R30476 vss.n13196 vss.t1097 501.3
R30477 vss.t1097 vss.n728 501.3
R30478 vss.t1079 vss.n6203 501.3
R30479 vss.t1079 vss.n6195 501.3
R30480 vss.t1090 vss.n6195 501.3
R30481 vss.t1090 vss.n6197 501.3
R30482 vss.n6197 vss.t1089 501.3
R30483 vss.n9373 vss.t1089 501.3
R30484 vss.n9373 vss.t1092 501.3
R30485 vss.n9382 vss.t1092 501.3
R30486 vss.t1322 vss.n9967 501.3
R30487 vss.t1322 vss.n9961 501.3
R30488 vss.t518 vss.n9961 501.3
R30489 vss.t518 vss.n2636 501.3
R30490 vss.t520 vss.n2636 501.3
R30491 vss.t520 vss.n9986 501.3
R30492 vss.n9986 vss.t277 501.3
R30493 vss.n9955 vss.t277 501.3
R30494 vss.n12088 vss.n12087 498.046
R30495 vss.n12599 vss.n12598 498.046
R30496 vss.n11528 vss.n11527 498.046
R30497 vss.n12757 vss.n12756 498.046
R30498 vss.n13873 vss.n13336 498.046
R30499 vss.n13768 vss.n13416 498.046
R30500 vss.n13663 vss.n13496 498.046
R30501 vss.n14154 vss.n457 498.046
R30502 vss.n668 vss.n667 498.046
R30503 vss.n1749 vss.n1706 498.046
R30504 vss.n1853 vss.n1210 498.046
R30505 vss.n715 vss.n698 498.046
R30506 vss.n8283 vss.n7894 498.046
R30507 vss.n8645 vss.n8644 498.046
R30508 vss.n8558 vss.n8557 498.046
R30509 vss.n7256 vss.n7255 498.046
R30510 vss.n6785 vss.n6726 498.046
R30511 vss.n6880 vss.n6879 498.046
R30512 vss.n9141 vss.n9140 498.046
R30513 vss.n3281 vss.n2716 498.046
R30514 vss.n5583 vss.n5582 498.046
R30515 vss.n5497 vss.n5496 498.046
R30516 vss.n5411 vss.n5410 498.046
R30517 vss.n4557 vss.n4421 498.046
R30518 vss.n3827 vss.n3811 498.046
R30519 vss.n3923 vss.n3922 498.046
R30520 vss.n5735 vss.n5734 498.046
R30521 vss.n8153 vss.n8116 498.046
R30522 vss.n12152 vss.n11806 498.046
R30523 vss.n12548 vss.n11719 498.046
R30524 vss.n12831 vss.n10315 498.046
R30525 vss.n10042 vss.n10029 498.046
R30526 vss.n12044 vss.n12043 482.334
R30527 vss.n12007 vss.n12006 482.334
R30528 vss.n11614 vss.n11613 482.334
R30529 vss.n10858 vss.n10824 482.334
R30530 vss.n11479 vss.n11478 482.334
R30531 vss.n10927 vss.n10926 482.334
R30532 vss.n13844 vss.n13364 482.334
R30533 vss.n13819 vss.n13377 482.334
R30534 vss.n13739 vss.n13444 482.334
R30535 vss.n13714 vss.n13457 482.334
R30536 vss.n13634 vss.n13524 482.334
R30537 vss.n13609 vss.n13537 482.334
R30538 vss.n13967 vss.n569 482.334
R30539 vss.n778 vss.n762 482.334
R30540 vss.n1779 vss.n1756 482.334
R30541 vss.n1820 vss.n1263 482.334
R30542 vss.n1883 vss.n1860 482.334
R30543 vss.n1924 vss.n1145 482.334
R30544 vss.n8078 vss.n7275 482.334
R30545 vss.n9017 vss.n9016 482.334
R30546 vss.n8688 vss.n8687 482.334
R30547 vss.n8673 vss.n8672 482.334
R30548 vss.n8601 vss.n8600 482.334
R30549 vss.n8586 vss.n8585 482.334
R30550 vss.n9516 vss.n6109 482.334
R30551 vss.n7237 vss.n7236 482.334
R30552 vss.n7061 vss.n6792 482.334
R30553 vss.n7046 vss.n7045 482.334
R30554 vss.n9224 vss.n6503 482.334
R30555 vss.n9209 vss.n9208 482.334
R30556 vss.n4668 vss.n4667 482.334
R30557 vss.n5611 vss.n5610 482.334
R30558 vss.n5540 vss.n5539 482.334
R30559 vss.n5525 vss.n5524 482.334
R30560 vss.n5454 vss.n5453 482.334
R30561 vss.n5439 vss.n5438 482.334
R30562 vss.n4587 vss.n4564 482.334
R30563 vss.n3771 vss.n3639 482.334
R30564 vss.n4149 vss.n3834 482.334
R30565 vss.n4136 vss.n4135 482.334
R30566 vss.n5816 vss.n3557 482.334
R30567 vss.n5803 vss.n5802 482.334
R30568 vss.n12175 vss.n11786 482.334
R30569 vss.n12251 vss.n12183 482.334
R30570 vss.n12571 vss.n11699 482.334
R30571 vss.n11687 vss.n11686 482.334
R30572 vss.n12809 vss.n12791 482.334
R30573 vss.n12921 vss.n10083 482.334
R30574 vss.n12059 vss.n12058 467.584
R30575 vss.n10671 vss.n10633 467.584
R30576 vss.n11494 vss.n11493 467.584
R30577 vss.n12724 vss.n12723 467.584
R30578 vss.n13898 vss.n13325 467.584
R30579 vss.n13793 vss.n13405 467.584
R30580 vss.n13688 vss.n13485 467.584
R30581 vss.n13596 vss.n13583 467.584
R30582 vss.n14002 vss.n530 467.584
R30583 vss.n1727 vss.n750 467.584
R30584 vss.n1831 vss.n1231 467.584
R30585 vss.n1954 vss.n1931 467.584
R30586 vss.n8305 vss.n8304 467.584
R30587 vss.n8630 vss.n8629 467.584
R30588 vss.n8543 vss.n8542 467.584
R30589 vss.n9551 vss.n6070 467.584
R30590 vss.n6763 vss.n6747 467.584
R30591 vss.n6893 vss.n6843 467.584
R30592 vss.n9081 vss.n9065 467.584
R30593 vss.n9909 vss.n9908 467.584
R30594 vss.n5568 vss.n5567 467.584
R30595 vss.n5482 vss.n5481 467.584
R30596 vss.n5396 vss.n5395 467.584
R30597 vss.n4535 vss.n4443 467.584
R30598 vss.n4184 vss.n3778 467.584
R30599 vss.n3936 vss.n3886 467.584
R30600 vss.n5675 vss.n5659 467.584
R30601 vss.n12122 vss.n11826 467.584
R30602 vss.n12227 vss.n12209 467.584
R30603 vss.n11662 vss.n11660 467.584
R30604 vss.n12942 vss.n10058 467.584
R30605 vss.n14731 vss.n191 376
R30606 vss.n14685 vss.n14684 376
R30607 vss.n14536 vss.n250 376
R30608 vss.n14490 vss.n14489 376
R30609 vss.n14341 vss.n309 376
R30610 vss.n14295 vss.n14294 376
R30611 vss.n14222 vss.n432 376
R30612 vss.n9952 vss.n9951 376
R30613 vss.n9949 vss.n9948 376
R30614 vss.n9946 vss.n9945 376
R30615 vss.n9943 vss.n9942 376
R30616 vss.n9940 vss.n9939 376
R30617 vss.n9937 vss.n9936 376
R30618 vss.n9934 vss.n9933 376
R30619 vss.n9818 vss.n2935 376
R30620 vss.n9816 vss.n9815 376
R30621 vss.n9813 vss.n9812 376
R30622 vss.n9810 vss.n9809 376
R30623 vss.n9807 vss.n9806 376
R30624 vss.n9804 vss.n9803 376
R30625 vss.n9900 vss.n9899 376
R30626 vss.n9386 vss.n9385 376
R30627 vss.n9389 vss.n9388 376
R30628 vss.n9392 vss.n9391 376
R30629 vss.n9395 vss.n9394 376
R30630 vss.n9398 vss.n9397 376
R30631 vss.n9491 vss.n9490 376
R30632 vss.n9488 vss.n9487 376
R30633 vss.n8949 vss.n7537 376
R30634 vss.n8903 vss.n8902 376
R30635 vss.n8830 vss.n7680 376
R30636 vss.n8784 vss.n8783 376
R30637 vss.n8711 vss.n8710 376
R30638 vss.n9008 vss.n9007 376
R30639 vss.n13263 vss.n13262 376
R30640 vss.n13260 vss.n13259 376
R30641 vss.n13257 vss.n13256 376
R30642 vss.n13254 vss.n13253 376
R30643 vss.n13251 vss.n13250 376
R30644 vss.n13942 vss.n13941 376
R30645 vss.n13939 vss.n13938 376
R30646 vss.n12993 vss.n2305 376
R30647 vss.n12991 vss.n12990 376
R30648 vss.n12988 vss.n12987 376
R30649 vss.n12985 vss.n12984 376
R30650 vss.n12982 vss.n12981 376
R30651 vss.n12979 vss.n12978 376
R30652 vss.n12976 vss.n12975 376
R30653 vss.n13135 vss.n13134 376
R30654 vss.n13132 vss.n13131 376
R30655 vss.n13129 vss.n13128 376
R30656 vss.n13126 vss.n13125 376
R30657 vss.n13123 vss.n13122 376
R30658 vss.n13120 vss.n13119 376
R30659 vss.n13117 vss.n13116 376
R30660 vss.t876 vss.n13266 315.219
R30661 vss.t876 vss.n722 315.219
R30662 vss.t780 vss.n722 315.219
R30663 vss.t780 vss.n712 315.219
R30664 vss.t782 vss.n712 315.219
R30665 vss.t782 vss.n13285 315.219
R30666 vss.n13285 vss.t645 315.219
R30667 vss.n716 vss.t645 315.219
R30668 vss.t888 vss.n6184 315.219
R30669 vss.t888 vss.n9114 315.219
R30670 vss.t1436 vss.n9114 315.219
R30671 vss.t1436 vss.n9105 315.219
R30672 vss.t1435 vss.n9105 315.219
R30673 vss.t1435 vss.n9106 315.219
R30674 vss.n9106 vss.t1179 315.219
R30675 vss.n9139 vss.t1179 315.219
R30676 vss.t884 vss.n2639 315.219
R30677 vss.t884 vss.n5708 315.219
R30678 vss.t513 vss.n5708 315.219
R30679 vss.t513 vss.n5699 315.219
R30680 vss.t515 vss.n5699 315.219
R30681 vss.t515 vss.n5700 315.219
R30682 vss.n5700 vss.t1427 315.219
R30683 vss.n5733 vss.t1427 315.219
R30684 vss.t1020 vss.n2048 315.219
R30685 vss.t1020 vss.n11874 315.219
R30686 vss.t893 vss.n11874 315.219
R30687 vss.t893 vss.n11865 315.219
R30688 vss.t895 vss.n11865 315.219
R30689 vss.t895 vss.n11866 315.219
R30690 vss.n11866 vss.t628 315.219
R30691 vss.n12086 vss.t628 315.219
R30692 vss.n12591 vss.t232 270.964
R30693 vss.n11520 vss.t142 270.964
R30694 vss.n12766 vss.t1147 270.964
R30695 vss.t268 vss.n689 270.964
R30696 vss.t516 vss.n685 270.964
R30697 vss.t1128 vss.n681 270.964
R30698 vss.n678 vss.t1279 270.964
R30699 vss.t545 vss.n682 270.964
R30700 vss.t315 vss.n686 270.964
R30701 vss.t1054 vss.n6574 270.964
R30702 vss.t1223 vss.n6570 270.964
R30703 vss.t424 vss.n6556 270.964
R30704 vss.n7266 vss.t839 270.964
R30705 vss.t248 vss.n6573 270.964
R30706 vss.t343 vss.n6569 270.964
R30707 vss.t699 vss.n3630 270.964
R30708 vss.t812 vss.n3626 270.964
R30709 vss.t1265 vss.n3612 270.964
R30710 vss.t155 vss.n4422 270.964
R30711 vss.t1284 vss.n3629 270.964
R30712 vss.t629 vss.n3625 270.964
R30713 vss.t1057 vss.n11807 270.964
R30714 vss.t1132 vss.n10615 270.964
R30715 vss.n12832 vss.t32 270.964
R30716 vss.t958 vss.n2051 267.55
R30717 vss.t1046 vss.n2054 267.55
R30718 vss.t841 vss.n2057 267.55
R30719 vss.t950 vss.n2060 267.55
R30720 vss.t993 vss.n2063 267.55
R30721 vss.t954 vss.n2066 267.55
R30722 vss.t1001 vss.n2069 267.55
R30723 vss.t914 vss.n13899 267.55
R30724 vss.t1024 vss.n192 267.55
R30725 vss.t47 vss.n13794 267.55
R30726 vss.t1026 vss.n251 267.55
R30727 vss.t991 vss.n13689 267.55
R30728 vss.t1040 vss.n310 267.55
R30729 vss.t1018 vss.n13588 267.55
R30730 vss.t999 vss.n536 267.55
R30731 vss.t952 vss.n575 267.55
R30732 vss.n13249 vss.t890 267.55
R30733 vss.t1022 vss.n740 267.55
R30734 vss.t997 vss.n737 267.55
R30735 vss.t847 vss.n734 267.55
R30736 vss.t886 vss.n731 267.55
R30737 vss.n9009 vss.t946 267.55
R30738 vss.n8709 vss.t912 267.55
R30739 vss.t1032 vss.n7681 267.55
R30740 vss.n8622 vss.t956 267.55
R30741 vss.t1030 vss.n7538 267.55
R30742 vss.n8535 vss.t1028 267.55
R30743 vss.t1042 vss.n6076 267.55
R30744 vss.t989 vss.n6115 267.55
R30745 vss.t43 vss.n6169 267.55
R30746 vss.t995 vss.n6172 267.55
R30747 vss.t918 vss.n6175 267.55
R30748 vss.t57 vss.n6178 267.55
R30749 vss.t1034 vss.n6181 267.55
R30750 vss.n9901 vss.t1044 267.55
R30751 vss.t787 vss.n2992 267.55
R30752 vss.t845 vss.n2989 267.55
R30753 vss.t966 vss.n2986 267.55
R30754 vss.t878 vss.n2983 267.55
R30755 vss.t964 vss.n2980 267.55
R30756 vss.n5388 vss.t55 267.55
R30757 vss.t948 vss.n2704 267.55
R30758 vss.t916 vss.n2701 267.55
R30759 vss.t1036 vss.n2698 267.55
R30760 vss.t962 vss.n2695 267.55
R30761 vss.t849 vss.n2692 267.55
R30762 vss.t51 vss.n2689 267.55
R30763 vss.t1003 vss.n2686 267.55
R30764 vss.t1038 vss.n11828 267.55
R30765 vss.t872 vss.n2350 267.55
R30766 vss.t851 vss.n2353 267.55
R30767 vss.t874 vss.n2356 267.55
R30768 vss.t882 vss.n2359 267.55
R30769 vss.t843 vss.n2362 267.55
R30770 vss.t45 vss.n2365 267.55
R30771 vss.n12036 vss.t1191 264.219
R30772 vss.n11623 vss.t685 264.219
R30773 vss.t1459 vss.n10322 264.219
R30774 vss.t722 vss.n687 264.219
R30775 vss.t687 vss.n683 264.219
R30776 vss.t988 vss.n679 264.219
R30777 vss.t1148 vss.n680 264.219
R30778 vss.t1067 vss.n684 264.219
R30779 vss.t1397 vss.n688 264.219
R30780 vss.t272 vss.n6572 264.219
R30781 vss.t1115 vss.n6568 264.219
R30782 vss.n7247 vss.t910 264.219
R30783 vss.t557 vss.n6571 264.219
R30784 vss.n6567 vss.t285 264.219
R30785 vss.n5631 vss.t752 264.219
R30786 vss.t938 vss.n3628 264.219
R30787 vss.t1438 vss.n3624 264.219
R30788 vss.n4627 vss.t465 264.219
R30789 vss.t423 vss.n3627 264.219
R30790 vss.n3623 vss.t1093 264.219
R30791 vss.n9037 vss.t1382 264.219
R30792 vss.n12252 vss.t1258 264.219
R30793 vss.n12586 vss.t757 264.219
R30794 vss.t1426 vss.n10084 264.219
R30795 vss.n120 vss.n119 263.154
R30796 vss.n409 vss.n408 263.154
R30797 vss.n286 vss.n285 263.154
R30798 vss.n14443 vss.n14442 263.154
R30799 vss.n227 vss.n226 263.154
R30800 vss.n14638 vss.n14637 263.154
R30801 vss.n150 vss.n149 263.154
R30802 vss.n14776 vss.n69 263.154
R30803 vss.n14048 vss.n14047 263.154
R30804 vss.n14055 vss.n507 263.154
R30805 vss.n14038 vss.n14034 263.154
R30806 vss.n1597 vss.n1594 263.154
R30807 vss.n1584 vss.n1581 263.154
R30808 vss.n1605 vss.n1604 263.154
R30809 vss.n1302 vss.n1299 263.154
R30810 vss.n1289 vss.n1286 263.154
R30811 vss.n1310 vss.n1309 263.154
R30812 vss.n1041 vss.n1038 263.154
R30813 vss.n1028 vss.n1025 263.154
R30814 vss.n1049 vss.n1048 263.154
R30815 vss.n1434 vss.n1431 263.154
R30816 vss.n1421 vss.n1418 263.154
R30817 vss.n1442 vss.n1441 263.154
R30818 vss.n1514 vss.n1511 263.154
R30819 vss.n1501 vss.n1498 263.154
R30820 vss.n1522 vss.n1521 263.154
R30821 vss.n956 vss.n953 263.154
R30822 vss.n966 vss.n937 263.154
R30823 vss.n964 vss.n963 263.154
R30824 vss.n1008 vss.n1005 263.154
R30825 vss.n13206 vss.n989 263.154
R30826 vss.n13204 vss.n1015 263.154
R30827 vss.n7368 vss.n7346 263.154
R30828 vss.n7844 vss.n7843 263.154
R30829 vss.n7657 vss.n7656 263.154
R30830 vss.n7468 vss.n7467 263.154
R30831 vss.n7434 vss.n7433 263.154
R30832 vss.n7622 vss.n7621 263.154
R30833 vss.n7765 vss.n7764 263.154
R30834 vss.n7986 vss.n7985 263.154
R30835 vss.n6248 vss.n6247 263.154
R30836 vss.n6254 vss.n6228 263.154
R30837 vss.n6237 vss.n6007 263.154
R30838 vss.n6603 vss.n6602 263.154
R30839 vss.n6608 vss.n6607 263.154
R30840 vss.n6628 vss.n6627 263.154
R30841 vss.n6376 vss.n6375 263.154
R30842 vss.n6381 vss.n6380 263.154
R30843 vss.n6401 vss.n6400 263.154
R30844 vss.n9277 vss.n9276 263.154
R30845 vss.n9283 vss.n6323 263.154
R30846 vss.n9266 vss.n9257 263.154
R30847 vss.n6912 vss.n6911 263.154
R30848 vss.n6917 vss.n6916 263.154
R30849 vss.n6937 vss.n6936 263.154
R30850 vss.n7101 vss.n7100 263.154
R30851 vss.n7106 vss.n7105 263.154
R30852 vss.n7126 vss.n7125 263.154
R30853 vss.n6286 vss.n6285 263.154
R30854 vss.n6292 vss.n6265 263.154
R30855 vss.n6275 vss.n6266 263.154
R30856 vss.n9300 vss.n9299 263.154
R30857 vss.n9313 vss.n9312 263.154
R30858 vss.n9319 vss.n9318 263.154
R30859 vss.n3319 vss.n3318 263.154
R30860 vss.n3332 vss.n3329 263.154
R30861 vss.n5888 vss.n5887 263.154
R30862 vss.n3230 vss.n3228 263.154
R30863 vss.n3073 vss.n3071 263.154
R30864 vss.n5047 vss.n5045 263.154
R30865 vss.n2839 vss.n2837 263.154
R30866 vss.n9862 vss.n9861 263.154
R30867 vss.n4970 vss.n4968 263.154
R30868 vss.n5172 vss.n5170 263.154
R30869 vss.n3153 vss.n3151 263.154
R30870 vss.n4301 vss.n4297 263.154
R30871 vss.n4312 vss.n4308 263.154
R30872 vss.n4320 vss.n4319 263.154
R30873 vss.n3656 vss.n3652 263.154
R30874 vss.n3667 vss.n3663 263.154
R30875 vss.n3675 vss.n3674 263.154
R30876 vss.n3436 vss.n3432 263.154
R30877 vss.n3447 vss.n3443 263.154
R30878 vss.n3455 vss.n3454 263.154
R30879 vss.n5874 vss.n5870 263.154
R30880 vss.n9996 vss.n2627 263.154
R30881 vss.n9994 vss.n2629 263.154
R30882 vss.n3373 vss.n3369 263.154
R30883 vss.n5854 vss.n5851 263.154
R30884 vss.n5849 vss.n3380 263.154
R30885 vss.n3958 vss.n3954 263.154
R30886 vss.n3969 vss.n3965 263.154
R30887 vss.n3977 vss.n3976 263.154
R30888 vss.n4225 vss.n4221 263.154
R30889 vss.n4236 vss.n4232 263.154
R30890 vss.n4244 vss.n4243 263.154
R30891 vss.n14047 vss.n14044 252.988
R30892 vss.n14056 vss.n14055 252.988
R30893 vss.n14039 vss.n14038 252.988
R30894 vss.n1598 vss.n1597 252.988
R30895 vss.n1585 vss.n1584 252.988
R30896 vss.n1604 vss.n1574 252.988
R30897 vss.n1303 vss.n1302 252.988
R30898 vss.n1290 vss.n1289 252.988
R30899 vss.n1309 vss.n1279 252.988
R30900 vss.n1042 vss.n1041 252.988
R30901 vss.n1029 vss.n1028 252.988
R30902 vss.n1048 vss.n1018 252.988
R30903 vss.n1435 vss.n1434 252.988
R30904 vss.n1422 vss.n1421 252.988
R30905 vss.n1441 vss.n1411 252.988
R30906 vss.n1515 vss.n1514 252.988
R30907 vss.n1502 vss.n1501 252.988
R30908 vss.n1521 vss.n1491 252.988
R30909 vss.n957 vss.n956 252.988
R30910 vss.n944 vss.n937 252.988
R30911 vss.n963 vss.n939 252.988
R30912 vss.n1009 vss.n1008 252.988
R30913 vss.n996 vss.n989 252.988
R30914 vss.n1015 vss.n991 252.988
R30915 vss.n6247 vss.n6246 252.988
R30916 vss.n6236 vss.n6228 252.988
R30917 vss.n6238 vss.n6237 252.988
R30918 vss.n6602 vss.n6601 252.988
R30919 vss.n6607 vss.n6599 252.988
R30920 vss.n6627 vss.n6626 252.988
R30921 vss.n6375 vss.n6374 252.988
R30922 vss.n6380 vss.n6372 252.988
R30923 vss.n6400 vss.n6399 252.988
R30924 vss.n9276 vss.n9275 252.988
R30925 vss.n9265 vss.n6323 252.988
R30926 vss.n9267 vss.n9266 252.988
R30927 vss.n6911 vss.n6910 252.988
R30928 vss.n6916 vss.n6908 252.988
R30929 vss.n6936 vss.n6935 252.988
R30930 vss.n7100 vss.n7099 252.988
R30931 vss.n7105 vss.n7097 252.988
R30932 vss.n7125 vss.n7124 252.988
R30933 vss.n6285 vss.n6284 252.988
R30934 vss.n6274 vss.n6265 252.988
R30935 vss.n6276 vss.n6275 252.988
R30936 vss.n9300 vss.n9293 252.988
R30937 vss.n9312 vss.n9311 252.988
R30938 vss.n9318 vss.n6216 252.988
R30939 vss.n3318 vss.n3315 252.988
R30940 vss.n3333 vss.n3332 252.988
R30941 vss.n5887 vss.n3310 252.988
R30942 vss.n4302 vss.n4301 252.988
R30943 vss.n4313 vss.n4312 252.988
R30944 vss.n4319 vss.n4315 252.988
R30945 vss.n3657 vss.n3656 252.988
R30946 vss.n3668 vss.n3667 252.988
R30947 vss.n3674 vss.n3670 252.988
R30948 vss.n3437 vss.n3436 252.988
R30949 vss.n3448 vss.n3447 252.988
R30950 vss.n3454 vss.n3450 252.988
R30951 vss.n5875 vss.n5874 252.988
R30952 vss.n5879 vss.n2627 252.988
R30953 vss.n5877 vss.n2629 252.988
R30954 vss.n3374 vss.n3373 252.988
R30955 vss.n5855 vss.n5854 252.988
R30956 vss.n3380 vss.n3376 252.988
R30957 vss.n3959 vss.n3958 252.988
R30958 vss.n3970 vss.n3969 252.988
R30959 vss.n3976 vss.n3972 252.988
R30960 vss.n4226 vss.n4225 252.988
R30961 vss.n4237 vss.n4236 252.988
R30962 vss.n4243 vss.n4239 252.988
R30963 vss.n11335 vss.n10458 239.812
R30964 vss.n12668 vss.n10458 239.812
R30965 vss.n11331 vss.n11330 239.812
R30966 vss.n11330 vss.n10459 239.812
R30967 vss.n11088 vss.n11087 239.812
R30968 vss.n11102 vss.n11087 239.812
R30969 vss.n11094 vss.n11086 239.812
R30970 vss.n11104 vss.n11086 239.812
R30971 vss.n11090 vss.n11085 239.812
R30972 vss.n11152 vss.n11085 239.812
R30973 vss.n11163 vss.n11045 239.812
R30974 vss.n11354 vss.n11045 239.812
R30975 vss.n11160 vss.n11044 239.812
R30976 vss.n11356 vss.n11044 239.812
R30977 vss.n11170 vss.n11169 239.812
R30978 vss.n11171 vss.n11170 239.812
R30979 vss.n11214 vss.n11213 239.812
R30980 vss.n11228 vss.n11213 239.812
R30981 vss.n11220 vss.n11212 239.812
R30982 vss.n11230 vss.n11212 239.812
R30983 vss.n11216 vss.n11211 239.812
R30984 vss.n11233 vss.n11211 239.812
R30985 vss.n11275 vss.n11274 239.812
R30986 vss.n11289 vss.n11274 239.812
R30987 vss.n11281 vss.n11273 239.812
R30988 vss.n11291 vss.n11273 239.812
R30989 vss.n11277 vss.n11272 239.812
R30990 vss.n11294 vss.n11272 239.812
R30991 vss.n13026 vss.n13025 239.812
R30992 vss.n13027 vss.n13026 239.812
R30993 vss.n13040 vss.n13039 239.812
R30994 vss.n13039 vss.n13038 239.812
R30995 vss.n376 vss.n368 239.812
R30996 vss.n372 vss.n368 239.812
R30997 vss.n378 vss.n364 239.812
R30998 vss.n370 vss.n364 239.812
R30999 vss.n14763 vss.n108 239.812
R31000 vss.n110 vss.n108 239.812
R31001 vss.n119 vss.n115 239.812
R31002 vss.n14768 vss.n14765 239.812
R31003 vss.n14769 vss.n14768 239.812
R31004 vss.n392 vss.n390 239.812
R31005 vss.n397 vss.n390 239.812
R31006 vss.n386 vss.n381 239.812
R31007 vss.n399 vss.n386 239.812
R31008 vss.n408 vss.n404 239.812
R31009 vss.n269 vss.n267 239.812
R31010 vss.n274 vss.n267 239.812
R31011 vss.n263 vss.n258 239.812
R31012 vss.n276 vss.n263 239.812
R31013 vss.n285 vss.n281 239.812
R31014 vss.n14426 vss.n14424 239.812
R31015 vss.n14431 vss.n14424 239.812
R31016 vss.n14420 vss.n14415 239.812
R31017 vss.n14433 vss.n14420 239.812
R31018 vss.n14442 vss.n14438 239.812
R31019 vss.n210 vss.n208 239.812
R31020 vss.n215 vss.n208 239.812
R31021 vss.n204 vss.n199 239.812
R31022 vss.n217 vss.n204 239.812
R31023 vss.n226 vss.n222 239.812
R31024 vss.n14621 vss.n14619 239.812
R31025 vss.n14626 vss.n14619 239.812
R31026 vss.n14615 vss.n14610 239.812
R31027 vss.n14628 vss.n14615 239.812
R31028 vss.n14637 vss.n14633 239.812
R31029 vss.n133 vss.n131 239.812
R31030 vss.n138 vss.n131 239.812
R31031 vss.n127 vss.n122 239.812
R31032 vss.n140 vss.n127 239.812
R31033 vss.n149 vss.n145 239.812
R31034 vss.n14777 vss.n14776 239.812
R31035 vss.n7376 vss.n7344 239.812
R31036 vss.n7356 vss.n7344 239.812
R31037 vss.n7374 vss.n7345 239.812
R31038 vss.n7350 vss.n7345 239.812
R31039 vss.n7368 vss.n7367 239.812
R31040 vss.n7829 vss.n7828 239.812
R31041 vss.n7829 vss.n7820 239.812
R31042 vss.n7819 vss.n7812 239.812
R31043 vss.n7834 vss.n7819 239.812
R31044 vss.n7843 vss.n7814 239.812
R31045 vss.n7642 vss.n7641 239.812
R31046 vss.n7642 vss.n7633 239.812
R31047 vss.n7632 vss.n7625 239.812
R31048 vss.n7647 vss.n7632 239.812
R31049 vss.n7656 vss.n7627 239.812
R31050 vss.n7453 vss.n7452 239.812
R31051 vss.n7453 vss.n7444 239.812
R31052 vss.n7443 vss.n7436 239.812
R31053 vss.n7458 vss.n7443 239.812
R31054 vss.n7467 vss.n7438 239.812
R31055 vss.n8982 vss.n7409 239.812
R31056 vss.n7417 vss.n7409 239.812
R31057 vss.n8980 vss.n7410 239.812
R31058 vss.n7424 vss.n7410 239.812
R31059 vss.n7433 vss.n7412 239.812
R31060 vss.n7607 vss.n7606 239.812
R31061 vss.n7607 vss.n7598 239.812
R31062 vss.n7597 vss.n7590 239.812
R31063 vss.n7612 vss.n7597 239.812
R31064 vss.n7621 vss.n7592 239.812
R31065 vss.n7750 vss.n7749 239.812
R31066 vss.n7750 vss.n7741 239.812
R31067 vss.n7740 vss.n7733 239.812
R31068 vss.n7755 vss.n7740 239.812
R31069 vss.n7764 vss.n7735 239.812
R31070 vss.n7971 vss.n7970 239.812
R31071 vss.n7971 vss.n7962 239.812
R31072 vss.n7961 vss.n7954 239.812
R31073 vss.n7976 vss.n7961 239.812
R31074 vss.n7985 vss.n7956 239.812
R31075 vss.n3236 vss.n3235 239.812
R31076 vss.n3235 vss.n3234 239.812
R31077 vss.n3233 vss.n3227 239.812
R31078 vss.n3248 vss.n3233 239.812
R31079 vss.n3231 vss.n3230 239.812
R31080 vss.n3079 vss.n3078 239.812
R31081 vss.n3078 vss.n3077 239.812
R31082 vss.n3076 vss.n3070 239.812
R31083 vss.n3091 vss.n3076 239.812
R31084 vss.n3074 vss.n3073 239.812
R31085 vss.n5053 vss.n5052 239.812
R31086 vss.n5052 vss.n5051 239.812
R31087 vss.n5050 vss.n5044 239.812
R31088 vss.n5065 vss.n5050 239.812
R31089 vss.n5048 vss.n5047 239.812
R31090 vss.n2845 vss.n2844 239.812
R31091 vss.n2844 vss.n2843 239.812
R31092 vss.n2842 vss.n2836 239.812
R31093 vss.n2857 vss.n2842 239.812
R31094 vss.n2840 vss.n2839 239.812
R31095 vss.n9851 vss.n2828 239.812
R31096 vss.n9869 vss.n2828 239.812
R31097 vss.n9853 vss.n9852 239.812
R31098 vss.n9852 vss.n2829 239.812
R31099 vss.n9863 vss.n9862 239.812
R31100 vss.n4976 vss.n4975 239.812
R31101 vss.n4975 vss.n4974 239.812
R31102 vss.n4973 vss.n4967 239.812
R31103 vss.n4988 vss.n4973 239.812
R31104 vss.n4971 vss.n4970 239.812
R31105 vss.n5178 vss.n5177 239.812
R31106 vss.n5177 vss.n5176 239.812
R31107 vss.n5175 vss.n5169 239.812
R31108 vss.n5190 vss.n5175 239.812
R31109 vss.n5173 vss.n5172 239.812
R31110 vss.n3159 vss.n3158 239.812
R31111 vss.n3158 vss.n3157 239.812
R31112 vss.n3156 vss.n3150 239.812
R31113 vss.n3171 vss.n3156 239.812
R31114 vss.n3154 vss.n3153 239.812
R31115 vss.n10195 vss.n10194 239.812
R31116 vss.n10194 vss.n10193 239.812
R31117 vss.n10192 vss.n10186 239.812
R31118 vss.n10207 vss.n10192 239.812
R31119 vss.n10189 vss.n10187 239.812
R31120 vss.n10190 vss.n10189 239.812
R31121 vss.n12506 vss.n12505 239.812
R31122 vss.n12505 vss.n12504 239.812
R31123 vss.n12503 vss.n12497 239.812
R31124 vss.n12518 vss.n12503 239.812
R31125 vss.n12500 vss.n12498 239.812
R31126 vss.n12501 vss.n12500 239.812
R31127 vss.n2214 vss.n2213 239.812
R31128 vss.n2213 vss.n2212 239.812
R31129 vss.n2211 vss.n2205 239.812
R31130 vss.n2226 vss.n2211 239.812
R31131 vss.n2208 vss.n2206 239.812
R31132 vss.n2209 vss.n2208 239.812
R31133 vss.n12377 vss.n12376 239.812
R31134 vss.n12376 vss.n12375 239.812
R31135 vss.n12374 vss.n12368 239.812
R31136 vss.n12389 vss.n12374 239.812
R31137 vss.n12371 vss.n12369 239.812
R31138 vss.n12372 vss.n12371 239.812
R31139 vss.n10273 vss.n10272 239.812
R31140 vss.n10272 vss.n10271 239.812
R31141 vss.n10270 vss.n10264 239.812
R31142 vss.n10285 vss.n10270 239.812
R31143 vss.n10267 vss.n10265 239.812
R31144 vss.n10268 vss.n10267 239.812
R31145 vss.n2453 vss.n2452 239.812
R31146 vss.n2452 vss.n2451 239.812
R31147 vss.n2450 vss.n2444 239.812
R31148 vss.n2465 vss.n2450 239.812
R31149 vss.n2447 vss.n2445 239.812
R31150 vss.n2448 vss.n2447 239.812
R31151 vss.n2532 vss.n2531 239.812
R31152 vss.n2531 vss.n2530 239.812
R31153 vss.n2529 vss.n2523 239.812
R31154 vss.n2544 vss.n2529 239.812
R31155 vss.n2526 vss.n2524 239.812
R31156 vss.n2527 vss.n2526 239.812
R31157 vss.n13046 vss.n2202 239.812
R31158 vss.n2204 vss.n2202 239.812
R31159 vss.n11315 vss.n11306 239.812
R31160 vss.n11310 vss.n11306 239.812
R31161 vss.n11307 vss.n11303 239.812
R31162 vss.n11308 vss.n11307 239.812
R31163 vss.n11322 vss.n11321 239.812
R31164 vss.n11324 vss.n11322 239.812
R31165 vss.n11254 vss.n11245 239.812
R31166 vss.n11249 vss.n11245 239.812
R31167 vss.n11246 vss.n11242 239.812
R31168 vss.n11247 vss.n11246 239.812
R31169 vss.n11261 vss.n11260 239.812
R31170 vss.n11263 vss.n11261 239.812
R31171 vss.n11183 vss.n11182 239.812
R31172 vss.n11197 vss.n11182 239.812
R31173 vss.n11189 vss.n11181 239.812
R31174 vss.n11199 vss.n11181 239.812
R31175 vss.n11185 vss.n11180 239.812
R31176 vss.n11202 vss.n11180 239.812
R31177 vss.n11348 vss.n11341 239.812
R31178 vss.n11348 vss.n11347 239.812
R31179 vss.n8152 vss.t1219 231.517
R31180 vss.t1387 vss.n3282 231.517
R31181 vss.t1387 vss.n3275 231.517
R31182 vss.t1199 vss.n3275 231.517
R31183 vss.t1199 vss.n3268 231.517
R31184 vss.t1197 vss.n3268 231.517
R31185 vss.t49 vss.n3296 231.517
R31186 vss.t49 vss.n2742 231.517
R31187 vss.t293 vss.n14155 231.517
R31188 vss.t293 vss.n451 231.517
R31189 vss.t972 vss.n451 231.517
R31190 vss.t972 vss.n441 231.517
R31191 vss.t973 vss.n441 231.517
R31192 vss.n444 vss.t880 231.517
R31193 vss.n14175 vss.t880 231.517
R31194 vss.n10041 vss.t1087 231.517
R31195 vss.n3296 vss.n3269 223.119
R31196 vss.n444 vss.n442 223.119
R31197 vss.n8174 vss.n8099 219.322
R31198 vss.n8174 vss.t960 217.061
R31199 vss.n9703 vss.n2591 208.036
R31200 vss.n9649 vss.n9648 193.368
R31201 vss.n13093 vss.n13092 193.368
R31202 vss.n12060 vss.n12059 189.903
R31203 vss.n10671 vss.n10670 189.903
R31204 vss.n11495 vss.n11494 189.903
R31205 vss.n12725 vss.n12724 189.903
R31206 vss.n13898 vss.n13897 189.903
R31207 vss.n13793 vss.n13792 189.903
R31208 vss.n13688 vss.n13687 189.903
R31209 vss.n13583 vss.n13582 189.903
R31210 vss.n14002 vss.n14001 189.903
R31211 vss.n1728 vss.n1727 189.903
R31212 vss.n1832 vss.n1831 189.903
R31213 vss.n1954 vss.n1953 189.903
R31214 vss.n8304 vss.n8303 189.903
R31215 vss.n8631 vss.n8630 189.903
R31216 vss.n8544 vss.n8543 189.903
R31217 vss.n9551 vss.n9550 189.903
R31218 vss.n6764 vss.n6763 189.903
R31219 vss.n6893 vss.n6892 189.903
R31220 vss.n9082 vss.n9081 189.903
R31221 vss.n9910 vss.n9909 189.903
R31222 vss.n5569 vss.n5568 189.903
R31223 vss.n5483 vss.n5482 189.903
R31224 vss.n5397 vss.n5396 189.903
R31225 vss.n4536 vss.n4535 189.903
R31226 vss.n4184 vss.n4183 189.903
R31227 vss.n3936 vss.n3935 189.903
R31228 vss.n5676 vss.n5675 189.903
R31229 vss.n12123 vss.n12122 189.903
R31230 vss.n12227 vss.n12226 189.903
R31231 vss.n11662 vss.n11661 189.903
R31232 vss.n12943 vss.n12942 189.903
R31233 vss.t718 vss.n14114 188.209
R31234 vss.t718 vss.n14108 188.209
R31235 vss.t1224 vss.n14108 188.209
R31236 vss.t1224 vss.n14101 188.209
R31237 vss.t1225 vss.n14101 188.209
R31238 vss.t1225 vss.n14102 188.209
R31239 vss.t393 vss.n14102 188.209
R31240 vss.t393 vss.n26 188.209
R31241 vss.n8051 vss.t94 188.209
R31242 vss.t94 vss.n8012 188.209
R31243 vss.t1528 vss.n8012 188.209
R31244 vss.t1528 vss.n8019 188.209
R31245 vss.t1529 vss.n8019 188.209
R31246 vss.n8027 vss.t1529 188.209
R31247 vss.n8027 vss.t635 188.209
R31248 vss.t635 vss.n7323 188.209
R31249 vss.n9895 vss.t322 188.209
R31250 vss.n2751 vss.t322 188.209
R31251 vss.t129 vss.n2751 188.209
R31252 vss.t129 vss.n2752 188.209
R31253 vss.t130 vss.n2752 188.209
R31254 vss.t130 vss.n9883 188.209
R31255 vss.n9883 vss.t217 188.209
R31256 vss.n9876 vss.t217 188.209
R31257 vss.n13076 vss.t1149 188.209
R31258 vss.n2127 vss.t1149 188.209
R31259 vss.t854 vss.n2127 188.209
R31260 vss.t854 vss.n2128 188.209
R31261 vss.t855 vss.n2128 188.209
R31262 vss.t855 vss.n13064 188.209
R31263 vss.n13064 vss.t619 188.209
R31264 vss.n13057 vss.t619 188.209
R31265 vss.n13301 vss.t1412 186.228
R31266 vss.t351 vss.n9050 186.228
R31267 vss.t688 vss.n5644 186.228
R31268 vss.n12097 vss.t530 186.228
R31269 vss.n9648 vss.t1219 184.733
R31270 vss.n13092 vss.t1087 184.733
R31271 vss.n12672 vss.n10410 183.912
R31272 vss.n13136 vss.n2049 183.912
R31273 vss.n12673 vss.n12672 183.912
R31274 vss.n13117 vss.n2068 183.912
R31275 vss.n12672 vss.n10411 183.912
R31276 vss.n13120 vss.n2065 183.912
R31277 vss.n12672 vss.n10412 183.912
R31278 vss.n13118 vss.n2067 183.912
R31279 vss.n12672 vss.n10413 183.912
R31280 vss.n13123 vss.n2062 183.912
R31281 vss.n12672 vss.n10414 183.912
R31282 vss.n13126 vss.n2059 183.912
R31283 vss.n12672 vss.n10415 183.912
R31284 vss.n13124 vss.n2061 183.912
R31285 vss.n12672 vss.n10416 183.912
R31286 vss.n13129 vss.n2056 183.912
R31287 vss.n12672 vss.n10417 183.912
R31288 vss.n13132 vss.n2053 183.912
R31289 vss.n12672 vss.n10418 183.912
R31290 vss.n13130 vss.n2055 183.912
R31291 vss.n12672 vss.n10419 183.912
R31292 vss.n13135 vss.n2050 183.912
R31293 vss.n12008 vss.n12007 183.912
R31294 vss.n12600 vss.n12599 183.912
R31295 vss.n10858 vss.n10857 183.912
R31296 vss.n11529 vss.n11528 183.912
R31297 vss.n10928 vss.n10927 183.912
R31298 vss.n12756 vss.n12755 183.912
R31299 vss.n2304 vss.n2303 183.912
R31300 vss.n13056 vss.n2143 183.912
R31301 vss.n12994 vss.n12993 183.912
R31302 vss.n13056 vss.n2144 183.912
R31303 vss.n13873 vss.n13872 183.912
R31304 vss.n13844 vss.n13843 183.912
R31305 vss.n13768 vss.n13767 183.912
R31306 vss.n13739 vss.n13738 183.912
R31307 vss.n13663 vss.n13662 183.912
R31308 vss.n13634 vss.n13633 183.912
R31309 vss.n14732 vss.n14731 183.912
R31310 vss.n14783 vss.n19 183.912
R31311 vss.n14684 vss.n14683 183.912
R31312 vss.n14783 vss.n20 183.912
R31313 vss.n14537 vss.n14536 183.912
R31314 vss.n14783 vss.n21 183.912
R31315 vss.n14489 vss.n14488 183.912
R31316 vss.n14783 vss.n22 183.912
R31317 vss.n14342 vss.n14341 183.912
R31318 vss.n14783 vss.n23 183.912
R31319 vss.n14294 vss.n14293 183.912
R31320 vss.n14783 vss.n24 183.912
R31321 vss.n14223 vss.n14222 183.912
R31322 vss.n14783 vss.n25 183.912
R31323 vss.n14221 vss.n14220 183.912
R31324 vss.n14783 vss.n27 183.912
R31325 vss.n335 vss.n311 183.912
R31326 vss.n14783 vss.n28 183.912
R31327 vss.n14340 vss.n14339 183.912
R31328 vss.n14783 vss.n29 183.912
R31329 vss.n14388 vss.n252 183.912
R31330 vss.n14783 vss.n30 183.912
R31331 vss.n14535 vss.n14534 183.912
R31332 vss.n14783 vss.n31 183.912
R31333 vss.n14583 vss.n193 183.912
R31334 vss.n14783 vss.n32 183.912
R31335 vss.n14730 vss.n14729 183.912
R31336 vss.n14783 vss.n33 183.912
R31337 vss.n190 vss.n189 183.912
R31338 vss.n14784 vss.n14783 183.912
R31339 vss.n667 vss.n666 183.912
R31340 vss.n13967 vss.n13966 183.912
R31341 vss.n1750 vss.n1749 183.912
R31342 vss.n1779 vss.n1778 183.912
R31343 vss.n1854 vss.n1853 183.912
R31344 vss.n1883 vss.n1882 183.912
R31345 vss.n13210 vss.n813 183.912
R31346 vss.n13263 vss.n730 183.912
R31347 vss.n13210 vss.n814 183.912
R31348 vss.n13260 vss.n733 183.912
R31349 vss.n13210 vss.n815 183.912
R31350 vss.n13257 vss.n736 183.912
R31351 vss.n13210 vss.n816 183.912
R31352 vss.n13254 vss.n739 183.912
R31353 vss.n13211 vss.n13210 183.912
R31354 vss.n13251 vss.n742 183.912
R31355 vss.n13210 vss.n833 183.912
R31356 vss.n13943 vss.n13942 183.912
R31357 vss.n13210 vss.n874 183.912
R31358 vss.n13939 vss.n613 183.912
R31359 vss.n13210 vss.n918 183.912
R31360 vss.n13940 vss.n612 183.912
R31361 vss.n13210 vss.n919 183.912
R31362 vss.n1555 vss.n611 183.912
R31363 vss.n13210 vss.n920 183.912
R31364 vss.n13252 vss.n741 183.912
R31365 vss.n13210 vss.n921 183.912
R31366 vss.n13255 vss.n738 183.912
R31367 vss.n13210 vss.n922 183.912
R31368 vss.n13258 vss.n735 183.912
R31369 vss.n13210 vss.n923 183.912
R31370 vss.n13261 vss.n732 183.912
R31371 vss.n13210 vss.n924 183.912
R31372 vss.n13264 vss.n729 183.912
R31373 vss.n9018 vss.n9017 183.912
R31374 vss.n8283 vss.n8282 183.912
R31375 vss.n8674 vss.n8673 183.912
R31376 vss.n8646 vss.n8645 183.912
R31377 vss.n8587 vss.n8586 183.912
R31378 vss.n8559 vss.n8558 183.912
R31379 vss.n7255 vss.n7254 183.912
R31380 vss.n9516 vss.n9515 183.912
R31381 vss.n6786 vss.n6785 183.912
R31382 vss.n7061 vss.n7060 183.912
R31383 vss.n6879 vss.n6878 183.912
R31384 vss.n9224 vss.n9223 183.912
R31385 vss.n9168 vss.n5971 183.912
R31386 vss.n9385 vss.n6182 183.912
R31387 vss.n6465 vss.n5971 183.912
R31388 vss.n9388 vss.n6179 183.912
R31389 vss.n7005 vss.n5971 183.912
R31390 vss.n9391 vss.n6176 183.912
R31391 vss.n6691 vss.n5971 183.912
R31392 vss.n9394 vss.n6173 183.912
R31393 vss.n7196 vss.n5971 183.912
R31394 vss.n9397 vss.n6170 183.912
R31395 vss.n6153 vss.n5971 183.912
R31396 vss.n9492 vss.n9491 183.912
R31397 vss.n9462 vss.n5971 183.912
R31398 vss.n9488 vss.n9486 183.912
R31399 vss.n6026 vss.n5971 183.912
R31400 vss.n6041 vss.n5972 183.912
R31401 vss.n9418 vss.n5971 183.912
R31402 vss.n9489 vss.n9444 183.912
R31403 vss.n7145 vss.n5971 183.912
R31404 vss.n9399 vss.n6168 183.912
R31405 vss.n6647 vss.n5971 183.912
R31406 vss.n9396 vss.n6171 183.912
R31407 vss.n6956 vss.n5971 183.912
R31408 vss.n9393 vss.n6174 183.912
R31409 vss.n6420 vss.n5971 183.912
R31410 vss.n9390 vss.n6177 183.912
R31411 vss.n6342 vss.n5971 183.912
R31412 vss.n9387 vss.n6180 183.912
R31413 vss.n9338 vss.n5971 183.912
R31414 vss.n9384 vss.n6183 183.912
R31415 vss.n9899 vss.n2740 183.912
R31416 vss.n9875 vss.n2768 183.912
R31417 vss.n9898 vss.n2741 183.912
R31418 vss.n9875 vss.n2769 183.912
R31419 vss.n9803 vss.n9802 183.912
R31420 vss.n9875 vss.n2770 183.912
R31421 vss.n9806 vss.n2990 183.912
R31422 vss.n9875 vss.n2771 183.912
R31423 vss.n9805 vss.n2991 183.912
R31424 vss.n9875 vss.n2772 183.912
R31425 vss.n9809 vss.n2987 183.912
R31426 vss.n9875 vss.n2773 183.912
R31427 vss.n9812 vss.n2984 183.912
R31428 vss.n9875 vss.n2774 183.912
R31429 vss.n9811 vss.n2985 183.912
R31430 vss.n9875 vss.n2775 183.912
R31431 vss.n9815 vss.n2981 183.912
R31432 vss.n9875 vss.n2776 183.912
R31433 vss.n5612 vss.n5611 183.912
R31434 vss.n5584 vss.n5583 183.912
R31435 vss.n5526 vss.n5525 183.912
R31436 vss.n5498 vss.n5497 183.912
R31437 vss.n5440 vss.n5439 183.912
R31438 vss.n5412 vss.n5411 183.912
R31439 vss.n9819 vss.n9818 183.912
R31440 vss.n9875 vss.n2777 183.912
R31441 vss.n9817 vss.n2979 183.912
R31442 vss.n9875 vss.n2778 183.912
R31443 vss.n2934 vss.n2933 183.912
R31444 vss.n9875 vss.n2779 183.912
R31445 vss.n9814 vss.n2982 183.912
R31446 vss.n9875 vss.n2780 183.912
R31447 vss.n9808 vss.n2988 183.912
R31448 vss.n9875 vss.n2781 183.912
R31449 vss.n3122 vss.n2739 183.912
R31450 vss.n9875 vss.n2782 183.912
R31451 vss.n4480 vss.n2600 183.912
R31452 vss.n9934 vss.n2703 183.912
R31453 vss.n4388 vss.n2600 183.912
R31454 vss.n9937 vss.n2700 183.912
R31455 vss.n4340 vss.n2600 183.912
R31456 vss.n9935 vss.n2702 183.912
R31457 vss.n3740 vss.n2600 183.912
R31458 vss.n9940 vss.n2697 183.912
R31459 vss.n4042 vss.n2600 183.912
R31460 vss.n9943 vss.n2694 183.912
R31461 vss.n3695 vss.n2600 183.912
R31462 vss.n9941 vss.n2696 183.912
R31463 vss.n4096 vss.n2600 183.912
R31464 vss.n9946 vss.n2691 183.912
R31465 vss.n3520 vss.n2600 183.912
R31466 vss.n9949 vss.n2688 183.912
R31467 vss.n3475 vss.n2600 183.912
R31468 vss.n9947 vss.n2690 183.912
R31469 vss.n5763 vss.n2600 183.912
R31470 vss.n9952 vss.n2685 183.912
R31471 vss.n4558 vss.n4557 183.912
R31472 vss.n4587 vss.n4586 183.912
R31473 vss.n3828 vss.n3827 183.912
R31474 vss.n4149 vss.n4148 183.912
R31475 vss.n3922 vss.n3921 183.912
R31476 vss.n5816 vss.n5815 183.912
R31477 vss.n2662 vss.n2600 183.912
R31478 vss.n9953 vss.n2684 183.912
R31479 vss.n3400 vss.n2600 183.912
R31480 vss.n9950 vss.n2687 183.912
R31481 vss.n3997 vss.n2600 183.912
R31482 vss.n9944 vss.n2693 183.912
R31483 vss.n4264 vss.n2600 183.912
R31484 vss.n9938 vss.n2699 183.912
R31485 vss.n5907 vss.n2600 183.912
R31486 vss.n9932 vss.n2705 183.912
R31487 vss.n8950 vss.n8949 183.912
R31488 vss.n8986 vss.n7325 183.912
R31489 vss.n8902 vss.n8901 183.912
R31490 vss.n8986 vss.n7326 183.912
R31491 vss.n8831 vss.n8830 183.912
R31492 vss.n8986 vss.n7327 183.912
R31493 vss.n8783 vss.n8782 183.912
R31494 vss.n8986 vss.n7328 183.912
R31495 vss.n8712 vss.n8711 183.912
R31496 vss.n8986 vss.n7329 183.912
R31497 vss.n9007 vss.n9006 183.912
R31498 vss.n8987 vss.n8986 183.912
R31499 vss.n8221 vss.n8220 183.912
R31500 vss.n8986 vss.n7330 183.912
R31501 vss.n8986 vss.n7331 183.912
R31502 vss.n7927 vss.n7299 183.912
R31503 vss.n8986 vss.n7333 183.912
R31504 vss.n7786 vss.n7298 183.912
R31505 vss.n8986 vss.n7334 183.912
R31506 vss.n7706 vss.n7682 183.912
R31507 vss.n8986 vss.n7335 183.912
R31508 vss.n8829 vss.n8828 183.912
R31509 vss.n8986 vss.n7336 183.912
R31510 vss.n7563 vss.n7539 183.912
R31511 vss.n8986 vss.n7337 183.912
R31512 vss.n8948 vss.n8947 183.912
R31513 vss.n8986 vss.n7338 183.912
R31514 vss.n7536 vss.n7535 183.912
R31515 vss.n8986 vss.n7339 183.912
R31516 vss.n13937 vss.n658 183.912
R31517 vss.n12978 vss.n2363 183.912
R31518 vss.n13056 vss.n2146 183.912
R31519 vss.n12981 vss.n2360 183.912
R31520 vss.n13056 vss.n2147 183.912
R31521 vss.n12980 vss.n2361 183.912
R31522 vss.n13056 vss.n2148 183.912
R31523 vss.n12984 vss.n2357 183.912
R31524 vss.n13056 vss.n2149 183.912
R31525 vss.n12987 vss.n2354 183.912
R31526 vss.n13056 vss.n2150 183.912
R31527 vss.n12986 vss.n2355 183.912
R31528 vss.n13056 vss.n2151 183.912
R31529 vss.n12992 vss.n2349 183.912
R31530 vss.n13056 vss.n2152 183.912
R31531 vss.n12990 vss.n2351 183.912
R31532 vss.n13056 vss.n2153 183.912
R31533 vss.n12989 vss.n2352 183.912
R31534 vss.n13056 vss.n2154 183.912
R31535 vss.n12983 vss.n2358 183.912
R31536 vss.n13056 vss.n2155 183.912
R31537 vss.n12977 vss.n2364 183.912
R31538 vss.n13056 vss.n2156 183.912
R31539 vss.n12975 vss.n12974 183.912
R31540 vss.n13056 vss.n2157 183.912
R31541 vss.n2496 vss.n2119 183.912
R31542 vss.n13056 vss.n2158 183.912
R31543 vss.n12153 vss.n12152 183.912
R31544 vss.n12176 vss.n12175 183.912
R31545 vss.n12549 vss.n12548 183.912
R31546 vss.n12572 vss.n12571 183.912
R31547 vss.n12831 vss.n12830 183.912
R31548 vss.n12809 vss.n12808 183.912
R31549 vss.n12672 vss.n10420 183.912
R31550 vss.n13133 vss.n2052 183.912
R31551 vss.n12672 vss.n10421 183.912
R31552 vss.n13127 vss.n2058 183.912
R31553 vss.n12672 vss.n10422 183.912
R31554 vss.n13121 vss.n2064 183.912
R31555 vss.n12672 vss.n10423 183.912
R31556 vss.n13115 vss.n2070 183.912
R31557 vss.n12045 vss.n12044 178.287
R31558 vss.n11613 vss.n11612 178.287
R31559 vss.n11480 vss.n11479 178.287
R31560 vss.n13819 vss.n13818 178.287
R31561 vss.n13714 vss.n13713 178.287
R31562 vss.n13609 vss.n13608 178.287
R31563 vss.n779 vss.n778 178.287
R31564 vss.n1821 vss.n1820 178.287
R31565 vss.n1925 vss.n1924 178.287
R31566 vss.n8689 vss.n8688 178.287
R31567 vss.n8602 vss.n8601 178.287
R31568 vss.n7236 vss.n7235 178.287
R31569 vss.n7045 vss.n7044 178.287
R31570 vss.n9208 vss.n9207 178.287
R31571 vss.n4667 vss.n4666 178.287
R31572 vss.n5541 vss.n5540 178.287
R31573 vss.n5455 vss.n5454 178.287
R31574 vss.n3772 vss.n3771 178.287
R31575 vss.n4135 vss.n4134 178.287
R31576 vss.n5802 vss.n5801 178.287
R31577 vss.n8079 vss.n8078 178.287
R31578 vss.n12251 vss.n12250 178.287
R31579 vss.n11686 vss.n11685 178.287
R31580 vss.n12922 vss.n12921 178.287
R31581 vss.n9647 vss.t691 154.065
R31582 vss.n8129 vss.t691 154.065
R31583 vss.t689 vss.n8129 154.065
R31584 vss.t689 vss.n8130 154.065
R31585 vss.t1005 vss.n8130 154.065
R31586 vss.t1005 vss.n8052 154.065
R31587 vss.n13091 vss.t678 154.065
R31588 vss.n2104 vss.t678 154.065
R31589 vss.t676 vss.n2104 154.065
R31590 vss.t676 vss.n2105 154.065
R31591 vss.t53 vss.n2105 154.065
R31592 vss.t53 vss.n13078 154.065
R31593 vss.t1061 vss.n8123 153.452
R31594 vss.n9929 vss.t339 153.452
R31595 vss.t1275 vss.n458 153.452
R31596 vss.t318 vss.n10035 153.452
R31597 vss.n11154 vss.n11084 146.834
R31598 vss.n11100 vss.n11099 146.834
R31599 vss.n11173 vss.n11159 146.834
R31600 vss.n11352 vss.n11046 146.834
R31601 vss.n11235 vss.n11210 146.834
R31602 vss.n11226 vss.n11225 146.834
R31603 vss.n11296 vss.n11271 146.834
R31604 vss.n11287 vss.n11286 146.834
R31605 vss.n114 vss.n113 146.834
R31606 vss.n14770 vss.n102 146.834
R31607 vss.n403 vss.n402 146.834
R31608 vss.n396 vss.n395 146.834
R31609 vss.n280 vss.n279 146.834
R31610 vss.n273 vss.n272 146.834
R31611 vss.n14437 vss.n14436 146.834
R31612 vss.n14430 vss.n14429 146.834
R31613 vss.n221 vss.n220 146.834
R31614 vss.n214 vss.n213 146.834
R31615 vss.n14632 vss.n14631 146.834
R31616 vss.n14625 vss.n14624 146.834
R31617 vss.n144 vss.n143 146.834
R31618 vss.n137 vss.n136 146.834
R31619 vss.n14779 vss.n14778 146.834
R31620 vss.n374 vss.n373 146.834
R31621 vss.n14043 vss.n14042 146.834
R31622 vss.n14057 vss.n505 146.834
R31623 vss.n1592 vss.n1589 146.834
R31624 vss.n1579 vss.n1576 146.834
R31625 vss.n1297 vss.n1294 146.834
R31626 vss.n1284 vss.n1281 146.834
R31627 vss.n1036 vss.n1033 146.834
R31628 vss.n1023 vss.n1020 146.834
R31629 vss.n1429 vss.n1426 146.834
R31630 vss.n1416 vss.n1413 146.834
R31631 vss.n1509 vss.n1506 146.834
R31632 vss.n1496 vss.n1493 146.834
R31633 vss.n951 vss.n948 146.834
R31634 vss.n943 vss.n936 146.834
R31635 vss.n1003 vss.n1000 146.834
R31636 vss.n995 vss.n988 146.834
R31637 vss.n7366 vss.n7363 146.834
R31638 vss.n7355 vss.n7343 146.834
R31639 vss.n7839 vss.n7838 146.834
R31640 vss.n7825 vss.n7823 146.834
R31641 vss.n7652 vss.n7651 146.834
R31642 vss.n7638 vss.n7636 146.834
R31643 vss.n7463 vss.n7462 146.834
R31644 vss.n7449 vss.n7447 146.834
R31645 vss.n7429 vss.n7428 146.834
R31646 vss.n7418 vss.n7408 146.834
R31647 vss.n7617 vss.n7616 146.834
R31648 vss.n7603 vss.n7601 146.834
R31649 vss.n7760 vss.n7759 146.834
R31650 vss.n7746 vss.n7744 146.834
R31651 vss.n7981 vss.n7980 146.834
R31652 vss.n7967 vss.n7965 146.834
R31653 vss.n6245 vss.n6234 146.834
R31654 vss.n6256 vss.n6227 146.834
R31655 vss.n6619 vss.n6618 146.834
R31656 vss.n6606 vss.n6605 146.834
R31657 vss.n6392 vss.n6391 146.834
R31658 vss.n6379 vss.n6378 146.834
R31659 vss.n9274 vss.n9263 146.834
R31660 vss.n9285 vss.n6322 146.834
R31661 vss.n6928 vss.n6927 146.834
R31662 vss.n6915 vss.n6914 146.834
R31663 vss.n7117 vss.n7116 146.834
R31664 vss.n7104 vss.n7103 146.834
R31665 vss.n6283 vss.n6272 146.834
R31666 vss.n6294 vss.n6264 146.834
R31667 vss.n9297 vss.n9296 146.834
R31668 vss.n9315 vss.n9307 146.834
R31669 vss.n3322 vss.n3321 146.834
R31670 vss.n3334 vss.n3326 146.834
R31671 vss.n3254 vss.n3253 146.834
R31672 vss.n3243 vss.n3242 146.834
R31673 vss.n3097 vss.n3096 146.834
R31674 vss.n3086 vss.n3085 146.834
R31675 vss.n5071 vss.n5070 146.834
R31676 vss.n5060 vss.n5059 146.834
R31677 vss.n2863 vss.n2862 146.834
R31678 vss.n2852 vss.n2851 146.834
R31679 vss.n2834 vss.n2833 146.834
R31680 vss.n9871 vss.n9870 146.834
R31681 vss.n4994 vss.n4993 146.834
R31682 vss.n4983 vss.n4982 146.834
R31683 vss.n5196 vss.n5195 146.834
R31684 vss.n5185 vss.n5184 146.834
R31685 vss.n3177 vss.n3176 146.834
R31686 vss.n3166 vss.n3165 146.834
R31687 vss.n4295 vss.n4293 146.834
R31688 vss.n4306 vss.n4304 146.834
R31689 vss.n3650 vss.n3648 146.834
R31690 vss.n3661 vss.n3659 146.834
R31691 vss.n3430 vss.n3428 146.834
R31692 vss.n3441 vss.n3439 146.834
R31693 vss.n5868 vss.n5866 146.834
R31694 vss.n5880 vss.n2626 146.834
R31695 vss.n3367 vss.n3365 146.834
R31696 vss.n5856 vss.n3361 146.834
R31697 vss.n3952 vss.n3950 146.834
R31698 vss.n3963 vss.n3961 146.834
R31699 vss.n4219 vss.n4217 146.834
R31700 vss.n4230 vss.n4228 146.834
R31701 vss.n10202 vss.n10201 146.834
R31702 vss.n10213 vss.n10212 146.834
R31703 vss.n12513 vss.n12512 146.834
R31704 vss.n12524 vss.n12523 146.834
R31705 vss.n2221 vss.n2220 146.834
R31706 vss.n2232 vss.n2231 146.834
R31707 vss.n12384 vss.n12383 146.834
R31708 vss.n12395 vss.n12394 146.834
R31709 vss.n10280 vss.n10279 146.834
R31710 vss.n10291 vss.n10290 146.834
R31711 vss.n2460 vss.n2459 146.834
R31712 vss.n2471 vss.n2470 146.834
R31713 vss.n2539 vss.n2538 146.834
R31714 vss.n2550 vss.n2549 146.834
R31715 vss.n13031 vss.n13030 146.834
R31716 vss.n13050 vss.n13049 146.834
R31717 vss.n11326 vss.n11302 146.834
R31718 vss.n11314 vss.n11312 146.834
R31719 vss.n11265 vss.n11241 146.834
R31720 vss.n11253 vss.n11251 146.834
R31721 vss.n11204 vss.n11179 146.834
R31722 vss.n11195 vss.n11194 146.834
R31723 vss.n11334 vss.n10457 146.834
R31724 vss.n11345 vss.n11344 146.834
R31725 vss.n113 vss.n109 141.34
R31726 vss.n402 vss.n382 141.34
R31727 vss.n279 vss.n259 141.34
R31728 vss.n14436 vss.n14416 141.34
R31729 vss.n220 vss.n200 141.34
R31730 vss.n14631 vss.n14611 141.34
R31731 vss.n143 vss.n123 141.34
R31732 vss.n14779 vss.n66 141.34
R31733 vss.n14042 vss.n14035 141.34
R31734 vss.n508 vss.n505 141.34
R31735 vss.n1593 vss.n1592 141.34
R31736 vss.n1580 vss.n1579 141.34
R31737 vss.n1298 vss.n1297 141.34
R31738 vss.n1285 vss.n1284 141.34
R31739 vss.n1037 vss.n1036 141.34
R31740 vss.n1024 vss.n1023 141.34
R31741 vss.n1430 vss.n1429 141.34
R31742 vss.n1417 vss.n1416 141.34
R31743 vss.n1510 vss.n1509 141.34
R31744 vss.n1497 vss.n1496 141.34
R31745 vss.n952 vss.n951 141.34
R31746 vss.n967 vss.n936 141.34
R31747 vss.n1004 vss.n1003 141.34
R31748 vss.n13207 vss.n988 141.34
R31749 vss.n7363 vss.n7362 141.34
R31750 vss.n7838 vss.n7813 141.34
R31751 vss.n7651 vss.n7626 141.34
R31752 vss.n7462 vss.n7437 141.34
R31753 vss.n7428 vss.n7411 141.34
R31754 vss.n7616 vss.n7591 141.34
R31755 vss.n7759 vss.n7734 141.34
R31756 vss.n7980 vss.n7955 141.34
R31757 vss.n6234 vss.n6232 141.34
R31758 vss.n6256 vss.n6255 141.34
R31759 vss.n6618 vss.n6617 141.34
R31760 vss.n6609 vss.n6606 141.34
R31761 vss.n6391 vss.n6390 141.34
R31762 vss.n6382 vss.n6379 141.34
R31763 vss.n9263 vss.n9261 141.34
R31764 vss.n9285 vss.n9284 141.34
R31765 vss.n6927 vss.n6926 141.34
R31766 vss.n6918 vss.n6915 141.34
R31767 vss.n7116 vss.n7115 141.34
R31768 vss.n7107 vss.n7104 141.34
R31769 vss.n6272 vss.n6270 141.34
R31770 vss.n6294 vss.n6293 141.34
R31771 vss.n9298 vss.n9297 141.34
R31772 vss.n9315 vss.n9314 141.34
R31773 vss.n3321 vss.n3320 141.34
R31774 vss.n3328 vss.n3326 141.34
R31775 vss.n3255 vss.n3254 141.34
R31776 vss.n3098 vss.n3097 141.34
R31777 vss.n5072 vss.n5071 141.34
R31778 vss.n2864 vss.n2863 141.34
R31779 vss.n2835 vss.n2834 141.34
R31780 vss.n4995 vss.n4994 141.34
R31781 vss.n5197 vss.n5196 141.34
R31782 vss.n3178 vss.n3177 141.34
R31783 vss.n4296 vss.n4295 141.34
R31784 vss.n4307 vss.n4306 141.34
R31785 vss.n3651 vss.n3650 141.34
R31786 vss.n3662 vss.n3661 141.34
R31787 vss.n3431 vss.n3430 141.34
R31788 vss.n3442 vss.n3441 141.34
R31789 vss.n5869 vss.n5868 141.34
R31790 vss.n9997 vss.n2626 141.34
R31791 vss.n3368 vss.n3367 141.34
R31792 vss.n3363 vss.n3361 141.34
R31793 vss.n3953 vss.n3952 141.34
R31794 vss.n3964 vss.n3963 141.34
R31795 vss.n4220 vss.n4219 141.34
R31796 vss.n4231 vss.n4230 141.34
R31797 vss.n10214 vss.n10213 141.34
R31798 vss.n12525 vss.n12524 141.34
R31799 vss.n2233 vss.n2232 141.34
R31800 vss.n12396 vss.n12395 141.34
R31801 vss.n10292 vss.n10291 141.34
R31802 vss.n2472 vss.n2471 141.34
R31803 vss.n2551 vss.n2550 141.34
R31804 vss.n13049 vss.n13048 141.34
R31805 vss.n12672 vss.n10409 137.662
R31806 vss.n13210 vss.n812 137.662
R31807 vss.n6203 vss.n5971 137.662
R31808 vss.n9967 vss.n2600 137.662
R31809 vss.n11154 vss.n11153 133.615
R31810 vss.n11101 vss.n11100 133.615
R31811 vss.n11173 vss.n11172 133.615
R31812 vss.n11353 vss.n11352 133.615
R31813 vss.n11235 vss.n11234 133.615
R31814 vss.n11227 vss.n11226 133.615
R31815 vss.n11296 vss.n11295 133.615
R31816 vss.n11288 vss.n11287 133.615
R31817 vss.n104 vss.n102 133.615
R31818 vss.n395 vss.n393 133.615
R31819 vss.n272 vss.n270 133.615
R31820 vss.n14429 vss.n14427 133.615
R31821 vss.n213 vss.n211 133.615
R31822 vss.n14624 vss.n14622 133.615
R31823 vss.n136 vss.n134 133.615
R31824 vss.n375 vss.n374 133.615
R31825 vss.n7377 vss.n7343 133.615
R31826 vss.n7826 vss.n7825 133.615
R31827 vss.n7639 vss.n7638 133.615
R31828 vss.n7450 vss.n7449 133.615
R31829 vss.n8983 vss.n7408 133.615
R31830 vss.n7604 vss.n7603 133.615
R31831 vss.n7747 vss.n7746 133.615
R31832 vss.n7968 vss.n7967 133.615
R31833 vss.n3242 vss.n3241 133.615
R31834 vss.n3085 vss.n3084 133.615
R31835 vss.n5059 vss.n5058 133.615
R31836 vss.n2851 vss.n2850 133.615
R31837 vss.n9871 vss.n2827 133.615
R31838 vss.n4982 vss.n4981 133.615
R31839 vss.n5184 vss.n5183 133.615
R31840 vss.n3165 vss.n3164 133.615
R31841 vss.n10201 vss.n10200 133.615
R31842 vss.n12512 vss.n12511 133.615
R31843 vss.n2220 vss.n2219 133.615
R31844 vss.n12383 vss.n12382 133.615
R31845 vss.n10279 vss.n10278 133.615
R31846 vss.n2459 vss.n2458 133.615
R31847 vss.n2538 vss.n2537 133.615
R31848 vss.n13030 vss.n13029 133.615
R31849 vss.n11326 vss.n11325 133.615
R31850 vss.n11312 vss.n11311 133.615
R31851 vss.n11265 vss.n11264 133.615
R31852 vss.n11251 vss.n11250 133.615
R31853 vss.n11204 vss.n11203 133.615
R31854 vss.n11196 vss.n11195 133.615
R31855 vss.n12669 vss.n10457 133.615
R31856 vss.n11346 vss.n11345 133.615
R31857 vss.n8099 vss.n8010 119.837
R31858 vss.n8985 vss.t25 99.1734
R31859 vss.t25 vss.n496 99.1734
R31860 vss.t83 vss.n497 99.1734
R31861 vss.n13209 vss.t83 99.1734
R31862 vss.n6219 vss.n2793 94.4601
R31863 vss.n5882 vss.n2171 94.4601
R31864 vss.t79 vss.n11048 93.0605
R31865 vss.t77 vss.n2793 87.5028
R31866 vss.t27 vss.n6219 87.5028
R31867 vss.t27 vss.n6220 87.5028
R31868 vss.t76 vss.n2171 87.5028
R31869 vss.n5882 vss.t90 87.5028
R31870 vss.n13266 vss.n13265 86.5632
R31871 vss.n716 vss.n715 86.5632
R31872 vss.n9383 vss.n6184 86.5632
R31873 vss.n9140 vss.n9139 86.5632
R31874 vss.n9954 vss.n2639 86.5632
R31875 vss.n5734 vss.n5733 86.5632
R31876 vss.n13137 vss.n2048 86.5632
R31877 vss.n12087 vss.n12086 86.5632
R31878 vss.n14782 vss.t26 82.8568
R31879 vss.n14772 vss.t26 82.8568
R31880 vss.n8986 vss.n8985 81.7347
R31881 vss.n13210 vss.n13209 81.7347
R31882 vss.n12672 vss.n12671 76.6967
R31883 vss.n12599 vss.t232 75.8142
R31884 vss.n11528 vss.t142 75.8142
R31885 vss.n12756 vss.t1147 75.8142
R31886 vss.t268 vss.n13873 75.8142
R31887 vss.t516 vss.n13768 75.8142
R31888 vss.t1128 vss.n13663 75.8142
R31889 vss.n667 vss.t1279 75.8142
R31890 vss.n1749 vss.t545 75.8142
R31891 vss.n1853 vss.t315 75.8142
R31892 vss.t1054 vss.n8283 75.8142
R31893 vss.n8645 vss.t1223 75.8142
R31894 vss.n8558 vss.t424 75.8142
R31895 vss.n7255 vss.t839 75.8142
R31896 vss.n6785 vss.t248 75.8142
R31897 vss.n6879 vss.t343 75.8142
R31898 vss.n5583 vss.t699 75.8142
R31899 vss.n5497 vss.t812 75.8142
R31900 vss.n5411 vss.t1265 75.8142
R31901 vss.n4557 vss.t155 75.8142
R31902 vss.n3827 vss.t1284 75.8142
R31903 vss.n3922 vss.t629 75.8142
R31904 vss.n12152 vss.t1057 75.8142
R31905 vss.n12548 vss.t1132 75.8142
R31906 vss.t32 vss.n12831 75.8142
R31907 vss.n10000 vss.t90 75.3274
R31908 vss.n12059 vss.t958 74.8587
R31909 vss.n12007 vss.t1046 74.8587
R31910 vss.t841 vss.n10671 74.8587
R31911 vss.t950 vss.n10858 74.8587
R31912 vss.n11494 vss.t993 74.8587
R31913 vss.n10927 vss.t954 74.8587
R31914 vss.n12724 vss.t1001 74.8587
R31915 vss.t914 vss.n13898 74.8587
R31916 vss.t1024 vss.n13844 74.8587
R31917 vss.t47 vss.n13793 74.8587
R31918 vss.t1026 vss.n13739 74.8587
R31919 vss.t991 vss.n13688 74.8587
R31920 vss.t1040 vss.n13634 74.8587
R31921 vss.t1018 vss.n13583 74.8587
R31922 vss.t999 vss.n14002 74.8587
R31923 vss.t952 vss.n13967 74.8587
R31924 vss.n1727 vss.t890 74.8587
R31925 vss.t1022 vss.n1779 74.8587
R31926 vss.n1831 vss.t997 74.8587
R31927 vss.t847 vss.n1883 74.8587
R31928 vss.t886 vss.n1954 74.8587
R31929 vss.n9017 vss.t946 74.8587
R31930 vss.n8304 vss.t912 74.8587
R31931 vss.n8673 vss.t1032 74.8587
R31932 vss.n8630 vss.t956 74.8587
R31933 vss.n8586 vss.t1030 74.8587
R31934 vss.n8543 vss.t1028 74.8587
R31935 vss.t1042 vss.n9551 74.8587
R31936 vss.t989 vss.n9516 74.8587
R31937 vss.n6763 vss.t43 74.8587
R31938 vss.t995 vss.n7061 74.8587
R31939 vss.t918 vss.n6893 74.8587
R31940 vss.t57 vss.n9224 74.8587
R31941 vss.n9081 vss.t1034 74.8587
R31942 vss.n9909 vss.t1044 74.8587
R31943 vss.n5611 vss.t787 74.8587
R31944 vss.n5568 vss.t845 74.8587
R31945 vss.n5525 vss.t966 74.8587
R31946 vss.n5482 vss.t878 74.8587
R31947 vss.n5439 vss.t964 74.8587
R31948 vss.n5396 vss.t55 74.8587
R31949 vss.n4535 vss.t948 74.8587
R31950 vss.t916 vss.n4587 74.8587
R31951 vss.t1036 vss.n4184 74.8587
R31952 vss.t962 vss.n4149 74.8587
R31953 vss.t849 vss.n3936 74.8587
R31954 vss.t51 vss.n5816 74.8587
R31955 vss.n5675 vss.t1003 74.8587
R31956 vss.n12122 vss.t1038 74.8587
R31957 vss.n12175 vss.t872 74.8587
R31958 vss.t851 vss.n12227 74.8587
R31959 vss.n12571 vss.t874 74.8587
R31960 vss.t882 vss.n11662 74.8587
R31961 vss.t843 vss.n12809 74.8587
R31962 vss.n12942 vss.t45 74.8587
R31963 vss.n12591 vss.n12590 74.4102
R31964 vss.n11520 vss.n10321 74.4102
R31965 vss.n12767 vss.n12766 74.4102
R31966 vss.n13923 vss.n689 74.4102
R31967 vss.n13927 vss.n685 74.4102
R31968 vss.n13931 vss.n681 74.4102
R31969 vss.n13934 vss.n678 74.4102
R31970 vss.n13930 vss.n682 74.4102
R31971 vss.n13926 vss.n686 74.4102
R31972 vss.n9040 vss.n6574 74.4102
R31973 vss.n9044 vss.n6570 74.4102
R31974 vss.n9048 vss.n6556 74.4102
R31975 vss.n7267 vss.n7266 74.4102
R31976 vss.n9041 vss.n6573 74.4102
R31977 vss.n9045 vss.n6569 74.4102
R31978 vss.n5634 vss.n3630 74.4102
R31979 vss.n5638 vss.n3626 74.4102
R31980 vss.n5642 vss.n3612 74.4102
R31981 vss.n4422 vss.n2708 74.4102
R31982 vss.n5635 vss.n3629 74.4102
R31983 vss.n5639 vss.n3625 74.4102
R31984 vss.n11850 vss.n11807 74.4102
R31985 vss.n12589 vss.n10615 74.4102
R31986 vss.n12832 vss.n12770 74.4102
R31987 vss.n12044 vss.t1191 73.9271
R31988 vss.n11613 vss.t685 73.9271
R31989 vss.n11479 vss.t1459 73.9271
R31990 vss.t722 vss.n13819 73.9271
R31991 vss.t687 vss.n13714 73.9271
R31992 vss.t988 vss.n13609 73.9271
R31993 vss.n778 vss.t1148 73.9271
R31994 vss.n1820 vss.t1067 73.9271
R31995 vss.n1924 vss.t1397 73.9271
R31996 vss.n8688 vss.t272 73.9271
R31997 vss.n8601 vss.t1115 73.9271
R31998 vss.n7236 vss.t910 73.9271
R31999 vss.n7045 vss.t557 73.9271
R32000 vss.n9208 vss.t285 73.9271
R32001 vss.n4667 vss.t752 73.9271
R32002 vss.n5540 vss.t938 73.9271
R32003 vss.n5454 vss.t1438 73.9271
R32004 vss.n3771 vss.t465 73.9271
R32005 vss.n4135 vss.t423 73.9271
R32006 vss.n5802 vss.t1093 73.9271
R32007 vss.n8078 vss.t1382 73.9271
R32008 vss.t1258 vss.n12251 73.9271
R32009 vss.n11686 vss.t757 73.9271
R32010 vss.n12921 vss.t1426 73.9271
R32011 vss.n13134 vss.n2051 73.4725
R32012 vss.n13131 vss.n2054 73.4725
R32013 vss.n13128 vss.n2057 73.4725
R32014 vss.n13125 vss.n2060 73.4725
R32015 vss.n13122 vss.n2063 73.4725
R32016 vss.n13119 vss.n2066 73.4725
R32017 vss.n13116 vss.n2069 73.4725
R32018 vss.n13899 vss.n191 73.4725
R32019 vss.n14685 vss.n192 73.4725
R32020 vss.n13794 vss.n250 73.4725
R32021 vss.n14490 vss.n251 73.4725
R32022 vss.n13689 vss.n309 73.4725
R32023 vss.n14295 vss.n310 73.4725
R32024 vss.n13588 vss.n432 73.4725
R32025 vss.n13938 vss.n536 73.4725
R32026 vss.n13941 vss.n575 73.4725
R32027 vss.n13250 vss.n13249 73.4725
R32028 vss.n13253 vss.n740 73.4725
R32029 vss.n13256 vss.n737 73.4725
R32030 vss.n13259 vss.n734 73.4725
R32031 vss.n13262 vss.n731 73.4725
R32032 vss.n9009 vss.n9008 73.4725
R32033 vss.n8710 vss.n8709 73.4725
R32034 vss.n8784 vss.n7681 73.4725
R32035 vss.n8622 vss.n7680 73.4725
R32036 vss.n8903 vss.n7538 73.4725
R32037 vss.n8535 vss.n7537 73.4725
R32038 vss.n9487 vss.n6076 73.4725
R32039 vss.n9490 vss.n6115 73.4725
R32040 vss.n9398 vss.n6169 73.4725
R32041 vss.n9395 vss.n6172 73.4725
R32042 vss.n9392 vss.n6175 73.4725
R32043 vss.n9389 vss.n6178 73.4725
R32044 vss.n9386 vss.n6181 73.4725
R32045 vss.n9901 vss.n9900 73.4725
R32046 vss.n9804 vss.n2992 73.4725
R32047 vss.n9807 vss.n2989 73.4725
R32048 vss.n9810 vss.n2986 73.4725
R32049 vss.n9813 vss.n2983 73.4725
R32050 vss.n9816 vss.n2980 73.4725
R32051 vss.n5388 vss.n2935 73.4725
R32052 vss.n9933 vss.n2704 73.4725
R32053 vss.n9936 vss.n2701 73.4725
R32054 vss.n9939 vss.n2698 73.4725
R32055 vss.n9942 vss.n2695 73.4725
R32056 vss.n9945 vss.n2692 73.4725
R32057 vss.n9948 vss.n2689 73.4725
R32058 vss.n9951 vss.n2686 73.4725
R32059 vss.n11828 vss.n2305 73.4725
R32060 vss.n12991 vss.n2350 73.4725
R32061 vss.n12988 vss.n2353 73.4725
R32062 vss.n12985 vss.n2356 73.4725
R32063 vss.n12982 vss.n2359 73.4725
R32064 vss.n12979 vss.n2362 73.4725
R32065 vss.n12976 vss.n2365 73.4725
R32066 vss.n12036 vss.n12035 72.5581
R32067 vss.n12588 vss.n11623 72.5581
R32068 vss.n12769 vss.n10322 72.5581
R32069 vss.n13925 vss.n687 72.5581
R32070 vss.n13929 vss.n683 72.5581
R32071 vss.n13933 vss.n679 72.5581
R32072 vss.n13932 vss.n680 72.5581
R32073 vss.n13928 vss.n684 72.5581
R32074 vss.n13924 vss.n688 72.5581
R32075 vss.n9042 vss.n6572 72.5581
R32076 vss.n9046 vss.n6568 72.5581
R32077 vss.n9039 vss.n7247 72.5581
R32078 vss.n9043 vss.n6571 72.5581
R32079 vss.n9047 vss.n6567 72.5581
R32080 vss.n5632 vss.n5631 72.5581
R32081 vss.n5636 vss.n3628 72.5581
R32082 vss.n5640 vss.n3624 72.5581
R32083 vss.n5633 vss.n4627 72.5581
R32084 vss.n5637 vss.n3627 72.5581
R32085 vss.n5641 vss.n3623 72.5581
R32086 vss.n9038 vss.n9037 72.5581
R32087 vss.n12252 vss.n10614 72.5581
R32088 vss.n12587 vss.n12586 72.5581
R32089 vss.n12768 vss.n10084 72.5581
R32090 vss.n9999 vss.n2600 72.1163
R32091 vss.n13141 vss.n2045 71.8634
R32092 vss.n10407 vss.n10406 71.8634
R32093 vss.n12655 vss.n12650 71.8634
R32094 vss.n12640 vss.n12639 71.8634
R32095 vss.n12688 vss.n12687 71.8634
R32096 vss.n12675 vss.n12674 71.8634
R32097 vss.n11438 vss.n11437 71.8634
R32098 vss.n11425 vss.n11424 71.8634
R32099 vss.n11391 vss.n11390 71.8634
R32100 vss.n11378 vss.n11377 71.8634
R32101 vss.n10966 vss.n10965 71.8634
R32102 vss.n10953 vss.n10952 71.8634
R32103 vss.n10803 vss.n10802 71.8634
R32104 vss.n10790 vss.n10789 71.8634
R32105 vss.n10759 vss.n10758 71.8634
R32106 vss.n10746 vss.n10745 71.8634
R32107 vss.n11585 vss.n11584 71.8634
R32108 vss.n11572 vss.n11571 71.8634
R32109 vss.n10582 vss.n10581 71.8634
R32110 vss.n10569 vss.n10568 71.8634
R32111 vss.n10538 vss.n10537 71.8634
R32112 vss.n10525 vss.n10524 71.8634
R32113 vss.n11959 vss.n11958 71.8634
R32114 vss.n11946 vss.n11945 71.8634
R32115 vss.n12095 vss.n12094 71.8634
R32116 vss.n12065 vss.n11902 71.8634
R32117 vss.n12048 vss.n11918 71.8634
R32118 vss.n11912 vss.n11907 71.8634
R32119 vss.n12039 vss.n12032 71.8634
R32120 vss.n12025 vss.n11989 71.8634
R32121 vss.n12603 vss.n10604 71.8634
R32122 vss.n12000 vss.n11995 71.8634
R32123 vss.n12594 vss.n10611 71.8634
R32124 vss.n10668 vss.n10667 71.8634
R32125 vss.n11610 vss.n11609 71.8634
R32126 vss.n10673 vss.n10639 71.8634
R32127 vss.n11621 vss.n11620 71.8634
R32128 vss.n10855 vss.n10854 71.8634
R32129 vss.n11532 vss.n10870 71.8634
R32130 vss.n10860 vss.n10859 71.8634
R32131 vss.n11523 vss.n11517 71.8634
R32132 vss.n11510 vss.n10881 71.8634
R32133 vss.n11483 vss.n10897 71.8634
R32134 vss.n10891 vss.n10886 71.8634
R32135 vss.n11474 vss.n11469 71.8634
R32136 vss.n11462 vss.n10907 71.8634
R32137 vss.n12753 vss.n12752 71.8634
R32138 vss.n10920 vss.n10915 71.8634
R32139 vss.n12764 vss.n12763 71.8634
R32140 vss.n12730 vss.n10351 71.8634
R32141 vss.n12713 vss.n10367 71.8634
R32142 vss.n10361 vss.n10356 71.8634
R32143 vss.n12996 vss.n12995 71.8634
R32144 vss.n13011 vss.n13006 71.8634
R32145 vss.n2301 vss.n2261 71.8634
R32146 vss.n2283 vss.n2282 71.8634
R32147 vss.n13110 vss.n2075 71.8634
R32148 vss.n2094 vss.n2093 71.8634
R32149 vss.n1129 vss.n1124 71.8634
R32150 vss.n1114 vss.n1113 71.8634
R32151 vss.n863 vss.n845 71.8634
R32152 vss.n872 vss.n871 71.8634
R32153 vss.n14156 vss.n455 71.8634
R32154 vss.n14173 vss.n436 71.8634
R32155 vss.n187 vss.n175 71.8634
R32156 vss.n14786 vss.n14 71.8634
R32157 vss.n337 vss.n336 71.8634
R32158 vss.n352 vss.n347 71.8634
R32159 vss.n14218 vss.n14179 71.8634
R32160 vss.n14200 vss.n14199 71.8634
R32161 vss.n14116 vss.n14115 71.8634
R32162 vss.n14131 vss.n14126 71.8634
R32163 vss.n14225 vss.n14224 71.8634
R32164 vss.n14240 vss.n14235 71.8634
R32165 vss.n14152 vss.n462 71.8634
R32166 vss.n13580 vss.n13568 71.8634
R32167 vss.n13606 vss.n13547 71.8634
R32168 vss.n13589 vss.n13586 71.8634
R32169 vss.n14681 vss.n196 71.8634
R32170 vss.n14663 vss.n14662 71.8634
R32171 vss.n14539 vss.n14538 71.8634
R32172 vss.n14554 vss.n14549 71.8634
R32173 vss.n14486 vss.n255 71.8634
R32174 vss.n14468 vss.n14467 71.8634
R32175 vss.n14344 vss.n14343 71.8634
R32176 vss.n14359 vss.n14354 71.8634
R32177 vss.n14291 vss.n314 71.8634
R32178 vss.n14273 vss.n14272 71.8634
R32179 vss.n14337 vss.n14298 71.8634
R32180 vss.n14319 vss.n14318 71.8634
R32181 vss.n14390 vss.n14389 71.8634
R32182 vss.n14405 vss.n14400 71.8634
R32183 vss.n14532 vss.n14493 71.8634
R32184 vss.n14514 vss.n14513 71.8634
R32185 vss.n14585 vss.n14584 71.8634
R32186 vss.n14600 vss.n14595 71.8634
R32187 vss.n14727 vss.n14688 71.8634
R32188 vss.n14709 vss.n14708 71.8634
R32189 vss.n14734 vss.n14733 71.8634
R32190 vss.n14749 vss.n14744 71.8634
R32191 vss.n13918 vss.n13306 71.8634
R32192 vss.n13906 vss.n13905 71.8634
R32193 vss.n13874 vss.n13342 71.8634
R32194 vss.n13895 vss.n13328 71.8634
R32195 vss.n13870 vss.n13348 71.8634
R32196 vss.n13851 vss.n13850 71.8634
R32197 vss.n13820 vss.n13383 71.8634
R32198 vss.n13841 vss.n13367 71.8634
R32199 vss.n13816 vss.n13389 71.8634
R32200 vss.n13801 vss.n13800 71.8634
R32201 vss.n13769 vss.n13422 71.8634
R32202 vss.n13790 vss.n13408 71.8634
R32203 vss.n13765 vss.n13428 71.8634
R32204 vss.n13746 vss.n13745 71.8634
R32205 vss.n13715 vss.n13463 71.8634
R32206 vss.n13736 vss.n13447 71.8634
R32207 vss.n13711 vss.n13469 71.8634
R32208 vss.n13696 vss.n13695 71.8634
R32209 vss.n13664 vss.n13502 71.8634
R32210 vss.n13685 vss.n13488 71.8634
R32211 vss.n13660 vss.n13508 71.8634
R32212 vss.n13641 vss.n13640 71.8634
R32213 vss.n13610 vss.n13543 71.8634
R32214 vss.n13631 vss.n13527 71.8634
R32215 vss.n656 vss.n655 71.8634
R32216 vss.n635 vss.n630 71.8634
R32217 vss.n13228 vss.n13223 71.8634
R32218 vss.n13213 vss.n13212 71.8634
R32219 vss.n1687 vss.n1682 71.8634
R32220 vss.n1672 vss.n1671 71.8634
R32221 vss.n1640 vss.n1635 71.8634
R32222 vss.n1625 vss.n1624 71.8634
R32223 vss.n1392 vss.n1387 71.8634
R32224 vss.n1377 vss.n1376 71.8634
R32225 vss.n1193 vss.n1188 71.8634
R32226 vss.n1178 vss.n1177 71.8634
R32227 vss.n1345 vss.n1340 71.8634
R32228 vss.n1330 vss.n1329 71.8634
R32229 vss.n1084 vss.n1079 71.8634
R32230 vss.n1069 vss.n1068 71.8634
R32231 vss.n1477 vss.n1472 71.8634
R32232 vss.n1462 vss.n1461 71.8634
R32233 vss.n1558 vss.n1552 71.8634
R32234 vss.n1542 vss.n1541 71.8634
R32235 vss.n13946 vss.n608 71.8634
R32236 vss.n831 vss.n830 71.8634
R32237 vss.n907 vss.n885 71.8634
R32238 vss.n916 vss.n915 71.8634
R32239 vss.n14017 vss.n14016 71.8634
R32240 vss.n14004 vss.n14003 71.8634
R32241 vss.n676 vss.n675 71.8634
R32242 vss.n13999 vss.n13998 71.8634
R32243 vss.n13982 vss.n13981 71.8634
R32244 vss.n13969 vss.n13968 71.8634
R32245 vss.n775 vss.n774 71.8634
R32246 vss.n13964 vss.n13963 71.8634
R32247 vss.n786 vss.n785 71.8634
R32248 vss.n13247 vss.n13246 71.8634
R32249 vss.n1746 vss.n1745 71.8634
R32250 vss.n1732 vss.n1725 71.8634
R32251 vss.n1794 vss.n1793 71.8634
R32252 vss.n1781 vss.n1780 71.8634
R32253 vss.n1817 vss.n1816 71.8634
R32254 vss.n1776 vss.n1775 71.8634
R32255 vss.n1261 vss.n1247 71.8634
R32256 vss.n1255 vss.n1254 71.8634
R32257 vss.n1850 vss.n1849 71.8634
R32258 vss.n1836 vss.n1229 71.8634
R32259 vss.n1898 vss.n1897 71.8634
R32260 vss.n1885 vss.n1884 71.8634
R32261 vss.n1921 vss.n1920 71.8634
R32262 vss.n1880 vss.n1879 71.8634
R32263 vss.n1969 vss.n1968 71.8634
R32264 vss.n1956 vss.n1955 71.8634
R32265 vss.n13299 vss.n13298 71.8634
R32266 vss.n1951 vss.n1950 71.8634
R32267 vss.n13281 vss.n13280 71.8634
R32268 vss.n13268 vss.n13267 71.8634
R32269 vss.n2019 vss.n2014 71.8634
R32270 vss.n2004 vss.n2003 71.8634
R32271 vss.n13178 vss.n13177 71.8634
R32272 vss.n13192 vss.n13187 71.8634
R32273 vss.n9606 vss.n9605 71.8634
R32274 vss.n9621 vss.n9616 71.8634
R32275 vss.n9185 vss.n9180 71.8634
R32276 vss.n9170 vss.n9169 71.8634
R32277 vss.n9484 vss.n9483 71.8634
R32278 vss.n9467 vss.n9460 71.8634
R32279 vss.n8049 vss.n8015 71.8634
R32280 vss.n8033 vss.n8026 71.8634
R32281 vss.n9666 vss.n5976 71.8634
R32282 vss.n5995 vss.n5994 71.8634
R32283 vss.n8150 vss.n8148 71.8634
R32284 vss.n8138 vss.n8137 71.8634
R32285 vss.n8154 vss.n8120 71.8634
R32286 vss.n8171 vss.n8102 71.8634
R32287 vss.n8080 vss.n8076 71.8634
R32288 vss.n8097 vss.n8055 71.8634
R32289 vss.n8223 vss.n8222 71.8634
R32290 vss.n8238 vss.n8233 71.8634
R32291 vss.n8216 vss.n8177 71.8634
R32292 vss.n8198 vss.n8197 71.8634
R32293 vss.n9004 vss.n7302 71.8634
R32294 vss.n7321 vss.n7320 71.8634
R32295 vss.n8714 vss.n8713 71.8634
R32296 vss.n8729 vss.n8724 71.8634
R32297 vss.n7788 vss.n7787 71.8634
R32298 vss.n7803 vss.n7798 71.8634
R32299 vss.n8780 vss.n7685 71.8634
R32300 vss.n8762 vss.n8761 71.8634
R32301 vss.n8833 vss.n8832 71.8634
R32302 vss.n8848 vss.n8843 71.8634
R32303 vss.n8826 vss.n8787 71.8634
R32304 vss.n8808 vss.n8807 71.8634
R32305 vss.n8899 vss.n7542 71.8634
R32306 vss.n8881 vss.n8880 71.8634
R32307 vss.n9035 vss.n7270 71.8634
R32308 vss.n7289 vss.n7288 71.8634
R32309 vss.n8280 vss.n7902 71.8634
R32310 vss.n7296 vss.n7295 71.8634
R32311 vss.n8284 vss.n7898 71.8634
R32312 vss.n8301 vss.n7880 71.8634
R32313 vss.n8690 vss.n8317 71.8634
R32314 vss.n8707 vss.n7869 71.8634
R32315 vss.n8323 vss.n8322 71.8634
R32316 vss.n8676 vss.n8344 71.8634
R32317 vss.n8651 vss.n8362 71.8634
R32318 vss.n8664 vss.n8663 71.8634
R32319 vss.n8368 vss.n8367 71.8634
R32320 vss.n8633 vss.n8394 71.8634
R32321 vss.n8607 vss.n8415 71.8634
R32322 vss.n8620 vss.n8619 71.8634
R32323 vss.n8421 vss.n8420 71.8634
R32324 vss.n8589 vss.n8442 71.8634
R32325 vss.n8564 vss.n8460 71.8634
R32326 vss.n8577 vss.n8576 71.8634
R32327 vss.n8466 vss.n8465 71.8634
R32328 vss.n8546 vss.n8492 71.8634
R32329 vss.n8522 vss.n8508 71.8634
R32330 vss.n8533 vss.n8532 71.8634
R32331 vss.n8952 vss.n8951 71.8634
R32332 vss.n8967 vss.n8962 71.8634
R32333 vss.n8945 vss.n8906 71.8634
R32334 vss.n8927 vss.n8926 71.8634
R32335 vss.n7533 vss.n7493 71.8634
R32336 vss.n7515 vss.n7514 71.8634
R32337 vss.n7565 vss.n7564 71.8634
R32338 vss.n7580 vss.n7575 71.8634
R32339 vss.n7708 vss.n7707 71.8634
R32340 vss.n7723 vss.n7718 71.8634
R32341 vss.n7929 vss.n7928 71.8634
R32342 vss.n7944 vss.n7939 71.8634
R32343 vss.n6044 vss.n6038 71.8634
R32344 vss.n6028 vss.n6027 71.8634
R32345 vss.n7213 vss.n7208 71.8634
R32346 vss.n7198 vss.n7197 71.8634
R32347 vss.n6708 vss.n6703 71.8634
R32348 vss.n6693 vss.n6692 71.8634
R32349 vss.n6664 vss.n6659 71.8634
R32350 vss.n6649 vss.n6648 71.8634
R32351 vss.n7022 vss.n7017 71.8634
R32352 vss.n7007 vss.n7006 71.8634
R32353 vss.n6482 vss.n6477 71.8634
R32354 vss.n6467 vss.n6466 71.8634
R32355 vss.n6437 vss.n6432 71.8634
R32356 vss.n6422 vss.n6421 71.8634
R32357 vss.n6359 vss.n6354 71.8634
R32358 vss.n6344 vss.n6343 71.8634
R32359 vss.n6973 vss.n6968 71.8634
R32360 vss.n6958 vss.n6957 71.8634
R32361 vss.n7162 vss.n7157 71.8634
R32362 vss.n7147 vss.n7146 71.8634
R32363 vss.n9495 vss.n6165 71.8634
R32364 vss.n6155 vss.n6154 71.8634
R32365 vss.n9442 vss.n9441 71.8634
R32366 vss.n9422 vss.n9416 71.8634
R32367 vss.n9566 vss.n9565 71.8634
R32368 vss.n9553 vss.n9552 71.8634
R32369 vss.n7264 vss.n7263 71.8634
R32370 vss.n9548 vss.n9547 71.8634
R32371 vss.n9531 vss.n9530 71.8634
R32372 vss.n9518 vss.n9517 71.8634
R32373 vss.n7245 vss.n7244 71.8634
R32374 vss.n9513 vss.n9512 71.8634
R32375 vss.n7233 vss.n7232 71.8634
R32376 vss.n6756 vss.n6755 71.8634
R32377 vss.n6782 vss.n6781 71.8634
R32378 vss.n6768 vss.n6745 71.8634
R32379 vss.n7076 vss.n7075 71.8634
R32380 vss.n7063 vss.n7062 71.8634
R32381 vss.n6824 vss.n6823 71.8634
R32382 vss.n7058 vss.n7057 71.8634
R32383 vss.n7042 vss.n7041 71.8634
R32384 vss.n6897 vss.n6847 71.8634
R32385 vss.n6875 vss.n6874 71.8634
R32386 vss.n6890 vss.n6889 71.8634
R32387 vss.n9239 vss.n9238 71.8634
R32388 vss.n9226 vss.n9225 71.8634
R32389 vss.n6565 vss.n6564 71.8634
R32390 vss.n9221 vss.n9220 71.8634
R32391 vss.n9205 vss.n9204 71.8634
R32392 vss.n9074 vss.n9073 71.8634
R32393 vss.n9095 vss.n9094 71.8634
R32394 vss.n9084 vss.n9083 71.8634
R32395 vss.n9137 vss.n9136 71.8634
R32396 vss.n9123 vss.n9118 71.8634
R32397 vss.n9355 vss.n9350 71.8634
R32398 vss.n9340 vss.n9339 71.8634
R32399 vss.n9380 vss.n9379 71.8634
R32400 vss.n6207 vss.n6201 71.8634
R32401 vss.n5956 vss.n5955 71.8634
R32402 vss.n9675 vss.n5966 71.8634
R32403 vss.n9706 vss.n9705 71.8634
R32404 vss.n9722 vss.n9716 71.8634
R32405 vss.n2577 vss.n2576 71.8634
R32406 vss.n10003 vss.n2587 71.8634
R32407 vss.n9893 vss.n2746 71.8634
R32408 vss.n2765 vss.n2764 71.8634
R32409 vss.n3284 vss.n3283 71.8634
R32410 vss.n3300 vss.n3293 71.8634
R32411 vss.n9763 vss.n9762 71.8634
R32412 vss.n9778 vss.n9777 71.8634
R32413 vss.n3203 vss.n3202 71.8634
R32414 vss.n3218 vss.n3217 71.8634
R32415 vss.n9800 vss.n2997 71.8634
R32416 vss.n3020 vss.n3019 71.8634
R32417 vss.n5233 vss.n5232 71.8634
R32418 vss.n5248 vss.n5247 71.8634
R32419 vss.n3046 vss.n3045 71.8634
R32420 vss.n3061 vss.n3060 71.8634
R32421 vss.n5103 vss.n5102 71.8634
R32422 vss.n5118 vss.n5117 71.8634
R32423 vss.n5292 vss.n5291 71.8634
R32424 vss.n5307 vss.n5306 71.8634
R32425 vss.n5020 vss.n5019 71.8634
R32426 vss.n5035 vss.n5034 71.8634
R32427 vss.n4901 vss.n4900 71.8634
R32428 vss.n4916 vss.n4915 71.8634
R32429 vss.n9927 vss.n2711 71.8634
R32430 vss.n2730 vss.n2729 71.8634
R32431 vss.n4664 vss.n4639 71.8634
R32432 vss.n2737 vss.n2736 71.8634
R32433 vss.n5629 vss.n4630 71.8634
R32434 vss.n4682 vss.n4681 71.8634
R32435 vss.n5589 vss.n4697 71.8634
R32436 vss.n5602 vss.n5601 71.8634
R32437 vss.n4703 vss.n4702 71.8634
R32438 vss.n5571 vss.n4722 71.8634
R32439 vss.n5546 vss.n4740 71.8634
R32440 vss.n5559 vss.n5558 71.8634
R32441 vss.n4746 vss.n4745 71.8634
R32442 vss.n5528 vss.n4765 71.8634
R32443 vss.n5503 vss.n4783 71.8634
R32444 vss.n5516 vss.n5515 71.8634
R32445 vss.n4789 vss.n4788 71.8634
R32446 vss.n5485 vss.n4808 71.8634
R32447 vss.n5460 vss.n4826 71.8634
R32448 vss.n5473 vss.n5472 71.8634
R32449 vss.n4832 vss.n4831 71.8634
R32450 vss.n5442 vss.n4851 71.8634
R32451 vss.n5417 vss.n4869 71.8634
R32452 vss.n5430 vss.n5429 71.8634
R32453 vss.n4875 vss.n4874 71.8634
R32454 vss.n5399 vss.n5345 71.8634
R32455 vss.n5375 vss.n5361 71.8634
R32456 vss.n5386 vss.n5385 71.8634
R32457 vss.n9822 vss.n9821 71.8634
R32458 vss.n9837 vss.n9836 71.8634
R32459 vss.n2977 vss.n2940 71.8634
R32460 vss.n2963 vss.n2962 71.8634
R32461 vss.n2931 vss.n2893 71.8634
R32462 vss.n2916 vss.n2915 71.8634
R32463 vss.n4942 vss.n4941 71.8634
R32464 vss.n4957 vss.n4956 71.8634
R32465 vss.n5144 vss.n5143 71.8634
R32466 vss.n5159 vss.n5158 71.8634
R32467 vss.n3125 vss.n3124 71.8634
R32468 vss.n3140 vss.n3139 71.8634
R32469 vss.n4495 vss.n4494 71.8634
R32470 vss.n4482 vss.n4481 71.8634
R32471 vss.n4403 vss.n4402 71.8634
R32472 vss.n4390 vss.n4389 71.8634
R32473 vss.n4355 vss.n4354 71.8634
R32474 vss.n4342 vss.n4341 71.8634
R32475 vss.n3755 vss.n3754 71.8634
R32476 vss.n3742 vss.n3741 71.8634
R32477 vss.n4057 vss.n4056 71.8634
R32478 vss.n4044 vss.n4043 71.8634
R32479 vss.n3710 vss.n3709 71.8634
R32480 vss.n3697 vss.n3696 71.8634
R32481 vss.n4111 vss.n4110 71.8634
R32482 vss.n4098 vss.n4097 71.8634
R32483 vss.n3535 vss.n3534 71.8634
R32484 vss.n3522 vss.n3521 71.8634
R32485 vss.n3490 vss.n3489 71.8634
R32486 vss.n3477 vss.n3476 71.8634
R32487 vss.n5778 vss.n5777 71.8634
R32488 vss.n5765 vss.n5764 71.8634
R32489 vss.n4524 vss.n4510 71.8634
R32490 vss.n4518 vss.n4517 71.8634
R32491 vss.n4554 vss.n4553 71.8634
R32492 vss.n4540 vss.n4441 71.8634
R32493 vss.n4602 vss.n4601 71.8634
R32494 vss.n4589 vss.n4588 71.8634
R32495 vss.n4625 vss.n4624 71.8634
R32496 vss.n4584 vss.n4583 71.8634
R32497 vss.n4199 vss.n4198 71.8634
R32498 vss.n4186 vss.n4185 71.8634
R32499 vss.n3824 vss.n3823 71.8634
R32500 vss.n4181 vss.n4180 71.8634
R32501 vss.n4164 vss.n4163 71.8634
R32502 vss.n4151 vss.n4150 71.8634
R32503 vss.n3867 vss.n3866 71.8634
R32504 vss.n4146 vss.n4145 71.8634
R32505 vss.n4132 vss.n4131 71.8634
R32506 vss.n3940 vss.n3890 71.8634
R32507 vss.n3918 vss.n3917 71.8634
R32508 vss.n3933 vss.n3932 71.8634
R32509 vss.n5831 vss.n5830 71.8634
R32510 vss.n5818 vss.n5817 71.8634
R32511 vss.n3621 vss.n3620 71.8634
R32512 vss.n5813 vss.n5812 71.8634
R32513 vss.n5799 vss.n5798 71.8634
R32514 vss.n5668 vss.n5667 71.8634
R32515 vss.n5689 vss.n5688 71.8634
R32516 vss.n5678 vss.n5677 71.8634
R32517 vss.n5731 vss.n5730 71.8634
R32518 vss.n5717 vss.n5712 71.8634
R32519 vss.n9982 vss.n9981 71.8634
R32520 vss.n9969 vss.n9968 71.8634
R32521 vss.n2682 vss.n2681 71.8634
R32522 vss.n2666 vss.n2660 71.8634
R32523 vss.n3415 vss.n3414 71.8634
R32524 vss.n3402 vss.n3401 71.8634
R32525 vss.n4012 vss.n4011 71.8634
R32526 vss.n3999 vss.n3998 71.8634
R32527 vss.n4279 vss.n4278 71.8634
R32528 vss.n4266 vss.n4265 71.8634
R32529 vss.n5924 vss.n5919 71.8634
R32530 vss.n5909 vss.n5908 71.8634
R32531 vss.n14066 vss.n14065 71.8634
R32532 vss.n14081 vss.n14080 71.8634
R32533 vss.n10121 vss.n10120 71.8634
R32534 vss.n10136 vss.n10135 71.8634
R32535 vss.n12879 vss.n12878 71.8634
R32536 vss.n12894 vss.n12893 71.8634
R32537 vss.n10162 vss.n10161 71.8634
R32538 vss.n10177 vss.n10176 71.8634
R32539 vss.n12428 vss.n12427 71.8634
R32540 vss.n12443 vss.n12442 71.8634
R32541 vss.n11757 vss.n11756 71.8634
R32542 vss.n11772 vss.n11771 71.8634
R32543 vss.n12473 vss.n12472 71.8634
R32544 vss.n12488 vss.n12487 71.8634
R32545 vss.n2347 vss.n2310 71.8634
R32546 vss.n2333 vss.n2332 71.8634
R32547 vss.n12298 vss.n12297 71.8634
R32548 vss.n12313 vss.n12312 71.8634
R32549 vss.n12343 vss.n12342 71.8634
R32550 vss.n12358 vss.n12357 71.8634
R32551 vss.n10239 vss.n10238 71.8634
R32552 vss.n10254 vss.n10253 71.8634
R32553 vss.n2419 vss.n2418 71.8634
R32554 vss.n2434 vss.n2433 71.8634
R32555 vss.n12972 vss.n2370 71.8634
R32556 vss.n2393 vss.n2392 71.8634
R32557 vss.n10044 vss.n10043 71.8634
R32558 vss.n12945 vss.n10054 71.8634
R32559 vss.n10039 vss.n10038 71.8634
R32560 vss.n13080 vss.n2114 71.8634
R32561 vss.n12923 vss.n10081 71.8634
R32562 vss.n12940 vss.n12939 71.8634
R32563 vss.n2499 vss.n2498 71.8634
R32564 vss.n2514 vss.n2513 71.8634
R32565 vss.n13074 vss.n2122 71.8634
R32566 vss.n2141 vss.n2140 71.8634
R32567 vss.n12101 vss.n11848 71.8634
R32568 vss.n12120 vss.n12119 71.8634
R32569 vss.n12150 vss.n11811 71.8634
R32570 vss.n12132 vss.n12131 71.8634
R32571 vss.n12154 vss.n11804 71.8634
R32572 vss.n12173 vss.n12172 71.8634
R32573 vss.n12254 vss.n12187 71.8634
R32574 vss.n12269 vss.n12268 71.8634
R32575 vss.n12248 vss.n12193 71.8634
R32576 vss.n12234 vss.n12233 71.8634
R32577 vss.n12546 vss.n11723 71.8634
R32578 vss.n12224 vss.n12212 71.8634
R32579 vss.n12550 vss.n11717 71.8634
R32580 vss.n12569 vss.n12568 71.8634
R32581 vss.n12584 vss.n11626 71.8634
R32582 vss.n11697 vss.n11634 71.8634
R32583 vss.n11683 vss.n11644 71.8634
R32584 vss.n11669 vss.n11668 71.8634
R32585 vss.n12834 vss.n10319 71.8634
R32586 vss.n12849 vss.n12848 71.8634
R32587 vss.n12828 vss.n12775 71.8634
R32588 vss.n12816 vss.n12815 71.8634
R32589 vss.n12919 vss.n10088 71.8634
R32590 vss.n12806 vss.n12794 71.8634
R32591 vss.n12084 vss.n12083 71.8634
R32592 vss.n11883 vss.n11878 71.8634
R32593 vss.n10494 vss.n10493 71.8634
R32594 vss.n10481 vss.n10480 71.8634
R32595 vss.n10715 vss.n10714 71.8634
R32596 vss.n10702 vss.n10701 71.8634
R32597 vss.n11029 vss.n11028 71.8634
R32598 vss.n11016 vss.n11015 71.8634
R32599 vss.n11139 vss.n11134 71.8634
R32600 vss.n11124 vss.n11123 71.8634
R32601 vss.n10397 vss.n10396 68.5181
R32602 vss.n10405 vss.n10397 68.5181
R32603 vss.n13147 vss.n2032 68.5181
R32604 vss.n2042 vss.n2032 68.5181
R32605 vss.n2044 vss.n2034 68.5181
R32606 vss.n13142 vss.n2044 68.5181
R32607 vss.n12637 vss.n12636 68.5181
R32608 vss.n12636 vss.n12631 68.5181
R32609 vss.n12661 vss.n12621 68.5181
R32610 vss.n12647 vss.n12621 68.5181
R32611 vss.n12649 vss.n12623 68.5181
R32612 vss.n12656 vss.n12649 68.5181
R32613 vss.n10381 vss.n10376 68.5181
R32614 vss.n12684 vss.n10381 68.5181
R32615 vss.n12695 vss.n10374 68.5181
R32616 vss.n12682 vss.n10374 68.5181
R32617 vss.n10391 vss.n10390 68.5181
R32618 vss.n10390 vss.n10383 68.5181
R32619 vss.n11412 vss.n11407 68.5181
R32620 vss.n11434 vss.n11412 68.5181
R32621 vss.n11445 vss.n11405 68.5181
R32622 vss.n11432 vss.n11405 68.5181
R32623 vss.n11422 vss.n11421 68.5181
R32624 vss.n11421 vss.n11414 68.5181
R32625 vss.n11365 vss.n11360 68.5181
R32626 vss.n11387 vss.n11365 68.5181
R32627 vss.n11398 vss.n11358 68.5181
R32628 vss.n11385 vss.n11358 68.5181
R32629 vss.n11375 vss.n11374 68.5181
R32630 vss.n11374 vss.n11367 68.5181
R32631 vss.n10940 vss.n10935 68.5181
R32632 vss.n10962 vss.n10940 68.5181
R32633 vss.n10973 vss.n10933 68.5181
R32634 vss.n10960 vss.n10933 68.5181
R32635 vss.n10950 vss.n10949 68.5181
R32636 vss.n10949 vss.n10942 68.5181
R32637 vss.n10777 vss.n10772 68.5181
R32638 vss.n10799 vss.n10777 68.5181
R32639 vss.n10810 vss.n10770 68.5181
R32640 vss.n10797 vss.n10770 68.5181
R32641 vss.n10787 vss.n10786 68.5181
R32642 vss.n10786 vss.n10779 68.5181
R32643 vss.n10733 vss.n10728 68.5181
R32644 vss.n10755 vss.n10733 68.5181
R32645 vss.n10766 vss.n10726 68.5181
R32646 vss.n10753 vss.n10726 68.5181
R32647 vss.n10743 vss.n10742 68.5181
R32648 vss.n10742 vss.n10735 68.5181
R32649 vss.n11559 vss.n11554 68.5181
R32650 vss.n11581 vss.n11559 68.5181
R32651 vss.n11592 vss.n11552 68.5181
R32652 vss.n11579 vss.n11552 68.5181
R32653 vss.n11569 vss.n11568 68.5181
R32654 vss.n11568 vss.n11561 68.5181
R32655 vss.n10556 vss.n10551 68.5181
R32656 vss.n10578 vss.n10556 68.5181
R32657 vss.n10589 vss.n10549 68.5181
R32658 vss.n10576 vss.n10549 68.5181
R32659 vss.n10566 vss.n10565 68.5181
R32660 vss.n10565 vss.n10558 68.5181
R32661 vss.n10512 vss.n10507 68.5181
R32662 vss.n10534 vss.n10512 68.5181
R32663 vss.n10545 vss.n10505 68.5181
R32664 vss.n10532 vss.n10505 68.5181
R32665 vss.n10522 vss.n10521 68.5181
R32666 vss.n10521 vss.n10514 68.5181
R32667 vss.n11933 vss.n11928 68.5181
R32668 vss.n11955 vss.n11933 68.5181
R32669 vss.n11966 vss.n11926 68.5181
R32670 vss.n11953 vss.n11926 68.5181
R32671 vss.n11943 vss.n11942 68.5181
R32672 vss.n11942 vss.n11935 68.5181
R32673 vss.n12077 vss.n11861 68.5181
R32674 vss.n12082 vss.n11861 68.5181
R32675 vss.n12076 vss.n11871 68.5181
R32676 vss.n11871 vss.n11862 68.5181
R32677 vss.n12061 vss.n11901 68.5181
R32678 vss.n12066 vss.n11901 68.5181
R32679 vss.n12073 vss.n11892 68.5181
R32680 vss.n11892 vss.n11855 68.5181
R32681 vss.n11894 vss.n11854 68.5181
R32682 vss.n12093 vss.n11854 68.5181
R32683 vss.n12056 vss.n11906 68.5181
R32684 vss.n12056 vss.n12055 68.5181
R32685 vss.n11972 vss.n11922 68.5181
R32686 vss.n11922 vss.n11913 68.5181
R32687 vss.n11978 vss.n11917 68.5181
R32688 vss.n12049 vss.n11917 68.5181
R32689 vss.n12021 vss.n11988 68.5181
R32690 vss.n12026 vss.n11988 68.5181
R32691 vss.n12015 vss.n12012 68.5181
R32692 vss.n12012 vss.n11984 68.5181
R32693 vss.n12041 vss.n11983 68.5181
R32694 vss.n12041 vss.n12040 68.5181
R32695 vss.n12004 vss.n11994 68.5181
R32696 vss.n12004 vss.n12003 68.5181
R32697 vss.n12609 vss.n10591 68.5181
R32698 vss.n10601 vss.n10591 68.5181
R32699 vss.n10603 vss.n10593 68.5181
R32700 vss.n12604 vss.n10603 68.5181
R32701 vss.n10650 vss.n10646 68.5181
R32702 vss.n10666 vss.n10646 68.5181
R32703 vss.n10659 vss.n10658 68.5181
R32704 vss.n10659 vss.n10647 68.5181
R32705 vss.n12596 vss.n10609 68.5181
R32706 vss.n12596 vss.n12595 68.5181
R32707 vss.n10638 vss.n10631 68.5181
R32708 vss.n10674 vss.n10638 68.5181
R32709 vss.n11598 vss.n10630 68.5181
R32710 vss.n10630 vss.n10627 68.5181
R32711 vss.n11599 vss.n10626 68.5181
R32712 vss.n11608 vss.n10626 68.5181
R32713 vss.n10840 vss.n10833 68.5181
R32714 vss.n10853 vss.n10833 68.5181
R32715 vss.n10848 vss.n10842 68.5181
R32716 vss.n10842 vss.n10620 68.5181
R32717 vss.n10845 vss.n10619 68.5181
R32718 vss.n11619 vss.n10619 68.5181
R32719 vss.n10828 vss.n10827 68.5181
R32720 vss.n10827 vss.n10822 68.5181
R32721 vss.n11538 vss.n10812 68.5181
R32722 vss.n10867 vss.n10812 68.5181
R32723 vss.n10869 vss.n10814 68.5181
R32724 vss.n11533 vss.n10869 68.5181
R32725 vss.n11506 vss.n10880 68.5181
R32726 vss.n11511 vss.n10880 68.5181
R32727 vss.n11500 vss.n11499 68.5181
R32728 vss.n11499 vss.n10876 68.5181
R32729 vss.n11525 vss.n10875 68.5181
R32730 vss.n11525 vss.n11524 68.5181
R32731 vss.n11491 vss.n10885 68.5181
R32732 vss.n11491 vss.n11490 68.5181
R32733 vss.n10987 vss.n10976 68.5181
R32734 vss.n10976 vss.n10892 68.5181
R32735 vss.n10979 vss.n10896 68.5181
R32736 vss.n11484 vss.n10896 68.5181
R32737 vss.n11458 vss.n10906 68.5181
R32738 vss.n11463 vss.n10906 68.5181
R32739 vss.n11452 vss.n10932 68.5181
R32740 vss.n10932 vss.n10902 68.5181
R32741 vss.n11476 vss.n10901 68.5181
R32742 vss.n11476 vss.n11475 68.5181
R32743 vss.n10924 vss.n10914 68.5181
R32744 vss.n10924 vss.n10923 68.5181
R32745 vss.n12741 vss.n10337 68.5181
R32746 vss.n10337 vss.n10334 68.5181
R32747 vss.n12742 vss.n10333 68.5181
R32748 vss.n12751 vss.n10333 68.5181
R32749 vss.n12726 vss.n10350 68.5181
R32750 vss.n12731 vss.n10350 68.5181
R32751 vss.n12738 vss.n10341 68.5181
R32752 vss.n10341 vss.n10327 68.5181
R32753 vss.n10343 vss.n10326 68.5181
R32754 vss.n12762 vss.n10326 68.5181
R32755 vss.n12721 vss.n10355 68.5181
R32756 vss.n12721 vss.n12720 68.5181
R32757 vss.n12701 vss.n10371 68.5181
R32758 vss.n10371 vss.n10362 68.5181
R32759 vss.n12707 vss.n10366 68.5181
R32760 vss.n12714 vss.n10366 68.5181
R32761 vss.n12803 vss.n12795 68.5181
R32762 vss.n12804 vss.n12803 68.5181
R32763 vss.n12814 vss.n12811 68.5181
R32764 vss.n12811 vss.n12787 68.5181
R32765 vss.n12786 vss.n12777 68.5181
R32766 vss.n12822 vss.n12786 68.5181
R32767 vss.n10311 vss.n10310 68.5181
R32768 vss.n10310 vss.n10305 68.5181
R32769 vss.n11667 vss.n11664 68.5181
R32770 vss.n11664 vss.n11656 68.5181
R32771 vss.n11655 vss.n11646 68.5181
R32772 vss.n11677 vss.n11655 68.5181
R32773 vss.n11696 vss.n11633 68.5181
R32774 vss.n12576 vss.n11633 68.5181
R32775 vss.n11704 vss.n11703 68.5181
R32776 vss.n12566 vss.n11704 68.5181
R32777 vss.n12559 vss.n11710 68.5181
R32778 vss.n11710 vss.n11705 68.5181
R32779 vss.n12221 vss.n12213 68.5181
R32780 vss.n12222 vss.n12221 68.5181
R32781 vss.n12232 vss.n12229 68.5181
R32782 vss.n12229 vss.n12205 68.5181
R32783 vss.n12204 vss.n12195 68.5181
R32784 vss.n12242 vss.n12204 68.5181
R32785 vss.n12179 vss.n12178 68.5181
R32786 vss.n12178 vss.n11782 68.5181
R32787 vss.n11791 vss.n11790 68.5181
R32788 vss.n12170 vss.n11791 68.5181
R32789 vss.n12163 vss.n11797 68.5181
R32790 vss.n11797 vss.n11792 68.5181
R32791 vss.n12126 vss.n12125 68.5181
R32792 vss.n12125 vss.n11823 68.5181
R32793 vss.n13012 vss.n13005 68.5181
R32794 vss.n13005 vss.n2243 68.5181
R32795 vss.n13003 vss.n2241 68.5181
R32796 vss.n13017 vss.n2241 68.5181
R32797 vss.n2256 vss.n2251 68.5181
R32798 vss.n2257 vss.n2256 68.5181
R32799 vss.n2289 vss.n2277 68.5181
R32800 vss.n2289 vss.n2288 68.5181
R32801 vss.n2294 vss.n2276 68.5181
R32802 vss.n2276 vss.n2266 68.5181
R32803 vss.n2274 vss.n2262 68.5181
R32804 vss.n2299 vss.n2262 68.5181
R32805 vss.n13098 vss.n2088 68.5181
R32806 vss.n13098 vss.n13097 68.5181
R32807 vss.n13103 vss.n2087 68.5181
R32808 vss.n2087 vss.n2077 68.5181
R32809 vss.n2085 vss.n2076 68.5181
R32810 vss.n13108 vss.n2076 68.5181
R32811 vss.n485 vss.n484 68.5181
R32812 vss.n484 vss.n477 68.5181
R32813 vss.n14075 vss.n475 68.5181
R32814 vss.n14087 vss.n475 68.5181
R32815 vss.n13199 vss.n13159 68.5181
R32816 vss.n13185 vss.n13159 68.5181
R32817 vss.n1111 vss.n1110 68.5181
R32818 vss.n1110 vss.n1105 68.5181
R32819 vss.n1135 vss.n1095 68.5181
R32820 vss.n1121 vss.n1095 68.5181
R32821 vss.n1123 vss.n1097 68.5181
R32822 vss.n1130 vss.n1123 68.5181
R32823 vss.n714 vss.n709 68.5181
R32824 vss.n13277 vss.n714 68.5181
R32825 vss.n13288 vss.n707 68.5181
R32826 vss.n13275 vss.n707 68.5181
R32827 vss.n13291 vss.n703 68.5181
R32828 vss.n703 vss.n694 68.5181
R32829 vss.n1144 vss.n1139 68.5181
R32830 vss.n1965 vss.n1144 68.5181
R32831 vss.n1976 vss.n1137 68.5181
R32832 vss.n1963 vss.n1137 68.5181
R32833 vss.n1913 vss.n1157 68.5181
R32834 vss.n1157 vss.n1150 68.5181
R32835 vss.n1209 vss.n1204 68.5181
R32836 vss.n1894 vss.n1209 68.5181
R32837 vss.n1905 vss.n1202 68.5181
R32838 vss.n1892 vss.n1202 68.5181
R32839 vss.n1842 vss.n1222 68.5181
R32840 vss.n1222 vss.n1215 68.5181
R32841 vss.n1824 vss.n1246 68.5181
R32842 vss.n1260 vss.n1246 68.5181
R32843 vss.n1251 vss.n1245 68.5181
R32844 vss.n1258 vss.n1251 68.5181
R32845 vss.n1809 vss.n1275 68.5181
R32846 vss.n1275 vss.n1268 68.5181
R32847 vss.n1705 vss.n1700 68.5181
R32848 vss.n1790 vss.n1705 68.5181
R32849 vss.n1801 vss.n1698 68.5181
R32850 vss.n1788 vss.n1698 68.5181
R32851 vss.n1738 vss.n1718 68.5181
R32852 vss.n1718 vss.n1711 68.5181
R32853 vss.n761 vss.n758 68.5181
R32854 vss.n782 vss.n761 68.5181
R32855 vss.n13240 vss.n757 68.5181
R32856 vss.n757 vss.n747 68.5181
R32857 vss.n13957 vss.n590 68.5181
R32858 vss.n590 vss.n580 68.5181
R32859 vss.n563 vss.n558 68.5181
R32860 vss.n13978 vss.n563 68.5181
R32861 vss.n13989 vss.n556 68.5181
R32862 vss.n13976 vss.n556 68.5181
R32863 vss.n13992 vss.n551 68.5181
R32864 vss.n551 vss.n541 68.5181
R32865 vss.n852 vss.n837 68.5181
R32866 vss.n870 vss.n837 68.5181
R32867 vss.n840 vss.n516 68.5181
R32868 vss.n840 vss.n838 68.5181
R32869 vss.n858 vss.n844 68.5181
R32870 vss.n864 vss.n844 68.5181
R32871 vss.n14166 vss.n437 68.5181
R32872 vss.n14171 vss.n437 68.5181
R32873 vss.n14165 vss.n448 68.5181
R32874 vss.n448 vss.n438 68.5181
R32875 vss.n454 vss.n449 68.5181
R32876 vss.n14160 vss.n454 68.5181
R32877 vss.n14787 vss.n13 68.5181
R32878 vss.n13 vss.n3 68.5181
R32879 vss.n11 vss.n1 68.5181
R32880 vss.n14792 vss.n1 68.5181
R32881 vss.n184 vss.n176 68.5181
R32882 vss.n185 vss.n184 68.5181
R32883 vss.n353 vss.n346 68.5181
R32884 vss.n346 vss.n319 68.5181
R32885 vss.n344 vss.n317 68.5181
R32886 vss.n358 vss.n317 68.5181
R32887 vss.n332 vss.n327 68.5181
R32888 vss.n333 vss.n332 68.5181
R32889 vss.n14206 vss.n14194 68.5181
R32890 vss.n14206 vss.n14205 68.5181
R32891 vss.n14211 vss.n14193 68.5181
R32892 vss.n14193 vss.n14183 68.5181
R32893 vss.n14191 vss.n14180 68.5181
R32894 vss.n14216 vss.n14180 68.5181
R32895 vss.n14132 vss.n14125 68.5181
R32896 vss.n14125 vss.n14098 68.5181
R32897 vss.n14123 vss.n14096 68.5181
R32898 vss.n14137 vss.n14096 68.5181
R32899 vss.n14111 vss.n14106 68.5181
R32900 vss.n14112 vss.n14111 68.5181
R32901 vss.n14241 vss.n14234 68.5181
R32902 vss.n14234 vss.n416 68.5181
R32903 vss.n14232 vss.n414 68.5181
R32904 vss.n14246 vss.n414 68.5181
R32905 vss.n429 vss.n424 68.5181
R32906 vss.n430 vss.n429 68.5181
R32907 vss.n13577 vss.n13569 68.5181
R32908 vss.n13578 vss.n13577 68.5181
R32909 vss.n473 vss.n464 68.5181
R32910 vss.n14146 vss.n473 68.5181
R32911 vss.n14151 vss.n463 68.5181
R32912 vss.n471 vss.n463 68.5181
R32913 vss.n13594 vss.n13563 68.5181
R32914 vss.n13594 vss.n13593 68.5181
R32915 vss.n13599 vss.n13562 68.5181
R32916 vss.n13562 vss.n13552 68.5181
R32917 vss.n13560 vss.n13548 68.5181
R32918 vss.n13604 vss.n13548 68.5181
R32919 vss.n13620 vss.n13528 68.5181
R32920 vss.n13629 vss.n13528 68.5181
R32921 vss.n13639 vss.n13636 68.5181
R32922 vss.n13636 vss.n13520 68.5181
R32923 vss.n13519 vss.n13510 68.5181
R32924 vss.n13654 vss.n13519 68.5181
R32925 vss.n13674 vss.n13489 68.5181
R32926 vss.n13683 vss.n13489 68.5181
R32927 vss.n13694 vss.n13691 68.5181
R32928 vss.n13691 vss.n13481 68.5181
R32929 vss.n13480 vss.n13471 68.5181
R32930 vss.n13705 vss.n13480 68.5181
R32931 vss.n13725 vss.n13448 68.5181
R32932 vss.n13734 vss.n13448 68.5181
R32933 vss.n13744 vss.n13741 68.5181
R32934 vss.n13741 vss.n13440 68.5181
R32935 vss.n13439 vss.n13430 68.5181
R32936 vss.n13759 vss.n13439 68.5181
R32937 vss.n13779 vss.n13409 68.5181
R32938 vss.n13788 vss.n13409 68.5181
R32939 vss.n13799 vss.n13796 68.5181
R32940 vss.n13796 vss.n13401 68.5181
R32941 vss.n13400 vss.n13391 68.5181
R32942 vss.n13810 vss.n13400 68.5181
R32943 vss.n13830 vss.n13368 68.5181
R32944 vss.n13839 vss.n13368 68.5181
R32945 vss.n13849 vss.n13846 68.5181
R32946 vss.n13846 vss.n13360 68.5181
R32947 vss.n13359 vss.n13350 68.5181
R32948 vss.n13864 vss.n13359 68.5181
R32949 vss.n13884 vss.n13329 68.5181
R32950 vss.n13893 vss.n13329 68.5181
R32951 vss.n14669 vss.n14657 68.5181
R32952 vss.n14669 vss.n14668 68.5181
R32953 vss.n14674 vss.n14656 68.5181
R32954 vss.n14656 vss.n14646 68.5181
R32955 vss.n14654 vss.n197 68.5181
R32956 vss.n14679 vss.n197 68.5181
R32957 vss.n14555 vss.n14548 68.5181
R32958 vss.n14548 vss.n234 68.5181
R32959 vss.n14546 vss.n232 68.5181
R32960 vss.n14560 vss.n232 68.5181
R32961 vss.n247 vss.n242 68.5181
R32962 vss.n248 vss.n247 68.5181
R32963 vss.n14474 vss.n14462 68.5181
R32964 vss.n14474 vss.n14473 68.5181
R32965 vss.n14479 vss.n14461 68.5181
R32966 vss.n14461 vss.n14451 68.5181
R32967 vss.n14459 vss.n256 68.5181
R32968 vss.n14484 vss.n256 68.5181
R32969 vss.n14360 vss.n14353 68.5181
R32970 vss.n14353 vss.n293 68.5181
R32971 vss.n14351 vss.n291 68.5181
R32972 vss.n14365 vss.n291 68.5181
R32973 vss.n306 vss.n301 68.5181
R32974 vss.n307 vss.n306 68.5181
R32975 vss.n14279 vss.n14267 68.5181
R32976 vss.n14279 vss.n14278 68.5181
R32977 vss.n14284 vss.n14266 68.5181
R32978 vss.n14266 vss.n14256 68.5181
R32979 vss.n14264 vss.n315 68.5181
R32980 vss.n14289 vss.n315 68.5181
R32981 vss.n14325 vss.n14313 68.5181
R32982 vss.n14325 vss.n14324 68.5181
R32983 vss.n14330 vss.n14312 68.5181
R32984 vss.n14312 vss.n14302 68.5181
R32985 vss.n14310 vss.n14299 68.5181
R32986 vss.n14335 vss.n14299 68.5181
R32987 vss.n14406 vss.n14399 68.5181
R32988 vss.n14399 vss.n14372 68.5181
R32989 vss.n14397 vss.n14370 68.5181
R32990 vss.n14411 vss.n14370 68.5181
R32991 vss.n14385 vss.n14380 68.5181
R32992 vss.n14386 vss.n14385 68.5181
R32993 vss.n14520 vss.n14508 68.5181
R32994 vss.n14520 vss.n14519 68.5181
R32995 vss.n14525 vss.n14507 68.5181
R32996 vss.n14507 vss.n14497 68.5181
R32997 vss.n14505 vss.n14494 68.5181
R32998 vss.n14530 vss.n14494 68.5181
R32999 vss.n14601 vss.n14594 68.5181
R33000 vss.n14594 vss.n14567 68.5181
R33001 vss.n14592 vss.n14565 68.5181
R33002 vss.n14606 vss.n14565 68.5181
R33003 vss.n14580 vss.n14575 68.5181
R33004 vss.n14581 vss.n14580 68.5181
R33005 vss.n14715 vss.n14703 68.5181
R33006 vss.n14715 vss.n14714 68.5181
R33007 vss.n14720 vss.n14702 68.5181
R33008 vss.n14702 vss.n14692 68.5181
R33009 vss.n14700 vss.n14689 68.5181
R33010 vss.n14725 vss.n14689 68.5181
R33011 vss.n14750 vss.n14743 68.5181
R33012 vss.n14743 vss.n157 68.5181
R33013 vss.n14741 vss.n155 68.5181
R33014 vss.n14755 vss.n155 68.5181
R33015 vss.n170 vss.n165 68.5181
R33016 vss.n171 vss.n170 68.5181
R33017 vss.n13904 vss.n13901 68.5181
R33018 vss.n13901 vss.n13321 68.5181
R33019 vss.n13317 vss.n13308 68.5181
R33020 vss.n13912 vss.n13317 68.5181
R33021 vss.n13917 vss.n13307 68.5181
R33022 vss.n13315 vss.n13307 68.5181
R33023 vss.n13883 vss.n13333 68.5181
R33024 vss.n13333 vss.n13330 68.5181
R33025 vss.n13341 vss.n13334 68.5181
R33026 vss.n13878 vss.n13341 68.5181
R33027 vss.n13869 vss.n13349 68.5181
R33028 vss.n13357 vss.n13349 68.5181
R33029 vss.n13829 vss.n13374 68.5181
R33030 vss.n13374 vss.n13371 68.5181
R33031 vss.n13382 vss.n13375 68.5181
R33032 vss.n13824 vss.n13382 68.5181
R33033 vss.n13815 vss.n13390 68.5181
R33034 vss.n13398 vss.n13390 68.5181
R33035 vss.n13778 vss.n13413 68.5181
R33036 vss.n13413 vss.n13410 68.5181
R33037 vss.n13421 vss.n13414 68.5181
R33038 vss.n13773 vss.n13421 68.5181
R33039 vss.n13764 vss.n13429 68.5181
R33040 vss.n13437 vss.n13429 68.5181
R33041 vss.n13724 vss.n13454 68.5181
R33042 vss.n13454 vss.n13451 68.5181
R33043 vss.n13462 vss.n13455 68.5181
R33044 vss.n13719 vss.n13462 68.5181
R33045 vss.n13710 vss.n13470 68.5181
R33046 vss.n13478 vss.n13470 68.5181
R33047 vss.n13673 vss.n13493 68.5181
R33048 vss.n13493 vss.n13490 68.5181
R33049 vss.n13501 vss.n13494 68.5181
R33050 vss.n13668 vss.n13501 68.5181
R33051 vss.n13659 vss.n13509 68.5181
R33052 vss.n13517 vss.n13509 68.5181
R33053 vss.n13619 vss.n13534 68.5181
R33054 vss.n13534 vss.n13531 68.5181
R33055 vss.n13542 vss.n13535 68.5181
R33056 vss.n13614 vss.n13542 68.5181
R33057 vss.n629 vss.n622 68.5181
R33058 vss.n636 vss.n629 68.5181
R33059 vss.n644 vss.n621 68.5181
R33060 vss.n621 vss.n618 68.5181
R33061 vss.n645 vss.n617 68.5181
R33062 vss.n654 vss.n617 68.5181
R33063 vss.n810 vss.n809 68.5181
R33064 vss.n809 vss.n804 68.5181
R33065 vss.n13234 vss.n794 68.5181
R33066 vss.n13220 vss.n794 68.5181
R33067 vss.n13222 vss.n796 68.5181
R33068 vss.n13229 vss.n13222 68.5181
R33069 vss.n1669 vss.n1668 68.5181
R33070 vss.n1668 vss.n1663 68.5181
R33071 vss.n1693 vss.n1653 68.5181
R33072 vss.n1679 vss.n1653 68.5181
R33073 vss.n1681 vss.n1655 68.5181
R33074 vss.n1688 vss.n1681 68.5181
R33075 vss.n1622 vss.n1621 68.5181
R33076 vss.n1621 vss.n1616 68.5181
R33077 vss.n1646 vss.n1606 68.5181
R33078 vss.n1632 vss.n1606 68.5181
R33079 vss.n1634 vss.n1608 68.5181
R33080 vss.n1641 vss.n1634 68.5181
R33081 vss.n1374 vss.n1373 68.5181
R33082 vss.n1373 vss.n1368 68.5181
R33083 vss.n1398 vss.n1358 68.5181
R33084 vss.n1384 vss.n1358 68.5181
R33085 vss.n1386 vss.n1360 68.5181
R33086 vss.n1393 vss.n1386 68.5181
R33087 vss.n1175 vss.n1174 68.5181
R33088 vss.n1174 vss.n1169 68.5181
R33089 vss.n1199 vss.n1159 68.5181
R33090 vss.n1185 vss.n1159 68.5181
R33091 vss.n1187 vss.n1161 68.5181
R33092 vss.n1194 vss.n1187 68.5181
R33093 vss.n1327 vss.n1326 68.5181
R33094 vss.n1326 vss.n1321 68.5181
R33095 vss.n1351 vss.n1311 68.5181
R33096 vss.n1337 vss.n1311 68.5181
R33097 vss.n1339 vss.n1313 68.5181
R33098 vss.n1346 vss.n1339 68.5181
R33099 vss.n1066 vss.n1065 68.5181
R33100 vss.n1065 vss.n1060 68.5181
R33101 vss.n1090 vss.n1050 68.5181
R33102 vss.n1076 vss.n1050 68.5181
R33103 vss.n1078 vss.n1052 68.5181
R33104 vss.n1085 vss.n1078 68.5181
R33105 vss.n1459 vss.n1458 68.5181
R33106 vss.n1458 vss.n1453 68.5181
R33107 vss.n1483 vss.n1443 68.5181
R33108 vss.n1469 vss.n1443 68.5181
R33109 vss.n1471 vss.n1445 68.5181
R33110 vss.n1478 vss.n1471 68.5181
R33111 vss.n1539 vss.n1538 68.5181
R33112 vss.n1538 vss.n1533 68.5181
R33113 vss.n1564 vss.n1523 68.5181
R33114 vss.n1549 vss.n1523 68.5181
R33115 vss.n1551 vss.n1525 68.5181
R33116 vss.n1559 vss.n1551 68.5181
R33117 vss.n821 vss.n820 68.5181
R33118 vss.n829 vss.n821 68.5181
R33119 vss.n13952 vss.n595 68.5181
R33120 vss.n605 vss.n595 68.5181
R33121 vss.n607 vss.n597 68.5181
R33122 vss.n13947 vss.n607 68.5181
R33123 vss.n896 vss.n878 68.5181
R33124 vss.n914 vss.n878 68.5181
R33125 vss.n892 vss.n889 68.5181
R33126 vss.n889 vss.n879 68.5181
R33127 vss.n902 vss.n884 68.5181
R33128 vss.n908 vss.n884 68.5181
R33129 vss.n524 vss.n519 68.5181
R33130 vss.n14013 vss.n524 68.5181
R33131 vss.n14024 vss.n517 68.5181
R33132 vss.n14011 vss.n517 68.5181
R33133 vss.n534 vss.n533 68.5181
R33134 vss.n533 vss.n526 68.5181
R33135 vss.n549 vss.n540 68.5181
R33136 vss.n13997 vss.n540 68.5181
R33137 vss.n664 vss.n663 68.5181
R33138 vss.n674 vss.n664 68.5181
R33139 vss.n573 vss.n572 68.5181
R33140 vss.n572 vss.n565 68.5181
R33141 vss.n588 vss.n579 68.5181
R33142 vss.n13962 vss.n579 68.5181
R33143 vss.n767 vss.n766 68.5181
R33144 vss.n773 vss.n767 68.5181
R33145 vss.n755 vss.n746 68.5181
R33146 vss.n13245 vss.n746 68.5181
R33147 vss.n1724 vss.n1719 68.5181
R33148 vss.n1733 vss.n1724 68.5181
R33149 vss.n1739 vss.n1710 68.5181
R33150 vss.n1744 vss.n1710 68.5181
R33151 vss.n1760 vss.n1759 68.5181
R33152 vss.n1759 vss.n1752 68.5181
R33153 vss.n1766 vss.n1765 68.5181
R33154 vss.n1774 vss.n1766 68.5181
R33155 vss.n1810 vss.n1267 68.5181
R33156 vss.n1815 vss.n1267 68.5181
R33157 vss.n1253 vss.n1252 68.5181
R33158 vss.n1256 vss.n1253 68.5181
R33159 vss.n1228 vss.n1223 68.5181
R33160 vss.n1837 vss.n1228 68.5181
R33161 vss.n1843 vss.n1214 68.5181
R33162 vss.n1848 vss.n1214 68.5181
R33163 vss.n1864 vss.n1863 68.5181
R33164 vss.n1863 vss.n1856 68.5181
R33165 vss.n1870 vss.n1869 68.5181
R33166 vss.n1878 vss.n1870 68.5181
R33167 vss.n1914 vss.n1149 68.5181
R33168 vss.n1919 vss.n1149 68.5181
R33169 vss.n1935 vss.n1934 68.5181
R33170 vss.n1934 vss.n1927 68.5181
R33171 vss.n1941 vss.n1940 68.5181
R33172 vss.n1949 vss.n1941 68.5181
R33173 vss.n13292 vss.n693 68.5181
R33174 vss.n13297 vss.n693 68.5181
R33175 vss.n726 vss.n725 68.5181
R33176 vss.n725 vss.n718 68.5181
R33177 vss.n2001 vss.n2000 68.5181
R33178 vss.n2000 vss.n1995 68.5181
R33179 vss.n2025 vss.n1985 68.5181
R33180 vss.n2011 vss.n1985 68.5181
R33181 vss.n2013 vss.n1987 68.5181
R33182 vss.n2020 vss.n2013 68.5181
R33183 vss.n13194 vss.n13161 68.5181
R33184 vss.n13194 vss.n13193 68.5181
R33185 vss.n13175 vss.n13174 68.5181
R33186 vss.n13174 vss.n13167 68.5181
R33187 vss.n9622 vss.n9615 68.5181
R33188 vss.n9615 vss.n9588 68.5181
R33189 vss.n9613 vss.n9586 68.5181
R33190 vss.n9627 vss.n9586 68.5181
R33191 vss.n9601 vss.n9596 68.5181
R33192 vss.n9602 vss.n9601 68.5181
R33193 vss.n9166 vss.n9165 68.5181
R33194 vss.n9165 vss.n9160 68.5181
R33195 vss.n9191 vss.n9150 68.5181
R33196 vss.n9177 vss.n9150 68.5181
R33197 vss.n9179 vss.n9152 68.5181
R33198 vss.n9186 vss.n9179 68.5181
R33199 vss.n9130 vss.n9101 68.5181
R33200 vss.n9135 vss.n9101 68.5181
R33201 vss.n9129 vss.n9111 68.5181
R33202 vss.n9111 vss.n9102 68.5181
R33203 vss.n9144 vss.n6547 68.5181
R33204 vss.n9091 vss.n6547 68.5181
R33205 vss.n9198 vss.n6531 68.5181
R33206 vss.n9203 vss.n6531 68.5181
R33207 vss.n9197 vss.n6541 68.5181
R33208 vss.n6541 vss.n6532 68.5181
R33209 vss.n9214 vss.n6523 68.5181
R33210 vss.n6523 vss.n6513 68.5181
R33211 vss.n6497 vss.n6492 68.5181
R33212 vss.n9235 vss.n6497 68.5181
R33213 vss.n9246 vss.n6490 68.5181
R33214 vss.n9233 vss.n6490 68.5181
R33215 vss.n6883 vss.n6863 68.5181
R33216 vss.n6863 vss.n6853 68.5181
R33217 vss.n7035 vss.n6830 68.5181
R33218 vss.n7040 vss.n6830 68.5181
R33219 vss.n7034 vss.n6840 68.5181
R33220 vss.n6840 vss.n6831 68.5181
R33221 vss.n7051 vss.n6812 68.5181
R33222 vss.n6812 vss.n6802 68.5181
R33223 vss.n6725 vss.n6720 68.5181
R33224 vss.n7072 vss.n6725 68.5181
R33225 vss.n7083 vss.n6718 68.5181
R33226 vss.n7070 vss.n6718 68.5181
R33227 vss.n6774 vss.n6738 68.5181
R33228 vss.n6738 vss.n6731 68.5181
R33229 vss.n7226 vss.n6584 68.5181
R33230 vss.n7231 vss.n6584 68.5181
R33231 vss.n7225 vss.n6594 68.5181
R33232 vss.n6594 vss.n6585 68.5181
R33233 vss.n9506 vss.n6130 68.5181
R33234 vss.n6130 vss.n6120 68.5181
R33235 vss.n6103 vss.n6098 68.5181
R33236 vss.n9527 vss.n6103 68.5181
R33237 vss.n9538 vss.n6096 68.5181
R33238 vss.n9525 vss.n6096 68.5181
R33239 vss.n9541 vss.n6091 68.5181
R33240 vss.n6091 vss.n6081 68.5181
R33241 vss.n9463 vss.n9459 68.5181
R33242 vss.n9468 vss.n9459 68.5181
R33243 vss.n9451 vss.n6055 68.5181
R33244 vss.n9451 vss.n9449 68.5181
R33245 vss.n9473 vss.n9448 68.5181
R33246 vss.n9482 vss.n9448 68.5181
R33247 vss.n8032 vss.n8025 68.5181
R33248 vss.n8038 vss.n8025 68.5181
R33249 vss.n8022 vss.n8017 68.5181
R33250 vss.n8022 vss.n6005 68.5181
R33251 vss.n8048 vss.n8016 68.5181
R33252 vss.n8043 vss.n8016 68.5181
R33253 vss.n8135 vss.n8134 68.5181
R33254 vss.n8134 vss.n8133 68.5181
R33255 vss.n8125 vss.n6002 68.5181
R33256 vss.n9642 vss.n6002 68.5181
R33257 vss.n9654 vss.n5989 68.5181
R33258 vss.n9654 vss.n9653 68.5181
R33259 vss.n9659 vss.n5988 68.5181
R33260 vss.n5988 vss.n5978 68.5181
R33261 vss.n5986 vss.n5977 68.5181
R33262 vss.n9664 vss.n5977 68.5181
R33263 vss.n8147 vss.n5998 68.5181
R33264 vss.n6001 vss.n5998 68.5181
R33265 vss.n8164 vss.n8103 68.5181
R33266 vss.n8169 vss.n8103 68.5181
R33267 vss.n8163 vss.n8113 68.5181
R33268 vss.n8113 vss.n8104 68.5181
R33269 vss.n8119 vss.n8114 68.5181
R33270 vss.n8158 vss.n8119 68.5181
R33271 vss.n8090 vss.n8056 68.5181
R33272 vss.n8095 vss.n8056 68.5181
R33273 vss.n8089 vss.n8069 68.5181
R33274 vss.n8069 vss.n8060 68.5181
R33275 vss.n8075 vss.n8070 68.5181
R33276 vss.n8084 vss.n8075 68.5181
R33277 vss.n8239 vss.n8232 68.5181
R33278 vss.n8232 vss.n7994 68.5181
R33279 vss.n8230 vss.n7992 68.5181
R33280 vss.n8244 vss.n7992 68.5181
R33281 vss.n8007 vss.n8002 68.5181
R33282 vss.n8008 vss.n8007 68.5181
R33283 vss.n8204 vss.n8192 68.5181
R33284 vss.n8204 vss.n8203 68.5181
R33285 vss.n8209 vss.n8191 68.5181
R33286 vss.n8191 vss.n8181 68.5181
R33287 vss.n8189 vss.n8178 68.5181
R33288 vss.n8214 vss.n8178 68.5181
R33289 vss.n8992 vss.n7315 68.5181
R33290 vss.n8992 vss.n8991 68.5181
R33291 vss.n8997 vss.n7314 68.5181
R33292 vss.n7314 vss.n7304 68.5181
R33293 vss.n7312 vss.n7303 68.5181
R33294 vss.n9002 vss.n7303 68.5181
R33295 vss.n8730 vss.n8723 68.5181
R33296 vss.n8723 vss.n7851 68.5181
R33297 vss.n8721 vss.n7849 68.5181
R33298 vss.n8735 vss.n7849 68.5181
R33299 vss.n7864 vss.n7859 68.5181
R33300 vss.n7865 vss.n7864 68.5181
R33301 vss.n7804 vss.n7797 68.5181
R33302 vss.n7797 vss.n7770 68.5181
R33303 vss.n7795 vss.n7768 68.5181
R33304 vss.n7809 vss.n7768 68.5181
R33305 vss.n7783 vss.n7778 68.5181
R33306 vss.n7784 vss.n7783 68.5181
R33307 vss.n8768 vss.n8756 68.5181
R33308 vss.n8768 vss.n8767 68.5181
R33309 vss.n8773 vss.n8755 68.5181
R33310 vss.n8755 vss.n8745 68.5181
R33311 vss.n8753 vss.n7686 68.5181
R33312 vss.n8778 vss.n7686 68.5181
R33313 vss.n8849 vss.n8842 68.5181
R33314 vss.n8842 vss.n7664 68.5181
R33315 vss.n8840 vss.n7662 68.5181
R33316 vss.n8854 vss.n7662 68.5181
R33317 vss.n7677 vss.n7672 68.5181
R33318 vss.n7678 vss.n7677 68.5181
R33319 vss.n8814 vss.n8802 68.5181
R33320 vss.n8814 vss.n8813 68.5181
R33321 vss.n8819 vss.n8801 68.5181
R33322 vss.n8801 vss.n8791 68.5181
R33323 vss.n8799 vss.n8788 68.5181
R33324 vss.n8824 vss.n8788 68.5181
R33325 vss.n8887 vss.n8875 68.5181
R33326 vss.n8887 vss.n8886 68.5181
R33327 vss.n8892 vss.n8874 68.5181
R33328 vss.n8874 vss.n8864 68.5181
R33329 vss.n8872 vss.n7543 68.5181
R33330 vss.n8897 vss.n7543 68.5181
R33331 vss.n8540 vss.n8499 68.5181
R33332 vss.n8540 vss.n8539 68.5181
R33333 vss.n8515 vss.n8514 68.5181
R33334 vss.n8514 vss.n8503 68.5181
R33335 vss.n9023 vss.n7283 68.5181
R33336 vss.n9023 vss.n9022 68.5181
R33337 vss.n9028 vss.n7282 68.5181
R33338 vss.n7282 vss.n7272 68.5181
R33339 vss.n7280 vss.n7271 68.5181
R33340 vss.n9033 vss.n7271 68.5181
R33341 vss.n9014 vss.n7293 68.5181
R33342 vss.n9014 vss.n9013 68.5181
R33343 vss.n8273 vss.n8270 68.5181
R33344 vss.n8270 vss.n8259 68.5181
R33345 vss.n8268 vss.n7903 68.5181
R33346 vss.n8278 vss.n7903 68.5181
R33347 vss.n8294 vss.n7881 68.5181
R33348 vss.n8299 vss.n7881 68.5181
R33349 vss.n8293 vss.n7891 68.5181
R33350 vss.n7891 vss.n7882 68.5181
R33351 vss.n7897 vss.n7892 68.5181
R33352 vss.n8288 vss.n7897 68.5181
R33353 vss.n8700 vss.n7870 68.5181
R33354 vss.n8705 vss.n7870 68.5181
R33355 vss.n8699 vss.n8310 68.5181
R33356 vss.n8310 vss.n7874 68.5181
R33357 vss.n8316 vss.n8311 68.5181
R33358 vss.n8694 vss.n8316 68.5181
R33359 vss.n8677 vss.n8343 68.5181
R33360 vss.n8346 vss.n8343 68.5181
R33361 vss.n8341 vss.n8338 68.5181
R33362 vss.n8338 vss.n8330 68.5181
R33363 vss.n8685 vss.n8321 68.5181
R33364 vss.n8685 vss.n8684 68.5181
R33365 vss.n8670 vss.n8351 68.5181
R33366 vss.n8670 vss.n8669 68.5181
R33367 vss.n8656 vss.n8653 68.5181
R33368 vss.n8653 vss.n8352 68.5181
R33369 vss.n8652 vss.n8361 68.5181
R33370 vss.n8647 vss.n8361 68.5181
R33371 vss.n8634 vss.n8393 68.5181
R33372 vss.n8396 vss.n8393 68.5181
R33373 vss.n8391 vss.n8388 68.5181
R33374 vss.n8388 vss.n8380 68.5181
R33375 vss.n8642 vss.n8366 68.5181
R33376 vss.n8642 vss.n8641 68.5181
R33377 vss.n8627 vss.n8401 68.5181
R33378 vss.n8627 vss.n8626 68.5181
R33379 vss.n8612 vss.n8609 68.5181
R33380 vss.n8609 vss.n8405 68.5181
R33381 vss.n8608 vss.n8414 68.5181
R33382 vss.n8603 vss.n8414 68.5181
R33383 vss.n8590 vss.n8441 68.5181
R33384 vss.n8444 vss.n8441 68.5181
R33385 vss.n8439 vss.n8436 68.5181
R33386 vss.n8436 vss.n8428 68.5181
R33387 vss.n8598 vss.n8419 68.5181
R33388 vss.n8598 vss.n8597 68.5181
R33389 vss.n8583 vss.n8449 68.5181
R33390 vss.n8583 vss.n8582 68.5181
R33391 vss.n8569 vss.n8566 68.5181
R33392 vss.n8566 vss.n8450 68.5181
R33393 vss.n8565 vss.n8459 68.5181
R33394 vss.n8560 vss.n8459 68.5181
R33395 vss.n8547 vss.n8491 68.5181
R33396 vss.n8494 vss.n8491 68.5181
R33397 vss.n8489 vss.n8486 68.5181
R33398 vss.n8486 vss.n8478 68.5181
R33399 vss.n8555 vss.n8464 68.5181
R33400 vss.n8555 vss.n8554 68.5181
R33401 vss.n8521 vss.n8507 68.5181
R33402 vss.n8526 vss.n8507 68.5181
R33403 vss.n8968 vss.n8961 68.5181
R33404 vss.n8961 vss.n7475 68.5181
R33405 vss.n8959 vss.n7473 68.5181
R33406 vss.n8973 vss.n7473 68.5181
R33407 vss.n7488 vss.n7483 68.5181
R33408 vss.n7489 vss.n7488 68.5181
R33409 vss.n8933 vss.n8921 68.5181
R33410 vss.n8933 vss.n8932 68.5181
R33411 vss.n8938 vss.n8920 68.5181
R33412 vss.n8920 vss.n8910 68.5181
R33413 vss.n8918 vss.n8907 68.5181
R33414 vss.n8943 vss.n8907 68.5181
R33415 vss.n7521 vss.n7509 68.5181
R33416 vss.n7521 vss.n7520 68.5181
R33417 vss.n7526 vss.n7508 68.5181
R33418 vss.n7508 vss.n7498 68.5181
R33419 vss.n7506 vss.n7494 68.5181
R33420 vss.n7531 vss.n7494 68.5181
R33421 vss.n7581 vss.n7574 68.5181
R33422 vss.n7574 vss.n7547 68.5181
R33423 vss.n7572 vss.n7545 68.5181
R33424 vss.n7586 vss.n7545 68.5181
R33425 vss.n7560 vss.n7555 68.5181
R33426 vss.n7561 vss.n7560 68.5181
R33427 vss.n7724 vss.n7717 68.5181
R33428 vss.n7717 vss.n7690 68.5181
R33429 vss.n7715 vss.n7688 68.5181
R33430 vss.n7729 vss.n7688 68.5181
R33431 vss.n7703 vss.n7698 68.5181
R33432 vss.n7704 vss.n7703 68.5181
R33433 vss.n7945 vss.n7938 68.5181
R33434 vss.n7938 vss.n7911 68.5181
R33435 vss.n7936 vss.n7909 68.5181
R33436 vss.n7950 vss.n7909 68.5181
R33437 vss.n7924 vss.n7919 68.5181
R33438 vss.n7925 vss.n7924 68.5181
R33439 vss.n6024 vss.n6023 68.5181
R33440 vss.n6023 vss.n6018 68.5181
R33441 vss.n6050 vss.n6008 68.5181
R33442 vss.n6035 vss.n6008 68.5181
R33443 vss.n6037 vss.n6010 68.5181
R33444 vss.n6045 vss.n6037 68.5181
R33445 vss.n7194 vss.n7193 68.5181
R33446 vss.n7193 vss.n7188 68.5181
R33447 vss.n7219 vss.n7178 68.5181
R33448 vss.n7205 vss.n7178 68.5181
R33449 vss.n7207 vss.n7180 68.5181
R33450 vss.n7214 vss.n7207 68.5181
R33451 vss.n6689 vss.n6688 68.5181
R33452 vss.n6688 vss.n6683 68.5181
R33453 vss.n6714 vss.n6673 68.5181
R33454 vss.n6700 vss.n6673 68.5181
R33455 vss.n6702 vss.n6675 68.5181
R33456 vss.n6709 vss.n6702 68.5181
R33457 vss.n6645 vss.n6644 68.5181
R33458 vss.n6644 vss.n6639 68.5181
R33459 vss.n6670 vss.n6629 68.5181
R33460 vss.n6656 vss.n6629 68.5181
R33461 vss.n6658 vss.n6631 68.5181
R33462 vss.n6665 vss.n6658 68.5181
R33463 vss.n7003 vss.n7002 68.5181
R33464 vss.n7002 vss.n6997 68.5181
R33465 vss.n7028 vss.n6987 68.5181
R33466 vss.n7014 vss.n6987 68.5181
R33467 vss.n7016 vss.n6989 68.5181
R33468 vss.n7023 vss.n7016 68.5181
R33469 vss.n6463 vss.n6462 68.5181
R33470 vss.n6462 vss.n6457 68.5181
R33471 vss.n6488 vss.n6447 68.5181
R33472 vss.n6474 vss.n6447 68.5181
R33473 vss.n6476 vss.n6449 68.5181
R33474 vss.n6483 vss.n6476 68.5181
R33475 vss.n6418 vss.n6417 68.5181
R33476 vss.n6417 vss.n6412 68.5181
R33477 vss.n6443 vss.n6402 68.5181
R33478 vss.n6429 vss.n6402 68.5181
R33479 vss.n6431 vss.n6404 68.5181
R33480 vss.n6438 vss.n6431 68.5181
R33481 vss.n6340 vss.n6339 68.5181
R33482 vss.n6339 vss.n6334 68.5181
R33483 vss.n6365 vss.n6324 68.5181
R33484 vss.n6351 vss.n6324 68.5181
R33485 vss.n6353 vss.n6326 68.5181
R33486 vss.n6360 vss.n6353 68.5181
R33487 vss.n6954 vss.n6953 68.5181
R33488 vss.n6953 vss.n6948 68.5181
R33489 vss.n6979 vss.n6938 68.5181
R33490 vss.n6965 vss.n6938 68.5181
R33491 vss.n6967 vss.n6940 68.5181
R33492 vss.n6974 vss.n6967 68.5181
R33493 vss.n7143 vss.n7142 68.5181
R33494 vss.n7142 vss.n7137 68.5181
R33495 vss.n7168 vss.n7127 68.5181
R33496 vss.n7154 vss.n7127 68.5181
R33497 vss.n7156 vss.n7129 68.5181
R33498 vss.n7163 vss.n7156 68.5181
R33499 vss.n6151 vss.n6150 68.5181
R33500 vss.n6150 vss.n6145 68.5181
R33501 vss.n9501 vss.n6135 68.5181
R33502 vss.n6162 vss.n6135 68.5181
R33503 vss.n6164 vss.n6137 68.5181
R33504 vss.n9496 vss.n6164 68.5181
R33505 vss.n9415 vss.n9408 68.5181
R33506 vss.n9423 vss.n9415 68.5181
R33507 vss.n9430 vss.n9407 68.5181
R33508 vss.n9407 vss.n9404 68.5181
R33509 vss.n9431 vss.n9403 68.5181
R33510 vss.n9440 vss.n9403 68.5181
R33511 vss.n6063 vss.n6058 68.5181
R33512 vss.n9562 vss.n6063 68.5181
R33513 vss.n9573 vss.n6056 68.5181
R33514 vss.n9560 vss.n6056 68.5181
R33515 vss.n6074 vss.n6073 68.5181
R33516 vss.n6073 vss.n6066 68.5181
R33517 vss.n6089 vss.n6080 68.5181
R33518 vss.n9546 vss.n6080 68.5181
R33519 vss.n7252 vss.n7251 68.5181
R33520 vss.n7262 vss.n7252 68.5181
R33521 vss.n6113 vss.n6112 68.5181
R33522 vss.n6112 vss.n6105 68.5181
R33523 vss.n6128 vss.n6119 68.5181
R33524 vss.n9511 vss.n6119 68.5181
R33525 vss.n6579 vss.n6578 68.5181
R33526 vss.n7243 vss.n6579 68.5181
R33527 vss.n6754 vss.n6753 68.5181
R33528 vss.n6757 vss.n6754 68.5181
R33529 vss.n6744 vss.n6739 68.5181
R33530 vss.n6769 vss.n6744 68.5181
R33531 vss.n6775 vss.n6730 68.5181
R33532 vss.n6780 vss.n6730 68.5181
R33533 vss.n6796 vss.n6795 68.5181
R33534 vss.n6795 vss.n6788 68.5181
R33535 vss.n6810 vss.n6801 68.5181
R33536 vss.n7056 vss.n6801 68.5181
R33537 vss.n6820 vss.n6813 68.5181
R33538 vss.n6822 vss.n6820 68.5181
R33539 vss.n6846 vss.n6841 68.5181
R33540 vss.n6898 vss.n6846 68.5181
R33541 vss.n6861 vss.n6852 68.5181
R33542 vss.n6888 vss.n6852 68.5181
R33543 vss.n6871 vss.n6864 68.5181
R33544 vss.n6873 vss.n6871 68.5181
R33545 vss.n6507 vss.n6506 68.5181
R33546 vss.n6506 vss.n6499 68.5181
R33547 vss.n6521 vss.n6512 68.5181
R33548 vss.n9219 vss.n6512 68.5181
R33549 vss.n6561 vss.n6524 68.5181
R33550 vss.n6563 vss.n6561 68.5181
R33551 vss.n9072 vss.n9071 68.5181
R33552 vss.n9075 vss.n9072 68.5181
R33553 vss.n9063 vss.n9062 68.5181
R33554 vss.n9062 vss.n9055 68.5181
R33555 vss.n9054 vss.n6549 68.5181
R33556 vss.n9093 vss.n9054 68.5181
R33557 vss.n9117 vss.n9112 68.5181
R33558 vss.n9124 vss.n9117 68.5181
R33559 vss.n9336 vss.n9335 68.5181
R33560 vss.n9335 vss.n9330 68.5181
R33561 vss.n9361 vss.n9320 68.5181
R33562 vss.n9347 vss.n9320 68.5181
R33563 vss.n9349 vss.n9322 68.5181
R33564 vss.n9356 vss.n9349 68.5181
R33565 vss.n6200 vss.n6193 68.5181
R33566 vss.n6208 vss.n6200 68.5181
R33567 vss.n9368 vss.n6192 68.5181
R33568 vss.n6192 vss.n6189 68.5181
R33569 vss.n9369 vss.n6188 68.5181
R33570 vss.n9378 vss.n6188 68.5181
R33571 vss.n9676 vss.n5965 68.5181
R33572 vss.n5965 vss.n5939 68.5181
R33573 vss.n5963 vss.n5937 68.5181
R33574 vss.n9681 vss.n5937 68.5181
R33575 vss.n5952 vss.n5947 68.5181
R33576 vss.n5953 vss.n5952 68.5181
R33577 vss.n9723 vss.n9715 68.5181
R33578 vss.n9715 vss.n9687 68.5181
R33579 vss.n9713 vss.n9685 68.5181
R33580 vss.n9728 vss.n9685 68.5181
R33581 vss.n9700 vss.n9695 68.5181
R33582 vss.n9701 vss.n9700 68.5181
R33583 vss.n10004 vss.n2586 68.5181
R33584 vss.n2586 vss.n2560 68.5181
R33585 vss.n2584 vss.n2558 68.5181
R33586 vss.n10009 vss.n2558 68.5181
R33587 vss.n2573 vss.n2568 68.5181
R33588 vss.n2574 vss.n2573 68.5181
R33589 vss.n9881 vss.n2759 68.5181
R33590 vss.n9881 vss.n9880 68.5181
R33591 vss.n9886 vss.n2758 68.5181
R33592 vss.n2758 vss.n2748 68.5181
R33593 vss.n2756 vss.n2747 68.5181
R33594 vss.n9891 vss.n2747 68.5181
R33595 vss.n3301 vss.n3292 68.5181
R33596 vss.n3292 vss.n3265 68.5181
R33597 vss.n3291 vss.n3263 68.5181
R33598 vss.n3306 vss.n3263 68.5181
R33599 vss.n3278 vss.n3273 68.5181
R33600 vss.n3279 vss.n3278 68.5181
R33601 vss.n9752 vss.n9751 68.5181
R33602 vss.n9751 vss.n9746 68.5181
R33603 vss.n9772 vss.n9744 68.5181
R33604 vss.n9784 vss.n9744 68.5181
R33605 vss.n9764 vss.n9754 68.5181
R33606 vss.n9765 vss.n9764 68.5181
R33607 vss.n3192 vss.n3191 68.5181
R33608 vss.n3191 vss.n3186 68.5181
R33609 vss.n3212 vss.n3184 68.5181
R33610 vss.n3224 vss.n3184 68.5181
R33611 vss.n3204 vss.n3194 68.5181
R33612 vss.n3205 vss.n3204 68.5181
R33613 vss.n3014 vss.n3013 68.5181
R33614 vss.n3013 vss.n3009 68.5181
R33615 vss.n3008 vss.n2999 68.5181
R33616 vss.n9794 vss.n3008 68.5181
R33617 vss.n9799 vss.n2998 68.5181
R33618 vss.n3006 vss.n2998 68.5181
R33619 vss.n5222 vss.n5221 68.5181
R33620 vss.n5221 vss.n5216 68.5181
R33621 vss.n5242 vss.n5214 68.5181
R33622 vss.n5254 vss.n5214 68.5181
R33623 vss.n5234 vss.n5224 68.5181
R33624 vss.n5235 vss.n5234 68.5181
R33625 vss.n3035 vss.n3034 68.5181
R33626 vss.n3034 vss.n3029 68.5181
R33627 vss.n3055 vss.n3027 68.5181
R33628 vss.n3067 vss.n3027 68.5181
R33629 vss.n3047 vss.n3037 68.5181
R33630 vss.n3048 vss.n3047 68.5181
R33631 vss.n5092 vss.n5091 68.5181
R33632 vss.n5091 vss.n5086 68.5181
R33633 vss.n5112 vss.n5084 68.5181
R33634 vss.n5124 vss.n5084 68.5181
R33635 vss.n5104 vss.n5094 68.5181
R33636 vss.n5105 vss.n5104 68.5181
R33637 vss.n5281 vss.n5280 68.5181
R33638 vss.n5280 vss.n5275 68.5181
R33639 vss.n5301 vss.n5273 68.5181
R33640 vss.n5313 vss.n5273 68.5181
R33641 vss.n5293 vss.n5283 68.5181
R33642 vss.n5294 vss.n5293 68.5181
R33643 vss.n5009 vss.n5008 68.5181
R33644 vss.n5008 vss.n5003 68.5181
R33645 vss.n5029 vss.n5001 68.5181
R33646 vss.n5041 vss.n5001 68.5181
R33647 vss.n5021 vss.n5011 68.5181
R33648 vss.n5022 vss.n5021 68.5181
R33649 vss.n4890 vss.n4889 68.5181
R33650 vss.n4889 vss.n4884 68.5181
R33651 vss.n4910 vss.n4882 68.5181
R33652 vss.n4922 vss.n4882 68.5181
R33653 vss.n4902 vss.n4892 68.5181
R33654 vss.n4903 vss.n4902 68.5181
R33655 vss.n5393 vss.n5352 68.5181
R33656 vss.n5393 vss.n5392 68.5181
R33657 vss.n5368 vss.n5367 68.5181
R33658 vss.n5367 vss.n5356 68.5181
R33659 vss.n9915 vss.n2724 68.5181
R33660 vss.n9915 vss.n9914 68.5181
R33661 vss.n9920 vss.n2723 68.5181
R33662 vss.n2723 vss.n2713 68.5181
R33663 vss.n2721 vss.n2712 68.5181
R33664 vss.n9925 vss.n2712 68.5181
R33665 vss.n9906 vss.n2734 68.5181
R33666 vss.n9906 vss.n9905 68.5181
R33667 vss.n4657 vss.n4654 68.5181
R33668 vss.n4654 vss.n4643 68.5181
R33669 vss.n4652 vss.n4640 68.5181
R33670 vss.n4662 vss.n4640 68.5181
R33671 vss.n5617 vss.n4676 68.5181
R33672 vss.n5617 vss.n5616 68.5181
R33673 vss.n5622 vss.n4675 68.5181
R33674 vss.n4675 vss.n4634 68.5181
R33675 vss.n4673 vss.n4631 68.5181
R33676 vss.n5627 vss.n4631 68.5181
R33677 vss.n5608 vss.n4686 68.5181
R33678 vss.n5608 vss.n5607 68.5181
R33679 vss.n5594 vss.n5591 68.5181
R33680 vss.n5591 vss.n4687 68.5181
R33681 vss.n5590 vss.n4696 68.5181
R33682 vss.n5585 vss.n4696 68.5181
R33683 vss.n5572 vss.n4721 68.5181
R33684 vss.n4724 vss.n4721 68.5181
R33685 vss.n4719 vss.n4716 68.5181
R33686 vss.n4716 vss.n4708 68.5181
R33687 vss.n5580 vss.n4701 68.5181
R33688 vss.n5580 vss.n5579 68.5181
R33689 vss.n5565 vss.n4729 68.5181
R33690 vss.n5565 vss.n5564 68.5181
R33691 vss.n5551 vss.n5548 68.5181
R33692 vss.n5548 vss.n4730 68.5181
R33693 vss.n5547 vss.n4739 68.5181
R33694 vss.n5542 vss.n4739 68.5181
R33695 vss.n5529 vss.n4764 68.5181
R33696 vss.n4767 vss.n4764 68.5181
R33697 vss.n4762 vss.n4759 68.5181
R33698 vss.n4759 vss.n4751 68.5181
R33699 vss.n5537 vss.n4744 68.5181
R33700 vss.n5537 vss.n5536 68.5181
R33701 vss.n5522 vss.n4772 68.5181
R33702 vss.n5522 vss.n5521 68.5181
R33703 vss.n5508 vss.n5505 68.5181
R33704 vss.n5505 vss.n4773 68.5181
R33705 vss.n5504 vss.n4782 68.5181
R33706 vss.n5499 vss.n4782 68.5181
R33707 vss.n5486 vss.n4807 68.5181
R33708 vss.n4810 vss.n4807 68.5181
R33709 vss.n4805 vss.n4802 68.5181
R33710 vss.n4802 vss.n4794 68.5181
R33711 vss.n5494 vss.n4787 68.5181
R33712 vss.n5494 vss.n5493 68.5181
R33713 vss.n5479 vss.n4815 68.5181
R33714 vss.n5479 vss.n5478 68.5181
R33715 vss.n5465 vss.n5462 68.5181
R33716 vss.n5462 vss.n4816 68.5181
R33717 vss.n5461 vss.n4825 68.5181
R33718 vss.n5456 vss.n4825 68.5181
R33719 vss.n5443 vss.n4850 68.5181
R33720 vss.n4853 vss.n4850 68.5181
R33721 vss.n4848 vss.n4845 68.5181
R33722 vss.n4845 vss.n4837 68.5181
R33723 vss.n5451 vss.n4830 68.5181
R33724 vss.n5451 vss.n5450 68.5181
R33725 vss.n5436 vss.n4858 68.5181
R33726 vss.n5436 vss.n5435 68.5181
R33727 vss.n5422 vss.n5419 68.5181
R33728 vss.n5419 vss.n4859 68.5181
R33729 vss.n5418 vss.n4868 68.5181
R33730 vss.n5413 vss.n4868 68.5181
R33731 vss.n5400 vss.n5344 68.5181
R33732 vss.n5347 vss.n5344 68.5181
R33733 vss.n5342 vss.n5339 68.5181
R33734 vss.n5339 vss.n5331 68.5181
R33735 vss.n5408 vss.n4873 68.5181
R33736 vss.n5408 vss.n5407 68.5181
R33737 vss.n5374 vss.n5360 68.5181
R33738 vss.n5379 vss.n5360 68.5181
R33739 vss.n2880 vss.n2879 68.5181
R33740 vss.n2879 vss.n2874 68.5181
R33741 vss.n9831 vss.n2872 68.5181
R33742 vss.n9843 vss.n2872 68.5181
R33743 vss.n9823 vss.n2882 68.5181
R33744 vss.n9824 vss.n9823 68.5181
R33745 vss.n2957 vss.n2956 68.5181
R33746 vss.n2956 vss.n2952 68.5181
R33747 vss.n2951 vss.n2942 68.5181
R33748 vss.n2971 vss.n2951 68.5181
R33749 vss.n2976 vss.n2941 68.5181
R33750 vss.n2949 vss.n2941 68.5181
R33751 vss.n2910 vss.n2909 68.5181
R33752 vss.n2909 vss.n2905 68.5181
R33753 vss.n2904 vss.n2895 68.5181
R33754 vss.n2925 vss.n2904 68.5181
R33755 vss.n2930 vss.n2894 68.5181
R33756 vss.n2902 vss.n2894 68.5181
R33757 vss.n4931 vss.n4930 68.5181
R33758 vss.n4930 vss.n4925 68.5181
R33759 vss.n4951 vss.n4923 68.5181
R33760 vss.n4963 vss.n4923 68.5181
R33761 vss.n4943 vss.n4933 68.5181
R33762 vss.n4944 vss.n4943 68.5181
R33763 vss.n5133 vss.n5132 68.5181
R33764 vss.n5132 vss.n5127 68.5181
R33765 vss.n5153 vss.n5125 68.5181
R33766 vss.n5165 vss.n5125 68.5181
R33767 vss.n5145 vss.n5135 68.5181
R33768 vss.n5146 vss.n5145 68.5181
R33769 vss.n3113 vss.n3112 68.5181
R33770 vss.n3112 vss.n3107 68.5181
R33771 vss.n3134 vss.n3105 68.5181
R33772 vss.n3146 vss.n3105 68.5181
R33773 vss.n3126 vss.n3115 68.5181
R33774 vss.n3127 vss.n3126 68.5181
R33775 vss.n4468 vss.n4463 68.5181
R33776 vss.n4491 vss.n4468 68.5181
R33777 vss.n4502 vss.n4461 68.5181
R33778 vss.n4489 vss.n4461 68.5181
R33779 vss.n4478 vss.n4477 68.5181
R33780 vss.n4477 vss.n4470 68.5181
R33781 vss.n4376 vss.n4371 68.5181
R33782 vss.n4399 vss.n4376 68.5181
R33783 vss.n4410 vss.n4369 68.5181
R33784 vss.n4397 vss.n4369 68.5181
R33785 vss.n4386 vss.n4385 68.5181
R33786 vss.n4385 vss.n4378 68.5181
R33787 vss.n4328 vss.n4323 68.5181
R33788 vss.n4351 vss.n4328 68.5181
R33789 vss.n4362 vss.n4321 68.5181
R33790 vss.n4349 vss.n4321 68.5181
R33791 vss.n4338 vss.n4337 68.5181
R33792 vss.n4337 vss.n4330 68.5181
R33793 vss.n3728 vss.n3723 68.5181
R33794 vss.n3751 vss.n3728 68.5181
R33795 vss.n3762 vss.n3721 68.5181
R33796 vss.n3749 vss.n3721 68.5181
R33797 vss.n3738 vss.n3737 68.5181
R33798 vss.n3737 vss.n3730 68.5181
R33799 vss.n4030 vss.n4025 68.5181
R33800 vss.n4053 vss.n4030 68.5181
R33801 vss.n4064 vss.n4023 68.5181
R33802 vss.n4051 vss.n4023 68.5181
R33803 vss.n4040 vss.n4039 68.5181
R33804 vss.n4039 vss.n4032 68.5181
R33805 vss.n3683 vss.n3678 68.5181
R33806 vss.n3706 vss.n3683 68.5181
R33807 vss.n3717 vss.n3676 68.5181
R33808 vss.n3704 vss.n3676 68.5181
R33809 vss.n3693 vss.n3692 68.5181
R33810 vss.n3692 vss.n3685 68.5181
R33811 vss.n4084 vss.n4079 68.5181
R33812 vss.n4107 vss.n4084 68.5181
R33813 vss.n4118 vss.n4077 68.5181
R33814 vss.n4105 vss.n4077 68.5181
R33815 vss.n4094 vss.n4093 68.5181
R33816 vss.n4093 vss.n4086 68.5181
R33817 vss.n3508 vss.n3503 68.5181
R33818 vss.n3531 vss.n3508 68.5181
R33819 vss.n3542 vss.n3501 68.5181
R33820 vss.n3529 vss.n3501 68.5181
R33821 vss.n3518 vss.n3517 68.5181
R33822 vss.n3517 vss.n3510 68.5181
R33823 vss.n3463 vss.n3458 68.5181
R33824 vss.n3486 vss.n3463 68.5181
R33825 vss.n3497 vss.n3456 68.5181
R33826 vss.n3484 vss.n3456 68.5181
R33827 vss.n3473 vss.n3472 68.5181
R33828 vss.n3472 vss.n3465 68.5181
R33829 vss.n5751 vss.n5746 68.5181
R33830 vss.n5774 vss.n5751 68.5181
R33831 vss.n5785 vss.n5744 68.5181
R33832 vss.n5772 vss.n5744 68.5181
R33833 vss.n5761 vss.n5760 68.5181
R33834 vss.n5760 vss.n5753 68.5181
R33835 vss.n5724 vss.n5695 68.5181
R33836 vss.n5729 vss.n5695 68.5181
R33837 vss.n5723 vss.n5705 68.5181
R33838 vss.n5705 vss.n5696 68.5181
R33839 vss.n5738 vss.n3603 68.5181
R33840 vss.n5685 vss.n3603 68.5181
R33841 vss.n5792 vss.n3587 68.5181
R33842 vss.n5797 vss.n3587 68.5181
R33843 vss.n5791 vss.n3597 68.5181
R33844 vss.n3597 vss.n3588 68.5181
R33845 vss.n5806 vss.n3577 68.5181
R33846 vss.n3577 vss.n3567 68.5181
R33847 vss.n3551 vss.n3546 68.5181
R33848 vss.n5827 vss.n3551 68.5181
R33849 vss.n5838 vss.n3544 68.5181
R33850 vss.n5825 vss.n3544 68.5181
R33851 vss.n3926 vss.n3906 68.5181
R33852 vss.n3906 vss.n3896 68.5181
R33853 vss.n4125 vss.n3873 68.5181
R33854 vss.n4130 vss.n3873 68.5181
R33855 vss.n4124 vss.n3883 68.5181
R33856 vss.n3883 vss.n3874 68.5181
R33857 vss.n4139 vss.n3854 68.5181
R33858 vss.n3854 vss.n3844 68.5181
R33859 vss.n3810 vss.n3805 68.5181
R33860 vss.n4160 vss.n3810 68.5181
R33861 vss.n4171 vss.n3803 68.5181
R33862 vss.n4158 vss.n3803 68.5181
R33863 vss.n4174 vss.n3798 68.5181
R33864 vss.n3798 vss.n3788 68.5181
R33865 vss.n3770 vss.n3765 68.5181
R33866 vss.n4195 vss.n3770 68.5181
R33867 vss.n4206 vss.n3763 68.5181
R33868 vss.n4193 vss.n3763 68.5181
R33869 vss.n4617 vss.n3644 68.5181
R33870 vss.n3644 vss.n3635 68.5181
R33871 vss.n4420 vss.n4415 68.5181
R33872 vss.n4598 vss.n4420 68.5181
R33873 vss.n4609 vss.n4413 68.5181
R33874 vss.n4596 vss.n4413 68.5181
R33875 vss.n4546 vss.n4434 68.5181
R33876 vss.n4434 vss.n4427 68.5181
R33877 vss.n4528 vss.n4509 68.5181
R33878 vss.n4523 vss.n4509 68.5181
R33879 vss.n4514 vss.n4508 68.5181
R33880 vss.n4521 vss.n4514 68.5181
R33881 vss.n4516 vss.n4515 68.5181
R33882 vss.n4519 vss.n4516 68.5181
R33883 vss.n4440 vss.n4435 68.5181
R33884 vss.n4541 vss.n4440 68.5181
R33885 vss.n4547 vss.n4426 68.5181
R33886 vss.n4552 vss.n4426 68.5181
R33887 vss.n4568 vss.n4567 68.5181
R33888 vss.n4567 vss.n4560 68.5181
R33889 vss.n4574 vss.n4573 68.5181
R33890 vss.n4582 vss.n4574 68.5181
R33891 vss.n4618 vss.n3634 68.5181
R33892 vss.n4623 vss.n3634 68.5181
R33893 vss.n3782 vss.n3781 68.5181
R33894 vss.n3781 vss.n3774 68.5181
R33895 vss.n3796 vss.n3787 68.5181
R33896 vss.n4179 vss.n3787 68.5181
R33897 vss.n3816 vss.n3815 68.5181
R33898 vss.n3822 vss.n3816 68.5181
R33899 vss.n3838 vss.n3837 68.5181
R33900 vss.n3837 vss.n3830 68.5181
R33901 vss.n3852 vss.n3843 68.5181
R33902 vss.n4144 vss.n3843 68.5181
R33903 vss.n3863 vss.n3856 68.5181
R33904 vss.n3865 vss.n3863 68.5181
R33905 vss.n3889 vss.n3884 68.5181
R33906 vss.n3941 vss.n3889 68.5181
R33907 vss.n3904 vss.n3895 68.5181
R33908 vss.n3931 vss.n3895 68.5181
R33909 vss.n3914 vss.n3907 68.5181
R33910 vss.n3916 vss.n3914 68.5181
R33911 vss.n3561 vss.n3560 68.5181
R33912 vss.n3560 vss.n3553 68.5181
R33913 vss.n3575 vss.n3566 68.5181
R33914 vss.n5811 vss.n3566 68.5181
R33915 vss.n3617 vss.n3580 68.5181
R33916 vss.n3619 vss.n3617 68.5181
R33917 vss.n5666 vss.n5665 68.5181
R33918 vss.n5669 vss.n5666 68.5181
R33919 vss.n5657 vss.n5656 68.5181
R33920 vss.n5656 vss.n5649 68.5181
R33921 vss.n5648 vss.n3605 68.5181
R33922 vss.n5687 vss.n5648 68.5181
R33923 vss.n5711 vss.n5706 68.5181
R33924 vss.n5718 vss.n5711 68.5181
R33925 vss.n2638 vss.n2633 68.5181
R33926 vss.n9978 vss.n2638 68.5181
R33927 vss.n9989 vss.n2631 68.5181
R33928 vss.n9976 vss.n2631 68.5181
R33929 vss.n9965 vss.n9964 68.5181
R33930 vss.n9964 vss.n9957 68.5181
R33931 vss.n2675 vss.n2643 68.5181
R33932 vss.n2680 vss.n2643 68.5181
R33933 vss.n2674 vss.n2653 68.5181
R33934 vss.n2653 vss.n2644 68.5181
R33935 vss.n2659 vss.n2654 68.5181
R33936 vss.n2667 vss.n2659 68.5181
R33937 vss.n3388 vss.n3383 68.5181
R33938 vss.n3411 vss.n3388 68.5181
R33939 vss.n3422 vss.n3381 68.5181
R33940 vss.n3409 vss.n3381 68.5181
R33941 vss.n3398 vss.n3397 68.5181
R33942 vss.n3397 vss.n3390 68.5181
R33943 vss.n3985 vss.n3980 68.5181
R33944 vss.n4008 vss.n3985 68.5181
R33945 vss.n4019 vss.n3978 68.5181
R33946 vss.n4006 vss.n3978 68.5181
R33947 vss.n3995 vss.n3994 68.5181
R33948 vss.n3994 vss.n3987 68.5181
R33949 vss.n4252 vss.n4247 68.5181
R33950 vss.n4275 vss.n4252 68.5181
R33951 vss.n4286 vss.n4245 68.5181
R33952 vss.n4273 vss.n4245 68.5181
R33953 vss.n4262 vss.n4261 68.5181
R33954 vss.n4261 vss.n4254 68.5181
R33955 vss.n5905 vss.n5904 68.5181
R33956 vss.n5904 vss.n5899 68.5181
R33957 vss.n5930 vss.n5889 68.5181
R33958 vss.n5916 vss.n5889 68.5181
R33959 vss.n5918 vss.n5891 68.5181
R33960 vss.n5925 vss.n5918 68.5181
R33961 vss.n14067 vss.n487 68.5181
R33962 vss.n14068 vss.n14067 68.5181
R33963 vss.n10110 vss.n10109 68.5181
R33964 vss.n10109 vss.n10104 68.5181
R33965 vss.n10130 vss.n10102 68.5181
R33966 vss.n10142 vss.n10102 68.5181
R33967 vss.n10122 vss.n10112 68.5181
R33968 vss.n10123 vss.n10122 68.5181
R33969 vss.n12868 vss.n12867 68.5181
R33970 vss.n12867 vss.n12862 68.5181
R33971 vss.n12888 vss.n12860 68.5181
R33972 vss.n12900 vss.n12860 68.5181
R33973 vss.n12880 vss.n12870 68.5181
R33974 vss.n12881 vss.n12880 68.5181
R33975 vss.n10151 vss.n10150 68.5181
R33976 vss.n10150 vss.n10145 68.5181
R33977 vss.n10171 vss.n10143 68.5181
R33978 vss.n10183 vss.n10143 68.5181
R33979 vss.n10163 vss.n10153 68.5181
R33980 vss.n10164 vss.n10163 68.5181
R33981 vss.n12417 vss.n12416 68.5181
R33982 vss.n12416 vss.n12411 68.5181
R33983 vss.n12437 vss.n12409 68.5181
R33984 vss.n12449 vss.n12409 68.5181
R33985 vss.n12429 vss.n12419 68.5181
R33986 vss.n12430 vss.n12429 68.5181
R33987 vss.n11746 vss.n11745 68.5181
R33988 vss.n11745 vss.n11740 68.5181
R33989 vss.n11766 vss.n11738 68.5181
R33990 vss.n11778 vss.n11738 68.5181
R33991 vss.n11758 vss.n11748 68.5181
R33992 vss.n11759 vss.n11758 68.5181
R33993 vss.n12462 vss.n12461 68.5181
R33994 vss.n12461 vss.n12456 68.5181
R33995 vss.n12482 vss.n12454 68.5181
R33996 vss.n12494 vss.n12454 68.5181
R33997 vss.n12474 vss.n12464 68.5181
R33998 vss.n12475 vss.n12474 68.5181
R33999 vss.n2327 vss.n2326 68.5181
R34000 vss.n2326 vss.n2322 68.5181
R34001 vss.n2321 vss.n2312 68.5181
R34002 vss.n2341 vss.n2321 68.5181
R34003 vss.n2346 vss.n2311 68.5181
R34004 vss.n2319 vss.n2311 68.5181
R34005 vss.n12287 vss.n12286 68.5181
R34006 vss.n12286 vss.n12281 68.5181
R34007 vss.n12307 vss.n12279 68.5181
R34008 vss.n12319 vss.n12279 68.5181
R34009 vss.n12299 vss.n12289 68.5181
R34010 vss.n12300 vss.n12299 68.5181
R34011 vss.n12332 vss.n12331 68.5181
R34012 vss.n12331 vss.n12326 68.5181
R34013 vss.n12352 vss.n12324 68.5181
R34014 vss.n12364 vss.n12324 68.5181
R34015 vss.n12344 vss.n12334 68.5181
R34016 vss.n12345 vss.n12344 68.5181
R34017 vss.n10228 vss.n10227 68.5181
R34018 vss.n10227 vss.n10222 68.5181
R34019 vss.n10248 vss.n10220 68.5181
R34020 vss.n10260 vss.n10220 68.5181
R34021 vss.n10240 vss.n10230 68.5181
R34022 vss.n10241 vss.n10240 68.5181
R34023 vss.n2408 vss.n2407 68.5181
R34024 vss.n2407 vss.n2402 68.5181
R34025 vss.n2428 vss.n2400 68.5181
R34026 vss.n2440 vss.n2400 68.5181
R34027 vss.n2420 vss.n2410 68.5181
R34028 vss.n2421 vss.n2420 68.5181
R34029 vss.n2387 vss.n2386 68.5181
R34030 vss.n2386 vss.n2382 68.5181
R34031 vss.n2381 vss.n2372 68.5181
R34032 vss.n12966 vss.n2381 68.5181
R34033 vss.n12971 vss.n2371 68.5181
R34034 vss.n2379 vss.n2371 68.5181
R34035 vss.n13081 vss.n2113 68.5181
R34036 vss.n2116 vss.n2113 68.5181
R34037 vss.n2111 vss.n2108 68.5181
R34038 vss.n2108 vss.n2100 68.5181
R34039 vss.n13089 vss.n2098 68.5181
R34040 vss.n13089 vss.n13088 68.5181
R34041 vss.n12946 vss.n10053 68.5181
R34042 vss.n10053 vss.n10019 68.5181
R34043 vss.n10051 vss.n10017 68.5181
R34044 vss.n12951 vss.n10017 68.5181
R34045 vss.n10032 vss.n10027 68.5181
R34046 vss.n10033 vss.n10032 68.5181
R34047 vss.n10063 vss.n10062 68.5181
R34048 vss.n12937 vss.n10063 68.5181
R34049 vss.n12932 vss.n10074 68.5181
R34050 vss.n10074 vss.n10067 68.5181
R34051 vss.n10080 vss.n10075 68.5181
R34052 vss.n12927 vss.n10080 68.5181
R34053 vss.n2487 vss.n2486 68.5181
R34054 vss.n2486 vss.n2481 68.5181
R34055 vss.n2508 vss.n2479 68.5181
R34056 vss.n2520 vss.n2479 68.5181
R34057 vss.n2500 vss.n2489 68.5181
R34058 vss.n2501 vss.n2500 68.5181
R34059 vss.n13062 vss.n2135 68.5181
R34060 vss.n13062 vss.n13061 68.5181
R34061 vss.n13067 vss.n2134 68.5181
R34062 vss.n2134 vss.n2124 68.5181
R34063 vss.n2132 vss.n2123 68.5181
R34064 vss.n13072 vss.n2123 68.5181
R34065 vss.n11832 vss.n11831 68.5181
R34066 vss.n12117 vss.n11832 68.5181
R34067 vss.n12110 vss.n11841 68.5181
R34068 vss.n11841 vss.n11836 68.5181
R34069 vss.n11847 vss.n11842 68.5181
R34070 vss.n12105 vss.n11847 68.5181
R34071 vss.n11822 vss.n11813 68.5181
R34072 vss.n12144 vss.n11822 68.5181
R34073 vss.n12149 vss.n11812 68.5181
R34074 vss.n11820 vss.n11812 68.5181
R34075 vss.n11803 vss.n11798 68.5181
R34076 vss.n12158 vss.n11803 68.5181
R34077 vss.n12263 vss.n11780 68.5181
R34078 vss.n12275 vss.n11780 68.5181
R34079 vss.n12257 vss.n12181 68.5181
R34080 vss.n12257 vss.n12256 68.5181
R34081 vss.n12247 vss.n12194 68.5181
R34082 vss.n12202 vss.n12194 68.5181
R34083 vss.n11734 vss.n11725 68.5181
R34084 vss.n12540 vss.n11734 68.5181
R34085 vss.n12545 vss.n11724 68.5181
R34086 vss.n11732 vss.n11724 68.5181
R34087 vss.n11716 vss.n11711 68.5181
R34088 vss.n12554 vss.n11716 68.5181
R34089 vss.n11639 vss.n11638 68.5181
R34090 vss.n11638 vss.n11628 68.5181
R34091 vss.n11690 vss.n11627 68.5181
R34092 vss.n12582 vss.n11627 68.5181
R34093 vss.n11682 vss.n11645 68.5181
R34094 vss.n11653 vss.n11645 68.5181
R34095 vss.n12843 vss.n10303 68.5181
R34096 vss.n12855 vss.n10303 68.5181
R34097 vss.n12837 vss.n10313 68.5181
R34098 vss.n12837 vss.n12836 68.5181
R34099 vss.n12827 vss.n12776 68.5181
R34100 vss.n12784 vss.n12776 68.5181
R34101 vss.n10099 vss.n10090 68.5181
R34102 vss.n12913 vss.n10099 68.5181
R34103 vss.n12918 vss.n10089 68.5181
R34104 vss.n10097 vss.n10089 68.5181
R34105 vss.n11877 vss.n11872 68.5181
R34106 vss.n11884 vss.n11877 68.5181
R34107 vss.n10468 vss.n10463 68.5181
R34108 vss.n10490 vss.n10468 68.5181
R34109 vss.n10501 vss.n10461 68.5181
R34110 vss.n10488 vss.n10461 68.5181
R34111 vss.n10478 vss.n10477 68.5181
R34112 vss.n10477 vss.n10470 68.5181
R34113 vss.n10689 vss.n10684 68.5181
R34114 vss.n10711 vss.n10689 68.5181
R34115 vss.n10722 vss.n10682 68.5181
R34116 vss.n10709 vss.n10682 68.5181
R34117 vss.n10699 vss.n10698 68.5181
R34118 vss.n10698 vss.n10691 68.5181
R34119 vss.n11003 vss.n10998 68.5181
R34120 vss.n11025 vss.n11003 68.5181
R34121 vss.n11036 vss.n10996 68.5181
R34122 vss.n11023 vss.n10996 68.5181
R34123 vss.n11013 vss.n11012 68.5181
R34124 vss.n11012 vss.n11005 68.5181
R34125 vss.n11121 vss.n11120 68.5181
R34126 vss.n11120 vss.n11115 68.5181
R34127 vss.n11145 vss.n11105 68.5181
R34128 vss.n11131 vss.n11105 68.5181
R34129 vss.n11133 vss.n11107 68.5181
R34130 vss.n11140 vss.n11133 68.5181
R34131 vss.n13056 vss.n13055 68.2878
R34132 vss.n9875 vss.n9874 68.2878
R34133 vss.n14783 vss.n14782 68.2873
R34134 vss.n5971 vss.n5970 68.2362
R34135 vss.n8153 vss.n8152 63.5774
R34136 vss.n3282 vss.n3281 63.5774
R34137 vss.n9897 vss.n2742 63.5774
R34138 vss.n14155 vss.n14154 63.5774
R34139 vss.n14176 vss.n14175 63.5774
R34140 vss.n10042 vss.n10041 63.5774
R34141 vss.n13054 vss.t76 59.9409
R34142 vss.n12671 vss.n2072 58.4831
R34143 vss.n14060 vss.n496 53.5296
R34144 vss.n14060 vss.n497 53.5296
R34145 vss.n715 vss.t1412 52.1058
R34146 vss.n9140 vss.t351 52.1058
R34147 vss.n5734 vss.t688 52.1058
R34148 vss.n12087 vss.t530 52.1058
R34149 vss.n14114 vss.n433 51.6849
R34150 vss.n14783 vss.n26 51.6849
R34151 vss.n8986 vss.n7323 51.6849
R34152 vss.n9896 vss.n9895 51.6849
R34153 vss.n9876 vss.n9875 51.6849
R34154 vss.n13057 vss.n13056 51.6849
R34155 vss.n13922 vss.n13301 51.1409
R34156 vss.n9050 vss.n9049 51.1409
R34157 vss.n5644 vss.n5643 51.1409
R34158 vss.n12098 vss.n12097 51.1409
R34159 vss.n2046 vss.n2045 51.0489
R34160 vss.n10407 vss.n10395 51.0489
R34161 vss.n12651 vss.n12650 51.0489
R34162 vss.n12639 vss.n12638 51.0489
R34163 vss.n12687 vss.n12686 51.0489
R34164 vss.n12674 vss.n10392 51.0489
R34165 vss.n11437 vss.n11436 51.0489
R34166 vss.n11424 vss.n11423 51.0489
R34167 vss.n11390 vss.n11389 51.0489
R34168 vss.n11377 vss.n11376 51.0489
R34169 vss.n10965 vss.n10964 51.0489
R34170 vss.n10952 vss.n10951 51.0489
R34171 vss.n10802 vss.n10801 51.0489
R34172 vss.n10789 vss.n10788 51.0489
R34173 vss.n10758 vss.n10757 51.0489
R34174 vss.n10745 vss.n10744 51.0489
R34175 vss.n11584 vss.n11583 51.0489
R34176 vss.n11571 vss.n11570 51.0489
R34177 vss.n10581 vss.n10580 51.0489
R34178 vss.n10568 vss.n10567 51.0489
R34179 vss.n10537 vss.n10536 51.0489
R34180 vss.n10524 vss.n10523 51.0489
R34181 vss.n11958 vss.n11957 51.0489
R34182 vss.n11945 vss.n11944 51.0489
R34183 vss.n12095 vss.n11853 51.0489
R34184 vss.n12062 vss.n11902 51.0489
R34185 vss.n11979 vss.n11918 51.0489
R34186 vss.n11908 vss.n11907 51.0489
R34187 vss.n12033 vss.n12032 51.0489
R34188 vss.n12022 vss.n11989 51.0489
R34189 vss.n10605 vss.n10604 51.0489
R34190 vss.n11996 vss.n11995 51.0489
R34191 vss.n10612 vss.n10611 51.0489
R34192 vss.n10668 vss.n10645 51.0489
R34193 vss.n11610 vss.n10625 51.0489
R34194 vss.n10641 vss.n10639 51.0489
R34195 vss.n11621 vss.n10618 51.0489
R34196 vss.n10855 vss.n10832 51.0489
R34197 vss.n10871 vss.n10870 51.0489
R34198 vss.n10859 vss.n10829 51.0489
R34199 vss.n11518 vss.n11517 51.0489
R34200 vss.n11507 vss.n10881 51.0489
R34201 vss.n10978 vss.n10897 51.0489
R34202 vss.n10887 vss.n10886 51.0489
R34203 vss.n11470 vss.n11469 51.0489
R34204 vss.n11459 vss.n10907 51.0489
R34205 vss.n12753 vss.n10332 51.0489
R34206 vss.n10916 vss.n10915 51.0489
R34207 vss.n12764 vss.n10325 51.0489
R34208 vss.n12727 vss.n10351 51.0489
R34209 vss.n12708 vss.n10367 51.0489
R34210 vss.n10357 vss.n10356 51.0489
R34211 vss.n12995 vss.n2258 51.0489
R34212 vss.n13008 vss.n13006 51.0489
R34213 vss.n2301 vss.n2300 51.0489
R34214 vss.n2287 vss.n2282 51.0489
R34215 vss.n13110 vss.n13109 51.0489
R34216 vss.n13096 vss.n2093 51.0489
R34217 vss.n1125 vss.n1124 51.0489
R34218 vss.n1113 vss.n1112 51.0489
R34219 vss.n859 vss.n845 51.0489
R34220 vss.n872 vss.n836 51.0489
R34221 vss.n14159 vss.n455 51.0489
R34222 vss.n14173 vss.n14172 51.0489
R34223 vss.n187 vss.n186 51.0489
R34224 vss.n16 vss.n14 51.0489
R34225 vss.n336 vss.n334 51.0489
R34226 vss.n349 vss.n347 51.0489
R34227 vss.n14218 vss.n14217 51.0489
R34228 vss.n14204 vss.n14199 51.0489
R34229 vss.n14115 vss.n14113 51.0489
R34230 vss.n14128 vss.n14126 51.0489
R34231 vss.n14224 vss.n431 51.0489
R34232 vss.n14237 vss.n14235 51.0489
R34233 vss.n470 vss.n462 51.0489
R34234 vss.n13580 vss.n13579 51.0489
R34235 vss.n13606 vss.n13605 51.0489
R34236 vss.n13592 vss.n13586 51.0489
R34237 vss.n14681 vss.n14680 51.0489
R34238 vss.n14667 vss.n14662 51.0489
R34239 vss.n14538 vss.n249 51.0489
R34240 vss.n14551 vss.n14549 51.0489
R34241 vss.n14486 vss.n14485 51.0489
R34242 vss.n14472 vss.n14467 51.0489
R34243 vss.n14343 vss.n308 51.0489
R34244 vss.n14356 vss.n14354 51.0489
R34245 vss.n14291 vss.n14290 51.0489
R34246 vss.n14277 vss.n14272 51.0489
R34247 vss.n14337 vss.n14336 51.0489
R34248 vss.n14323 vss.n14318 51.0489
R34249 vss.n14389 vss.n14387 51.0489
R34250 vss.n14402 vss.n14400 51.0489
R34251 vss.n14532 vss.n14531 51.0489
R34252 vss.n14518 vss.n14513 51.0489
R34253 vss.n14584 vss.n14582 51.0489
R34254 vss.n14597 vss.n14595 51.0489
R34255 vss.n14727 vss.n14726 51.0489
R34256 vss.n14713 vss.n14708 51.0489
R34257 vss.n14733 vss.n172 51.0489
R34258 vss.n14746 vss.n14744 51.0489
R34259 vss.n13314 vss.n13306 51.0489
R34260 vss.n13905 vss.n13323 51.0489
R34261 vss.n13877 vss.n13342 51.0489
R34262 vss.n13895 vss.n13894 51.0489
R34263 vss.n13356 vss.n13348 51.0489
R34264 vss.n13850 vss.n13362 51.0489
R34265 vss.n13823 vss.n13383 51.0489
R34266 vss.n13841 vss.n13840 51.0489
R34267 vss.n13397 vss.n13389 51.0489
R34268 vss.n13800 vss.n13403 51.0489
R34269 vss.n13772 vss.n13422 51.0489
R34270 vss.n13790 vss.n13789 51.0489
R34271 vss.n13436 vss.n13428 51.0489
R34272 vss.n13745 vss.n13442 51.0489
R34273 vss.n13718 vss.n13463 51.0489
R34274 vss.n13736 vss.n13735 51.0489
R34275 vss.n13477 vss.n13469 51.0489
R34276 vss.n13695 vss.n13483 51.0489
R34277 vss.n13667 vss.n13502 51.0489
R34278 vss.n13685 vss.n13684 51.0489
R34279 vss.n13516 vss.n13508 51.0489
R34280 vss.n13640 vss.n13522 51.0489
R34281 vss.n13613 vss.n13543 51.0489
R34282 vss.n13631 vss.n13630 51.0489
R34283 vss.n656 vss.n616 51.0489
R34284 vss.n632 vss.n630 51.0489
R34285 vss.n13224 vss.n13223 51.0489
R34286 vss.n13212 vss.n811 51.0489
R34287 vss.n1683 vss.n1682 51.0489
R34288 vss.n1671 vss.n1670 51.0489
R34289 vss.n1636 vss.n1635 51.0489
R34290 vss.n1624 vss.n1623 51.0489
R34291 vss.n1388 vss.n1387 51.0489
R34292 vss.n1376 vss.n1375 51.0489
R34293 vss.n1189 vss.n1188 51.0489
R34294 vss.n1177 vss.n1176 51.0489
R34295 vss.n1341 vss.n1340 51.0489
R34296 vss.n1329 vss.n1328 51.0489
R34297 vss.n1080 vss.n1079 51.0489
R34298 vss.n1068 vss.n1067 51.0489
R34299 vss.n1473 vss.n1472 51.0489
R34300 vss.n1461 vss.n1460 51.0489
R34301 vss.n1553 vss.n1552 51.0489
R34302 vss.n1541 vss.n1540 51.0489
R34303 vss.n609 vss.n608 51.0489
R34304 vss.n831 vss.n819 51.0489
R34305 vss.n903 vss.n885 51.0489
R34306 vss.n916 vss.n877 51.0489
R34307 vss.n14016 vss.n14015 51.0489
R34308 vss.n14003 vss.n535 51.0489
R34309 vss.n676 vss.n662 51.0489
R34310 vss.n13999 vss.n539 51.0489
R34311 vss.n13981 vss.n13980 51.0489
R34312 vss.n13968 vss.n574 51.0489
R34313 vss.n775 vss.n765 51.0489
R34314 vss.n13964 vss.n578 51.0489
R34315 vss.n785 vss.n784 51.0489
R34316 vss.n13247 vss.n745 51.0489
R34317 vss.n1746 vss.n1709 51.0489
R34318 vss.n1729 vss.n1725 51.0489
R34319 vss.n1793 vss.n1792 51.0489
R34320 vss.n1780 vss.n1761 51.0489
R34321 vss.n1817 vss.n1266 51.0489
R34322 vss.n1776 vss.n1764 51.0489
R34323 vss.n1823 vss.n1247 51.0489
R34324 vss.n1254 vss.n1234 51.0489
R34325 vss.n1850 vss.n1213 51.0489
R34326 vss.n1833 vss.n1229 51.0489
R34327 vss.n1897 vss.n1896 51.0489
R34328 vss.n1884 vss.n1865 51.0489
R34329 vss.n1921 vss.n1148 51.0489
R34330 vss.n1880 vss.n1868 51.0489
R34331 vss.n1968 vss.n1967 51.0489
R34332 vss.n1955 vss.n1936 51.0489
R34333 vss.n13299 vss.n692 51.0489
R34334 vss.n1951 vss.n1939 51.0489
R34335 vss.n13280 vss.n13279 51.0489
R34336 vss.n13267 vss.n727 51.0489
R34337 vss.n2015 vss.n2014 51.0489
R34338 vss.n2003 vss.n2002 51.0489
R34339 vss.n13177 vss.n13176 51.0489
R34340 vss.n13188 vss.n13187 51.0489
R34341 vss.n9605 vss.n9603 51.0489
R34342 vss.n9618 vss.n9616 51.0489
R34343 vss.n9181 vss.n9180 51.0489
R34344 vss.n9169 vss.n9167 51.0489
R34345 vss.n9484 vss.n9447 51.0489
R34346 vss.n9464 vss.n9460 51.0489
R34347 vss.n8042 vss.n8015 51.0489
R34348 vss.n8037 vss.n8026 51.0489
R34349 vss.n9666 vss.n9665 51.0489
R34350 vss.n9652 vss.n5994 51.0489
R34351 vss.n8150 vss.n8149 51.0489
R34352 vss.n8139 vss.n8138 51.0489
R34353 vss.n8157 vss.n8120 51.0489
R34354 vss.n8171 vss.n8170 51.0489
R34355 vss.n8083 vss.n8076 51.0489
R34356 vss.n8097 vss.n8096 51.0489
R34357 vss.n8222 vss.n8009 51.0489
R34358 vss.n8235 vss.n8233 51.0489
R34359 vss.n8216 vss.n8215 51.0489
R34360 vss.n8202 vss.n8197 51.0489
R34361 vss.n9004 vss.n9003 51.0489
R34362 vss.n8990 vss.n7320 51.0489
R34363 vss.n8713 vss.n7866 51.0489
R34364 vss.n8726 vss.n8724 51.0489
R34365 vss.n7787 vss.n7785 51.0489
R34366 vss.n7800 vss.n7798 51.0489
R34367 vss.n8780 vss.n8779 51.0489
R34368 vss.n8766 vss.n8761 51.0489
R34369 vss.n8832 vss.n7679 51.0489
R34370 vss.n8845 vss.n8843 51.0489
R34371 vss.n8826 vss.n8825 51.0489
R34372 vss.n8812 vss.n8807 51.0489
R34373 vss.n8899 vss.n8898 51.0489
R34374 vss.n8885 vss.n8880 51.0489
R34375 vss.n9035 vss.n9034 51.0489
R34376 vss.n9021 vss.n7288 51.0489
R34377 vss.n8280 vss.n8279 51.0489
R34378 vss.n9012 vss.n7295 51.0489
R34379 vss.n8287 vss.n7898 51.0489
R34380 vss.n8301 vss.n8300 51.0489
R34381 vss.n8693 vss.n8317 51.0489
R34382 vss.n8707 vss.n8706 51.0489
R34383 vss.n8327 vss.n8322 51.0489
R34384 vss.n8347 vss.n8344 51.0489
R34385 vss.n8648 vss.n8362 51.0489
R34386 vss.n8668 vss.n8663 51.0489
R34387 vss.n8372 vss.n8367 51.0489
R34388 vss.n8397 vss.n8394 51.0489
R34389 vss.n8604 vss.n8415 51.0489
R34390 vss.n8625 vss.n8619 51.0489
R34391 vss.n8425 vss.n8420 51.0489
R34392 vss.n8445 vss.n8442 51.0489
R34393 vss.n8561 vss.n8460 51.0489
R34394 vss.n8581 vss.n8576 51.0489
R34395 vss.n8470 vss.n8465 51.0489
R34396 vss.n8495 vss.n8492 51.0489
R34397 vss.n8525 vss.n8508 51.0489
R34398 vss.n8538 vss.n8532 51.0489
R34399 vss.n8951 vss.n7490 51.0489
R34400 vss.n8964 vss.n8962 51.0489
R34401 vss.n8945 vss.n8944 51.0489
R34402 vss.n8931 vss.n8926 51.0489
R34403 vss.n7533 vss.n7532 51.0489
R34404 vss.n7519 vss.n7514 51.0489
R34405 vss.n7564 vss.n7562 51.0489
R34406 vss.n7577 vss.n7575 51.0489
R34407 vss.n7707 vss.n7705 51.0489
R34408 vss.n7720 vss.n7718 51.0489
R34409 vss.n7928 vss.n7926 51.0489
R34410 vss.n7941 vss.n7939 51.0489
R34411 vss.n6039 vss.n6038 51.0489
R34412 vss.n6027 vss.n6025 51.0489
R34413 vss.n7209 vss.n7208 51.0489
R34414 vss.n7197 vss.n7195 51.0489
R34415 vss.n6704 vss.n6703 51.0489
R34416 vss.n6692 vss.n6690 51.0489
R34417 vss.n6660 vss.n6659 51.0489
R34418 vss.n6648 vss.n6646 51.0489
R34419 vss.n7018 vss.n7017 51.0489
R34420 vss.n7006 vss.n7004 51.0489
R34421 vss.n6478 vss.n6477 51.0489
R34422 vss.n6466 vss.n6464 51.0489
R34423 vss.n6433 vss.n6432 51.0489
R34424 vss.n6421 vss.n6419 51.0489
R34425 vss.n6355 vss.n6354 51.0489
R34426 vss.n6343 vss.n6341 51.0489
R34427 vss.n6969 vss.n6968 51.0489
R34428 vss.n6957 vss.n6955 51.0489
R34429 vss.n7158 vss.n7157 51.0489
R34430 vss.n7146 vss.n7144 51.0489
R34431 vss.n6166 vss.n6165 51.0489
R34432 vss.n6154 vss.n6152 51.0489
R34433 vss.n9442 vss.n9402 51.0489
R34434 vss.n9419 vss.n9416 51.0489
R34435 vss.n9565 vss.n9564 51.0489
R34436 vss.n9552 vss.n6075 51.0489
R34437 vss.n7264 vss.n7250 51.0489
R34438 vss.n9548 vss.n6079 51.0489
R34439 vss.n9530 vss.n9529 51.0489
R34440 vss.n9517 vss.n6114 51.0489
R34441 vss.n7245 vss.n6577 51.0489
R34442 vss.n9513 vss.n6118 51.0489
R34443 vss.n7233 vss.n6583 51.0489
R34444 vss.n6755 vss.n6750 51.0489
R34445 vss.n6782 vss.n6729 51.0489
R34446 vss.n6765 vss.n6745 51.0489
R34447 vss.n7075 vss.n7074 51.0489
R34448 vss.n7062 vss.n6797 51.0489
R34449 vss.n6824 vss.n6819 51.0489
R34450 vss.n7058 vss.n6800 51.0489
R34451 vss.n7042 vss.n6829 51.0489
R34452 vss.n6894 vss.n6847 51.0489
R34453 vss.n6875 vss.n6870 51.0489
R34454 vss.n6890 vss.n6851 51.0489
R34455 vss.n9238 vss.n9237 51.0489
R34456 vss.n9225 vss.n6508 51.0489
R34457 vss.n6565 vss.n6560 51.0489
R34458 vss.n9221 vss.n6511 51.0489
R34459 vss.n9205 vss.n6530 51.0489
R34460 vss.n9073 vss.n9068 51.0489
R34461 vss.n9095 vss.n9053 51.0489
R34462 vss.n9083 vss.n9064 51.0489
R34463 vss.n9137 vss.n9100 51.0489
R34464 vss.n9120 vss.n9118 51.0489
R34465 vss.n9351 vss.n9350 51.0489
R34466 vss.n9339 vss.n9337 51.0489
R34467 vss.n9380 vss.n6187 51.0489
R34468 vss.n6204 vss.n6201 51.0489
R34469 vss.n5955 vss.n5954 51.0489
R34470 vss.n5968 vss.n5966 51.0489
R34471 vss.n9705 vss.n9702 51.0489
R34472 vss.n9718 vss.n9716 51.0489
R34473 vss.n2576 vss.n2575 51.0489
R34474 vss.n2589 vss.n2587 51.0489
R34475 vss.n9893 vss.n9892 51.0489
R34476 vss.n9879 vss.n2764 51.0489
R34477 vss.n3283 vss.n3280 51.0489
R34478 vss.n3297 vss.n3293 51.0489
R34479 vss.n9766 vss.n9763 51.0489
R34480 vss.n9779 vss.n9778 51.0489
R34481 vss.n3206 vss.n3203 51.0489
R34482 vss.n3219 vss.n3218 51.0489
R34483 vss.n3005 vss.n2997 51.0489
R34484 vss.n3021 vss.n3020 51.0489
R34485 vss.n5236 vss.n5233 51.0489
R34486 vss.n5249 vss.n5248 51.0489
R34487 vss.n3049 vss.n3046 51.0489
R34488 vss.n3062 vss.n3061 51.0489
R34489 vss.n5106 vss.n5103 51.0489
R34490 vss.n5119 vss.n5118 51.0489
R34491 vss.n5295 vss.n5292 51.0489
R34492 vss.n5308 vss.n5307 51.0489
R34493 vss.n5023 vss.n5020 51.0489
R34494 vss.n5036 vss.n5035 51.0489
R34495 vss.n4904 vss.n4901 51.0489
R34496 vss.n4917 vss.n4916 51.0489
R34497 vss.n9927 vss.n9926 51.0489
R34498 vss.n9913 vss.n2729 51.0489
R34499 vss.n4664 vss.n4663 51.0489
R34500 vss.n9904 vss.n2736 51.0489
R34501 vss.n5629 vss.n5628 51.0489
R34502 vss.n5615 vss.n4681 51.0489
R34503 vss.n5586 vss.n4697 51.0489
R34504 vss.n5606 vss.n5601 51.0489
R34505 vss.n4707 vss.n4702 51.0489
R34506 vss.n4725 vss.n4722 51.0489
R34507 vss.n5543 vss.n4740 51.0489
R34508 vss.n5563 vss.n5558 51.0489
R34509 vss.n4750 vss.n4745 51.0489
R34510 vss.n4768 vss.n4765 51.0489
R34511 vss.n5500 vss.n4783 51.0489
R34512 vss.n5520 vss.n5515 51.0489
R34513 vss.n4793 vss.n4788 51.0489
R34514 vss.n4811 vss.n4808 51.0489
R34515 vss.n5457 vss.n4826 51.0489
R34516 vss.n5477 vss.n5472 51.0489
R34517 vss.n4836 vss.n4831 51.0489
R34518 vss.n4854 vss.n4851 51.0489
R34519 vss.n5414 vss.n4869 51.0489
R34520 vss.n5434 vss.n5429 51.0489
R34521 vss.n4879 vss.n4874 51.0489
R34522 vss.n5348 vss.n5345 51.0489
R34523 vss.n5378 vss.n5361 51.0489
R34524 vss.n5391 vss.n5385 51.0489
R34525 vss.n9825 vss.n9822 51.0489
R34526 vss.n9838 vss.n9837 51.0489
R34527 vss.n2948 vss.n2940 51.0489
R34528 vss.n2964 vss.n2963 51.0489
R34529 vss.n2901 vss.n2893 51.0489
R34530 vss.n2917 vss.n2916 51.0489
R34531 vss.n4945 vss.n4942 51.0489
R34532 vss.n4958 vss.n4957 51.0489
R34533 vss.n5147 vss.n5144 51.0489
R34534 vss.n5160 vss.n5159 51.0489
R34535 vss.n3128 vss.n3125 51.0489
R34536 vss.n3141 vss.n3140 51.0489
R34537 vss.n4494 vss.n4493 51.0489
R34538 vss.n4481 vss.n4479 51.0489
R34539 vss.n4402 vss.n4401 51.0489
R34540 vss.n4389 vss.n4387 51.0489
R34541 vss.n4354 vss.n4353 51.0489
R34542 vss.n4341 vss.n4339 51.0489
R34543 vss.n3754 vss.n3753 51.0489
R34544 vss.n3741 vss.n3739 51.0489
R34545 vss.n4056 vss.n4055 51.0489
R34546 vss.n4043 vss.n4041 51.0489
R34547 vss.n3709 vss.n3708 51.0489
R34548 vss.n3696 vss.n3694 51.0489
R34549 vss.n4110 vss.n4109 51.0489
R34550 vss.n4097 vss.n4095 51.0489
R34551 vss.n3534 vss.n3533 51.0489
R34552 vss.n3521 vss.n3519 51.0489
R34553 vss.n3489 vss.n3488 51.0489
R34554 vss.n3476 vss.n3474 51.0489
R34555 vss.n5777 vss.n5776 51.0489
R34556 vss.n5764 vss.n5762 51.0489
R34557 vss.n4527 vss.n4510 51.0489
R34558 vss.n4517 vss.n4446 51.0489
R34559 vss.n4554 vss.n4425 51.0489
R34560 vss.n4537 vss.n4441 51.0489
R34561 vss.n4601 vss.n4600 51.0489
R34562 vss.n4588 vss.n4569 51.0489
R34563 vss.n4625 vss.n3633 51.0489
R34564 vss.n4584 vss.n4572 51.0489
R34565 vss.n4198 vss.n4197 51.0489
R34566 vss.n4185 vss.n3783 51.0489
R34567 vss.n3824 vss.n3814 51.0489
R34568 vss.n4181 vss.n3786 51.0489
R34569 vss.n4163 vss.n4162 51.0489
R34570 vss.n4150 vss.n3839 51.0489
R34571 vss.n3867 vss.n3862 51.0489
R34572 vss.n4146 vss.n3842 51.0489
R34573 vss.n4132 vss.n3872 51.0489
R34574 vss.n3937 vss.n3890 51.0489
R34575 vss.n3918 vss.n3913 51.0489
R34576 vss.n3933 vss.n3894 51.0489
R34577 vss.n5830 vss.n5829 51.0489
R34578 vss.n5817 vss.n3562 51.0489
R34579 vss.n3621 vss.n3616 51.0489
R34580 vss.n5813 vss.n3565 51.0489
R34581 vss.n5799 vss.n3586 51.0489
R34582 vss.n5667 vss.n5662 51.0489
R34583 vss.n5689 vss.n5647 51.0489
R34584 vss.n5677 vss.n5658 51.0489
R34585 vss.n5731 vss.n5694 51.0489
R34586 vss.n5714 vss.n5712 51.0489
R34587 vss.n9981 vss.n9980 51.0489
R34588 vss.n9968 vss.n9966 51.0489
R34589 vss.n2682 vss.n2642 51.0489
R34590 vss.n2663 vss.n2660 51.0489
R34591 vss.n3414 vss.n3413 51.0489
R34592 vss.n3401 vss.n3399 51.0489
R34593 vss.n4011 vss.n4010 51.0489
R34594 vss.n3998 vss.n3996 51.0489
R34595 vss.n4278 vss.n4277 51.0489
R34596 vss.n4265 vss.n4263 51.0489
R34597 vss.n5920 vss.n5919 51.0489
R34598 vss.n5908 vss.n5906 51.0489
R34599 vss.n14069 vss.n14066 51.0489
R34600 vss.n14082 vss.n14081 51.0489
R34601 vss.n10124 vss.n10121 51.0489
R34602 vss.n10137 vss.n10136 51.0489
R34603 vss.n12882 vss.n12879 51.0489
R34604 vss.n12895 vss.n12894 51.0489
R34605 vss.n10165 vss.n10162 51.0489
R34606 vss.n10178 vss.n10177 51.0489
R34607 vss.n12431 vss.n12428 51.0489
R34608 vss.n12444 vss.n12443 51.0489
R34609 vss.n11760 vss.n11757 51.0489
R34610 vss.n11773 vss.n11772 51.0489
R34611 vss.n12476 vss.n12473 51.0489
R34612 vss.n12489 vss.n12488 51.0489
R34613 vss.n2318 vss.n2310 51.0489
R34614 vss.n2334 vss.n2333 51.0489
R34615 vss.n12301 vss.n12298 51.0489
R34616 vss.n12314 vss.n12313 51.0489
R34617 vss.n12346 vss.n12343 51.0489
R34618 vss.n12359 vss.n12358 51.0489
R34619 vss.n10242 vss.n10239 51.0489
R34620 vss.n10255 vss.n10254 51.0489
R34621 vss.n2422 vss.n2419 51.0489
R34622 vss.n2435 vss.n2434 51.0489
R34623 vss.n2378 vss.n2370 51.0489
R34624 vss.n2394 vss.n2393 51.0489
R34625 vss.n10043 vss.n10034 51.0489
R34626 vss.n10056 vss.n10054 51.0489
R34627 vss.n10039 vss.n2099 51.0489
R34628 vss.n2117 vss.n2114 51.0489
R34629 vss.n12926 vss.n10081 51.0489
R34630 vss.n12939 vss.n12938 51.0489
R34631 vss.n2502 vss.n2499 51.0489
R34632 vss.n2515 vss.n2514 51.0489
R34633 vss.n13074 vss.n13073 51.0489
R34634 vss.n13060 vss.n2140 51.0489
R34635 vss.n12104 vss.n11848 51.0489
R34636 vss.n12119 vss.n12118 51.0489
R34637 vss.n11819 vss.n11811 51.0489
R34638 vss.n12133 vss.n12132 51.0489
R34639 vss.n12157 vss.n11804 51.0489
R34640 vss.n12172 vss.n12171 51.0489
R34641 vss.n12255 vss.n12254 51.0489
R34642 vss.n12270 vss.n12269 51.0489
R34643 vss.n12201 vss.n12193 51.0489
R34644 vss.n12233 vss.n12207 51.0489
R34645 vss.n11731 vss.n11723 51.0489
R34646 vss.n12224 vss.n12223 51.0489
R34647 vss.n12553 vss.n11717 51.0489
R34648 vss.n12568 vss.n12567 51.0489
R34649 vss.n12584 vss.n12583 51.0489
R34650 vss.n12575 vss.n11634 51.0489
R34651 vss.n11652 vss.n11644 51.0489
R34652 vss.n11668 vss.n11658 51.0489
R34653 vss.n12835 vss.n12834 51.0489
R34654 vss.n12850 vss.n12849 51.0489
R34655 vss.n12783 vss.n12775 51.0489
R34656 vss.n12815 vss.n12789 51.0489
R34657 vss.n10096 vss.n10088 51.0489
R34658 vss.n12806 vss.n12805 51.0489
R34659 vss.n12084 vss.n11860 51.0489
R34660 vss.n11880 vss.n11878 51.0489
R34661 vss.n10493 vss.n10492 51.0489
R34662 vss.n10480 vss.n10479 51.0489
R34663 vss.n10714 vss.n10713 51.0489
R34664 vss.n10701 vss.n10700 51.0489
R34665 vss.n11028 vss.n11027 51.0489
R34666 vss.n11015 vss.n11014 51.0489
R34667 vss.n11135 vss.n11134 51.0489
R34668 vss.n11123 vss.n11122 51.0489
R34669 vss.n9873 vss.t77 43.8854
R34670 vss.t1061 vss.n8153 42.9351
R34671 vss.n3281 vss.t339 42.9351
R34672 vss.n14154 vss.t1275 42.9351
R34673 vss.t318 vss.n10042 42.9351
R34674 vss.n8219 vss.n8052 42.3082
R34675 vss.n13078 vss.n13077 42.3082
R34676 vss.n8123 vss.n8122 42.14
R34677 vss.n9930 vss.n9929 42.14
R34678 vss.n13935 vss.n458 42.14
R34679 vss.n10035 vss.n2071 42.14
R34680 vss.n0 vss.t1110 41.7571
R34681 vss.n14760 vss.t1082 41.7571
R34682 vss.n2031 vss.t1461 41.7571
R34683 vss.n12664 vss.t1345 41.7571
R34684 vss.n11399 vss.t421 41.7571
R34685 vss.n11400 vss.t20 41.7571
R34686 vss.n10767 vss.t320 41.7571
R34687 vss.n10768 vss.t577 41.7571
R34688 vss.n10546 vss.t1389 41.7571
R34689 vss.n10547 vss.t12 41.7571
R34690 vss.n11971 vss.t306 41.7571
R34691 vss.n11970 vss.t959 41.7571
R34692 vss.n12014 vss.t701 41.7571
R34693 vss.n12013 vss.t1472 41.7571
R34694 vss.n11597 vss.t1246 41.7571
R34695 vss.n11596 vss.t842 41.7571
R34696 vss.n10844 vss.t684 41.7571
R34697 vss.n10843 vss.t1394 41.7571
R34698 vss.n10988 vss.t694 41.7571
R34699 vss.n10989 vss.t994 41.7571
R34700 vss.n11451 vss.t1100 41.7571
R34701 vss.n11450 vss.t594 41.7571
R34702 vss.n12700 vss.t1251 41.7571
R34703 vss.n12699 vss.t1002 41.7571
R34704 vss.n11835 vss.t539 41.7571
R34705 vss.n11834 vss.t1039 41.7571
R34706 vss.n13019 vss.t643 41.7571
R34707 vss.n13020 vss.t501 41.7571
R34708 vss.n12958 vss.t856 41.7571
R34709 vss.n12959 vss.t620 41.7571
R34710 vss.n13201 vss.t349 41.7571
R34711 vss.n13202 vss.t1496 41.7571
R34712 vss.n1977 vss.t366 41.7571
R34713 vss.n1978 vss.t887 41.7571
R34714 vss.n14144 vss.t1274 41.7571
R34715 vss.n14143 vss.t817 41.7571
R34716 vss.n14248 vss.t1190 41.7571
R34717 vss.n14249 vss.t1333 41.7571
R34718 vss.n14182 vss.t1523 41.7571
R34719 vss.n14181 vss.t1317 41.7571
R34720 vss.n13551 vss.t1263 41.7571
R34721 vss.n13550 vss.t1019 41.7571
R34722 vss.n13320 vss.t251 41.7571
R34723 vss.n13319 vss.t915 41.7571
R34724 vss.n13858 vss.t680 41.7571
R34725 vss.n13857 vss.t821 41.7571
R34726 vss.n13862 vss.t808 41.7571
R34727 vss.n13861 vss.t1025 41.7571
R34728 vss.n13370 vss.t1414 41.7571
R34729 vss.n13369 vss.t112 41.7571
R34730 vss.n14644 vss.t1051 41.7571
R34731 vss.n14643 vss.t1498 41.7571
R34732 vss.n13753 vss.t309 41.7571
R34733 vss.n13752 vss.t796 41.7571
R34734 vss.n13757 vss.t1418 41.7571
R34735 vss.n13756 vss.t1027 41.7571
R34736 vss.n13450 vss.t1434 41.7571
R34737 vss.n13449 vss.t1392 41.7571
R34738 vss.n14449 vss.t835 41.7571
R34739 vss.n14448 vss.t382 41.7571
R34740 vss.n13648 vss.t270 41.7571
R34741 vss.n13647 vss.t827 41.7571
R34742 vss.n13652 vss.t632 41.7571
R34743 vss.n13651 vss.t1041 41.7571
R34744 vss.n13530 vss.t1385 41.7571
R34745 vss.n13529 vss.t108 41.7571
R34746 vss.n14254 vss.t157 41.7571
R34747 vss.n14253 vss.t503 41.7571
R34748 vss.n14301 vss.t755 41.7571
R34749 vss.n14300 vss.t1478 41.7571
R34750 vss.n13704 vss.t1290 41.7571
R34751 vss.n13703 vss.t992 41.7571
R34752 vss.n14367 vss.t1103 41.7571
R34753 vss.n14368 vss.t1351 41.7571
R34754 vss.n14413 vss.t1209 41.7571
R34755 vss.n14414 vss.t467 41.7571
R34756 vss.n14496 vss.t267 41.7571
R34757 vss.n14495 vss.t1078 41.7571
R34758 vss.n13809 vss.t717 41.7571
R34759 vss.n13808 vss.t48 41.7571
R34760 vss.n14562 vss.t363 41.7571
R34761 vss.n14563 vss.t1325 41.7571
R34762 vss.n14608 vss.t75 41.7571
R34763 vss.n14609 vss.t1337 41.7571
R34764 vss.n14691 vss.t347 41.7571
R34765 vss.n14690 vss.t475 41.7571
R34766 vss.n14757 vss.t1113 41.7571
R34767 vss.n14758 vss.t614 41.7571
R34768 vss.n360 vss.t1405 41.7571
R34769 vss.n361 vss.t1353 41.7571
R34770 vss.n14141 vss.t974 41.7571
R34771 vss.n14140 vss.t881 41.7571
R34772 vss.n14095 vss.t1226 41.7571
R34773 vss.n14094 vss.t394 41.7571
R34774 vss.n642 vss.t137 41.7571
R34775 vss.n641 vss.t24 41.7571
R34776 vss.n13239 vss.t528 41.7571
R34777 vss.n13238 vss.t891 41.7571
R34778 vss.n1808 vss.t418 41.7571
R34779 vss.n1807 vss.t1160 41.7571
R34780 vss.n1647 vss.t584 41.7571
R34781 vss.n1648 vss.t622 41.7571
R34782 vss.n1401 vss.t280 41.7571
R34783 vss.n1402 vss.t998 41.7571
R34784 vss.n1912 vss.t151 41.7571
R34785 vss.n1911 vss.t600 41.7571
R34786 vss.n1352 vss.t765 41.7571
R34787 vss.n1353 vss.t1084 41.7571
R34788 vss.n1092 vss.t924 41.7571
R34789 vss.n1093 vss.t1373 41.7571
R34790 vss.n1354 vss.t543 41.7571
R34791 vss.n1355 vss.t14 41.7571
R34792 vss.n1907 vss.t1277 41.7571
R34793 vss.n1908 vss.t848 41.7571
R34794 vss.n1399 vss.t1456 41.7571
R34795 vss.n1400 vss.t175 41.7571
R34796 vss.n1406 vss.t1408 41.7571
R34797 vss.n1407 vss.t616 41.7571
R34798 vss.n1485 vss.t172 41.7571
R34799 vss.n1486 vss.t499 41.7571
R34800 vss.n1652 vss.t1532 41.7571
R34801 vss.n1651 vss.t1361 41.7571
R34802 vss.n1803 vss.t290 41.7571
R34803 vss.n1804 vss.t1023 41.7571
R34804 vss.n1696 vss.t909 41.7571
R34805 vss.n1695 vss.t658 41.7571
R34806 vss.n793 vss.t1175 41.7571
R34807 vss.n1488 vss.t507 41.7571
R34808 vss.n1566 vss.t1430 41.7571
R34809 vss.n1567 vss.t398 41.7571
R34810 vss.n554 vss.t674 41.7571
R34811 vss.n553 vss.t654 41.7571
R34812 vss.n555 vss.t302 41.7571
R34813 vss.n592 vss.t953 41.7571
R34814 vss.n13956 vss.t768 41.7571
R34815 vss.n13955 vss.t110 41.7571
R34816 vss.n594 vss.t359 41.7571
R34817 vss.n1568 vss.t18 41.7571
R34818 vss.n891 vss.t936 41.7571
R34819 vss.n890 vss.t505 41.7571
R34820 vss.n14030 vss.t763 41.7571
R34821 vss.n14031 vss.t396 41.7571
R34822 vss.n14025 vss.t295 41.7571
R34823 vss.n14026 vss.t1000 41.7571
R34824 vss.n706 vss.t781 41.7571
R34825 vss.n13156 vss.t877 41.7571
R34826 vss.n705 vss.t115 41.7571
R34827 vss.n1136 vss.t825 41.7571
R34828 vss.n1982 vss.t324 41.7571
R34829 vss.n1983 vss.t579 41.7571
R34830 vss.n2026 vss.t522 41.7571
R34831 vss.n2027 vss.t1321 41.7571
R34832 vss.n9366 vss.t1091 41.7571
R34833 vss.n9365 vss.t1080 41.7571
R34834 vss.n9196 vss.t1205 41.7571
R34835 vss.n9195 vss.t1035 41.7571
R34836 vss.n7989 vss.t1060 41.7571
R34837 vss.n7990 vss.t864 41.7571
R34838 vss.n8059 vss.t184 41.7571
R34839 vss.n8058 vss.t961 41.7571
R34840 vss.n8246 vss.t560 41.7571
R34841 vss.n8247 vss.t1508 41.7571
R34842 vss.n8180 vss.t372 41.7571
R34843 vss.n8179 vss.t1347 41.7571
R34844 vss.n7905 vss.t810 41.7571
R34845 vss.n7904 vss.t66 41.7571
R34846 vss.n8737 vss.t1297 41.7571
R34847 vss.n8738 vss.t612 41.7571
R34848 vss.n7810 vss.t164 41.7571
R34849 vss.n7811 vss.t497 41.7571
R34850 vss.n8378 vss.t607 41.7571
R34851 vss.n8377 vss.t866 41.7571
R34852 vss.n8856 vss.t785 41.7571
R34853 vss.n8857 vss.t1074 41.7571
R34854 vss.n8790 vss.t1012 41.7571
R34855 vss.n8789 vss.t206 41.7571
R34856 vss.n8476 vss.t793 41.7571
R34857 vss.n8475 vss.t179 41.7571
R34858 vss.n7907 vss.t721 41.7571
R34859 vss.n7908 vss.t586 41.7571
R34860 vss.n7873 vss.t96 41.7571
R34861 vss.n7872 vss.t913 41.7571
R34862 vss.n8329 vss.t1229 41.7571
R34863 vss.n8328 vss.t1154 41.7571
R34864 vss.n8404 vss.t149 41.7571
R34865 vss.n8403 vss.t957 41.7571
R34866 vss.n8427 vss.t99 41.7571
R34867 vss.n8426 vss.t596 41.7571
R34868 vss.n8502 vss.t1107 41.7571
R34869 vss.n8501 vss.t1029 41.7571
R34870 vss.n8975 vss.t263 41.7571
R34871 vss.n8976 vss.t1506 41.7571
R34872 vss.n8909 vss.t311 41.7571
R34873 vss.n8908 vss.t10 41.7571
R34874 vss.n7496 vss.t1469 41.7571
R34875 vss.n7495 vss.t216 41.7571
R34876 vss.n8473 vss.t945 41.7571
R34877 vss.n8472 vss.t1031 41.7571
R34878 vss.n8862 vss.t196 41.7571
R34879 vss.n8861 vss.t573 41.7571
R34880 vss.n7588 vss.t837 41.7571
R34881 vss.n7589 vss.t634 41.7571
R34882 vss.n8375 vss.t668 41.7571
R34883 vss.n8374 vss.t1033 41.7571
R34884 vss.n8743 vss.t1536 41.7571
R34885 vss.n8742 vss.t1377 41.7571
R34886 vss.n7731 vss.t224 41.7571
R34887 vss.n7732 vss.t6 41.7571
R34888 vss.n8257 vss.t774 41.7571
R34889 vss.n8256 vss.t947 41.7571
R34890 vss.n8252 vss.t413 41.7571
R34891 vss.n8251 vss.t384 41.7571
R34892 vss.n7952 vss.t652 41.7571
R34893 vss.n7953 vss.t485 41.7571
R34894 vss.n9640 vss.t690 41.7571
R34895 vss.n9639 vss.t1006 41.7571
R34896 vss.n9636 vss.t1530 41.7571
R34897 vss.n9635 vss.t636 41.7571
R34898 vss.n6052 vss.t732 41.7571
R34899 vss.n6053 vss.t212 41.7571
R34900 vss.n7224 vss.t533 41.7571
R34901 vss.n7223 vss.t44 41.7571
R34902 vss.n7050 vss.t556 41.7571
R34903 vss.n7049 vss.t1158 41.7571
R34904 vss.n6671 vss.t1119 41.7571
R34905 vss.n6672 vss.t1331 41.7571
R34906 vss.n7033 vss.t671 41.7571
R34907 vss.n7032 vss.t919 41.7571
R34908 vss.n9213 vss.t1411 41.7571
R34909 vss.n9212 vss.t590 41.7571
R34910 vss.n6444 vss.t901 41.7571
R34911 vss.n6445 vss.t1492 41.7571
R34912 vss.n6367 vss.t190 41.7571
R34913 vss.n6368 vss.t1357 41.7571
R34914 vss.n9253 vss.t1466 41.7571
R34915 vss.n9254 vss.t1335 41.7571
R34916 vss.n9248 vss.t256 41.7571
R34917 vss.n9249 vss.t58 41.7571
R34918 vss.n6903 vss.t141 41.7571
R34919 vss.n6904 vss.t798 41.7571
R34920 vss.n6986 vss.t334 41.7571
R34921 vss.n6985 vss.t1315 41.7571
R34922 vss.n6981 vss.t548 41.7571
R34923 vss.n6982 vss.t483 41.7571
R34924 vss.n7090 vss.t986 41.7571
R34925 vss.n7091 vss.t1371 41.7571
R34926 vss.n7085 vss.t328 41.7571
R34927 vss.n7086 vss.t996 41.7571
R34928 vss.n6716 vss.t247 41.7571
R34929 vss.n6715 vss.t447 41.7571
R34930 vss.n7177 vss.t86 41.7571
R34931 vss.n7176 vss.t214 41.7571
R34932 vss.n7170 vss.t1282 41.7571
R34933 vss.n7171 vss.t1502 41.7571
R34934 vss.n6094 vss.t904 41.7571
R34935 vss.n6093 vss.t823 41.7571
R34936 vss.n6095 vss.t259 41.7571
R34937 vss.n6132 vss.t990 41.7571
R34938 vss.n9505 vss.t454 41.7571
R34939 vss.n9504 vss.t106 41.7571
R34940 vss.n6134 vss.t1294 41.7571
R34941 vss.n7172 vss.t1341 41.7571
R34942 vss.n9429 vss.t942 41.7571
R34943 vss.n9428 vss.t1488 41.7571
R34944 vss.n9579 vss.t231 41.7571
R34945 vss.n9580 vss.t511 41.7571
R34946 vss.n9574 vss.t1301 41.7571
R34947 vss.n9575 vss.t1043 41.7571
R34948 vss.n6545 vss.t1437 41.7571
R34949 vss.n6544 vss.t889 41.7571
R34950 vss.n9146 vss.t461 41.7571
R34951 vss.n9147 vss.t860 41.7571
R34952 vss.n9149 vss.t898 41.7571
R34953 vss.n9148 vss.t473 41.7571
R34954 vss.n9362 vss.t536 41.7571
R34955 vss.n9363 vss.t610 41.7571
R34956 vss.n9741 vss.t779 41.7571
R34957 vss.n9742 vss.t70 41.7571
R34958 vss.n9786 vss.t714 41.7571
R34959 vss.n9787 vss.t477 41.7571
R34960 vss.n3225 vss.t493 41.7571
R34961 vss.n3226 vss.t1359 41.7571
R34962 vss.n5211 vss.t1234 41.7571
R34963 vss.n5212 vss.t68 41.7571
R34964 vss.n5256 vss.t1187 41.7571
R34965 vss.n5257 vss.t481 41.7571
R34966 vss.n3068 vss.t200 41.7571
R34967 vss.n3069 vss.t1367 41.7571
R34968 vss.n5270 vss.t1538 41.7571
R34969 vss.n5271 vss.t819 41.7571
R34970 vss.n5315 vss.t706 41.7571
R34971 vss.n5316 vss.t1349 41.7571
R34972 vss.n5042 vss.t1164 41.7571
R34973 vss.n5043 vss.t1381 41.7571
R34974 vss.n5329 vss.t193 41.7571
R34975 vss.n5328 vss.t181 41.7571
R34976 vss.n4642 vss.t29 41.7571
R34977 vss.n4641 vss.t1045 41.7571
R34978 vss.n4633 vss.t751 41.7571
R34979 vss.n4632 vss.t588 41.7571
R34980 vss.n5203 vss.t660 41.7571
R34981 vss.n5204 vss.t846 41.7571
R34982 vss.n5082 vss.t805 41.7571
R34983 vss.n5083 vss.t1156 41.7571
R34984 vss.n5079 vss.t338 41.7571
R34985 vss.n5080 vss.t879 41.7571
R34986 vss.n4880 vss.t1527 41.7571
R34987 vss.n4881 vss.t602 41.7571
R34988 vss.n5355 vss.t743 41.7571
R34989 vss.n5354 vss.t56 41.7571
R34990 vss.n9845 vss.t409 41.7571
R34991 vss.n9846 vss.t16 41.7571
R34992 vss.n2970 vss.t1424 41.7571
R34993 vss.n2969 vss.t1319 41.7571
R34994 vss.n2923 vss.t791 41.7571
R34995 vss.n2922 vss.t471 41.7571
R34996 vss.n5326 vss.t1244 41.7571
R34997 vss.n5325 vss.t965 41.7571
R34998 vss.n5321 vss.t605 41.7571
R34999 vss.n5320 vss.t1086 41.7571
R35000 vss.n4965 vss.t1236 41.7571
R35001 vss.n4966 vss.t1510 41.7571
R35002 vss.n5267 vss.t1222 41.7571
R35003 vss.n5266 vss.t967 41.7571
R35004 vss.n5262 vss.t2 41.7571
R35005 vss.n5261 vss.t1486 41.7571
R35006 vss.n5167 vss.t1309 41.7571
R35007 vss.n5168 vss.t509 41.7571
R35008 vss.n5208 vss.t1421 41.7571
R35009 vss.n5207 vss.t788 41.7571
R35010 vss.n9792 vss.t970 41.7571
R35011 vss.n9791 vss.t626 41.7571
R35012 vss.n3148 vss.t709 41.7571
R35013 vss.n3149 vss.t1343 41.7571
R35014 vss.n9738 vss.t1198 41.7571
R35015 vss.n9737 vss.t50 41.7571
R35016 vss.n9734 vss.t131 41.7571
R35017 vss.n9733 vss.t218 41.7571
R35018 vss.n4363 vss.t1260 41.7571
R35019 vss.n4364 vss.t1504 41.7571
R35020 vss.n3718 vss.t1442 41.7571
R35021 vss.n3719 vss.t1494 41.7571
R35022 vss.n3498 vss.t1213 41.7571
R35023 vss.n3499 vss.t618 41.7571
R35024 vss.n5790 vss.t1137 41.7571
R35025 vss.n5789 vss.t1004 41.7571
R35026 vss.n3579 vss.t739 41.7571
R35027 vss.n3578 vss.t1476 41.7571
R35028 vss.n4123 vss.t1195 41.7571
R35029 vss.n4122 vss.t850 41.7571
R35030 vss.n3855 vss.t427 41.7571
R35031 vss.n4065 vss.t1152 41.7571
R35032 vss.n4207 vss.t235 41.7571
R35033 vss.n4208 vss.t1037 41.7571
R35034 vss.n4616 vss.t1268 41.7571
R35035 vss.n4615 vss.t598 41.7571
R35036 vss.n4507 vss.t725 41.7571
R35037 vss.n4506 vss.t949 41.7571
R35038 vss.n9991 vss.t519 41.7571
R35039 vss.n9992 vss.t1323 41.7571
R35040 vss.n2673 vss.t406 41.7571
R35041 vss.n2672 vss.t1076 41.7571
R35042 vss.n3601 vss.t514 41.7571
R35043 vss.n3600 vss.t885 41.7571
R35044 vss.n5740 vss.t1514 41.7571
R35045 vss.n5741 vss.t64 41.7571
R35046 vss.n5743 vss.t747 41.7571
R35047 vss.n5742 vss.t380 41.7571
R35048 vss.n3424 vss.t648 41.7571
R35049 vss.n3425 vss.t4 41.7571
R35050 vss.n5845 vss.t728 41.7571
R35051 vss.n5846 vss.t567 41.7571
R35052 vss.n5840 vss.t330 41.7571
R35053 vss.n5841 vss.t52 41.7571
R35054 vss.n3946 vss.t118 41.7571
R35055 vss.n3947 vss.t449 41.7571
R35056 vss.n4076 vss.t353 41.7571
R35057 vss.n4075 vss.t1484 41.7571
R35058 vss.n4021 vss.t432 41.7571
R35059 vss.n4022 vss.t392 41.7571
R35060 vss.n4070 vss.t1127 41.7571
R35061 vss.n4071 vss.t624 41.7571
R35062 vss.n3802 vss.t526 41.7571
R35063 vss.n4066 vss.t963 41.7571
R35064 vss.n3801 vss.t374 41.7571
R35065 vss.n3800 vss.t868 41.7571
R35066 vss.n4212 vss.t1256 41.7571
R35067 vss.n4213 vss.t1072 41.7571
R35068 vss.n4288 vss.t1453 41.7571
R35069 vss.n4289 vss.t487 41.7571
R35070 vss.n4368 vss.t489 41.7571
R35071 vss.n4367 vss.t569 41.7571
R35072 vss.n4611 vss.t696 41.7571
R35073 vss.n4612 vss.t917 41.7571
R35074 vss.n4457 vss.t457 41.7571
R35075 vss.n4458 vss.t443 41.7571
R35076 vss.n4460 vss.t160 41.7571
R35077 vss.n4459 vss.t581 41.7571
R35078 vss.n5932 vss.t1065 41.7571
R35079 vss.n5933 vss.t479 41.7571
R35080 vss.n10012 vss.t1183 41.7571
R35081 vss.n10011 vss.t38 41.7571
R35082 vss.n2557 vss.t1202 41.7571
R35083 vss.n5935 vss.t1015 41.7571
R35084 vss.n9684 vss.t1446 41.7571
R35085 vss.n9683 vss.t40 41.7571
R35086 vss.n5936 vss.t565 41.7571
R35087 vss.n9583 vss.t1215 41.7571
R35088 vss.n9630 vss.t737 41.7571
R35089 vss.n9629 vss.t42 41.7571
R35090 vss.n9585 vss.t1141 41.7571
R35091 vss.n9584 vss.t1017 41.7571
R35092 vss.n14089 vss.t922 41.7571
R35093 vss.n14088 vss.t36 41.7571
R35094 vss.n12912 vss.t1449 41.7571
R35095 vss.n12911 vss.t1474 41.7571
R35096 vss.n12857 vss.t283 41.7571
R35097 vss.n12858 vss.t802 41.7571
R35098 vss.n11676 vss.t830 41.7571
R35099 vss.n11675 vss.t883 41.7571
R35100 vss.n12902 vss.t287 41.7571
R35101 vss.n12903 vss.t1480 41.7571
R35102 vss.n10184 vss.t298 41.7571
R35103 vss.n10185 vss.t386 41.7571
R35104 vss.n12406 vss.t640 41.7571
R35105 vss.n12407 vss.t1396 41.7571
R35106 vss.n12538 vss.t144 41.7571
R35107 vss.n12537 vss.t72 41.7571
R35108 vss.n12241 vss.t92 41.7571
R35109 vss.n12240 vss.t852 41.7571
R35110 vss.n12534 vss.t227 41.7571
R35111 vss.n12533 vss.t210 41.7571
R35112 vss.n12495 vss.t220 41.7571
R35113 vss.n12496 vss.t1500 41.7571
R35114 vss.n2340 vss.t980 41.7571
R35115 vss.n2339 vss.t1363 41.7571
R35116 vss.n12276 vss.t415 41.7571
R35117 vss.n12277 vss.t592 41.7571
R35118 vss.n12142 vss.t341 41.7571
R35119 vss.n12141 vss.t800 41.7571
R35120 vss.n12139 vss.t1123 41.7571
R35121 vss.n12138 vss.t873 41.7571
R35122 vss.n12321 vss.t1170 41.7571
R35123 vss.n12322 vss.t1339 41.7571
R35124 vss.n12366 vss.t932 41.7571
R35125 vss.n12367 vss.t1327 41.7571
R35126 vss.n12403 vss.t1401 41.7571
R35127 vss.n12404 vss.t875 41.7571
R35128 vss.n12451 vss.t463 41.7571
R35129 vss.n12452 vss.t8 41.7571
R35130 vss.n10262 vss.t438 41.7571
R35131 vss.n10263 vss.t1355 41.7571
R35132 vss.n10301 vss.t1239 41.7571
R35133 vss.n10300 vss.t844 41.7571
R35134 vss.n12908 vss.t1304 41.7571
R35135 vss.n12907 vss.t469 41.7571
R35136 vss.n2442 vss.t134 41.7571
R35137 vss.n2443 vss.t390 41.7571
R35138 vss.n10016 vss.t1519 41.7571
R35139 vss.n10015 vss.t858 41.7571
R35140 vss.n12954 vss.t677 41.7571
R35141 vss.n12955 vss.t54 41.7571
R35142 vss.n10066 vss.t274 41.7571
R35143 vss.n10065 vss.t46 41.7571
R35144 vss.n12964 vss.t1167 41.7571
R35145 vss.n12963 vss.t204 41.7571
R35146 vss.n2521 vss.t60 41.7571
R35147 vss.n2522 vss.t571 41.7571
R35148 vss.n2264 vss.t186 41.7571
R35149 vss.n2263 vss.t1512 41.7571
R35150 vss.n11890 vss.t894 41.7571
R35151 vss.n11889 vss.t1021 41.7571
R35152 vss.n11891 vss.t127 41.7571
R35153 vss.n11923 vss.t177 41.7571
R35154 vss.n11925 vss.t1069 41.7571
R35155 vss.n11924 vss.t1482 41.7571
R35156 vss.n10503 vss.t759 41.7571
R35157 vss.n10504 vss.t388 41.7571
R35158 vss.n12616 vss.t1144 41.7571
R35159 vss.n12617 vss.t202 41.7571
R35160 vss.n12611 vss.t238 41.7571
R35161 vss.n12612 vss.t1047 41.7571
R35162 vss.n10679 vss.t870 41.7571
R35163 vss.n10680 vss.t445 41.7571
R35164 vss.n11551 vss.t664 41.7571
R35165 vss.n11550 vss.t1365 41.7571
R35166 vss.n10724 vss.t1130 41.7571
R35167 vss.n10725 vss.t1490 41.7571
R35168 vss.n11545 vss.t169 41.7571
R35169 vss.n11546 vss.t22 41.7571
R35170 vss.n11540 vss.t402 41.7571
R35171 vss.n11541 vss.t951 41.7571
R35172 vss.n10974 vss.t377 41.7571
R35173 vss.n10975 vss.t862 41.7571
R35174 vss.n10993 vss.t814 41.7571
R35175 vss.n10994 vss.t1369 41.7571
R35176 vss.n11038 vss.t928 41.7571
R35177 vss.n11039 vss.t1329 41.7571
R35178 vss.n11404 vss.t103 41.7571
R35179 vss.n11403 vss.t208 41.7571
R35180 vss.n10339 vss.t977 41.7571
R35181 vss.n11447 vss.t955 41.7571
R35182 vss.n10340 vss.t1217 41.7571
R35183 vss.n10372 vss.t656 41.7571
R35184 vss.n10373 vss.t1096 41.7571
R35185 vss.n11041 vss.t575 41.7571
R35186 vss.n11147 vss.t356 41.7571
R35187 vss.n11148 vss.t1379 41.7571
R35188 vss.n12662 vss.t122 41.7571
R35189 vss.n12663 vss.t1375 41.7571
R35190 vss.n9874 vss.n9873 41.3025
R35191 vss.n10406 vss.n10405 35.2919
R35192 vss.n10405 vss.n10404 35.2919
R35193 vss.n10404 vss.n2042 35.2919
R35194 vss.n13143 vss.n2042 35.2919
R35195 vss.n13143 vss.n13142 35.2919
R35196 vss.n13142 vss.n13141 35.2919
R35197 vss.n12640 vss.n12631 35.2919
R35198 vss.n12646 vss.n12631 35.2919
R35199 vss.n12647 vss.n12646 35.2919
R35200 vss.n12657 vss.n12647 35.2919
R35201 vss.n12657 vss.n12656 35.2919
R35202 vss.n12656 vss.n12655 35.2919
R35203 vss.n12675 vss.n10383 35.2919
R35204 vss.n12681 vss.n10383 35.2919
R35205 vss.n12682 vss.n12681 35.2919
R35206 vss.n12683 vss.n12682 35.2919
R35207 vss.n12684 vss.n12683 35.2919
R35208 vss.n12688 vss.n12684 35.2919
R35209 vss.n11425 vss.n11414 35.2919
R35210 vss.n11431 vss.n11414 35.2919
R35211 vss.n11432 vss.n11431 35.2919
R35212 vss.n11433 vss.n11432 35.2919
R35213 vss.n11434 vss.n11433 35.2919
R35214 vss.n11438 vss.n11434 35.2919
R35215 vss.n11378 vss.n11367 35.2919
R35216 vss.n11384 vss.n11367 35.2919
R35217 vss.n11385 vss.n11384 35.2919
R35218 vss.n11386 vss.n11385 35.2919
R35219 vss.n11387 vss.n11386 35.2919
R35220 vss.n11391 vss.n11387 35.2919
R35221 vss.n10953 vss.n10942 35.2919
R35222 vss.n10959 vss.n10942 35.2919
R35223 vss.n10960 vss.n10959 35.2919
R35224 vss.n10961 vss.n10960 35.2919
R35225 vss.n10962 vss.n10961 35.2919
R35226 vss.n10966 vss.n10962 35.2919
R35227 vss.n10790 vss.n10779 35.2919
R35228 vss.n10796 vss.n10779 35.2919
R35229 vss.n10797 vss.n10796 35.2919
R35230 vss.n10798 vss.n10797 35.2919
R35231 vss.n10799 vss.n10798 35.2919
R35232 vss.n10803 vss.n10799 35.2919
R35233 vss.n10746 vss.n10735 35.2919
R35234 vss.n10752 vss.n10735 35.2919
R35235 vss.n10753 vss.n10752 35.2919
R35236 vss.n10754 vss.n10753 35.2919
R35237 vss.n10755 vss.n10754 35.2919
R35238 vss.n10759 vss.n10755 35.2919
R35239 vss.n11572 vss.n11561 35.2919
R35240 vss.n11578 vss.n11561 35.2919
R35241 vss.n11579 vss.n11578 35.2919
R35242 vss.n11580 vss.n11579 35.2919
R35243 vss.n11581 vss.n11580 35.2919
R35244 vss.n11585 vss.n11581 35.2919
R35245 vss.n10569 vss.n10558 35.2919
R35246 vss.n10575 vss.n10558 35.2919
R35247 vss.n10576 vss.n10575 35.2919
R35248 vss.n10577 vss.n10576 35.2919
R35249 vss.n10578 vss.n10577 35.2919
R35250 vss.n10582 vss.n10578 35.2919
R35251 vss.n10525 vss.n10514 35.2919
R35252 vss.n10531 vss.n10514 35.2919
R35253 vss.n10532 vss.n10531 35.2919
R35254 vss.n10533 vss.n10532 35.2919
R35255 vss.n10534 vss.n10533 35.2919
R35256 vss.n10538 vss.n10534 35.2919
R35257 vss.n11946 vss.n11935 35.2919
R35258 vss.n11952 vss.n11935 35.2919
R35259 vss.n11953 vss.n11952 35.2919
R35260 vss.n11954 vss.n11953 35.2919
R35261 vss.n11955 vss.n11954 35.2919
R35262 vss.n11959 vss.n11955 35.2919
R35263 vss.n12066 vss.n12065 35.2919
R35264 vss.n12067 vss.n12066 35.2919
R35265 vss.n12067 vss.n11855 35.2919
R35266 vss.n12092 vss.n11855 35.2919
R35267 vss.n12093 vss.n12092 35.2919
R35268 vss.n12094 vss.n12093 35.2919
R35269 vss.n12055 vss.n11912 35.2919
R35270 vss.n12055 vss.n12054 35.2919
R35271 vss.n12054 vss.n11913 35.2919
R35272 vss.n12050 vss.n11913 35.2919
R35273 vss.n12050 vss.n12049 35.2919
R35274 vss.n12049 vss.n12048 35.2919
R35275 vss.n12026 vss.n12025 35.2919
R35276 vss.n12027 vss.n12026 35.2919
R35277 vss.n12027 vss.n11984 35.2919
R35278 vss.n12031 vss.n11984 35.2919
R35279 vss.n12040 vss.n12031 35.2919
R35280 vss.n12040 vss.n12039 35.2919
R35281 vss.n12003 vss.n12000 35.2919
R35282 vss.n12003 vss.n12002 35.2919
R35283 vss.n12002 vss.n10601 35.2919
R35284 vss.n12605 vss.n10601 35.2919
R35285 vss.n12605 vss.n12604 35.2919
R35286 vss.n12604 vss.n12603 35.2919
R35287 vss.n10667 vss.n10666 35.2919
R35288 vss.n10666 vss.n10665 35.2919
R35289 vss.n10665 vss.n10647 35.2919
R35290 vss.n10647 vss.n10610 35.2919
R35291 vss.n12595 vss.n10610 35.2919
R35292 vss.n12595 vss.n12594 35.2919
R35293 vss.n10674 vss.n10673 35.2919
R35294 vss.n10675 vss.n10674 35.2919
R35295 vss.n10675 vss.n10627 35.2919
R35296 vss.n11607 vss.n10627 35.2919
R35297 vss.n11608 vss.n11607 35.2919
R35298 vss.n11609 vss.n11608 35.2919
R35299 vss.n10854 vss.n10853 35.2919
R35300 vss.n10853 vss.n10852 35.2919
R35301 vss.n10852 vss.n10620 35.2919
R35302 vss.n11618 vss.n10620 35.2919
R35303 vss.n11619 vss.n11618 35.2919
R35304 vss.n11620 vss.n11619 35.2919
R35305 vss.n10860 vss.n10822 35.2919
R35306 vss.n10866 vss.n10822 35.2919
R35307 vss.n10867 vss.n10866 35.2919
R35308 vss.n11534 vss.n10867 35.2919
R35309 vss.n11534 vss.n11533 35.2919
R35310 vss.n11533 vss.n11532 35.2919
R35311 vss.n11511 vss.n11510 35.2919
R35312 vss.n11512 vss.n11511 35.2919
R35313 vss.n11512 vss.n10876 35.2919
R35314 vss.n11516 vss.n10876 35.2919
R35315 vss.n11524 vss.n11516 35.2919
R35316 vss.n11524 vss.n11523 35.2919
R35317 vss.n11490 vss.n10891 35.2919
R35318 vss.n11490 vss.n11489 35.2919
R35319 vss.n11489 vss.n10892 35.2919
R35320 vss.n11485 vss.n10892 35.2919
R35321 vss.n11485 vss.n11484 35.2919
R35322 vss.n11484 vss.n11483 35.2919
R35323 vss.n11463 vss.n11462 35.2919
R35324 vss.n11464 vss.n11463 35.2919
R35325 vss.n11464 vss.n10902 35.2919
R35326 vss.n11468 vss.n10902 35.2919
R35327 vss.n11475 vss.n11468 35.2919
R35328 vss.n11475 vss.n11474 35.2919
R35329 vss.n10923 vss.n10920 35.2919
R35330 vss.n10923 vss.n10922 35.2919
R35331 vss.n10922 vss.n10334 35.2919
R35332 vss.n12750 vss.n10334 35.2919
R35333 vss.n12751 vss.n12750 35.2919
R35334 vss.n12752 vss.n12751 35.2919
R35335 vss.n12731 vss.n12730 35.2919
R35336 vss.n12732 vss.n12731 35.2919
R35337 vss.n12732 vss.n10327 35.2919
R35338 vss.n12761 vss.n10327 35.2919
R35339 vss.n12762 vss.n12761 35.2919
R35340 vss.n12763 vss.n12762 35.2919
R35341 vss.n12720 vss.n10361 35.2919
R35342 vss.n12720 vss.n12719 35.2919
R35343 vss.n12719 vss.n10362 35.2919
R35344 vss.n12715 vss.n10362 35.2919
R35345 vss.n12715 vss.n12714 35.2919
R35346 vss.n12714 vss.n12713 35.2919
R35347 vss.n12996 vss.n2251 35.2919
R35348 vss.n13002 vss.n2251 35.2919
R35349 vss.n13003 vss.n13002 35.2919
R35350 vss.n13013 vss.n13003 35.2919
R35351 vss.n13013 vss.n13012 35.2919
R35352 vss.n13012 vss.n13011 35.2919
R35353 vss.n2274 vss.n2261 35.2919
R35354 vss.n2295 vss.n2274 35.2919
R35355 vss.n2295 vss.n2294 35.2919
R35356 vss.n2294 vss.n2293 35.2919
R35357 vss.n2293 vss.n2277 35.2919
R35358 vss.n2283 vss.n2277 35.2919
R35359 vss.n2085 vss.n2075 35.2919
R35360 vss.n13104 vss.n2085 35.2919
R35361 vss.n13104 vss.n13103 35.2919
R35362 vss.n13103 vss.n13102 35.2919
R35363 vss.n13102 vss.n2088 35.2919
R35364 vss.n2094 vss.n2088 35.2919
R35365 vss.n1114 vss.n1105 35.2919
R35366 vss.n1120 vss.n1105 35.2919
R35367 vss.n1121 vss.n1120 35.2919
R35368 vss.n1131 vss.n1121 35.2919
R35369 vss.n1131 vss.n1130 35.2919
R35370 vss.n1130 vss.n1129 35.2919
R35371 vss.n871 vss.n870 35.2919
R35372 vss.n870 vss.n869 35.2919
R35373 vss.n869 vss.n838 35.2919
R35374 vss.n865 vss.n838 35.2919
R35375 vss.n865 vss.n864 35.2919
R35376 vss.n864 vss.n863 35.2919
R35377 vss.n14156 vss.n449 35.2919
R35378 vss.n14164 vss.n449 35.2919
R35379 vss.n14165 vss.n14164 35.2919
R35380 vss.n14167 vss.n14165 35.2919
R35381 vss.n14167 vss.n14166 35.2919
R35382 vss.n14166 vss.n436 35.2919
R35383 vss.n176 vss.n175 35.2919
R35384 vss.n180 vss.n176 35.2919
R35385 vss.n180 vss.n11 35.2919
R35386 vss.n14788 vss.n11 35.2919
R35387 vss.n14788 vss.n14787 35.2919
R35388 vss.n14787 vss.n14786 35.2919
R35389 vss.n337 vss.n327 35.2919
R35390 vss.n343 vss.n327 35.2919
R35391 vss.n344 vss.n343 35.2919
R35392 vss.n354 vss.n344 35.2919
R35393 vss.n354 vss.n353 35.2919
R35394 vss.n353 vss.n352 35.2919
R35395 vss.n14191 vss.n14179 35.2919
R35396 vss.n14212 vss.n14191 35.2919
R35397 vss.n14212 vss.n14211 35.2919
R35398 vss.n14211 vss.n14210 35.2919
R35399 vss.n14210 vss.n14194 35.2919
R35400 vss.n14200 vss.n14194 35.2919
R35401 vss.n14116 vss.n14106 35.2919
R35402 vss.n14122 vss.n14106 35.2919
R35403 vss.n14123 vss.n14122 35.2919
R35404 vss.n14133 vss.n14123 35.2919
R35405 vss.n14133 vss.n14132 35.2919
R35406 vss.n14132 vss.n14131 35.2919
R35407 vss.n14225 vss.n424 35.2919
R35408 vss.n14231 vss.n424 35.2919
R35409 vss.n14232 vss.n14231 35.2919
R35410 vss.n14242 vss.n14232 35.2919
R35411 vss.n14242 vss.n14241 35.2919
R35412 vss.n14241 vss.n14240 35.2919
R35413 vss.n14152 vss.n14151 35.2919
R35414 vss.n14151 vss.n14150 35.2919
R35415 vss.n14150 vss.n464 35.2919
R35416 vss.n13573 vss.n464 35.2919
R35417 vss.n13573 vss.n13569 35.2919
R35418 vss.n13569 vss.n13568 35.2919
R35419 vss.n13560 vss.n13547 35.2919
R35420 vss.n13600 vss.n13560 35.2919
R35421 vss.n13600 vss.n13599 35.2919
R35422 vss.n13599 vss.n13598 35.2919
R35423 vss.n13598 vss.n13563 35.2919
R35424 vss.n13589 vss.n13563 35.2919
R35425 vss.n14654 vss.n196 35.2919
R35426 vss.n14675 vss.n14654 35.2919
R35427 vss.n14675 vss.n14674 35.2919
R35428 vss.n14674 vss.n14673 35.2919
R35429 vss.n14673 vss.n14657 35.2919
R35430 vss.n14663 vss.n14657 35.2919
R35431 vss.n14539 vss.n242 35.2919
R35432 vss.n14545 vss.n242 35.2919
R35433 vss.n14546 vss.n14545 35.2919
R35434 vss.n14556 vss.n14546 35.2919
R35435 vss.n14556 vss.n14555 35.2919
R35436 vss.n14555 vss.n14554 35.2919
R35437 vss.n14459 vss.n255 35.2919
R35438 vss.n14480 vss.n14459 35.2919
R35439 vss.n14480 vss.n14479 35.2919
R35440 vss.n14479 vss.n14478 35.2919
R35441 vss.n14478 vss.n14462 35.2919
R35442 vss.n14468 vss.n14462 35.2919
R35443 vss.n14344 vss.n301 35.2919
R35444 vss.n14350 vss.n301 35.2919
R35445 vss.n14351 vss.n14350 35.2919
R35446 vss.n14361 vss.n14351 35.2919
R35447 vss.n14361 vss.n14360 35.2919
R35448 vss.n14360 vss.n14359 35.2919
R35449 vss.n14264 vss.n314 35.2919
R35450 vss.n14285 vss.n14264 35.2919
R35451 vss.n14285 vss.n14284 35.2919
R35452 vss.n14284 vss.n14283 35.2919
R35453 vss.n14283 vss.n14267 35.2919
R35454 vss.n14273 vss.n14267 35.2919
R35455 vss.n14310 vss.n14298 35.2919
R35456 vss.n14331 vss.n14310 35.2919
R35457 vss.n14331 vss.n14330 35.2919
R35458 vss.n14330 vss.n14329 35.2919
R35459 vss.n14329 vss.n14313 35.2919
R35460 vss.n14319 vss.n14313 35.2919
R35461 vss.n14390 vss.n14380 35.2919
R35462 vss.n14396 vss.n14380 35.2919
R35463 vss.n14397 vss.n14396 35.2919
R35464 vss.n14407 vss.n14397 35.2919
R35465 vss.n14407 vss.n14406 35.2919
R35466 vss.n14406 vss.n14405 35.2919
R35467 vss.n14505 vss.n14493 35.2919
R35468 vss.n14526 vss.n14505 35.2919
R35469 vss.n14526 vss.n14525 35.2919
R35470 vss.n14525 vss.n14524 35.2919
R35471 vss.n14524 vss.n14508 35.2919
R35472 vss.n14514 vss.n14508 35.2919
R35473 vss.n14585 vss.n14575 35.2919
R35474 vss.n14591 vss.n14575 35.2919
R35475 vss.n14592 vss.n14591 35.2919
R35476 vss.n14602 vss.n14592 35.2919
R35477 vss.n14602 vss.n14601 35.2919
R35478 vss.n14601 vss.n14600 35.2919
R35479 vss.n14700 vss.n14688 35.2919
R35480 vss.n14721 vss.n14700 35.2919
R35481 vss.n14721 vss.n14720 35.2919
R35482 vss.n14720 vss.n14719 35.2919
R35483 vss.n14719 vss.n14703 35.2919
R35484 vss.n14709 vss.n14703 35.2919
R35485 vss.n14734 vss.n165 35.2919
R35486 vss.n14740 vss.n165 35.2919
R35487 vss.n14741 vss.n14740 35.2919
R35488 vss.n14751 vss.n14741 35.2919
R35489 vss.n14751 vss.n14750 35.2919
R35490 vss.n14750 vss.n14749 35.2919
R35491 vss.n13918 vss.n13917 35.2919
R35492 vss.n13917 vss.n13916 35.2919
R35493 vss.n13916 vss.n13308 35.2919
R35494 vss.n13903 vss.n13308 35.2919
R35495 vss.n13904 vss.n13903 35.2919
R35496 vss.n13906 vss.n13904 35.2919
R35497 vss.n13874 vss.n13334 35.2919
R35498 vss.n13882 vss.n13334 35.2919
R35499 vss.n13883 vss.n13882 35.2919
R35500 vss.n13885 vss.n13883 35.2919
R35501 vss.n13885 vss.n13884 35.2919
R35502 vss.n13884 vss.n13328 35.2919
R35503 vss.n13870 vss.n13869 35.2919
R35504 vss.n13869 vss.n13868 35.2919
R35505 vss.n13868 vss.n13350 35.2919
R35506 vss.n13848 vss.n13350 35.2919
R35507 vss.n13849 vss.n13848 35.2919
R35508 vss.n13851 vss.n13849 35.2919
R35509 vss.n13820 vss.n13375 35.2919
R35510 vss.n13828 vss.n13375 35.2919
R35511 vss.n13829 vss.n13828 35.2919
R35512 vss.n13831 vss.n13829 35.2919
R35513 vss.n13831 vss.n13830 35.2919
R35514 vss.n13830 vss.n13367 35.2919
R35515 vss.n13816 vss.n13815 35.2919
R35516 vss.n13815 vss.n13814 35.2919
R35517 vss.n13814 vss.n13391 35.2919
R35518 vss.n13798 vss.n13391 35.2919
R35519 vss.n13799 vss.n13798 35.2919
R35520 vss.n13801 vss.n13799 35.2919
R35521 vss.n13769 vss.n13414 35.2919
R35522 vss.n13777 vss.n13414 35.2919
R35523 vss.n13778 vss.n13777 35.2919
R35524 vss.n13780 vss.n13778 35.2919
R35525 vss.n13780 vss.n13779 35.2919
R35526 vss.n13779 vss.n13408 35.2919
R35527 vss.n13765 vss.n13764 35.2919
R35528 vss.n13764 vss.n13763 35.2919
R35529 vss.n13763 vss.n13430 35.2919
R35530 vss.n13743 vss.n13430 35.2919
R35531 vss.n13744 vss.n13743 35.2919
R35532 vss.n13746 vss.n13744 35.2919
R35533 vss.n13715 vss.n13455 35.2919
R35534 vss.n13723 vss.n13455 35.2919
R35535 vss.n13724 vss.n13723 35.2919
R35536 vss.n13726 vss.n13724 35.2919
R35537 vss.n13726 vss.n13725 35.2919
R35538 vss.n13725 vss.n13447 35.2919
R35539 vss.n13711 vss.n13710 35.2919
R35540 vss.n13710 vss.n13709 35.2919
R35541 vss.n13709 vss.n13471 35.2919
R35542 vss.n13693 vss.n13471 35.2919
R35543 vss.n13694 vss.n13693 35.2919
R35544 vss.n13696 vss.n13694 35.2919
R35545 vss.n13664 vss.n13494 35.2919
R35546 vss.n13672 vss.n13494 35.2919
R35547 vss.n13673 vss.n13672 35.2919
R35548 vss.n13675 vss.n13673 35.2919
R35549 vss.n13675 vss.n13674 35.2919
R35550 vss.n13674 vss.n13488 35.2919
R35551 vss.n13660 vss.n13659 35.2919
R35552 vss.n13659 vss.n13658 35.2919
R35553 vss.n13658 vss.n13510 35.2919
R35554 vss.n13638 vss.n13510 35.2919
R35555 vss.n13639 vss.n13638 35.2919
R35556 vss.n13641 vss.n13639 35.2919
R35557 vss.n13610 vss.n13535 35.2919
R35558 vss.n13618 vss.n13535 35.2919
R35559 vss.n13619 vss.n13618 35.2919
R35560 vss.n13621 vss.n13619 35.2919
R35561 vss.n13621 vss.n13620 35.2919
R35562 vss.n13620 vss.n13527 35.2919
R35563 vss.n636 vss.n635 35.2919
R35564 vss.n637 vss.n636 35.2919
R35565 vss.n637 vss.n618 35.2919
R35566 vss.n653 vss.n618 35.2919
R35567 vss.n654 vss.n653 35.2919
R35568 vss.n655 vss.n654 35.2919
R35569 vss.n13213 vss.n804 35.2919
R35570 vss.n13219 vss.n804 35.2919
R35571 vss.n13220 vss.n13219 35.2919
R35572 vss.n13230 vss.n13220 35.2919
R35573 vss.n13230 vss.n13229 35.2919
R35574 vss.n13229 vss.n13228 35.2919
R35575 vss.n1672 vss.n1663 35.2919
R35576 vss.n1678 vss.n1663 35.2919
R35577 vss.n1679 vss.n1678 35.2919
R35578 vss.n1689 vss.n1679 35.2919
R35579 vss.n1689 vss.n1688 35.2919
R35580 vss.n1688 vss.n1687 35.2919
R35581 vss.n1625 vss.n1616 35.2919
R35582 vss.n1631 vss.n1616 35.2919
R35583 vss.n1632 vss.n1631 35.2919
R35584 vss.n1642 vss.n1632 35.2919
R35585 vss.n1642 vss.n1641 35.2919
R35586 vss.n1641 vss.n1640 35.2919
R35587 vss.n1377 vss.n1368 35.2919
R35588 vss.n1383 vss.n1368 35.2919
R35589 vss.n1384 vss.n1383 35.2919
R35590 vss.n1394 vss.n1384 35.2919
R35591 vss.n1394 vss.n1393 35.2919
R35592 vss.n1393 vss.n1392 35.2919
R35593 vss.n1178 vss.n1169 35.2919
R35594 vss.n1184 vss.n1169 35.2919
R35595 vss.n1185 vss.n1184 35.2919
R35596 vss.n1195 vss.n1185 35.2919
R35597 vss.n1195 vss.n1194 35.2919
R35598 vss.n1194 vss.n1193 35.2919
R35599 vss.n1330 vss.n1321 35.2919
R35600 vss.n1336 vss.n1321 35.2919
R35601 vss.n1337 vss.n1336 35.2919
R35602 vss.n1347 vss.n1337 35.2919
R35603 vss.n1347 vss.n1346 35.2919
R35604 vss.n1346 vss.n1345 35.2919
R35605 vss.n1069 vss.n1060 35.2919
R35606 vss.n1075 vss.n1060 35.2919
R35607 vss.n1076 vss.n1075 35.2919
R35608 vss.n1086 vss.n1076 35.2919
R35609 vss.n1086 vss.n1085 35.2919
R35610 vss.n1085 vss.n1084 35.2919
R35611 vss.n1462 vss.n1453 35.2919
R35612 vss.n1468 vss.n1453 35.2919
R35613 vss.n1469 vss.n1468 35.2919
R35614 vss.n1479 vss.n1469 35.2919
R35615 vss.n1479 vss.n1478 35.2919
R35616 vss.n1478 vss.n1477 35.2919
R35617 vss.n1542 vss.n1533 35.2919
R35618 vss.n1548 vss.n1533 35.2919
R35619 vss.n1549 vss.n1548 35.2919
R35620 vss.n1560 vss.n1549 35.2919
R35621 vss.n1560 vss.n1559 35.2919
R35622 vss.n1559 vss.n1558 35.2919
R35623 vss.n830 vss.n829 35.2919
R35624 vss.n829 vss.n828 35.2919
R35625 vss.n828 vss.n605 35.2919
R35626 vss.n13948 vss.n605 35.2919
R35627 vss.n13948 vss.n13947 35.2919
R35628 vss.n13947 vss.n13946 35.2919
R35629 vss.n915 vss.n914 35.2919
R35630 vss.n914 vss.n913 35.2919
R35631 vss.n913 vss.n879 35.2919
R35632 vss.n909 vss.n879 35.2919
R35633 vss.n909 vss.n908 35.2919
R35634 vss.n908 vss.n907 35.2919
R35635 vss.n14004 vss.n526 35.2919
R35636 vss.n14010 vss.n526 35.2919
R35637 vss.n14011 vss.n14010 35.2919
R35638 vss.n14012 vss.n14011 35.2919
R35639 vss.n14013 vss.n14012 35.2919
R35640 vss.n14017 vss.n14013 35.2919
R35641 vss.n13998 vss.n13997 35.2919
R35642 vss.n13997 vss.n13996 35.2919
R35643 vss.n13996 vss.n541 35.2919
R35644 vss.n673 vss.n541 35.2919
R35645 vss.n674 vss.n673 35.2919
R35646 vss.n675 vss.n674 35.2919
R35647 vss.n13969 vss.n565 35.2919
R35648 vss.n13975 vss.n565 35.2919
R35649 vss.n13976 vss.n13975 35.2919
R35650 vss.n13977 vss.n13976 35.2919
R35651 vss.n13978 vss.n13977 35.2919
R35652 vss.n13982 vss.n13978 35.2919
R35653 vss.n13963 vss.n13962 35.2919
R35654 vss.n13962 vss.n13961 35.2919
R35655 vss.n13961 vss.n580 35.2919
R35656 vss.n772 vss.n580 35.2919
R35657 vss.n773 vss.n772 35.2919
R35658 vss.n774 vss.n773 35.2919
R35659 vss.n13246 vss.n13245 35.2919
R35660 vss.n13245 vss.n13244 35.2919
R35661 vss.n13244 vss.n747 35.2919
R35662 vss.n781 vss.n747 35.2919
R35663 vss.n782 vss.n781 35.2919
R35664 vss.n786 vss.n782 35.2919
R35665 vss.n1733 vss.n1732 35.2919
R35666 vss.n1734 vss.n1733 35.2919
R35667 vss.n1734 vss.n1711 35.2919
R35668 vss.n1743 vss.n1711 35.2919
R35669 vss.n1744 vss.n1743 35.2919
R35670 vss.n1745 vss.n1744 35.2919
R35671 vss.n1781 vss.n1752 35.2919
R35672 vss.n1787 vss.n1752 35.2919
R35673 vss.n1788 vss.n1787 35.2919
R35674 vss.n1789 vss.n1788 35.2919
R35675 vss.n1790 vss.n1789 35.2919
R35676 vss.n1794 vss.n1790 35.2919
R35677 vss.n1775 vss.n1774 35.2919
R35678 vss.n1774 vss.n1773 35.2919
R35679 vss.n1773 vss.n1268 35.2919
R35680 vss.n1814 vss.n1268 35.2919
R35681 vss.n1815 vss.n1814 35.2919
R35682 vss.n1816 vss.n1815 35.2919
R35683 vss.n1256 vss.n1255 35.2919
R35684 vss.n1257 vss.n1256 35.2919
R35685 vss.n1258 vss.n1257 35.2919
R35686 vss.n1259 vss.n1258 35.2919
R35687 vss.n1260 vss.n1259 35.2919
R35688 vss.n1261 vss.n1260 35.2919
R35689 vss.n1837 vss.n1836 35.2919
R35690 vss.n1838 vss.n1837 35.2919
R35691 vss.n1838 vss.n1215 35.2919
R35692 vss.n1847 vss.n1215 35.2919
R35693 vss.n1848 vss.n1847 35.2919
R35694 vss.n1849 vss.n1848 35.2919
R35695 vss.n1885 vss.n1856 35.2919
R35696 vss.n1891 vss.n1856 35.2919
R35697 vss.n1892 vss.n1891 35.2919
R35698 vss.n1893 vss.n1892 35.2919
R35699 vss.n1894 vss.n1893 35.2919
R35700 vss.n1898 vss.n1894 35.2919
R35701 vss.n1879 vss.n1878 35.2919
R35702 vss.n1878 vss.n1877 35.2919
R35703 vss.n1877 vss.n1150 35.2919
R35704 vss.n1918 vss.n1150 35.2919
R35705 vss.n1919 vss.n1918 35.2919
R35706 vss.n1920 vss.n1919 35.2919
R35707 vss.n1956 vss.n1927 35.2919
R35708 vss.n1962 vss.n1927 35.2919
R35709 vss.n1963 vss.n1962 35.2919
R35710 vss.n1964 vss.n1963 35.2919
R35711 vss.n1965 vss.n1964 35.2919
R35712 vss.n1969 vss.n1965 35.2919
R35713 vss.n1950 vss.n1949 35.2919
R35714 vss.n1949 vss.n1948 35.2919
R35715 vss.n1948 vss.n694 35.2919
R35716 vss.n13296 vss.n694 35.2919
R35717 vss.n13297 vss.n13296 35.2919
R35718 vss.n13298 vss.n13297 35.2919
R35719 vss.n13268 vss.n718 35.2919
R35720 vss.n13274 vss.n718 35.2919
R35721 vss.n13275 vss.n13274 35.2919
R35722 vss.n13276 vss.n13275 35.2919
R35723 vss.n13277 vss.n13276 35.2919
R35724 vss.n13281 vss.n13277 35.2919
R35725 vss.n2004 vss.n1995 35.2919
R35726 vss.n2010 vss.n1995 35.2919
R35727 vss.n2011 vss.n2010 35.2919
R35728 vss.n2021 vss.n2011 35.2919
R35729 vss.n2021 vss.n2020 35.2919
R35730 vss.n2020 vss.n2019 35.2919
R35731 vss.n13178 vss.n13167 35.2919
R35732 vss.n13184 vss.n13167 35.2919
R35733 vss.n13185 vss.n13184 35.2919
R35734 vss.n13186 vss.n13185 35.2919
R35735 vss.n13193 vss.n13186 35.2919
R35736 vss.n13193 vss.n13192 35.2919
R35737 vss.n9606 vss.n9596 35.2919
R35738 vss.n9612 vss.n9596 35.2919
R35739 vss.n9613 vss.n9612 35.2919
R35740 vss.n9623 vss.n9613 35.2919
R35741 vss.n9623 vss.n9622 35.2919
R35742 vss.n9622 vss.n9621 35.2919
R35743 vss.n9170 vss.n9160 35.2919
R35744 vss.n9176 vss.n9160 35.2919
R35745 vss.n9177 vss.n9176 35.2919
R35746 vss.n9187 vss.n9177 35.2919
R35747 vss.n9187 vss.n9186 35.2919
R35748 vss.n9186 vss.n9185 35.2919
R35749 vss.n9468 vss.n9467 35.2919
R35750 vss.n9469 vss.n9468 35.2919
R35751 vss.n9469 vss.n9449 35.2919
R35752 vss.n9481 vss.n9449 35.2919
R35753 vss.n9482 vss.n9481 35.2919
R35754 vss.n9483 vss.n9482 35.2919
R35755 vss.n8049 vss.n8048 35.2919
R35756 vss.n8048 vss.n8047 35.2919
R35757 vss.n8047 vss.n8017 35.2919
R35758 vss.n8031 vss.n8017 35.2919
R35759 vss.n8032 vss.n8031 35.2919
R35760 vss.n8033 vss.n8032 35.2919
R35761 vss.n5986 vss.n5976 35.2919
R35762 vss.n9660 vss.n5986 35.2919
R35763 vss.n9660 vss.n9659 35.2919
R35764 vss.n9659 vss.n9658 35.2919
R35765 vss.n9658 vss.n5989 35.2919
R35766 vss.n5995 vss.n5989 35.2919
R35767 vss.n8148 vss.n8147 35.2919
R35768 vss.n8147 vss.n8146 35.2919
R35769 vss.n8146 vss.n8125 35.2919
R35770 vss.n8128 vss.n8125 35.2919
R35771 vss.n8135 vss.n8128 35.2919
R35772 vss.n8137 vss.n8135 35.2919
R35773 vss.n8154 vss.n8114 35.2919
R35774 vss.n8162 vss.n8114 35.2919
R35775 vss.n8163 vss.n8162 35.2919
R35776 vss.n8165 vss.n8163 35.2919
R35777 vss.n8165 vss.n8164 35.2919
R35778 vss.n8164 vss.n8102 35.2919
R35779 vss.n8080 vss.n8070 35.2919
R35780 vss.n8088 vss.n8070 35.2919
R35781 vss.n8089 vss.n8088 35.2919
R35782 vss.n8091 vss.n8089 35.2919
R35783 vss.n8091 vss.n8090 35.2919
R35784 vss.n8090 vss.n8055 35.2919
R35785 vss.n8223 vss.n8002 35.2919
R35786 vss.n8229 vss.n8002 35.2919
R35787 vss.n8230 vss.n8229 35.2919
R35788 vss.n8240 vss.n8230 35.2919
R35789 vss.n8240 vss.n8239 35.2919
R35790 vss.n8239 vss.n8238 35.2919
R35791 vss.n8189 vss.n8177 35.2919
R35792 vss.n8210 vss.n8189 35.2919
R35793 vss.n8210 vss.n8209 35.2919
R35794 vss.n8209 vss.n8208 35.2919
R35795 vss.n8208 vss.n8192 35.2919
R35796 vss.n8198 vss.n8192 35.2919
R35797 vss.n7312 vss.n7302 35.2919
R35798 vss.n8998 vss.n7312 35.2919
R35799 vss.n8998 vss.n8997 35.2919
R35800 vss.n8997 vss.n8996 35.2919
R35801 vss.n8996 vss.n7315 35.2919
R35802 vss.n7321 vss.n7315 35.2919
R35803 vss.n8714 vss.n7859 35.2919
R35804 vss.n8720 vss.n7859 35.2919
R35805 vss.n8721 vss.n8720 35.2919
R35806 vss.n8731 vss.n8721 35.2919
R35807 vss.n8731 vss.n8730 35.2919
R35808 vss.n8730 vss.n8729 35.2919
R35809 vss.n7788 vss.n7778 35.2919
R35810 vss.n7794 vss.n7778 35.2919
R35811 vss.n7795 vss.n7794 35.2919
R35812 vss.n7805 vss.n7795 35.2919
R35813 vss.n7805 vss.n7804 35.2919
R35814 vss.n7804 vss.n7803 35.2919
R35815 vss.n8753 vss.n7685 35.2919
R35816 vss.n8774 vss.n8753 35.2919
R35817 vss.n8774 vss.n8773 35.2919
R35818 vss.n8773 vss.n8772 35.2919
R35819 vss.n8772 vss.n8756 35.2919
R35820 vss.n8762 vss.n8756 35.2919
R35821 vss.n8833 vss.n7672 35.2919
R35822 vss.n8839 vss.n7672 35.2919
R35823 vss.n8840 vss.n8839 35.2919
R35824 vss.n8850 vss.n8840 35.2919
R35825 vss.n8850 vss.n8849 35.2919
R35826 vss.n8849 vss.n8848 35.2919
R35827 vss.n8799 vss.n8787 35.2919
R35828 vss.n8820 vss.n8799 35.2919
R35829 vss.n8820 vss.n8819 35.2919
R35830 vss.n8819 vss.n8818 35.2919
R35831 vss.n8818 vss.n8802 35.2919
R35832 vss.n8808 vss.n8802 35.2919
R35833 vss.n8872 vss.n7542 35.2919
R35834 vss.n8893 vss.n8872 35.2919
R35835 vss.n8893 vss.n8892 35.2919
R35836 vss.n8892 vss.n8891 35.2919
R35837 vss.n8891 vss.n8875 35.2919
R35838 vss.n8881 vss.n8875 35.2919
R35839 vss.n7280 vss.n7270 35.2919
R35840 vss.n9029 vss.n7280 35.2919
R35841 vss.n9029 vss.n9028 35.2919
R35842 vss.n9028 vss.n9027 35.2919
R35843 vss.n9027 vss.n7283 35.2919
R35844 vss.n7289 vss.n7283 35.2919
R35845 vss.n8268 vss.n7902 35.2919
R35846 vss.n8274 vss.n8268 35.2919
R35847 vss.n8274 vss.n8273 35.2919
R35848 vss.n8273 vss.n8272 35.2919
R35849 vss.n8272 vss.n7293 35.2919
R35850 vss.n7296 vss.n7293 35.2919
R35851 vss.n8284 vss.n7892 35.2919
R35852 vss.n8292 vss.n7892 35.2919
R35853 vss.n8293 vss.n8292 35.2919
R35854 vss.n8295 vss.n8293 35.2919
R35855 vss.n8295 vss.n8294 35.2919
R35856 vss.n8294 vss.n7880 35.2919
R35857 vss.n8690 vss.n8311 35.2919
R35858 vss.n8698 vss.n8311 35.2919
R35859 vss.n8699 vss.n8698 35.2919
R35860 vss.n8701 vss.n8699 35.2919
R35861 vss.n8701 vss.n8700 35.2919
R35862 vss.n8700 vss.n7869 35.2919
R35863 vss.n8323 vss.n8321 35.2919
R35864 vss.n8340 vss.n8321 35.2919
R35865 vss.n8341 vss.n8340 35.2919
R35866 vss.n8678 vss.n8341 35.2919
R35867 vss.n8678 vss.n8677 35.2919
R35868 vss.n8677 vss.n8676 35.2919
R35869 vss.n8652 vss.n8651 35.2919
R35870 vss.n8657 vss.n8652 35.2919
R35871 vss.n8657 vss.n8656 35.2919
R35872 vss.n8656 vss.n8655 35.2919
R35873 vss.n8655 vss.n8351 35.2919
R35874 vss.n8664 vss.n8351 35.2919
R35875 vss.n8368 vss.n8366 35.2919
R35876 vss.n8390 vss.n8366 35.2919
R35877 vss.n8391 vss.n8390 35.2919
R35878 vss.n8635 vss.n8391 35.2919
R35879 vss.n8635 vss.n8634 35.2919
R35880 vss.n8634 vss.n8633 35.2919
R35881 vss.n8608 vss.n8607 35.2919
R35882 vss.n8613 vss.n8608 35.2919
R35883 vss.n8613 vss.n8612 35.2919
R35884 vss.n8612 vss.n8611 35.2919
R35885 vss.n8611 vss.n8401 35.2919
R35886 vss.n8620 vss.n8401 35.2919
R35887 vss.n8421 vss.n8419 35.2919
R35888 vss.n8438 vss.n8419 35.2919
R35889 vss.n8439 vss.n8438 35.2919
R35890 vss.n8591 vss.n8439 35.2919
R35891 vss.n8591 vss.n8590 35.2919
R35892 vss.n8590 vss.n8589 35.2919
R35893 vss.n8565 vss.n8564 35.2919
R35894 vss.n8570 vss.n8565 35.2919
R35895 vss.n8570 vss.n8569 35.2919
R35896 vss.n8569 vss.n8568 35.2919
R35897 vss.n8568 vss.n8449 35.2919
R35898 vss.n8577 vss.n8449 35.2919
R35899 vss.n8466 vss.n8464 35.2919
R35900 vss.n8488 vss.n8464 35.2919
R35901 vss.n8489 vss.n8488 35.2919
R35902 vss.n8548 vss.n8489 35.2919
R35903 vss.n8548 vss.n8547 35.2919
R35904 vss.n8547 vss.n8546 35.2919
R35905 vss.n8522 vss.n8521 35.2919
R35906 vss.n8521 vss.n8520 35.2919
R35907 vss.n8520 vss.n8515 35.2919
R35908 vss.n8516 vss.n8515 35.2919
R35909 vss.n8516 vss.n8499 35.2919
R35910 vss.n8533 vss.n8499 35.2919
R35911 vss.n8952 vss.n7483 35.2919
R35912 vss.n8958 vss.n7483 35.2919
R35913 vss.n8959 vss.n8958 35.2919
R35914 vss.n8969 vss.n8959 35.2919
R35915 vss.n8969 vss.n8968 35.2919
R35916 vss.n8968 vss.n8967 35.2919
R35917 vss.n8918 vss.n8906 35.2919
R35918 vss.n8939 vss.n8918 35.2919
R35919 vss.n8939 vss.n8938 35.2919
R35920 vss.n8938 vss.n8937 35.2919
R35921 vss.n8937 vss.n8921 35.2919
R35922 vss.n8927 vss.n8921 35.2919
R35923 vss.n7506 vss.n7493 35.2919
R35924 vss.n7527 vss.n7506 35.2919
R35925 vss.n7527 vss.n7526 35.2919
R35926 vss.n7526 vss.n7525 35.2919
R35927 vss.n7525 vss.n7509 35.2919
R35928 vss.n7515 vss.n7509 35.2919
R35929 vss.n7565 vss.n7555 35.2919
R35930 vss.n7571 vss.n7555 35.2919
R35931 vss.n7572 vss.n7571 35.2919
R35932 vss.n7582 vss.n7572 35.2919
R35933 vss.n7582 vss.n7581 35.2919
R35934 vss.n7581 vss.n7580 35.2919
R35935 vss.n7708 vss.n7698 35.2919
R35936 vss.n7714 vss.n7698 35.2919
R35937 vss.n7715 vss.n7714 35.2919
R35938 vss.n7725 vss.n7715 35.2919
R35939 vss.n7725 vss.n7724 35.2919
R35940 vss.n7724 vss.n7723 35.2919
R35941 vss.n7929 vss.n7919 35.2919
R35942 vss.n7935 vss.n7919 35.2919
R35943 vss.n7936 vss.n7935 35.2919
R35944 vss.n7946 vss.n7936 35.2919
R35945 vss.n7946 vss.n7945 35.2919
R35946 vss.n7945 vss.n7944 35.2919
R35947 vss.n6028 vss.n6018 35.2919
R35948 vss.n6034 vss.n6018 35.2919
R35949 vss.n6035 vss.n6034 35.2919
R35950 vss.n6046 vss.n6035 35.2919
R35951 vss.n6046 vss.n6045 35.2919
R35952 vss.n6045 vss.n6044 35.2919
R35953 vss.n7198 vss.n7188 35.2919
R35954 vss.n7204 vss.n7188 35.2919
R35955 vss.n7205 vss.n7204 35.2919
R35956 vss.n7215 vss.n7205 35.2919
R35957 vss.n7215 vss.n7214 35.2919
R35958 vss.n7214 vss.n7213 35.2919
R35959 vss.n6693 vss.n6683 35.2919
R35960 vss.n6699 vss.n6683 35.2919
R35961 vss.n6700 vss.n6699 35.2919
R35962 vss.n6710 vss.n6700 35.2919
R35963 vss.n6710 vss.n6709 35.2919
R35964 vss.n6709 vss.n6708 35.2919
R35965 vss.n6649 vss.n6639 35.2919
R35966 vss.n6655 vss.n6639 35.2919
R35967 vss.n6656 vss.n6655 35.2919
R35968 vss.n6666 vss.n6656 35.2919
R35969 vss.n6666 vss.n6665 35.2919
R35970 vss.n6665 vss.n6664 35.2919
R35971 vss.n7007 vss.n6997 35.2919
R35972 vss.n7013 vss.n6997 35.2919
R35973 vss.n7014 vss.n7013 35.2919
R35974 vss.n7024 vss.n7014 35.2919
R35975 vss.n7024 vss.n7023 35.2919
R35976 vss.n7023 vss.n7022 35.2919
R35977 vss.n6467 vss.n6457 35.2919
R35978 vss.n6473 vss.n6457 35.2919
R35979 vss.n6474 vss.n6473 35.2919
R35980 vss.n6484 vss.n6474 35.2919
R35981 vss.n6484 vss.n6483 35.2919
R35982 vss.n6483 vss.n6482 35.2919
R35983 vss.n6422 vss.n6412 35.2919
R35984 vss.n6428 vss.n6412 35.2919
R35985 vss.n6429 vss.n6428 35.2919
R35986 vss.n6439 vss.n6429 35.2919
R35987 vss.n6439 vss.n6438 35.2919
R35988 vss.n6438 vss.n6437 35.2919
R35989 vss.n6344 vss.n6334 35.2919
R35990 vss.n6350 vss.n6334 35.2919
R35991 vss.n6351 vss.n6350 35.2919
R35992 vss.n6361 vss.n6351 35.2919
R35993 vss.n6361 vss.n6360 35.2919
R35994 vss.n6360 vss.n6359 35.2919
R35995 vss.n6958 vss.n6948 35.2919
R35996 vss.n6964 vss.n6948 35.2919
R35997 vss.n6965 vss.n6964 35.2919
R35998 vss.n6975 vss.n6965 35.2919
R35999 vss.n6975 vss.n6974 35.2919
R36000 vss.n6974 vss.n6973 35.2919
R36001 vss.n7147 vss.n7137 35.2919
R36002 vss.n7153 vss.n7137 35.2919
R36003 vss.n7154 vss.n7153 35.2919
R36004 vss.n7164 vss.n7154 35.2919
R36005 vss.n7164 vss.n7163 35.2919
R36006 vss.n7163 vss.n7162 35.2919
R36007 vss.n6155 vss.n6145 35.2919
R36008 vss.n6161 vss.n6145 35.2919
R36009 vss.n6162 vss.n6161 35.2919
R36010 vss.n9497 vss.n6162 35.2919
R36011 vss.n9497 vss.n9496 35.2919
R36012 vss.n9496 vss.n9495 35.2919
R36013 vss.n9423 vss.n9422 35.2919
R36014 vss.n9424 vss.n9423 35.2919
R36015 vss.n9424 vss.n9404 35.2919
R36016 vss.n9439 vss.n9404 35.2919
R36017 vss.n9440 vss.n9439 35.2919
R36018 vss.n9441 vss.n9440 35.2919
R36019 vss.n9553 vss.n6066 35.2919
R36020 vss.n9559 vss.n6066 35.2919
R36021 vss.n9560 vss.n9559 35.2919
R36022 vss.n9561 vss.n9560 35.2919
R36023 vss.n9562 vss.n9561 35.2919
R36024 vss.n9566 vss.n9562 35.2919
R36025 vss.n9547 vss.n9546 35.2919
R36026 vss.n9546 vss.n9545 35.2919
R36027 vss.n9545 vss.n6081 35.2919
R36028 vss.n7261 vss.n6081 35.2919
R36029 vss.n7262 vss.n7261 35.2919
R36030 vss.n7263 vss.n7262 35.2919
R36031 vss.n9518 vss.n6105 35.2919
R36032 vss.n9524 vss.n6105 35.2919
R36033 vss.n9525 vss.n9524 35.2919
R36034 vss.n9526 vss.n9525 35.2919
R36035 vss.n9527 vss.n9526 35.2919
R36036 vss.n9531 vss.n9527 35.2919
R36037 vss.n9512 vss.n9511 35.2919
R36038 vss.n9511 vss.n9510 35.2919
R36039 vss.n9510 vss.n6120 35.2919
R36040 vss.n7242 vss.n6120 35.2919
R36041 vss.n7243 vss.n7242 35.2919
R36042 vss.n7244 vss.n7243 35.2919
R36043 vss.n6757 vss.n6756 35.2919
R36044 vss.n6758 vss.n6757 35.2919
R36045 vss.n6758 vss.n6585 35.2919
R36046 vss.n7230 vss.n6585 35.2919
R36047 vss.n7231 vss.n7230 35.2919
R36048 vss.n7232 vss.n7231 35.2919
R36049 vss.n6769 vss.n6768 35.2919
R36050 vss.n6770 vss.n6769 35.2919
R36051 vss.n6770 vss.n6731 35.2919
R36052 vss.n6779 vss.n6731 35.2919
R36053 vss.n6780 vss.n6779 35.2919
R36054 vss.n6781 vss.n6780 35.2919
R36055 vss.n7063 vss.n6788 35.2919
R36056 vss.n7069 vss.n6788 35.2919
R36057 vss.n7070 vss.n7069 35.2919
R36058 vss.n7071 vss.n7070 35.2919
R36059 vss.n7072 vss.n7071 35.2919
R36060 vss.n7076 vss.n7072 35.2919
R36061 vss.n7057 vss.n7056 35.2919
R36062 vss.n7056 vss.n7055 35.2919
R36063 vss.n7055 vss.n6802 35.2919
R36064 vss.n6821 vss.n6802 35.2919
R36065 vss.n6822 vss.n6821 35.2919
R36066 vss.n6823 vss.n6822 35.2919
R36067 vss.n6898 vss.n6897 35.2919
R36068 vss.n6899 vss.n6898 35.2919
R36069 vss.n6899 vss.n6831 35.2919
R36070 vss.n7039 vss.n6831 35.2919
R36071 vss.n7040 vss.n7039 35.2919
R36072 vss.n7041 vss.n7040 35.2919
R36073 vss.n6889 vss.n6888 35.2919
R36074 vss.n6888 vss.n6887 35.2919
R36075 vss.n6887 vss.n6853 35.2919
R36076 vss.n6872 vss.n6853 35.2919
R36077 vss.n6873 vss.n6872 35.2919
R36078 vss.n6874 vss.n6873 35.2919
R36079 vss.n9226 vss.n6499 35.2919
R36080 vss.n9232 vss.n6499 35.2919
R36081 vss.n9233 vss.n9232 35.2919
R36082 vss.n9234 vss.n9233 35.2919
R36083 vss.n9235 vss.n9234 35.2919
R36084 vss.n9239 vss.n9235 35.2919
R36085 vss.n9220 vss.n9219 35.2919
R36086 vss.n9219 vss.n9218 35.2919
R36087 vss.n9218 vss.n6513 35.2919
R36088 vss.n6562 vss.n6513 35.2919
R36089 vss.n6563 vss.n6562 35.2919
R36090 vss.n6564 vss.n6563 35.2919
R36091 vss.n9075 vss.n9074 35.2919
R36092 vss.n9076 vss.n9075 35.2919
R36093 vss.n9076 vss.n6532 35.2919
R36094 vss.n9202 vss.n6532 35.2919
R36095 vss.n9203 vss.n9202 35.2919
R36096 vss.n9204 vss.n9203 35.2919
R36097 vss.n9084 vss.n9055 35.2919
R36098 vss.n9090 vss.n9055 35.2919
R36099 vss.n9091 vss.n9090 35.2919
R36100 vss.n9092 vss.n9091 35.2919
R36101 vss.n9093 vss.n9092 35.2919
R36102 vss.n9094 vss.n9093 35.2919
R36103 vss.n9124 vss.n9123 35.2919
R36104 vss.n9125 vss.n9124 35.2919
R36105 vss.n9125 vss.n9102 35.2919
R36106 vss.n9134 vss.n9102 35.2919
R36107 vss.n9135 vss.n9134 35.2919
R36108 vss.n9136 vss.n9135 35.2919
R36109 vss.n9340 vss.n9330 35.2919
R36110 vss.n9346 vss.n9330 35.2919
R36111 vss.n9347 vss.n9346 35.2919
R36112 vss.n9357 vss.n9347 35.2919
R36113 vss.n9357 vss.n9356 35.2919
R36114 vss.n9356 vss.n9355 35.2919
R36115 vss.n6208 vss.n6207 35.2919
R36116 vss.n6209 vss.n6208 35.2919
R36117 vss.n6209 vss.n6189 35.2919
R36118 vss.n9377 vss.n6189 35.2919
R36119 vss.n9378 vss.n9377 35.2919
R36120 vss.n9379 vss.n9378 35.2919
R36121 vss.n5956 vss.n5947 35.2919
R36122 vss.n5962 vss.n5947 35.2919
R36123 vss.n5963 vss.n5962 35.2919
R36124 vss.n9677 vss.n5963 35.2919
R36125 vss.n9677 vss.n9676 35.2919
R36126 vss.n9676 vss.n9675 35.2919
R36127 vss.n9706 vss.n9695 35.2919
R36128 vss.n9712 vss.n9695 35.2919
R36129 vss.n9713 vss.n9712 35.2919
R36130 vss.n9724 vss.n9713 35.2919
R36131 vss.n9724 vss.n9723 35.2919
R36132 vss.n9723 vss.n9722 35.2919
R36133 vss.n2577 vss.n2568 35.2919
R36134 vss.n2583 vss.n2568 35.2919
R36135 vss.n2584 vss.n2583 35.2919
R36136 vss.n10005 vss.n2584 35.2919
R36137 vss.n10005 vss.n10004 35.2919
R36138 vss.n10004 vss.n10003 35.2919
R36139 vss.n2756 vss.n2746 35.2919
R36140 vss.n9887 vss.n2756 35.2919
R36141 vss.n9887 vss.n9886 35.2919
R36142 vss.n9886 vss.n9885 35.2919
R36143 vss.n9885 vss.n2759 35.2919
R36144 vss.n2765 vss.n2759 35.2919
R36145 vss.n3284 vss.n3273 35.2919
R36146 vss.n3290 vss.n3273 35.2919
R36147 vss.n3291 vss.n3290 35.2919
R36148 vss.n3302 vss.n3291 35.2919
R36149 vss.n3302 vss.n3301 35.2919
R36150 vss.n3301 vss.n3300 35.2919
R36151 vss.n9762 vss.n9754 35.2919
R36152 vss.n9771 vss.n9754 35.2919
R36153 vss.n9772 vss.n9771 35.2919
R36154 vss.n9773 vss.n9772 35.2919
R36155 vss.n9773 vss.n9752 35.2919
R36156 vss.n9777 vss.n9752 35.2919
R36157 vss.n3202 vss.n3194 35.2919
R36158 vss.n3211 vss.n3194 35.2919
R36159 vss.n3212 vss.n3211 35.2919
R36160 vss.n3213 vss.n3212 35.2919
R36161 vss.n3213 vss.n3192 35.2919
R36162 vss.n3217 vss.n3192 35.2919
R36163 vss.n9800 vss.n9799 35.2919
R36164 vss.n9799 vss.n9798 35.2919
R36165 vss.n9798 vss.n2999 35.2919
R36166 vss.n3015 vss.n2999 35.2919
R36167 vss.n3015 vss.n3014 35.2919
R36168 vss.n3019 vss.n3014 35.2919
R36169 vss.n5232 vss.n5224 35.2919
R36170 vss.n5241 vss.n5224 35.2919
R36171 vss.n5242 vss.n5241 35.2919
R36172 vss.n5243 vss.n5242 35.2919
R36173 vss.n5243 vss.n5222 35.2919
R36174 vss.n5247 vss.n5222 35.2919
R36175 vss.n3045 vss.n3037 35.2919
R36176 vss.n3054 vss.n3037 35.2919
R36177 vss.n3055 vss.n3054 35.2919
R36178 vss.n3056 vss.n3055 35.2919
R36179 vss.n3056 vss.n3035 35.2919
R36180 vss.n3060 vss.n3035 35.2919
R36181 vss.n5102 vss.n5094 35.2919
R36182 vss.n5111 vss.n5094 35.2919
R36183 vss.n5112 vss.n5111 35.2919
R36184 vss.n5113 vss.n5112 35.2919
R36185 vss.n5113 vss.n5092 35.2919
R36186 vss.n5117 vss.n5092 35.2919
R36187 vss.n5291 vss.n5283 35.2919
R36188 vss.n5300 vss.n5283 35.2919
R36189 vss.n5301 vss.n5300 35.2919
R36190 vss.n5302 vss.n5301 35.2919
R36191 vss.n5302 vss.n5281 35.2919
R36192 vss.n5306 vss.n5281 35.2919
R36193 vss.n5019 vss.n5011 35.2919
R36194 vss.n5028 vss.n5011 35.2919
R36195 vss.n5029 vss.n5028 35.2919
R36196 vss.n5030 vss.n5029 35.2919
R36197 vss.n5030 vss.n5009 35.2919
R36198 vss.n5034 vss.n5009 35.2919
R36199 vss.n4900 vss.n4892 35.2919
R36200 vss.n4909 vss.n4892 35.2919
R36201 vss.n4910 vss.n4909 35.2919
R36202 vss.n4911 vss.n4910 35.2919
R36203 vss.n4911 vss.n4890 35.2919
R36204 vss.n4915 vss.n4890 35.2919
R36205 vss.n2721 vss.n2711 35.2919
R36206 vss.n9921 vss.n2721 35.2919
R36207 vss.n9921 vss.n9920 35.2919
R36208 vss.n9920 vss.n9919 35.2919
R36209 vss.n9919 vss.n2724 35.2919
R36210 vss.n2730 vss.n2724 35.2919
R36211 vss.n4652 vss.n4639 35.2919
R36212 vss.n4658 vss.n4652 35.2919
R36213 vss.n4658 vss.n4657 35.2919
R36214 vss.n4657 vss.n4656 35.2919
R36215 vss.n4656 vss.n2734 35.2919
R36216 vss.n2737 vss.n2734 35.2919
R36217 vss.n4673 vss.n4630 35.2919
R36218 vss.n5623 vss.n4673 35.2919
R36219 vss.n5623 vss.n5622 35.2919
R36220 vss.n5622 vss.n5621 35.2919
R36221 vss.n5621 vss.n4676 35.2919
R36222 vss.n4682 vss.n4676 35.2919
R36223 vss.n5590 vss.n5589 35.2919
R36224 vss.n5595 vss.n5590 35.2919
R36225 vss.n5595 vss.n5594 35.2919
R36226 vss.n5594 vss.n5593 35.2919
R36227 vss.n5593 vss.n4686 35.2919
R36228 vss.n5602 vss.n4686 35.2919
R36229 vss.n4703 vss.n4701 35.2919
R36230 vss.n4718 vss.n4701 35.2919
R36231 vss.n4719 vss.n4718 35.2919
R36232 vss.n5573 vss.n4719 35.2919
R36233 vss.n5573 vss.n5572 35.2919
R36234 vss.n5572 vss.n5571 35.2919
R36235 vss.n5547 vss.n5546 35.2919
R36236 vss.n5552 vss.n5547 35.2919
R36237 vss.n5552 vss.n5551 35.2919
R36238 vss.n5551 vss.n5550 35.2919
R36239 vss.n5550 vss.n4729 35.2919
R36240 vss.n5559 vss.n4729 35.2919
R36241 vss.n4746 vss.n4744 35.2919
R36242 vss.n4761 vss.n4744 35.2919
R36243 vss.n4762 vss.n4761 35.2919
R36244 vss.n5530 vss.n4762 35.2919
R36245 vss.n5530 vss.n5529 35.2919
R36246 vss.n5529 vss.n5528 35.2919
R36247 vss.n5504 vss.n5503 35.2919
R36248 vss.n5509 vss.n5504 35.2919
R36249 vss.n5509 vss.n5508 35.2919
R36250 vss.n5508 vss.n5507 35.2919
R36251 vss.n5507 vss.n4772 35.2919
R36252 vss.n5516 vss.n4772 35.2919
R36253 vss.n4789 vss.n4787 35.2919
R36254 vss.n4804 vss.n4787 35.2919
R36255 vss.n4805 vss.n4804 35.2919
R36256 vss.n5487 vss.n4805 35.2919
R36257 vss.n5487 vss.n5486 35.2919
R36258 vss.n5486 vss.n5485 35.2919
R36259 vss.n5461 vss.n5460 35.2919
R36260 vss.n5466 vss.n5461 35.2919
R36261 vss.n5466 vss.n5465 35.2919
R36262 vss.n5465 vss.n5464 35.2919
R36263 vss.n5464 vss.n4815 35.2919
R36264 vss.n5473 vss.n4815 35.2919
R36265 vss.n4832 vss.n4830 35.2919
R36266 vss.n4847 vss.n4830 35.2919
R36267 vss.n4848 vss.n4847 35.2919
R36268 vss.n5444 vss.n4848 35.2919
R36269 vss.n5444 vss.n5443 35.2919
R36270 vss.n5443 vss.n5442 35.2919
R36271 vss.n5418 vss.n5417 35.2919
R36272 vss.n5423 vss.n5418 35.2919
R36273 vss.n5423 vss.n5422 35.2919
R36274 vss.n5422 vss.n5421 35.2919
R36275 vss.n5421 vss.n4858 35.2919
R36276 vss.n5430 vss.n4858 35.2919
R36277 vss.n4875 vss.n4873 35.2919
R36278 vss.n5341 vss.n4873 35.2919
R36279 vss.n5342 vss.n5341 35.2919
R36280 vss.n5401 vss.n5342 35.2919
R36281 vss.n5401 vss.n5400 35.2919
R36282 vss.n5400 vss.n5399 35.2919
R36283 vss.n5375 vss.n5374 35.2919
R36284 vss.n5374 vss.n5373 35.2919
R36285 vss.n5373 vss.n5368 35.2919
R36286 vss.n5369 vss.n5368 35.2919
R36287 vss.n5369 vss.n5352 35.2919
R36288 vss.n5386 vss.n5352 35.2919
R36289 vss.n9821 vss.n2882 35.2919
R36290 vss.n9830 vss.n2882 35.2919
R36291 vss.n9831 vss.n9830 35.2919
R36292 vss.n9832 vss.n9831 35.2919
R36293 vss.n9832 vss.n2880 35.2919
R36294 vss.n9836 vss.n2880 35.2919
R36295 vss.n2977 vss.n2976 35.2919
R36296 vss.n2976 vss.n2975 35.2919
R36297 vss.n2975 vss.n2942 35.2919
R36298 vss.n2958 vss.n2942 35.2919
R36299 vss.n2958 vss.n2957 35.2919
R36300 vss.n2962 vss.n2957 35.2919
R36301 vss.n2931 vss.n2930 35.2919
R36302 vss.n2930 vss.n2929 35.2919
R36303 vss.n2929 vss.n2895 35.2919
R36304 vss.n2911 vss.n2895 35.2919
R36305 vss.n2911 vss.n2910 35.2919
R36306 vss.n2915 vss.n2910 35.2919
R36307 vss.n4941 vss.n4933 35.2919
R36308 vss.n4950 vss.n4933 35.2919
R36309 vss.n4951 vss.n4950 35.2919
R36310 vss.n4952 vss.n4951 35.2919
R36311 vss.n4952 vss.n4931 35.2919
R36312 vss.n4956 vss.n4931 35.2919
R36313 vss.n5143 vss.n5135 35.2919
R36314 vss.n5152 vss.n5135 35.2919
R36315 vss.n5153 vss.n5152 35.2919
R36316 vss.n5154 vss.n5153 35.2919
R36317 vss.n5154 vss.n5133 35.2919
R36318 vss.n5158 vss.n5133 35.2919
R36319 vss.n3124 vss.n3115 35.2919
R36320 vss.n3133 vss.n3115 35.2919
R36321 vss.n3134 vss.n3133 35.2919
R36322 vss.n3135 vss.n3134 35.2919
R36323 vss.n3135 vss.n3113 35.2919
R36324 vss.n3139 vss.n3113 35.2919
R36325 vss.n4482 vss.n4470 35.2919
R36326 vss.n4488 vss.n4470 35.2919
R36327 vss.n4489 vss.n4488 35.2919
R36328 vss.n4490 vss.n4489 35.2919
R36329 vss.n4491 vss.n4490 35.2919
R36330 vss.n4495 vss.n4491 35.2919
R36331 vss.n4390 vss.n4378 35.2919
R36332 vss.n4396 vss.n4378 35.2919
R36333 vss.n4397 vss.n4396 35.2919
R36334 vss.n4398 vss.n4397 35.2919
R36335 vss.n4399 vss.n4398 35.2919
R36336 vss.n4403 vss.n4399 35.2919
R36337 vss.n4342 vss.n4330 35.2919
R36338 vss.n4348 vss.n4330 35.2919
R36339 vss.n4349 vss.n4348 35.2919
R36340 vss.n4350 vss.n4349 35.2919
R36341 vss.n4351 vss.n4350 35.2919
R36342 vss.n4355 vss.n4351 35.2919
R36343 vss.n3742 vss.n3730 35.2919
R36344 vss.n3748 vss.n3730 35.2919
R36345 vss.n3749 vss.n3748 35.2919
R36346 vss.n3750 vss.n3749 35.2919
R36347 vss.n3751 vss.n3750 35.2919
R36348 vss.n3755 vss.n3751 35.2919
R36349 vss.n4044 vss.n4032 35.2919
R36350 vss.n4050 vss.n4032 35.2919
R36351 vss.n4051 vss.n4050 35.2919
R36352 vss.n4052 vss.n4051 35.2919
R36353 vss.n4053 vss.n4052 35.2919
R36354 vss.n4057 vss.n4053 35.2919
R36355 vss.n3697 vss.n3685 35.2919
R36356 vss.n3703 vss.n3685 35.2919
R36357 vss.n3704 vss.n3703 35.2919
R36358 vss.n3705 vss.n3704 35.2919
R36359 vss.n3706 vss.n3705 35.2919
R36360 vss.n3710 vss.n3706 35.2919
R36361 vss.n4098 vss.n4086 35.2919
R36362 vss.n4104 vss.n4086 35.2919
R36363 vss.n4105 vss.n4104 35.2919
R36364 vss.n4106 vss.n4105 35.2919
R36365 vss.n4107 vss.n4106 35.2919
R36366 vss.n4111 vss.n4107 35.2919
R36367 vss.n3522 vss.n3510 35.2919
R36368 vss.n3528 vss.n3510 35.2919
R36369 vss.n3529 vss.n3528 35.2919
R36370 vss.n3530 vss.n3529 35.2919
R36371 vss.n3531 vss.n3530 35.2919
R36372 vss.n3535 vss.n3531 35.2919
R36373 vss.n3477 vss.n3465 35.2919
R36374 vss.n3483 vss.n3465 35.2919
R36375 vss.n3484 vss.n3483 35.2919
R36376 vss.n3485 vss.n3484 35.2919
R36377 vss.n3486 vss.n3485 35.2919
R36378 vss.n3490 vss.n3486 35.2919
R36379 vss.n5765 vss.n5753 35.2919
R36380 vss.n5771 vss.n5753 35.2919
R36381 vss.n5772 vss.n5771 35.2919
R36382 vss.n5773 vss.n5772 35.2919
R36383 vss.n5774 vss.n5773 35.2919
R36384 vss.n5778 vss.n5774 35.2919
R36385 vss.n4519 vss.n4518 35.2919
R36386 vss.n4520 vss.n4519 35.2919
R36387 vss.n4521 vss.n4520 35.2919
R36388 vss.n4522 vss.n4521 35.2919
R36389 vss.n4523 vss.n4522 35.2919
R36390 vss.n4524 vss.n4523 35.2919
R36391 vss.n4541 vss.n4540 35.2919
R36392 vss.n4542 vss.n4541 35.2919
R36393 vss.n4542 vss.n4427 35.2919
R36394 vss.n4551 vss.n4427 35.2919
R36395 vss.n4552 vss.n4551 35.2919
R36396 vss.n4553 vss.n4552 35.2919
R36397 vss.n4589 vss.n4560 35.2919
R36398 vss.n4595 vss.n4560 35.2919
R36399 vss.n4596 vss.n4595 35.2919
R36400 vss.n4597 vss.n4596 35.2919
R36401 vss.n4598 vss.n4597 35.2919
R36402 vss.n4602 vss.n4598 35.2919
R36403 vss.n4583 vss.n4582 35.2919
R36404 vss.n4582 vss.n4581 35.2919
R36405 vss.n4581 vss.n3635 35.2919
R36406 vss.n4622 vss.n3635 35.2919
R36407 vss.n4623 vss.n4622 35.2919
R36408 vss.n4624 vss.n4623 35.2919
R36409 vss.n4186 vss.n3774 35.2919
R36410 vss.n4192 vss.n3774 35.2919
R36411 vss.n4193 vss.n4192 35.2919
R36412 vss.n4194 vss.n4193 35.2919
R36413 vss.n4195 vss.n4194 35.2919
R36414 vss.n4199 vss.n4195 35.2919
R36415 vss.n4180 vss.n4179 35.2919
R36416 vss.n4179 vss.n4178 35.2919
R36417 vss.n4178 vss.n3788 35.2919
R36418 vss.n3821 vss.n3788 35.2919
R36419 vss.n3822 vss.n3821 35.2919
R36420 vss.n3823 vss.n3822 35.2919
R36421 vss.n4151 vss.n3830 35.2919
R36422 vss.n4157 vss.n3830 35.2919
R36423 vss.n4158 vss.n4157 35.2919
R36424 vss.n4159 vss.n4158 35.2919
R36425 vss.n4160 vss.n4159 35.2919
R36426 vss.n4164 vss.n4160 35.2919
R36427 vss.n4145 vss.n4144 35.2919
R36428 vss.n4144 vss.n4143 35.2919
R36429 vss.n4143 vss.n3844 35.2919
R36430 vss.n3864 vss.n3844 35.2919
R36431 vss.n3865 vss.n3864 35.2919
R36432 vss.n3866 vss.n3865 35.2919
R36433 vss.n3941 vss.n3940 35.2919
R36434 vss.n3942 vss.n3941 35.2919
R36435 vss.n3942 vss.n3874 35.2919
R36436 vss.n4129 vss.n3874 35.2919
R36437 vss.n4130 vss.n4129 35.2919
R36438 vss.n4131 vss.n4130 35.2919
R36439 vss.n3932 vss.n3931 35.2919
R36440 vss.n3931 vss.n3930 35.2919
R36441 vss.n3930 vss.n3896 35.2919
R36442 vss.n3915 vss.n3896 35.2919
R36443 vss.n3916 vss.n3915 35.2919
R36444 vss.n3917 vss.n3916 35.2919
R36445 vss.n5818 vss.n3553 35.2919
R36446 vss.n5824 vss.n3553 35.2919
R36447 vss.n5825 vss.n5824 35.2919
R36448 vss.n5826 vss.n5825 35.2919
R36449 vss.n5827 vss.n5826 35.2919
R36450 vss.n5831 vss.n5827 35.2919
R36451 vss.n5812 vss.n5811 35.2919
R36452 vss.n5811 vss.n5810 35.2919
R36453 vss.n5810 vss.n3567 35.2919
R36454 vss.n3618 vss.n3567 35.2919
R36455 vss.n3619 vss.n3618 35.2919
R36456 vss.n3620 vss.n3619 35.2919
R36457 vss.n5669 vss.n5668 35.2919
R36458 vss.n5670 vss.n5669 35.2919
R36459 vss.n5670 vss.n3588 35.2919
R36460 vss.n5796 vss.n3588 35.2919
R36461 vss.n5797 vss.n5796 35.2919
R36462 vss.n5798 vss.n5797 35.2919
R36463 vss.n5678 vss.n5649 35.2919
R36464 vss.n5684 vss.n5649 35.2919
R36465 vss.n5685 vss.n5684 35.2919
R36466 vss.n5686 vss.n5685 35.2919
R36467 vss.n5687 vss.n5686 35.2919
R36468 vss.n5688 vss.n5687 35.2919
R36469 vss.n5718 vss.n5717 35.2919
R36470 vss.n5719 vss.n5718 35.2919
R36471 vss.n5719 vss.n5696 35.2919
R36472 vss.n5728 vss.n5696 35.2919
R36473 vss.n5729 vss.n5728 35.2919
R36474 vss.n5730 vss.n5729 35.2919
R36475 vss.n9969 vss.n9957 35.2919
R36476 vss.n9975 vss.n9957 35.2919
R36477 vss.n9976 vss.n9975 35.2919
R36478 vss.n9977 vss.n9976 35.2919
R36479 vss.n9978 vss.n9977 35.2919
R36480 vss.n9982 vss.n9978 35.2919
R36481 vss.n2667 vss.n2666 35.2919
R36482 vss.n2668 vss.n2667 35.2919
R36483 vss.n2668 vss.n2644 35.2919
R36484 vss.n2679 vss.n2644 35.2919
R36485 vss.n2680 vss.n2679 35.2919
R36486 vss.n2681 vss.n2680 35.2919
R36487 vss.n3402 vss.n3390 35.2919
R36488 vss.n3408 vss.n3390 35.2919
R36489 vss.n3409 vss.n3408 35.2919
R36490 vss.n3410 vss.n3409 35.2919
R36491 vss.n3411 vss.n3410 35.2919
R36492 vss.n3415 vss.n3411 35.2919
R36493 vss.n3999 vss.n3987 35.2919
R36494 vss.n4005 vss.n3987 35.2919
R36495 vss.n4006 vss.n4005 35.2919
R36496 vss.n4007 vss.n4006 35.2919
R36497 vss.n4008 vss.n4007 35.2919
R36498 vss.n4012 vss.n4008 35.2919
R36499 vss.n4266 vss.n4254 35.2919
R36500 vss.n4272 vss.n4254 35.2919
R36501 vss.n4273 vss.n4272 35.2919
R36502 vss.n4274 vss.n4273 35.2919
R36503 vss.n4275 vss.n4274 35.2919
R36504 vss.n4279 vss.n4275 35.2919
R36505 vss.n5909 vss.n5899 35.2919
R36506 vss.n5915 vss.n5899 35.2919
R36507 vss.n5916 vss.n5915 35.2919
R36508 vss.n5926 vss.n5916 35.2919
R36509 vss.n5926 vss.n5925 35.2919
R36510 vss.n5925 vss.n5924 35.2919
R36511 vss.n14065 vss.n487 35.2919
R36512 vss.n14074 vss.n487 35.2919
R36513 vss.n14075 vss.n14074 35.2919
R36514 vss.n14076 vss.n14075 35.2919
R36515 vss.n14076 vss.n485 35.2919
R36516 vss.n14080 vss.n485 35.2919
R36517 vss.n10120 vss.n10112 35.2919
R36518 vss.n10129 vss.n10112 35.2919
R36519 vss.n10130 vss.n10129 35.2919
R36520 vss.n10131 vss.n10130 35.2919
R36521 vss.n10131 vss.n10110 35.2919
R36522 vss.n10135 vss.n10110 35.2919
R36523 vss.n12878 vss.n12870 35.2919
R36524 vss.n12887 vss.n12870 35.2919
R36525 vss.n12888 vss.n12887 35.2919
R36526 vss.n12889 vss.n12888 35.2919
R36527 vss.n12889 vss.n12868 35.2919
R36528 vss.n12893 vss.n12868 35.2919
R36529 vss.n10161 vss.n10153 35.2919
R36530 vss.n10170 vss.n10153 35.2919
R36531 vss.n10171 vss.n10170 35.2919
R36532 vss.n10172 vss.n10171 35.2919
R36533 vss.n10172 vss.n10151 35.2919
R36534 vss.n10176 vss.n10151 35.2919
R36535 vss.n12427 vss.n12419 35.2919
R36536 vss.n12436 vss.n12419 35.2919
R36537 vss.n12437 vss.n12436 35.2919
R36538 vss.n12438 vss.n12437 35.2919
R36539 vss.n12438 vss.n12417 35.2919
R36540 vss.n12442 vss.n12417 35.2919
R36541 vss.n11756 vss.n11748 35.2919
R36542 vss.n11765 vss.n11748 35.2919
R36543 vss.n11766 vss.n11765 35.2919
R36544 vss.n11767 vss.n11766 35.2919
R36545 vss.n11767 vss.n11746 35.2919
R36546 vss.n11771 vss.n11746 35.2919
R36547 vss.n12472 vss.n12464 35.2919
R36548 vss.n12481 vss.n12464 35.2919
R36549 vss.n12482 vss.n12481 35.2919
R36550 vss.n12483 vss.n12482 35.2919
R36551 vss.n12483 vss.n12462 35.2919
R36552 vss.n12487 vss.n12462 35.2919
R36553 vss.n2347 vss.n2346 35.2919
R36554 vss.n2346 vss.n2345 35.2919
R36555 vss.n2345 vss.n2312 35.2919
R36556 vss.n2328 vss.n2312 35.2919
R36557 vss.n2328 vss.n2327 35.2919
R36558 vss.n2332 vss.n2327 35.2919
R36559 vss.n12297 vss.n12289 35.2919
R36560 vss.n12306 vss.n12289 35.2919
R36561 vss.n12307 vss.n12306 35.2919
R36562 vss.n12308 vss.n12307 35.2919
R36563 vss.n12308 vss.n12287 35.2919
R36564 vss.n12312 vss.n12287 35.2919
R36565 vss.n12342 vss.n12334 35.2919
R36566 vss.n12351 vss.n12334 35.2919
R36567 vss.n12352 vss.n12351 35.2919
R36568 vss.n12353 vss.n12352 35.2919
R36569 vss.n12353 vss.n12332 35.2919
R36570 vss.n12357 vss.n12332 35.2919
R36571 vss.n10238 vss.n10230 35.2919
R36572 vss.n10247 vss.n10230 35.2919
R36573 vss.n10248 vss.n10247 35.2919
R36574 vss.n10249 vss.n10248 35.2919
R36575 vss.n10249 vss.n10228 35.2919
R36576 vss.n10253 vss.n10228 35.2919
R36577 vss.n2418 vss.n2410 35.2919
R36578 vss.n2427 vss.n2410 35.2919
R36579 vss.n2428 vss.n2427 35.2919
R36580 vss.n2429 vss.n2428 35.2919
R36581 vss.n2429 vss.n2408 35.2919
R36582 vss.n2433 vss.n2408 35.2919
R36583 vss.n12972 vss.n12971 35.2919
R36584 vss.n12971 vss.n12970 35.2919
R36585 vss.n12970 vss.n2372 35.2919
R36586 vss.n2388 vss.n2372 35.2919
R36587 vss.n2388 vss.n2387 35.2919
R36588 vss.n2392 vss.n2387 35.2919
R36589 vss.n10044 vss.n10027 35.2919
R36590 vss.n10050 vss.n10027 35.2919
R36591 vss.n10051 vss.n10050 35.2919
R36592 vss.n12947 vss.n10051 35.2919
R36593 vss.n12947 vss.n12946 35.2919
R36594 vss.n12946 vss.n12945 35.2919
R36595 vss.n10038 vss.n2098 35.2919
R36596 vss.n2110 vss.n2098 35.2919
R36597 vss.n2111 vss.n2110 35.2919
R36598 vss.n13082 vss.n2111 35.2919
R36599 vss.n13082 vss.n13081 35.2919
R36600 vss.n13081 vss.n13080 35.2919
R36601 vss.n12923 vss.n10075 35.2919
R36602 vss.n12931 vss.n10075 35.2919
R36603 vss.n12932 vss.n12931 35.2919
R36604 vss.n12933 vss.n12932 35.2919
R36605 vss.n12933 vss.n10062 35.2919
R36606 vss.n12940 vss.n10062 35.2919
R36607 vss.n2498 vss.n2489 35.2919
R36608 vss.n2507 vss.n2489 35.2919
R36609 vss.n2508 vss.n2507 35.2919
R36610 vss.n2509 vss.n2508 35.2919
R36611 vss.n2509 vss.n2487 35.2919
R36612 vss.n2513 vss.n2487 35.2919
R36613 vss.n2132 vss.n2122 35.2919
R36614 vss.n13068 vss.n2132 35.2919
R36615 vss.n13068 vss.n13067 35.2919
R36616 vss.n13067 vss.n13066 35.2919
R36617 vss.n13066 vss.n2135 35.2919
R36618 vss.n2141 vss.n2135 35.2919
R36619 vss.n12101 vss.n11842 35.2919
R36620 vss.n12109 vss.n11842 35.2919
R36621 vss.n12110 vss.n12109 35.2919
R36622 vss.n12111 vss.n12110 35.2919
R36623 vss.n12111 vss.n11831 35.2919
R36624 vss.n12120 vss.n11831 35.2919
R36625 vss.n12150 vss.n12149 35.2919
R36626 vss.n12149 vss.n12148 35.2919
R36627 vss.n12148 vss.n11813 35.2919
R36628 vss.n12127 vss.n11813 35.2919
R36629 vss.n12127 vss.n12126 35.2919
R36630 vss.n12131 vss.n12126 35.2919
R36631 vss.n12154 vss.n11798 35.2919
R36632 vss.n12162 vss.n11798 35.2919
R36633 vss.n12163 vss.n12162 35.2919
R36634 vss.n12164 vss.n12163 35.2919
R36635 vss.n12164 vss.n11790 35.2919
R36636 vss.n12173 vss.n11790 35.2919
R36637 vss.n12187 vss.n12181 35.2919
R36638 vss.n12262 vss.n12181 35.2919
R36639 vss.n12263 vss.n12262 35.2919
R36640 vss.n12264 vss.n12263 35.2919
R36641 vss.n12264 vss.n12179 35.2919
R36642 vss.n12268 vss.n12179 35.2919
R36643 vss.n12248 vss.n12247 35.2919
R36644 vss.n12247 vss.n12246 35.2919
R36645 vss.n12246 vss.n12195 35.2919
R36646 vss.n12231 vss.n12195 35.2919
R36647 vss.n12232 vss.n12231 35.2919
R36648 vss.n12234 vss.n12232 35.2919
R36649 vss.n12546 vss.n12545 35.2919
R36650 vss.n12545 vss.n12544 35.2919
R36651 vss.n12544 vss.n11725 35.2919
R36652 vss.n12217 vss.n11725 35.2919
R36653 vss.n12217 vss.n12213 35.2919
R36654 vss.n12213 vss.n12212 35.2919
R36655 vss.n12550 vss.n11711 35.2919
R36656 vss.n12558 vss.n11711 35.2919
R36657 vss.n12559 vss.n12558 35.2919
R36658 vss.n12560 vss.n12559 35.2919
R36659 vss.n12560 vss.n11703 35.2919
R36660 vss.n12569 vss.n11703 35.2919
R36661 vss.n11690 vss.n11626 35.2919
R36662 vss.n11691 vss.n11690 35.2919
R36663 vss.n11691 vss.n11639 35.2919
R36664 vss.n11695 vss.n11639 35.2919
R36665 vss.n11696 vss.n11695 35.2919
R36666 vss.n11697 vss.n11696 35.2919
R36667 vss.n11683 vss.n11682 35.2919
R36668 vss.n11682 vss.n11681 35.2919
R36669 vss.n11681 vss.n11646 35.2919
R36670 vss.n11666 vss.n11646 35.2919
R36671 vss.n11667 vss.n11666 35.2919
R36672 vss.n11669 vss.n11667 35.2919
R36673 vss.n10319 vss.n10313 35.2919
R36674 vss.n12842 vss.n10313 35.2919
R36675 vss.n12843 vss.n12842 35.2919
R36676 vss.n12844 vss.n12843 35.2919
R36677 vss.n12844 vss.n10311 35.2919
R36678 vss.n12848 vss.n10311 35.2919
R36679 vss.n12828 vss.n12827 35.2919
R36680 vss.n12827 vss.n12826 35.2919
R36681 vss.n12826 vss.n12777 35.2919
R36682 vss.n12813 vss.n12777 35.2919
R36683 vss.n12814 vss.n12813 35.2919
R36684 vss.n12816 vss.n12814 35.2919
R36685 vss.n12919 vss.n12918 35.2919
R36686 vss.n12918 vss.n12917 35.2919
R36687 vss.n12917 vss.n10090 35.2919
R36688 vss.n12799 vss.n10090 35.2919
R36689 vss.n12799 vss.n12795 35.2919
R36690 vss.n12795 vss.n12794 35.2919
R36691 vss.n11884 vss.n11883 35.2919
R36692 vss.n11885 vss.n11884 35.2919
R36693 vss.n11885 vss.n11862 35.2919
R36694 vss.n12081 vss.n11862 35.2919
R36695 vss.n12082 vss.n12081 35.2919
R36696 vss.n12083 vss.n12082 35.2919
R36697 vss.n10481 vss.n10470 35.2919
R36698 vss.n10487 vss.n10470 35.2919
R36699 vss.n10488 vss.n10487 35.2919
R36700 vss.n10489 vss.n10488 35.2919
R36701 vss.n10490 vss.n10489 35.2919
R36702 vss.n10494 vss.n10490 35.2919
R36703 vss.n10702 vss.n10691 35.2919
R36704 vss.n10708 vss.n10691 35.2919
R36705 vss.n10709 vss.n10708 35.2919
R36706 vss.n10710 vss.n10709 35.2919
R36707 vss.n10711 vss.n10710 35.2919
R36708 vss.n10715 vss.n10711 35.2919
R36709 vss.n11016 vss.n11005 35.2919
R36710 vss.n11022 vss.n11005 35.2919
R36711 vss.n11023 vss.n11022 35.2919
R36712 vss.n11024 vss.n11023 35.2919
R36713 vss.n11025 vss.n11024 35.2919
R36714 vss.n11029 vss.n11025 35.2919
R36715 vss.n11124 vss.n11115 35.2919
R36716 vss.n11130 vss.n11115 35.2919
R36717 vss.n11131 vss.n11130 35.2919
R36718 vss.n11141 vss.n11131 35.2919
R36719 vss.n11141 vss.n11140 35.2919
R36720 vss.n11140 vss.n11139 35.2919
R36721 vss.t79 vss.n2072 34.5778
R36722 vss.n9648 vss.n9647 31.1326
R36723 vss.n13092 vss.n13091 31.1326
R36724 vss.n11090 vss.n11084 27.0634
R36725 vss.n11093 vss.n11090 27.0634
R36726 vss.n11094 vss.n11093 27.0634
R36727 vss.n11095 vss.n11094 27.0634
R36728 vss.n11095 vss.n11088 27.0634
R36729 vss.n11099 vss.n11088 27.0634
R36730 vss.n11169 vss.n11159 27.0634
R36731 vss.n11169 vss.n11168 27.0634
R36732 vss.n11168 vss.n11160 27.0634
R36733 vss.n11164 vss.n11160 27.0634
R36734 vss.n11164 vss.n11163 27.0634
R36735 vss.n11163 vss.n11046 27.0634
R36736 vss.n11216 vss.n11210 27.0634
R36737 vss.n11219 vss.n11216 27.0634
R36738 vss.n11220 vss.n11219 27.0634
R36739 vss.n11221 vss.n11220 27.0634
R36740 vss.n11221 vss.n11214 27.0634
R36741 vss.n11225 vss.n11214 27.0634
R36742 vss.n11277 vss.n11271 27.0634
R36743 vss.n11280 vss.n11277 27.0634
R36744 vss.n11281 vss.n11280 27.0634
R36745 vss.n11282 vss.n11281 27.0634
R36746 vss.n11282 vss.n11275 27.0634
R36747 vss.n11286 vss.n11275 27.0634
R36748 vss.n14770 vss.n14769 27.0634
R36749 vss.n14769 vss.n103 27.0634
R36750 vss.n110 vss.n103 27.0634
R36751 vss.n111 vss.n110 27.0634
R36752 vss.n115 vss.n111 27.0634
R36753 vss.n115 vss.n114 27.0634
R36754 vss.n397 vss.n396 27.0634
R36755 vss.n398 vss.n397 27.0634
R36756 vss.n399 vss.n398 27.0634
R36757 vss.n400 vss.n399 27.0634
R36758 vss.n404 vss.n400 27.0634
R36759 vss.n404 vss.n403 27.0634
R36760 vss.n274 vss.n273 27.0634
R36761 vss.n275 vss.n274 27.0634
R36762 vss.n276 vss.n275 27.0634
R36763 vss.n277 vss.n276 27.0634
R36764 vss.n281 vss.n277 27.0634
R36765 vss.n281 vss.n280 27.0634
R36766 vss.n14431 vss.n14430 27.0634
R36767 vss.n14432 vss.n14431 27.0634
R36768 vss.n14433 vss.n14432 27.0634
R36769 vss.n14434 vss.n14433 27.0634
R36770 vss.n14438 vss.n14434 27.0634
R36771 vss.n14438 vss.n14437 27.0634
R36772 vss.n215 vss.n214 27.0634
R36773 vss.n216 vss.n215 27.0634
R36774 vss.n217 vss.n216 27.0634
R36775 vss.n218 vss.n217 27.0634
R36776 vss.n222 vss.n218 27.0634
R36777 vss.n222 vss.n221 27.0634
R36778 vss.n14626 vss.n14625 27.0634
R36779 vss.n14627 vss.n14626 27.0634
R36780 vss.n14628 vss.n14627 27.0634
R36781 vss.n14629 vss.n14628 27.0634
R36782 vss.n14633 vss.n14629 27.0634
R36783 vss.n14633 vss.n14632 27.0634
R36784 vss.n138 vss.n137 27.0634
R36785 vss.n139 vss.n138 27.0634
R36786 vss.n140 vss.n139 27.0634
R36787 vss.n141 vss.n140 27.0634
R36788 vss.n145 vss.n141 27.0634
R36789 vss.n145 vss.n144 27.0634
R36790 vss.n373 vss.n372 27.0634
R36791 vss.n372 vss.n371 27.0634
R36792 vss.n371 vss.n370 27.0634
R36793 vss.n370 vss.n68 27.0634
R36794 vss.n14777 vss.n68 27.0634
R36795 vss.n14778 vss.n14777 27.0634
R36796 vss.n7356 vss.n7355 27.0634
R36797 vss.n7357 vss.n7356 27.0634
R36798 vss.n7357 vss.n7350 27.0634
R36799 vss.n7361 vss.n7350 27.0634
R36800 vss.n7367 vss.n7361 27.0634
R36801 vss.n7367 vss.n7366 27.0634
R36802 vss.n7823 vss.n7820 27.0634
R36803 vss.n7833 vss.n7820 27.0634
R36804 vss.n7834 vss.n7833 27.0634
R36805 vss.n7835 vss.n7834 27.0634
R36806 vss.n7835 vss.n7814 27.0634
R36807 vss.n7839 vss.n7814 27.0634
R36808 vss.n7636 vss.n7633 27.0634
R36809 vss.n7646 vss.n7633 27.0634
R36810 vss.n7647 vss.n7646 27.0634
R36811 vss.n7648 vss.n7647 27.0634
R36812 vss.n7648 vss.n7627 27.0634
R36813 vss.n7652 vss.n7627 27.0634
R36814 vss.n7447 vss.n7444 27.0634
R36815 vss.n7457 vss.n7444 27.0634
R36816 vss.n7458 vss.n7457 27.0634
R36817 vss.n7459 vss.n7458 27.0634
R36818 vss.n7459 vss.n7438 27.0634
R36819 vss.n7463 vss.n7438 27.0634
R36820 vss.n7418 vss.n7417 27.0634
R36821 vss.n7423 vss.n7417 27.0634
R36822 vss.n7424 vss.n7423 27.0634
R36823 vss.n7425 vss.n7424 27.0634
R36824 vss.n7425 vss.n7412 27.0634
R36825 vss.n7429 vss.n7412 27.0634
R36826 vss.n7601 vss.n7598 27.0634
R36827 vss.n7611 vss.n7598 27.0634
R36828 vss.n7612 vss.n7611 27.0634
R36829 vss.n7613 vss.n7612 27.0634
R36830 vss.n7613 vss.n7592 27.0634
R36831 vss.n7617 vss.n7592 27.0634
R36832 vss.n7744 vss.n7741 27.0634
R36833 vss.n7754 vss.n7741 27.0634
R36834 vss.n7755 vss.n7754 27.0634
R36835 vss.n7756 vss.n7755 27.0634
R36836 vss.n7756 vss.n7735 27.0634
R36837 vss.n7760 vss.n7735 27.0634
R36838 vss.n7965 vss.n7962 27.0634
R36839 vss.n7975 vss.n7962 27.0634
R36840 vss.n7976 vss.n7975 27.0634
R36841 vss.n7977 vss.n7976 27.0634
R36842 vss.n7977 vss.n7956 27.0634
R36843 vss.n7981 vss.n7956 27.0634
R36844 vss.n3243 vss.n3234 27.0634
R36845 vss.n3247 vss.n3234 27.0634
R36846 vss.n3248 vss.n3247 27.0634
R36847 vss.n3249 vss.n3248 27.0634
R36848 vss.n3249 vss.n3231 27.0634
R36849 vss.n3253 vss.n3231 27.0634
R36850 vss.n3086 vss.n3077 27.0634
R36851 vss.n3090 vss.n3077 27.0634
R36852 vss.n3091 vss.n3090 27.0634
R36853 vss.n3092 vss.n3091 27.0634
R36854 vss.n3092 vss.n3074 27.0634
R36855 vss.n3096 vss.n3074 27.0634
R36856 vss.n5060 vss.n5051 27.0634
R36857 vss.n5064 vss.n5051 27.0634
R36858 vss.n5065 vss.n5064 27.0634
R36859 vss.n5066 vss.n5065 27.0634
R36860 vss.n5066 vss.n5048 27.0634
R36861 vss.n5070 vss.n5048 27.0634
R36862 vss.n2852 vss.n2843 27.0634
R36863 vss.n2856 vss.n2843 27.0634
R36864 vss.n2857 vss.n2856 27.0634
R36865 vss.n2858 vss.n2857 27.0634
R36866 vss.n2858 vss.n2840 27.0634
R36867 vss.n2862 vss.n2840 27.0634
R36868 vss.n9870 vss.n9869 27.0634
R36869 vss.n9869 vss.n9868 27.0634
R36870 vss.n9868 vss.n2829 27.0634
R36871 vss.n9864 vss.n2829 27.0634
R36872 vss.n9864 vss.n9863 27.0634
R36873 vss.n9863 vss.n2833 27.0634
R36874 vss.n4983 vss.n4974 27.0634
R36875 vss.n4987 vss.n4974 27.0634
R36876 vss.n4988 vss.n4987 27.0634
R36877 vss.n4989 vss.n4988 27.0634
R36878 vss.n4989 vss.n4971 27.0634
R36879 vss.n4993 vss.n4971 27.0634
R36880 vss.n5185 vss.n5176 27.0634
R36881 vss.n5189 vss.n5176 27.0634
R36882 vss.n5190 vss.n5189 27.0634
R36883 vss.n5191 vss.n5190 27.0634
R36884 vss.n5191 vss.n5173 27.0634
R36885 vss.n5195 vss.n5173 27.0634
R36886 vss.n3166 vss.n3157 27.0634
R36887 vss.n3170 vss.n3157 27.0634
R36888 vss.n3171 vss.n3170 27.0634
R36889 vss.n3172 vss.n3171 27.0634
R36890 vss.n3172 vss.n3154 27.0634
R36891 vss.n3176 vss.n3154 27.0634
R36892 vss.n10202 vss.n10193 27.0634
R36893 vss.n10206 vss.n10193 27.0634
R36894 vss.n10207 vss.n10206 27.0634
R36895 vss.n10208 vss.n10207 27.0634
R36896 vss.n10208 vss.n10190 27.0634
R36897 vss.n10212 vss.n10190 27.0634
R36898 vss.n12513 vss.n12504 27.0634
R36899 vss.n12517 vss.n12504 27.0634
R36900 vss.n12518 vss.n12517 27.0634
R36901 vss.n12519 vss.n12518 27.0634
R36902 vss.n12519 vss.n12501 27.0634
R36903 vss.n12523 vss.n12501 27.0634
R36904 vss.n2221 vss.n2212 27.0634
R36905 vss.n2225 vss.n2212 27.0634
R36906 vss.n2226 vss.n2225 27.0634
R36907 vss.n2227 vss.n2226 27.0634
R36908 vss.n2227 vss.n2209 27.0634
R36909 vss.n2231 vss.n2209 27.0634
R36910 vss.n12384 vss.n12375 27.0634
R36911 vss.n12388 vss.n12375 27.0634
R36912 vss.n12389 vss.n12388 27.0634
R36913 vss.n12390 vss.n12389 27.0634
R36914 vss.n12390 vss.n12372 27.0634
R36915 vss.n12394 vss.n12372 27.0634
R36916 vss.n10280 vss.n10271 27.0634
R36917 vss.n10284 vss.n10271 27.0634
R36918 vss.n10285 vss.n10284 27.0634
R36919 vss.n10286 vss.n10285 27.0634
R36920 vss.n10286 vss.n10268 27.0634
R36921 vss.n10290 vss.n10268 27.0634
R36922 vss.n2460 vss.n2451 27.0634
R36923 vss.n2464 vss.n2451 27.0634
R36924 vss.n2465 vss.n2464 27.0634
R36925 vss.n2466 vss.n2465 27.0634
R36926 vss.n2466 vss.n2448 27.0634
R36927 vss.n2470 vss.n2448 27.0634
R36928 vss.n2539 vss.n2530 27.0634
R36929 vss.n2543 vss.n2530 27.0634
R36930 vss.n2544 vss.n2543 27.0634
R36931 vss.n2545 vss.n2544 27.0634
R36932 vss.n2545 vss.n2527 27.0634
R36933 vss.n2549 vss.n2527 27.0634
R36934 vss.n13031 vss.n13027 27.0634
R36935 vss.n13036 vss.n13027 27.0634
R36936 vss.n13038 vss.n13036 27.0634
R36937 vss.n13038 vss.n13037 27.0634
R36938 vss.n13037 vss.n2204 27.0634
R36939 vss.n13050 vss.n2204 27.0634
R36940 vss.n11321 vss.n11302 27.0634
R36941 vss.n11321 vss.n11320 27.0634
R36942 vss.n11320 vss.n11303 27.0634
R36943 vss.n11316 vss.n11303 27.0634
R36944 vss.n11316 vss.n11315 27.0634
R36945 vss.n11315 vss.n11314 27.0634
R36946 vss.n11260 vss.n11241 27.0634
R36947 vss.n11260 vss.n11259 27.0634
R36948 vss.n11259 vss.n11242 27.0634
R36949 vss.n11255 vss.n11242 27.0634
R36950 vss.n11255 vss.n11254 27.0634
R36951 vss.n11254 vss.n11253 27.0634
R36952 vss.n11185 vss.n11179 27.0634
R36953 vss.n11188 vss.n11185 27.0634
R36954 vss.n11189 vss.n11188 27.0634
R36955 vss.n11190 vss.n11189 27.0634
R36956 vss.n11190 vss.n11183 27.0634
R36957 vss.n11194 vss.n11183 27.0634
R36958 vss.n11335 vss.n11334 27.0634
R36959 vss.n11336 vss.n11335 27.0634
R36960 vss.n11336 vss.n11331 27.0634
R36961 vss.n11340 vss.n11331 27.0634
R36962 vss.n11341 vss.n11340 27.0634
R36963 vss.n11344 vss.n11341 27.0634
R36964 vss.n13055 vss.n13054 26.0995
R36965 vss.n14040 vss.n14039 23.9548
R36966 vss.n14044 vss.n14040 23.9548
R36967 vss.n14044 vss.n14043 23.9548
R36968 vss.n14057 vss.n14056 23.9548
R36969 vss.n14056 vss.n506 23.9548
R36970 vss.n14039 vss.n506 23.9548
R36971 vss.n1599 vss.n1574 23.9548
R36972 vss.n1599 vss.n1598 23.9548
R36973 vss.n1598 vss.n1589 23.9548
R36974 vss.n1585 vss.n1576 23.9548
R36975 vss.n1586 vss.n1585 23.9548
R36976 vss.n1586 vss.n1574 23.9548
R36977 vss.n1304 vss.n1279 23.9548
R36978 vss.n1304 vss.n1303 23.9548
R36979 vss.n1303 vss.n1294 23.9548
R36980 vss.n1290 vss.n1281 23.9548
R36981 vss.n1291 vss.n1290 23.9548
R36982 vss.n1291 vss.n1279 23.9548
R36983 vss.n1043 vss.n1018 23.9548
R36984 vss.n1043 vss.n1042 23.9548
R36985 vss.n1042 vss.n1033 23.9548
R36986 vss.n1029 vss.n1020 23.9548
R36987 vss.n1030 vss.n1029 23.9548
R36988 vss.n1030 vss.n1018 23.9548
R36989 vss.n1436 vss.n1411 23.9548
R36990 vss.n1436 vss.n1435 23.9548
R36991 vss.n1435 vss.n1426 23.9548
R36992 vss.n1422 vss.n1413 23.9548
R36993 vss.n1423 vss.n1422 23.9548
R36994 vss.n1423 vss.n1411 23.9548
R36995 vss.n1516 vss.n1491 23.9548
R36996 vss.n1516 vss.n1515 23.9548
R36997 vss.n1515 vss.n1506 23.9548
R36998 vss.n1502 vss.n1493 23.9548
R36999 vss.n1503 vss.n1502 23.9548
R37000 vss.n1503 vss.n1491 23.9548
R37001 vss.n958 vss.n939 23.9548
R37002 vss.n958 vss.n957 23.9548
R37003 vss.n957 vss.n948 23.9548
R37004 vss.n944 vss.n943 23.9548
R37005 vss.n945 vss.n944 23.9548
R37006 vss.n945 vss.n939 23.9548
R37007 vss.n1010 vss.n991 23.9548
R37008 vss.n1010 vss.n1009 23.9548
R37009 vss.n1009 vss.n1000 23.9548
R37010 vss.n996 vss.n995 23.9548
R37011 vss.n997 vss.n996 23.9548
R37012 vss.n997 vss.n991 23.9548
R37013 vss.n6238 vss.n6233 23.9548
R37014 vss.n6246 vss.n6233 23.9548
R37015 vss.n6246 vss.n6245 23.9548
R37016 vss.n6236 vss.n6227 23.9548
R37017 vss.n6239 vss.n6236 23.9548
R37018 vss.n6239 vss.n6238 23.9548
R37019 vss.n6626 vss.n6598 23.9548
R37020 vss.n6601 vss.n6598 23.9548
R37021 vss.n6619 vss.n6601 23.9548
R37022 vss.n6605 vss.n6599 23.9548
R37023 vss.n6625 vss.n6599 23.9548
R37024 vss.n6626 vss.n6625 23.9548
R37025 vss.n6399 vss.n6371 23.9548
R37026 vss.n6374 vss.n6371 23.9548
R37027 vss.n6392 vss.n6374 23.9548
R37028 vss.n6378 vss.n6372 23.9548
R37029 vss.n6398 vss.n6372 23.9548
R37030 vss.n6399 vss.n6398 23.9548
R37031 vss.n9267 vss.n9262 23.9548
R37032 vss.n9275 vss.n9262 23.9548
R37033 vss.n9275 vss.n9274 23.9548
R37034 vss.n9265 vss.n6322 23.9548
R37035 vss.n9268 vss.n9265 23.9548
R37036 vss.n9268 vss.n9267 23.9548
R37037 vss.n6935 vss.n6907 23.9548
R37038 vss.n6910 vss.n6907 23.9548
R37039 vss.n6928 vss.n6910 23.9548
R37040 vss.n6914 vss.n6908 23.9548
R37041 vss.n6934 vss.n6908 23.9548
R37042 vss.n6935 vss.n6934 23.9548
R37043 vss.n7124 vss.n7096 23.9548
R37044 vss.n7099 vss.n7096 23.9548
R37045 vss.n7117 vss.n7099 23.9548
R37046 vss.n7103 vss.n7097 23.9548
R37047 vss.n7123 vss.n7097 23.9548
R37048 vss.n7124 vss.n7123 23.9548
R37049 vss.n6276 vss.n6271 23.9548
R37050 vss.n6284 vss.n6271 23.9548
R37051 vss.n6284 vss.n6283 23.9548
R37052 vss.n6274 vss.n6264 23.9548
R37053 vss.n6277 vss.n6274 23.9548
R37054 vss.n6277 vss.n6276 23.9548
R37055 vss.n9292 vss.n6216 23.9548
R37056 vss.n9293 vss.n9292 23.9548
R37057 vss.n9296 vss.n9293 23.9548
R37058 vss.n9311 vss.n9307 23.9548
R37059 vss.n9311 vss.n9310 23.9548
R37060 vss.n9310 vss.n6216 23.9548
R37061 vss.n3313 vss.n3310 23.9548
R37062 vss.n3315 vss.n3313 23.9548
R37063 vss.n3322 vss.n3315 23.9548
R37064 vss.n3334 vss.n3333 23.9548
R37065 vss.n3333 vss.n3327 23.9548
R37066 vss.n3327 vss.n3310 23.9548
R37067 vss.n4315 vss.n4303 23.9548
R37068 vss.n4303 vss.n4302 23.9548
R37069 vss.n4302 vss.n4293 23.9548
R37070 vss.n4313 vss.n4304 23.9548
R37071 vss.n4314 vss.n4313 23.9548
R37072 vss.n4315 vss.n4314 23.9548
R37073 vss.n3670 vss.n3658 23.9548
R37074 vss.n3658 vss.n3657 23.9548
R37075 vss.n3657 vss.n3648 23.9548
R37076 vss.n3668 vss.n3659 23.9548
R37077 vss.n3669 vss.n3668 23.9548
R37078 vss.n3670 vss.n3669 23.9548
R37079 vss.n3450 vss.n3438 23.9548
R37080 vss.n3438 vss.n3437 23.9548
R37081 vss.n3437 vss.n3428 23.9548
R37082 vss.n3448 vss.n3439 23.9548
R37083 vss.n3449 vss.n3448 23.9548
R37084 vss.n3450 vss.n3449 23.9548
R37085 vss.n5877 vss.n5876 23.9548
R37086 vss.n5876 vss.n5875 23.9548
R37087 vss.n5875 vss.n5866 23.9548
R37088 vss.n5880 vss.n5879 23.9548
R37089 vss.n5879 vss.n5878 23.9548
R37090 vss.n5878 vss.n5877 23.9548
R37091 vss.n3376 vss.n3375 23.9548
R37092 vss.n3375 vss.n3374 23.9548
R37093 vss.n3374 vss.n3365 23.9548
R37094 vss.n5856 vss.n5855 23.9548
R37095 vss.n5855 vss.n3362 23.9548
R37096 vss.n3376 vss.n3362 23.9548
R37097 vss.n3972 vss.n3960 23.9548
R37098 vss.n3960 vss.n3959 23.9548
R37099 vss.n3959 vss.n3950 23.9548
R37100 vss.n3970 vss.n3961 23.9548
R37101 vss.n3971 vss.n3970 23.9548
R37102 vss.n3972 vss.n3971 23.9548
R37103 vss.n4239 vss.n4227 23.9548
R37104 vss.n4227 vss.n4226 23.9548
R37105 vss.n4226 vss.n4217 23.9548
R37106 vss.n4237 vss.n4228 23.9548
R37107 vss.n4238 vss.n4237 23.9548
R37108 vss.n4239 vss.n4238 23.9548
R37109 vss.n10396 vss.n10395 16.2531
R37110 vss.n10396 vss.n2033 16.2531
R37111 vss.n13147 vss.n2033 16.2531
R37112 vss.n13147 vss.n13146 16.2531
R37113 vss.n13146 vss.n2034 16.2531
R37114 vss.n2046 vss.n2034 16.2531
R37115 vss.n12638 vss.n12637 16.2531
R37116 vss.n12637 vss.n12622 16.2531
R37117 vss.n12661 vss.n12622 16.2531
R37118 vss.n12661 vss.n12660 16.2531
R37119 vss.n12660 vss.n12623 16.2531
R37120 vss.n12651 vss.n12623 16.2531
R37121 vss.n10392 vss.n10391 16.2531
R37122 vss.n10391 vss.n10375 16.2531
R37123 vss.n12695 vss.n10375 16.2531
R37124 vss.n12695 vss.n12694 16.2531
R37125 vss.n12694 vss.n10376 16.2531
R37126 vss.n12686 vss.n10376 16.2531
R37127 vss.n11423 vss.n11422 16.2531
R37128 vss.n11422 vss.n11406 16.2531
R37129 vss.n11445 vss.n11406 16.2531
R37130 vss.n11445 vss.n11444 16.2531
R37131 vss.n11444 vss.n11407 16.2531
R37132 vss.n11436 vss.n11407 16.2531
R37133 vss.n11376 vss.n11375 16.2531
R37134 vss.n11375 vss.n11359 16.2531
R37135 vss.n11398 vss.n11359 16.2531
R37136 vss.n11398 vss.n11397 16.2531
R37137 vss.n11397 vss.n11360 16.2531
R37138 vss.n11389 vss.n11360 16.2531
R37139 vss.n10951 vss.n10950 16.2531
R37140 vss.n10950 vss.n10934 16.2531
R37141 vss.n10973 vss.n10934 16.2531
R37142 vss.n10973 vss.n10972 16.2531
R37143 vss.n10972 vss.n10935 16.2531
R37144 vss.n10964 vss.n10935 16.2531
R37145 vss.n10788 vss.n10787 16.2531
R37146 vss.n10787 vss.n10771 16.2531
R37147 vss.n10810 vss.n10771 16.2531
R37148 vss.n10810 vss.n10809 16.2531
R37149 vss.n10809 vss.n10772 16.2531
R37150 vss.n10801 vss.n10772 16.2531
R37151 vss.n10744 vss.n10743 16.2531
R37152 vss.n10743 vss.n10727 16.2531
R37153 vss.n10766 vss.n10727 16.2531
R37154 vss.n10766 vss.n10765 16.2531
R37155 vss.n10765 vss.n10728 16.2531
R37156 vss.n10757 vss.n10728 16.2531
R37157 vss.n11570 vss.n11569 16.2531
R37158 vss.n11569 vss.n11553 16.2531
R37159 vss.n11592 vss.n11553 16.2531
R37160 vss.n11592 vss.n11591 16.2531
R37161 vss.n11591 vss.n11554 16.2531
R37162 vss.n11583 vss.n11554 16.2531
R37163 vss.n10567 vss.n10566 16.2531
R37164 vss.n10566 vss.n10550 16.2531
R37165 vss.n10589 vss.n10550 16.2531
R37166 vss.n10589 vss.n10588 16.2531
R37167 vss.n10588 vss.n10551 16.2531
R37168 vss.n10580 vss.n10551 16.2531
R37169 vss.n10523 vss.n10522 16.2531
R37170 vss.n10522 vss.n10506 16.2531
R37171 vss.n10545 vss.n10506 16.2531
R37172 vss.n10545 vss.n10544 16.2531
R37173 vss.n10544 vss.n10507 16.2531
R37174 vss.n10536 vss.n10507 16.2531
R37175 vss.n11944 vss.n11943 16.2531
R37176 vss.n11943 vss.n11927 16.2531
R37177 vss.n11966 vss.n11927 16.2531
R37178 vss.n11966 vss.n11965 16.2531
R37179 vss.n11965 vss.n11928 16.2531
R37180 vss.n11957 vss.n11928 16.2531
R37181 vss.n12062 vss.n12061 16.2531
R37182 vss.n12061 vss.n11893 16.2531
R37183 vss.n12073 vss.n11893 16.2531
R37184 vss.n12073 vss.n12072 16.2531
R37185 vss.n12072 vss.n11894 16.2531
R37186 vss.n11894 vss.n11853 16.2531
R37187 vss.n11908 vss.n11906 16.2531
R37188 vss.n11973 vss.n11906 16.2531
R37189 vss.n11973 vss.n11972 16.2531
R37190 vss.n11977 vss.n11972 16.2531
R37191 vss.n11978 vss.n11977 16.2531
R37192 vss.n11979 vss.n11978 16.2531
R37193 vss.n12022 vss.n12021 16.2531
R37194 vss.n12021 vss.n12020 16.2531
R37195 vss.n12020 vss.n12015 16.2531
R37196 vss.n12016 vss.n12015 16.2531
R37197 vss.n12016 vss.n11983 16.2531
R37198 vss.n12033 vss.n11983 16.2531
R37199 vss.n11996 vss.n11994 16.2531
R37200 vss.n11994 vss.n10592 16.2531
R37201 vss.n12609 vss.n10592 16.2531
R37202 vss.n12609 vss.n12608 16.2531
R37203 vss.n12608 vss.n10593 16.2531
R37204 vss.n10605 vss.n10593 16.2531
R37205 vss.n10650 vss.n10645 16.2531
R37206 vss.n10655 vss.n10650 16.2531
R37207 vss.n10658 vss.n10655 16.2531
R37208 vss.n10658 vss.n10657 16.2531
R37209 vss.n10657 vss.n10609 16.2531
R37210 vss.n10612 vss.n10609 16.2531
R37211 vss.n10641 vss.n10631 16.2531
R37212 vss.n10678 vss.n10631 16.2531
R37213 vss.n11598 vss.n10678 16.2531
R37214 vss.n11600 vss.n11598 16.2531
R37215 vss.n11600 vss.n11599 16.2531
R37216 vss.n11599 vss.n10625 16.2531
R37217 vss.n10840 vss.n10832 16.2531
R37218 vss.n10849 vss.n10840 16.2531
R37219 vss.n10849 vss.n10848 16.2531
R37220 vss.n10848 vss.n10847 16.2531
R37221 vss.n10847 vss.n10845 16.2531
R37222 vss.n10845 vss.n10618 16.2531
R37223 vss.n10829 vss.n10828 16.2531
R37224 vss.n10828 vss.n10813 16.2531
R37225 vss.n11538 vss.n10813 16.2531
R37226 vss.n11538 vss.n11537 16.2531
R37227 vss.n11537 vss.n10814 16.2531
R37228 vss.n10871 vss.n10814 16.2531
R37229 vss.n11507 vss.n11506 16.2531
R37230 vss.n11506 vss.n11505 16.2531
R37231 vss.n11505 vss.n11500 16.2531
R37232 vss.n11501 vss.n11500 16.2531
R37233 vss.n11501 vss.n10875 16.2531
R37234 vss.n11518 vss.n10875 16.2531
R37235 vss.n10887 vss.n10885 16.2531
R37236 vss.n10977 vss.n10885 16.2531
R37237 vss.n10987 vss.n10977 16.2531
R37238 vss.n10987 vss.n10986 16.2531
R37239 vss.n10986 vss.n10979 16.2531
R37240 vss.n10979 vss.n10978 16.2531
R37241 vss.n11459 vss.n11458 16.2531
R37242 vss.n11458 vss.n11457 16.2531
R37243 vss.n11457 vss.n11452 16.2531
R37244 vss.n11453 vss.n11452 16.2531
R37245 vss.n11453 vss.n10901 16.2531
R37246 vss.n11470 vss.n10901 16.2531
R37247 vss.n10916 vss.n10914 16.2531
R37248 vss.n10914 vss.n10338 16.2531
R37249 vss.n12741 vss.n10338 16.2531
R37250 vss.n12743 vss.n12741 16.2531
R37251 vss.n12743 vss.n12742 16.2531
R37252 vss.n12742 vss.n10332 16.2531
R37253 vss.n12727 vss.n12726 16.2531
R37254 vss.n12726 vss.n10342 16.2531
R37255 vss.n12738 vss.n10342 16.2531
R37256 vss.n12738 vss.n12737 16.2531
R37257 vss.n12737 vss.n10343 16.2531
R37258 vss.n10343 vss.n10325 16.2531
R37259 vss.n10357 vss.n10355 16.2531
R37260 vss.n12702 vss.n10355 16.2531
R37261 vss.n12702 vss.n12701 16.2531
R37262 vss.n12706 vss.n12701 16.2531
R37263 vss.n12707 vss.n12706 16.2531
R37264 vss.n12708 vss.n12707 16.2531
R37265 vss.n2258 vss.n2257 16.2531
R37266 vss.n2257 vss.n2242 16.2531
R37267 vss.n13017 vss.n2242 16.2531
R37268 vss.n13017 vss.n13016 16.2531
R37269 vss.n13016 vss.n2243 16.2531
R37270 vss.n13008 vss.n2243 16.2531
R37271 vss.n2300 vss.n2299 16.2531
R37272 vss.n2299 vss.n2298 16.2531
R37273 vss.n2298 vss.n2266 16.2531
R37274 vss.n2281 vss.n2266 16.2531
R37275 vss.n2288 vss.n2281 16.2531
R37276 vss.n2288 vss.n2287 16.2531
R37277 vss.n13109 vss.n13108 16.2531
R37278 vss.n13108 vss.n13107 16.2531
R37279 vss.n13107 vss.n2077 16.2531
R37280 vss.n2092 vss.n2077 16.2531
R37281 vss.n13097 vss.n2092 16.2531
R37282 vss.n13097 vss.n13096 16.2531
R37283 vss.n1112 vss.n1111 16.2531
R37284 vss.n1111 vss.n1096 16.2531
R37285 vss.n1135 vss.n1096 16.2531
R37286 vss.n1135 vss.n1134 16.2531
R37287 vss.n1134 vss.n1097 16.2531
R37288 vss.n1125 vss.n1097 16.2531
R37289 vss.n852 vss.n836 16.2531
R37290 vss.n853 vss.n852 16.2531
R37291 vss.n853 vss.n516 16.2531
R37292 vss.n857 vss.n516 16.2531
R37293 vss.n858 vss.n857 16.2531
R37294 vss.n859 vss.n858 16.2531
R37295 vss.n14160 vss.n14159 16.2531
R37296 vss.n14161 vss.n14160 16.2531
R37297 vss.n14161 vss.n438 16.2531
R37298 vss.n14170 vss.n438 16.2531
R37299 vss.n14171 vss.n14170 16.2531
R37300 vss.n14172 vss.n14171 16.2531
R37301 vss.n186 vss.n185 16.2531
R37302 vss.n185 vss.n2 16.2531
R37303 vss.n14792 vss.n2 16.2531
R37304 vss.n14792 vss.n14791 16.2531
R37305 vss.n14791 vss.n3 16.2531
R37306 vss.n16 vss.n3 16.2531
R37307 vss.n334 vss.n333 16.2531
R37308 vss.n333 vss.n318 16.2531
R37309 vss.n358 vss.n318 16.2531
R37310 vss.n358 vss.n357 16.2531
R37311 vss.n357 vss.n319 16.2531
R37312 vss.n349 vss.n319 16.2531
R37313 vss.n14217 vss.n14216 16.2531
R37314 vss.n14216 vss.n14215 16.2531
R37315 vss.n14215 vss.n14183 16.2531
R37316 vss.n14198 vss.n14183 16.2531
R37317 vss.n14205 vss.n14198 16.2531
R37318 vss.n14205 vss.n14204 16.2531
R37319 vss.n14113 vss.n14112 16.2531
R37320 vss.n14112 vss.n14097 16.2531
R37321 vss.n14137 vss.n14097 16.2531
R37322 vss.n14137 vss.n14136 16.2531
R37323 vss.n14136 vss.n14098 16.2531
R37324 vss.n14128 vss.n14098 16.2531
R37325 vss.n431 vss.n430 16.2531
R37326 vss.n430 vss.n415 16.2531
R37327 vss.n14246 vss.n415 16.2531
R37328 vss.n14246 vss.n14245 16.2531
R37329 vss.n14245 vss.n416 16.2531
R37330 vss.n14237 vss.n416 16.2531
R37331 vss.n471 vss.n470 16.2531
R37332 vss.n14147 vss.n471 16.2531
R37333 vss.n14147 vss.n14146 16.2531
R37334 vss.n14146 vss.n474 16.2531
R37335 vss.n13578 vss.n474 16.2531
R37336 vss.n13579 vss.n13578 16.2531
R37337 vss.n13605 vss.n13604 16.2531
R37338 vss.n13604 vss.n13603 16.2531
R37339 vss.n13603 vss.n13552 16.2531
R37340 vss.n13585 vss.n13552 16.2531
R37341 vss.n13593 vss.n13585 16.2531
R37342 vss.n13593 vss.n13592 16.2531
R37343 vss.n14680 vss.n14679 16.2531
R37344 vss.n14679 vss.n14678 16.2531
R37345 vss.n14678 vss.n14646 16.2531
R37346 vss.n14661 vss.n14646 16.2531
R37347 vss.n14668 vss.n14661 16.2531
R37348 vss.n14668 vss.n14667 16.2531
R37349 vss.n249 vss.n248 16.2531
R37350 vss.n248 vss.n233 16.2531
R37351 vss.n14560 vss.n233 16.2531
R37352 vss.n14560 vss.n14559 16.2531
R37353 vss.n14559 vss.n234 16.2531
R37354 vss.n14551 vss.n234 16.2531
R37355 vss.n14485 vss.n14484 16.2531
R37356 vss.n14484 vss.n14483 16.2531
R37357 vss.n14483 vss.n14451 16.2531
R37358 vss.n14466 vss.n14451 16.2531
R37359 vss.n14473 vss.n14466 16.2531
R37360 vss.n14473 vss.n14472 16.2531
R37361 vss.n308 vss.n307 16.2531
R37362 vss.n307 vss.n292 16.2531
R37363 vss.n14365 vss.n292 16.2531
R37364 vss.n14365 vss.n14364 16.2531
R37365 vss.n14364 vss.n293 16.2531
R37366 vss.n14356 vss.n293 16.2531
R37367 vss.n14290 vss.n14289 16.2531
R37368 vss.n14289 vss.n14288 16.2531
R37369 vss.n14288 vss.n14256 16.2531
R37370 vss.n14271 vss.n14256 16.2531
R37371 vss.n14278 vss.n14271 16.2531
R37372 vss.n14278 vss.n14277 16.2531
R37373 vss.n14336 vss.n14335 16.2531
R37374 vss.n14335 vss.n14334 16.2531
R37375 vss.n14334 vss.n14302 16.2531
R37376 vss.n14317 vss.n14302 16.2531
R37377 vss.n14324 vss.n14317 16.2531
R37378 vss.n14324 vss.n14323 16.2531
R37379 vss.n14387 vss.n14386 16.2531
R37380 vss.n14386 vss.n14371 16.2531
R37381 vss.n14411 vss.n14371 16.2531
R37382 vss.n14411 vss.n14410 16.2531
R37383 vss.n14410 vss.n14372 16.2531
R37384 vss.n14402 vss.n14372 16.2531
R37385 vss.n14531 vss.n14530 16.2531
R37386 vss.n14530 vss.n14529 16.2531
R37387 vss.n14529 vss.n14497 16.2531
R37388 vss.n14512 vss.n14497 16.2531
R37389 vss.n14519 vss.n14512 16.2531
R37390 vss.n14519 vss.n14518 16.2531
R37391 vss.n14582 vss.n14581 16.2531
R37392 vss.n14581 vss.n14566 16.2531
R37393 vss.n14606 vss.n14566 16.2531
R37394 vss.n14606 vss.n14605 16.2531
R37395 vss.n14605 vss.n14567 16.2531
R37396 vss.n14597 vss.n14567 16.2531
R37397 vss.n14726 vss.n14725 16.2531
R37398 vss.n14725 vss.n14724 16.2531
R37399 vss.n14724 vss.n14692 16.2531
R37400 vss.n14707 vss.n14692 16.2531
R37401 vss.n14714 vss.n14707 16.2531
R37402 vss.n14714 vss.n14713 16.2531
R37403 vss.n172 vss.n171 16.2531
R37404 vss.n171 vss.n156 16.2531
R37405 vss.n14755 vss.n156 16.2531
R37406 vss.n14755 vss.n14754 16.2531
R37407 vss.n14754 vss.n157 16.2531
R37408 vss.n14746 vss.n157 16.2531
R37409 vss.n13315 vss.n13314 16.2531
R37410 vss.n13913 vss.n13315 16.2531
R37411 vss.n13913 vss.n13912 16.2531
R37412 vss.n13912 vss.n13911 16.2531
R37413 vss.n13911 vss.n13321 16.2531
R37414 vss.n13323 vss.n13321 16.2531
R37415 vss.n13878 vss.n13877 16.2531
R37416 vss.n13879 vss.n13878 16.2531
R37417 vss.n13879 vss.n13330 16.2531
R37418 vss.n13892 vss.n13330 16.2531
R37419 vss.n13893 vss.n13892 16.2531
R37420 vss.n13894 vss.n13893 16.2531
R37421 vss.n13357 vss.n13356 16.2531
R37422 vss.n13865 vss.n13357 16.2531
R37423 vss.n13865 vss.n13864 16.2531
R37424 vss.n13864 vss.n13856 16.2531
R37425 vss.n13856 vss.n13360 16.2531
R37426 vss.n13362 vss.n13360 16.2531
R37427 vss.n13824 vss.n13823 16.2531
R37428 vss.n13825 vss.n13824 16.2531
R37429 vss.n13825 vss.n13371 16.2531
R37430 vss.n13838 vss.n13371 16.2531
R37431 vss.n13839 vss.n13838 16.2531
R37432 vss.n13840 vss.n13839 16.2531
R37433 vss.n13398 vss.n13397 16.2531
R37434 vss.n13811 vss.n13398 16.2531
R37435 vss.n13811 vss.n13810 16.2531
R37436 vss.n13810 vss.n13806 16.2531
R37437 vss.n13806 vss.n13401 16.2531
R37438 vss.n13403 vss.n13401 16.2531
R37439 vss.n13773 vss.n13772 16.2531
R37440 vss.n13774 vss.n13773 16.2531
R37441 vss.n13774 vss.n13410 16.2531
R37442 vss.n13787 vss.n13410 16.2531
R37443 vss.n13788 vss.n13787 16.2531
R37444 vss.n13789 vss.n13788 16.2531
R37445 vss.n13437 vss.n13436 16.2531
R37446 vss.n13760 vss.n13437 16.2531
R37447 vss.n13760 vss.n13759 16.2531
R37448 vss.n13759 vss.n13751 16.2531
R37449 vss.n13751 vss.n13440 16.2531
R37450 vss.n13442 vss.n13440 16.2531
R37451 vss.n13719 vss.n13718 16.2531
R37452 vss.n13720 vss.n13719 16.2531
R37453 vss.n13720 vss.n13451 16.2531
R37454 vss.n13733 vss.n13451 16.2531
R37455 vss.n13734 vss.n13733 16.2531
R37456 vss.n13735 vss.n13734 16.2531
R37457 vss.n13478 vss.n13477 16.2531
R37458 vss.n13706 vss.n13478 16.2531
R37459 vss.n13706 vss.n13705 16.2531
R37460 vss.n13705 vss.n13701 16.2531
R37461 vss.n13701 vss.n13481 16.2531
R37462 vss.n13483 vss.n13481 16.2531
R37463 vss.n13668 vss.n13667 16.2531
R37464 vss.n13669 vss.n13668 16.2531
R37465 vss.n13669 vss.n13490 16.2531
R37466 vss.n13682 vss.n13490 16.2531
R37467 vss.n13683 vss.n13682 16.2531
R37468 vss.n13684 vss.n13683 16.2531
R37469 vss.n13517 vss.n13516 16.2531
R37470 vss.n13655 vss.n13517 16.2531
R37471 vss.n13655 vss.n13654 16.2531
R37472 vss.n13654 vss.n13646 16.2531
R37473 vss.n13646 vss.n13520 16.2531
R37474 vss.n13522 vss.n13520 16.2531
R37475 vss.n13614 vss.n13613 16.2531
R37476 vss.n13615 vss.n13614 16.2531
R37477 vss.n13615 vss.n13531 16.2531
R37478 vss.n13628 vss.n13531 16.2531
R37479 vss.n13629 vss.n13628 16.2531
R37480 vss.n13630 vss.n13629 16.2531
R37481 vss.n632 vss.n622 16.2531
R37482 vss.n640 vss.n622 16.2531
R37483 vss.n644 vss.n640 16.2531
R37484 vss.n646 vss.n644 16.2531
R37485 vss.n646 vss.n645 16.2531
R37486 vss.n645 vss.n616 16.2531
R37487 vss.n811 vss.n810 16.2531
R37488 vss.n810 vss.n795 16.2531
R37489 vss.n13234 vss.n795 16.2531
R37490 vss.n13234 vss.n13233 16.2531
R37491 vss.n13233 vss.n796 16.2531
R37492 vss.n13224 vss.n796 16.2531
R37493 vss.n1670 vss.n1669 16.2531
R37494 vss.n1669 vss.n1654 16.2531
R37495 vss.n1693 vss.n1654 16.2531
R37496 vss.n1693 vss.n1692 16.2531
R37497 vss.n1692 vss.n1655 16.2531
R37498 vss.n1683 vss.n1655 16.2531
R37499 vss.n1623 vss.n1622 16.2531
R37500 vss.n1622 vss.n1607 16.2531
R37501 vss.n1646 vss.n1607 16.2531
R37502 vss.n1646 vss.n1645 16.2531
R37503 vss.n1645 vss.n1608 16.2531
R37504 vss.n1636 vss.n1608 16.2531
R37505 vss.n1375 vss.n1374 16.2531
R37506 vss.n1374 vss.n1359 16.2531
R37507 vss.n1398 vss.n1359 16.2531
R37508 vss.n1398 vss.n1397 16.2531
R37509 vss.n1397 vss.n1360 16.2531
R37510 vss.n1388 vss.n1360 16.2531
R37511 vss.n1176 vss.n1175 16.2531
R37512 vss.n1175 vss.n1160 16.2531
R37513 vss.n1199 vss.n1160 16.2531
R37514 vss.n1199 vss.n1198 16.2531
R37515 vss.n1198 vss.n1161 16.2531
R37516 vss.n1189 vss.n1161 16.2531
R37517 vss.n1328 vss.n1327 16.2531
R37518 vss.n1327 vss.n1312 16.2531
R37519 vss.n1351 vss.n1312 16.2531
R37520 vss.n1351 vss.n1350 16.2531
R37521 vss.n1350 vss.n1313 16.2531
R37522 vss.n1341 vss.n1313 16.2531
R37523 vss.n1067 vss.n1066 16.2531
R37524 vss.n1066 vss.n1051 16.2531
R37525 vss.n1090 vss.n1051 16.2531
R37526 vss.n1090 vss.n1089 16.2531
R37527 vss.n1089 vss.n1052 16.2531
R37528 vss.n1080 vss.n1052 16.2531
R37529 vss.n1460 vss.n1459 16.2531
R37530 vss.n1459 vss.n1444 16.2531
R37531 vss.n1483 vss.n1444 16.2531
R37532 vss.n1483 vss.n1482 16.2531
R37533 vss.n1482 vss.n1445 16.2531
R37534 vss.n1473 vss.n1445 16.2531
R37535 vss.n1540 vss.n1539 16.2531
R37536 vss.n1539 vss.n1524 16.2531
R37537 vss.n1564 vss.n1524 16.2531
R37538 vss.n1564 vss.n1563 16.2531
R37539 vss.n1563 vss.n1525 16.2531
R37540 vss.n1553 vss.n1525 16.2531
R37541 vss.n820 vss.n819 16.2531
R37542 vss.n820 vss.n596 16.2531
R37543 vss.n13952 vss.n596 16.2531
R37544 vss.n13952 vss.n13951 16.2531
R37545 vss.n13951 vss.n597 16.2531
R37546 vss.n609 vss.n597 16.2531
R37547 vss.n896 vss.n877 16.2531
R37548 vss.n897 vss.n896 16.2531
R37549 vss.n897 vss.n892 16.2531
R37550 vss.n901 vss.n892 16.2531
R37551 vss.n902 vss.n901 16.2531
R37552 vss.n903 vss.n902 16.2531
R37553 vss.n535 vss.n534 16.2531
R37554 vss.n534 vss.n518 16.2531
R37555 vss.n14024 vss.n518 16.2531
R37556 vss.n14024 vss.n14023 16.2531
R37557 vss.n14023 vss.n519 16.2531
R37558 vss.n14015 vss.n519 16.2531
R37559 vss.n549 vss.n539 16.2531
R37560 vss.n13993 vss.n549 16.2531
R37561 vss.n13993 vss.n13992 16.2531
R37562 vss.n13992 vss.n552 16.2531
R37563 vss.n663 vss.n552 16.2531
R37564 vss.n663 vss.n662 16.2531
R37565 vss.n574 vss.n573 16.2531
R37566 vss.n573 vss.n557 16.2531
R37567 vss.n13989 vss.n557 16.2531
R37568 vss.n13989 vss.n13988 16.2531
R37569 vss.n13988 vss.n558 16.2531
R37570 vss.n13980 vss.n558 16.2531
R37571 vss.n588 vss.n578 16.2531
R37572 vss.n13958 vss.n588 16.2531
R37573 vss.n13958 vss.n13957 16.2531
R37574 vss.n13957 vss.n591 16.2531
R37575 vss.n766 vss.n591 16.2531
R37576 vss.n766 vss.n765 16.2531
R37577 vss.n755 vss.n745 16.2531
R37578 vss.n13241 vss.n755 16.2531
R37579 vss.n13241 vss.n13240 16.2531
R37580 vss.n13240 vss.n792 16.2531
R37581 vss.n792 vss.n758 16.2531
R37582 vss.n784 vss.n758 16.2531
R37583 vss.n1729 vss.n1719 16.2531
R37584 vss.n1737 vss.n1719 16.2531
R37585 vss.n1738 vss.n1737 16.2531
R37586 vss.n1740 vss.n1738 16.2531
R37587 vss.n1740 vss.n1739 16.2531
R37588 vss.n1739 vss.n1709 16.2531
R37589 vss.n1761 vss.n1760 16.2531
R37590 vss.n1760 vss.n1699 16.2531
R37591 vss.n1801 vss.n1699 16.2531
R37592 vss.n1801 vss.n1800 16.2531
R37593 vss.n1800 vss.n1700 16.2531
R37594 vss.n1792 vss.n1700 16.2531
R37595 vss.n1765 vss.n1764 16.2531
R37596 vss.n1765 vss.n1276 16.2531
R37597 vss.n1809 vss.n1276 16.2531
R37598 vss.n1811 vss.n1809 16.2531
R37599 vss.n1811 vss.n1810 16.2531
R37600 vss.n1810 vss.n1266 16.2531
R37601 vss.n1252 vss.n1234 16.2531
R37602 vss.n1252 vss.n1237 16.2531
R37603 vss.n1245 vss.n1237 16.2531
R37604 vss.n1825 vss.n1245 16.2531
R37605 vss.n1825 vss.n1824 16.2531
R37606 vss.n1824 vss.n1823 16.2531
R37607 vss.n1833 vss.n1223 16.2531
R37608 vss.n1841 vss.n1223 16.2531
R37609 vss.n1842 vss.n1841 16.2531
R37610 vss.n1844 vss.n1842 16.2531
R37611 vss.n1844 vss.n1843 16.2531
R37612 vss.n1843 vss.n1213 16.2531
R37613 vss.n1865 vss.n1864 16.2531
R37614 vss.n1864 vss.n1203 16.2531
R37615 vss.n1905 vss.n1203 16.2531
R37616 vss.n1905 vss.n1904 16.2531
R37617 vss.n1904 vss.n1204 16.2531
R37618 vss.n1896 vss.n1204 16.2531
R37619 vss.n1869 vss.n1868 16.2531
R37620 vss.n1869 vss.n1158 16.2531
R37621 vss.n1913 vss.n1158 16.2531
R37622 vss.n1915 vss.n1913 16.2531
R37623 vss.n1915 vss.n1914 16.2531
R37624 vss.n1914 vss.n1148 16.2531
R37625 vss.n1936 vss.n1935 16.2531
R37626 vss.n1935 vss.n1138 16.2531
R37627 vss.n1976 vss.n1138 16.2531
R37628 vss.n1976 vss.n1975 16.2531
R37629 vss.n1975 vss.n1139 16.2531
R37630 vss.n1967 vss.n1139 16.2531
R37631 vss.n1940 vss.n1939 16.2531
R37632 vss.n1940 vss.n704 16.2531
R37633 vss.n13291 vss.n704 16.2531
R37634 vss.n13293 vss.n13291 16.2531
R37635 vss.n13293 vss.n13292 16.2531
R37636 vss.n13292 vss.n692 16.2531
R37637 vss.n727 vss.n726 16.2531
R37638 vss.n726 vss.n708 16.2531
R37639 vss.n13288 vss.n708 16.2531
R37640 vss.n13288 vss.n13287 16.2531
R37641 vss.n13287 vss.n709 16.2531
R37642 vss.n13279 vss.n709 16.2531
R37643 vss.n2002 vss.n2001 16.2531
R37644 vss.n2001 vss.n1986 16.2531
R37645 vss.n2025 vss.n1986 16.2531
R37646 vss.n2025 vss.n2024 16.2531
R37647 vss.n2024 vss.n1987 16.2531
R37648 vss.n2015 vss.n1987 16.2531
R37649 vss.n13176 vss.n13175 16.2531
R37650 vss.n13175 vss.n13160 16.2531
R37651 vss.n13199 vss.n13160 16.2531
R37652 vss.n13199 vss.n13198 16.2531
R37653 vss.n13198 vss.n13161 16.2531
R37654 vss.n13188 vss.n13161 16.2531
R37655 vss.n9603 vss.n9602 16.2531
R37656 vss.n9602 vss.n9587 16.2531
R37657 vss.n9627 vss.n9587 16.2531
R37658 vss.n9627 vss.n9626 16.2531
R37659 vss.n9626 vss.n9588 16.2531
R37660 vss.n9618 vss.n9588 16.2531
R37661 vss.n9167 vss.n9166 16.2531
R37662 vss.n9166 vss.n9151 16.2531
R37663 vss.n9191 vss.n9151 16.2531
R37664 vss.n9191 vss.n9190 16.2531
R37665 vss.n9190 vss.n9152 16.2531
R37666 vss.n9181 vss.n9152 16.2531
R37667 vss.n9464 vss.n9463 16.2531
R37668 vss.n9463 vss.n9454 16.2531
R37669 vss.n9454 vss.n6055 16.2531
R37670 vss.n9474 vss.n6055 16.2531
R37671 vss.n9474 vss.n9473 16.2531
R37672 vss.n9473 vss.n9447 16.2531
R37673 vss.n8043 vss.n8042 16.2531
R37674 vss.n8044 vss.n8043 16.2531
R37675 vss.n8044 vss.n6005 16.2531
R37676 vss.n8039 vss.n6005 16.2531
R37677 vss.n8039 vss.n8038 16.2531
R37678 vss.n8038 vss.n8037 16.2531
R37679 vss.n9665 vss.n9664 16.2531
R37680 vss.n9664 vss.n9663 16.2531
R37681 vss.n9663 vss.n5978 16.2531
R37682 vss.n5993 vss.n5978 16.2531
R37683 vss.n9653 vss.n5993 16.2531
R37684 vss.n9653 vss.n9652 16.2531
R37685 vss.n8149 vss.n6001 16.2531
R37686 vss.n9643 vss.n6001 16.2531
R37687 vss.n9643 vss.n9642 16.2531
R37688 vss.n9642 vss.n6003 16.2531
R37689 vss.n8133 vss.n6003 16.2531
R37690 vss.n8139 vss.n8133 16.2531
R37691 vss.n8158 vss.n8157 16.2531
R37692 vss.n8159 vss.n8158 16.2531
R37693 vss.n8159 vss.n8104 16.2531
R37694 vss.n8168 vss.n8104 16.2531
R37695 vss.n8169 vss.n8168 16.2531
R37696 vss.n8170 vss.n8169 16.2531
R37697 vss.n8084 vss.n8083 16.2531
R37698 vss.n8085 vss.n8084 16.2531
R37699 vss.n8085 vss.n8060 16.2531
R37700 vss.n8094 vss.n8060 16.2531
R37701 vss.n8095 vss.n8094 16.2531
R37702 vss.n8096 vss.n8095 16.2531
R37703 vss.n8009 vss.n8008 16.2531
R37704 vss.n8008 vss.n7993 16.2531
R37705 vss.n8244 vss.n7993 16.2531
R37706 vss.n8244 vss.n8243 16.2531
R37707 vss.n8243 vss.n7994 16.2531
R37708 vss.n8235 vss.n7994 16.2531
R37709 vss.n8215 vss.n8214 16.2531
R37710 vss.n8214 vss.n8213 16.2531
R37711 vss.n8213 vss.n8181 16.2531
R37712 vss.n8196 vss.n8181 16.2531
R37713 vss.n8203 vss.n8196 16.2531
R37714 vss.n8203 vss.n8202 16.2531
R37715 vss.n9003 vss.n9002 16.2531
R37716 vss.n9002 vss.n9001 16.2531
R37717 vss.n9001 vss.n7304 16.2531
R37718 vss.n7319 vss.n7304 16.2531
R37719 vss.n8991 vss.n7319 16.2531
R37720 vss.n8991 vss.n8990 16.2531
R37721 vss.n7866 vss.n7865 16.2531
R37722 vss.n7865 vss.n7850 16.2531
R37723 vss.n8735 vss.n7850 16.2531
R37724 vss.n8735 vss.n8734 16.2531
R37725 vss.n8734 vss.n7851 16.2531
R37726 vss.n8726 vss.n7851 16.2531
R37727 vss.n7785 vss.n7784 16.2531
R37728 vss.n7784 vss.n7769 16.2531
R37729 vss.n7809 vss.n7769 16.2531
R37730 vss.n7809 vss.n7808 16.2531
R37731 vss.n7808 vss.n7770 16.2531
R37732 vss.n7800 vss.n7770 16.2531
R37733 vss.n8779 vss.n8778 16.2531
R37734 vss.n8778 vss.n8777 16.2531
R37735 vss.n8777 vss.n8745 16.2531
R37736 vss.n8760 vss.n8745 16.2531
R37737 vss.n8767 vss.n8760 16.2531
R37738 vss.n8767 vss.n8766 16.2531
R37739 vss.n7679 vss.n7678 16.2531
R37740 vss.n7678 vss.n7663 16.2531
R37741 vss.n8854 vss.n7663 16.2531
R37742 vss.n8854 vss.n8853 16.2531
R37743 vss.n8853 vss.n7664 16.2531
R37744 vss.n8845 vss.n7664 16.2531
R37745 vss.n8825 vss.n8824 16.2531
R37746 vss.n8824 vss.n8823 16.2531
R37747 vss.n8823 vss.n8791 16.2531
R37748 vss.n8806 vss.n8791 16.2531
R37749 vss.n8813 vss.n8806 16.2531
R37750 vss.n8813 vss.n8812 16.2531
R37751 vss.n8898 vss.n8897 16.2531
R37752 vss.n8897 vss.n8896 16.2531
R37753 vss.n8896 vss.n8864 16.2531
R37754 vss.n8879 vss.n8864 16.2531
R37755 vss.n8886 vss.n8879 16.2531
R37756 vss.n8886 vss.n8885 16.2531
R37757 vss.n9034 vss.n9033 16.2531
R37758 vss.n9033 vss.n9032 16.2531
R37759 vss.n9032 vss.n7272 16.2531
R37760 vss.n7287 vss.n7272 16.2531
R37761 vss.n9022 vss.n7287 16.2531
R37762 vss.n9022 vss.n9021 16.2531
R37763 vss.n8279 vss.n8278 16.2531
R37764 vss.n8278 vss.n8277 16.2531
R37765 vss.n8277 vss.n8259 16.2531
R37766 vss.n8259 vss.n7294 16.2531
R37767 vss.n9013 vss.n7294 16.2531
R37768 vss.n9013 vss.n9012 16.2531
R37769 vss.n8288 vss.n8287 16.2531
R37770 vss.n8289 vss.n8288 16.2531
R37771 vss.n8289 vss.n7882 16.2531
R37772 vss.n8298 vss.n7882 16.2531
R37773 vss.n8299 vss.n8298 16.2531
R37774 vss.n8300 vss.n8299 16.2531
R37775 vss.n8694 vss.n8693 16.2531
R37776 vss.n8695 vss.n8694 16.2531
R37777 vss.n8695 vss.n7874 16.2531
R37778 vss.n8704 vss.n7874 16.2531
R37779 vss.n8705 vss.n8704 16.2531
R37780 vss.n8706 vss.n8705 16.2531
R37781 vss.n8684 vss.n8327 16.2531
R37782 vss.n8684 vss.n8683 16.2531
R37783 vss.n8683 vss.n8330 16.2531
R37784 vss.n8333 vss.n8330 16.2531
R37785 vss.n8346 vss.n8333 16.2531
R37786 vss.n8347 vss.n8346 16.2531
R37787 vss.n8648 vss.n8647 16.2531
R37788 vss.n8647 vss.n8355 16.2531
R37789 vss.n8355 vss.n8352 16.2531
R37790 vss.n8662 vss.n8352 16.2531
R37791 vss.n8669 vss.n8662 16.2531
R37792 vss.n8669 vss.n8668 16.2531
R37793 vss.n8641 vss.n8372 16.2531
R37794 vss.n8641 vss.n8640 16.2531
R37795 vss.n8640 vss.n8380 16.2531
R37796 vss.n8383 vss.n8380 16.2531
R37797 vss.n8396 vss.n8383 16.2531
R37798 vss.n8397 vss.n8396 16.2531
R37799 vss.n8604 vss.n8603 16.2531
R37800 vss.n8603 vss.n8408 16.2531
R37801 vss.n8408 vss.n8405 16.2531
R37802 vss.n8618 vss.n8405 16.2531
R37803 vss.n8626 vss.n8618 16.2531
R37804 vss.n8626 vss.n8625 16.2531
R37805 vss.n8597 vss.n8425 16.2531
R37806 vss.n8597 vss.n8596 16.2531
R37807 vss.n8596 vss.n8428 16.2531
R37808 vss.n8431 vss.n8428 16.2531
R37809 vss.n8444 vss.n8431 16.2531
R37810 vss.n8445 vss.n8444 16.2531
R37811 vss.n8561 vss.n8560 16.2531
R37812 vss.n8560 vss.n8453 16.2531
R37813 vss.n8453 vss.n8450 16.2531
R37814 vss.n8575 vss.n8450 16.2531
R37815 vss.n8582 vss.n8575 16.2531
R37816 vss.n8582 vss.n8581 16.2531
R37817 vss.n8554 vss.n8470 16.2531
R37818 vss.n8554 vss.n8553 16.2531
R37819 vss.n8553 vss.n8478 16.2531
R37820 vss.n8481 vss.n8478 16.2531
R37821 vss.n8494 vss.n8481 16.2531
R37822 vss.n8495 vss.n8494 16.2531
R37823 vss.n8526 vss.n8525 16.2531
R37824 vss.n8527 vss.n8526 16.2531
R37825 vss.n8527 vss.n8503 16.2531
R37826 vss.n8531 vss.n8503 16.2531
R37827 vss.n8539 vss.n8531 16.2531
R37828 vss.n8539 vss.n8538 16.2531
R37829 vss.n7490 vss.n7489 16.2531
R37830 vss.n7489 vss.n7474 16.2531
R37831 vss.n8973 vss.n7474 16.2531
R37832 vss.n8973 vss.n8972 16.2531
R37833 vss.n8972 vss.n7475 16.2531
R37834 vss.n8964 vss.n7475 16.2531
R37835 vss.n8944 vss.n8943 16.2531
R37836 vss.n8943 vss.n8942 16.2531
R37837 vss.n8942 vss.n8910 16.2531
R37838 vss.n8925 vss.n8910 16.2531
R37839 vss.n8932 vss.n8925 16.2531
R37840 vss.n8932 vss.n8931 16.2531
R37841 vss.n7532 vss.n7531 16.2531
R37842 vss.n7531 vss.n7530 16.2531
R37843 vss.n7530 vss.n7498 16.2531
R37844 vss.n7513 vss.n7498 16.2531
R37845 vss.n7520 vss.n7513 16.2531
R37846 vss.n7520 vss.n7519 16.2531
R37847 vss.n7562 vss.n7561 16.2531
R37848 vss.n7561 vss.n7546 16.2531
R37849 vss.n7586 vss.n7546 16.2531
R37850 vss.n7586 vss.n7585 16.2531
R37851 vss.n7585 vss.n7547 16.2531
R37852 vss.n7577 vss.n7547 16.2531
R37853 vss.n7705 vss.n7704 16.2531
R37854 vss.n7704 vss.n7689 16.2531
R37855 vss.n7729 vss.n7689 16.2531
R37856 vss.n7729 vss.n7728 16.2531
R37857 vss.n7728 vss.n7690 16.2531
R37858 vss.n7720 vss.n7690 16.2531
R37859 vss.n7926 vss.n7925 16.2531
R37860 vss.n7925 vss.n7910 16.2531
R37861 vss.n7950 vss.n7910 16.2531
R37862 vss.n7950 vss.n7949 16.2531
R37863 vss.n7949 vss.n7911 16.2531
R37864 vss.n7941 vss.n7911 16.2531
R37865 vss.n6025 vss.n6024 16.2531
R37866 vss.n6024 vss.n6009 16.2531
R37867 vss.n6050 vss.n6009 16.2531
R37868 vss.n6050 vss.n6049 16.2531
R37869 vss.n6049 vss.n6010 16.2531
R37870 vss.n6039 vss.n6010 16.2531
R37871 vss.n7195 vss.n7194 16.2531
R37872 vss.n7194 vss.n7179 16.2531
R37873 vss.n7219 vss.n7179 16.2531
R37874 vss.n7219 vss.n7218 16.2531
R37875 vss.n7218 vss.n7180 16.2531
R37876 vss.n7209 vss.n7180 16.2531
R37877 vss.n6690 vss.n6689 16.2531
R37878 vss.n6689 vss.n6674 16.2531
R37879 vss.n6714 vss.n6674 16.2531
R37880 vss.n6714 vss.n6713 16.2531
R37881 vss.n6713 vss.n6675 16.2531
R37882 vss.n6704 vss.n6675 16.2531
R37883 vss.n6646 vss.n6645 16.2531
R37884 vss.n6645 vss.n6630 16.2531
R37885 vss.n6670 vss.n6630 16.2531
R37886 vss.n6670 vss.n6669 16.2531
R37887 vss.n6669 vss.n6631 16.2531
R37888 vss.n6660 vss.n6631 16.2531
R37889 vss.n7004 vss.n7003 16.2531
R37890 vss.n7003 vss.n6988 16.2531
R37891 vss.n7028 vss.n6988 16.2531
R37892 vss.n7028 vss.n7027 16.2531
R37893 vss.n7027 vss.n6989 16.2531
R37894 vss.n7018 vss.n6989 16.2531
R37895 vss.n6464 vss.n6463 16.2531
R37896 vss.n6463 vss.n6448 16.2531
R37897 vss.n6488 vss.n6448 16.2531
R37898 vss.n6488 vss.n6487 16.2531
R37899 vss.n6487 vss.n6449 16.2531
R37900 vss.n6478 vss.n6449 16.2531
R37901 vss.n6419 vss.n6418 16.2531
R37902 vss.n6418 vss.n6403 16.2531
R37903 vss.n6443 vss.n6403 16.2531
R37904 vss.n6443 vss.n6442 16.2531
R37905 vss.n6442 vss.n6404 16.2531
R37906 vss.n6433 vss.n6404 16.2531
R37907 vss.n6341 vss.n6340 16.2531
R37908 vss.n6340 vss.n6325 16.2531
R37909 vss.n6365 vss.n6325 16.2531
R37910 vss.n6365 vss.n6364 16.2531
R37911 vss.n6364 vss.n6326 16.2531
R37912 vss.n6355 vss.n6326 16.2531
R37913 vss.n6955 vss.n6954 16.2531
R37914 vss.n6954 vss.n6939 16.2531
R37915 vss.n6979 vss.n6939 16.2531
R37916 vss.n6979 vss.n6978 16.2531
R37917 vss.n6978 vss.n6940 16.2531
R37918 vss.n6969 vss.n6940 16.2531
R37919 vss.n7144 vss.n7143 16.2531
R37920 vss.n7143 vss.n7128 16.2531
R37921 vss.n7168 vss.n7128 16.2531
R37922 vss.n7168 vss.n7167 16.2531
R37923 vss.n7167 vss.n7129 16.2531
R37924 vss.n7158 vss.n7129 16.2531
R37925 vss.n6152 vss.n6151 16.2531
R37926 vss.n6151 vss.n6136 16.2531
R37927 vss.n9501 vss.n6136 16.2531
R37928 vss.n9501 vss.n9500 16.2531
R37929 vss.n9500 vss.n6137 16.2531
R37930 vss.n6166 vss.n6137 16.2531
R37931 vss.n9419 vss.n9408 16.2531
R37932 vss.n9427 vss.n9408 16.2531
R37933 vss.n9430 vss.n9427 16.2531
R37934 vss.n9432 vss.n9430 16.2531
R37935 vss.n9432 vss.n9431 16.2531
R37936 vss.n9431 vss.n9402 16.2531
R37937 vss.n6075 vss.n6074 16.2531
R37938 vss.n6074 vss.n6057 16.2531
R37939 vss.n9573 vss.n6057 16.2531
R37940 vss.n9573 vss.n9572 16.2531
R37941 vss.n9572 vss.n6058 16.2531
R37942 vss.n9564 vss.n6058 16.2531
R37943 vss.n6089 vss.n6079 16.2531
R37944 vss.n9542 vss.n6089 16.2531
R37945 vss.n9542 vss.n9541 16.2531
R37946 vss.n9541 vss.n6092 16.2531
R37947 vss.n7251 vss.n6092 16.2531
R37948 vss.n7251 vss.n7250 16.2531
R37949 vss.n6114 vss.n6113 16.2531
R37950 vss.n6113 vss.n6097 16.2531
R37951 vss.n9538 vss.n6097 16.2531
R37952 vss.n9538 vss.n9537 16.2531
R37953 vss.n9537 vss.n6098 16.2531
R37954 vss.n9529 vss.n6098 16.2531
R37955 vss.n6128 vss.n6118 16.2531
R37956 vss.n9507 vss.n6128 16.2531
R37957 vss.n9507 vss.n9506 16.2531
R37958 vss.n9506 vss.n6131 16.2531
R37959 vss.n6578 vss.n6131 16.2531
R37960 vss.n6578 vss.n6577 16.2531
R37961 vss.n6753 vss.n6750 16.2531
R37962 vss.n6753 vss.n6595 16.2531
R37963 vss.n7225 vss.n6595 16.2531
R37964 vss.n7227 vss.n7225 16.2531
R37965 vss.n7227 vss.n7226 16.2531
R37966 vss.n7226 vss.n6583 16.2531
R37967 vss.n6765 vss.n6739 16.2531
R37968 vss.n6773 vss.n6739 16.2531
R37969 vss.n6774 vss.n6773 16.2531
R37970 vss.n6776 vss.n6774 16.2531
R37971 vss.n6776 vss.n6775 16.2531
R37972 vss.n6775 vss.n6729 16.2531
R37973 vss.n6797 vss.n6796 16.2531
R37974 vss.n6796 vss.n6719 16.2531
R37975 vss.n7083 vss.n6719 16.2531
R37976 vss.n7083 vss.n7082 16.2531
R37977 vss.n7082 vss.n6720 16.2531
R37978 vss.n7074 vss.n6720 16.2531
R37979 vss.n6810 vss.n6800 16.2531
R37980 vss.n7052 vss.n6810 16.2531
R37981 vss.n7052 vss.n7051 16.2531
R37982 vss.n7051 vss.n7048 16.2531
R37983 vss.n7048 vss.n6813 16.2531
R37984 vss.n6819 vss.n6813 16.2531
R37985 vss.n6894 vss.n6841 16.2531
R37986 vss.n6902 vss.n6841 16.2531
R37987 vss.n7034 vss.n6902 16.2531
R37988 vss.n7036 vss.n7034 16.2531
R37989 vss.n7036 vss.n7035 16.2531
R37990 vss.n7035 vss.n6829 16.2531
R37991 vss.n6861 vss.n6851 16.2531
R37992 vss.n6884 vss.n6861 16.2531
R37993 vss.n6884 vss.n6883 16.2531
R37994 vss.n6883 vss.n6882 16.2531
R37995 vss.n6882 vss.n6864 16.2531
R37996 vss.n6870 vss.n6864 16.2531
R37997 vss.n6508 vss.n6507 16.2531
R37998 vss.n6507 vss.n6491 16.2531
R37999 vss.n9246 vss.n6491 16.2531
R38000 vss.n9246 vss.n9245 16.2531
R38001 vss.n9245 vss.n6492 16.2531
R38002 vss.n9237 vss.n6492 16.2531
R38003 vss.n6521 vss.n6511 16.2531
R38004 vss.n9215 vss.n6521 16.2531
R38005 vss.n9215 vss.n9214 16.2531
R38006 vss.n9214 vss.n9211 16.2531
R38007 vss.n9211 vss.n6524 16.2531
R38008 vss.n6560 vss.n6524 16.2531
R38009 vss.n9071 vss.n9068 16.2531
R38010 vss.n9071 vss.n6542 16.2531
R38011 vss.n9197 vss.n6542 16.2531
R38012 vss.n9199 vss.n9197 16.2531
R38013 vss.n9199 vss.n9198 16.2531
R38014 vss.n9198 vss.n6530 16.2531
R38015 vss.n9064 vss.n9063 16.2531
R38016 vss.n9063 vss.n6548 16.2531
R38017 vss.n9144 vss.n6548 16.2531
R38018 vss.n9144 vss.n9143 16.2531
R38019 vss.n9143 vss.n6549 16.2531
R38020 vss.n9053 vss.n6549 16.2531
R38021 vss.n9120 vss.n9112 16.2531
R38022 vss.n9128 vss.n9112 16.2531
R38023 vss.n9129 vss.n9128 16.2531
R38024 vss.n9131 vss.n9129 16.2531
R38025 vss.n9131 vss.n9130 16.2531
R38026 vss.n9130 vss.n9100 16.2531
R38027 vss.n9337 vss.n9336 16.2531
R38028 vss.n9336 vss.n9321 16.2531
R38029 vss.n9361 vss.n9321 16.2531
R38030 vss.n9361 vss.n9360 16.2531
R38031 vss.n9360 vss.n9322 16.2531
R38032 vss.n9351 vss.n9322 16.2531
R38033 vss.n6204 vss.n6193 16.2531
R38034 vss.n6212 vss.n6193 16.2531
R38035 vss.n9368 vss.n6212 16.2531
R38036 vss.n9370 vss.n9368 16.2531
R38037 vss.n9370 vss.n9369 16.2531
R38038 vss.n9369 vss.n6187 16.2531
R38039 vss.n5954 vss.n5953 16.2531
R38040 vss.n5953 vss.n5938 16.2531
R38041 vss.n9681 vss.n5938 16.2531
R38042 vss.n9681 vss.n9680 16.2531
R38043 vss.n9680 vss.n5939 16.2531
R38044 vss.n5968 vss.n5939 16.2531
R38045 vss.n9702 vss.n9701 16.2531
R38046 vss.n9701 vss.n9686 16.2531
R38047 vss.n9728 vss.n9686 16.2531
R38048 vss.n9728 vss.n9727 16.2531
R38049 vss.n9727 vss.n9687 16.2531
R38050 vss.n9718 vss.n9687 16.2531
R38051 vss.n2575 vss.n2574 16.2531
R38052 vss.n2574 vss.n2559 16.2531
R38053 vss.n10009 vss.n2559 16.2531
R38054 vss.n10009 vss.n10008 16.2531
R38055 vss.n10008 vss.n2560 16.2531
R38056 vss.n2589 vss.n2560 16.2531
R38057 vss.n9892 vss.n9891 16.2531
R38058 vss.n9891 vss.n9890 16.2531
R38059 vss.n9890 vss.n2748 16.2531
R38060 vss.n2763 vss.n2748 16.2531
R38061 vss.n9880 vss.n2763 16.2531
R38062 vss.n9880 vss.n9879 16.2531
R38063 vss.n3280 vss.n3279 16.2531
R38064 vss.n3279 vss.n3264 16.2531
R38065 vss.n3306 vss.n3264 16.2531
R38066 vss.n3306 vss.n3305 16.2531
R38067 vss.n3305 vss.n3265 16.2531
R38068 vss.n3297 vss.n3265 16.2531
R38069 vss.n9766 vss.n9765 16.2531
R38070 vss.n9765 vss.n9745 16.2531
R38071 vss.n9784 vss.n9745 16.2531
R38072 vss.n9784 vss.n9783 16.2531
R38073 vss.n9783 vss.n9746 16.2531
R38074 vss.n9779 vss.n9746 16.2531
R38075 vss.n3206 vss.n3205 16.2531
R38076 vss.n3205 vss.n3185 16.2531
R38077 vss.n3224 vss.n3185 16.2531
R38078 vss.n3224 vss.n3223 16.2531
R38079 vss.n3223 vss.n3186 16.2531
R38080 vss.n3219 vss.n3186 16.2531
R38081 vss.n3006 vss.n3005 16.2531
R38082 vss.n9795 vss.n3006 16.2531
R38083 vss.n9795 vss.n9794 16.2531
R38084 vss.n9794 vss.n3025 16.2531
R38085 vss.n3025 vss.n3009 16.2531
R38086 vss.n3021 vss.n3009 16.2531
R38087 vss.n5236 vss.n5235 16.2531
R38088 vss.n5235 vss.n5215 16.2531
R38089 vss.n5254 vss.n5215 16.2531
R38090 vss.n5254 vss.n5253 16.2531
R38091 vss.n5253 vss.n5216 16.2531
R38092 vss.n5249 vss.n5216 16.2531
R38093 vss.n3049 vss.n3048 16.2531
R38094 vss.n3048 vss.n3028 16.2531
R38095 vss.n3067 vss.n3028 16.2531
R38096 vss.n3067 vss.n3066 16.2531
R38097 vss.n3066 vss.n3029 16.2531
R38098 vss.n3062 vss.n3029 16.2531
R38099 vss.n5106 vss.n5105 16.2531
R38100 vss.n5105 vss.n5085 16.2531
R38101 vss.n5124 vss.n5085 16.2531
R38102 vss.n5124 vss.n5123 16.2531
R38103 vss.n5123 vss.n5086 16.2531
R38104 vss.n5119 vss.n5086 16.2531
R38105 vss.n5295 vss.n5294 16.2531
R38106 vss.n5294 vss.n5274 16.2531
R38107 vss.n5313 vss.n5274 16.2531
R38108 vss.n5313 vss.n5312 16.2531
R38109 vss.n5312 vss.n5275 16.2531
R38110 vss.n5308 vss.n5275 16.2531
R38111 vss.n5023 vss.n5022 16.2531
R38112 vss.n5022 vss.n5002 16.2531
R38113 vss.n5041 vss.n5002 16.2531
R38114 vss.n5041 vss.n5040 16.2531
R38115 vss.n5040 vss.n5003 16.2531
R38116 vss.n5036 vss.n5003 16.2531
R38117 vss.n4904 vss.n4903 16.2531
R38118 vss.n4903 vss.n4883 16.2531
R38119 vss.n4922 vss.n4883 16.2531
R38120 vss.n4922 vss.n4921 16.2531
R38121 vss.n4921 vss.n4884 16.2531
R38122 vss.n4917 vss.n4884 16.2531
R38123 vss.n9926 vss.n9925 16.2531
R38124 vss.n9925 vss.n9924 16.2531
R38125 vss.n9924 vss.n2713 16.2531
R38126 vss.n2728 vss.n2713 16.2531
R38127 vss.n9914 vss.n2728 16.2531
R38128 vss.n9914 vss.n9913 16.2531
R38129 vss.n4663 vss.n4662 16.2531
R38130 vss.n4662 vss.n4661 16.2531
R38131 vss.n4661 vss.n4643 16.2531
R38132 vss.n4643 vss.n2735 16.2531
R38133 vss.n9905 vss.n2735 16.2531
R38134 vss.n9905 vss.n9904 16.2531
R38135 vss.n5628 vss.n5627 16.2531
R38136 vss.n5627 vss.n5626 16.2531
R38137 vss.n5626 vss.n4634 16.2531
R38138 vss.n4680 vss.n4634 16.2531
R38139 vss.n5616 vss.n4680 16.2531
R38140 vss.n5616 vss.n5615 16.2531
R38141 vss.n5586 vss.n5585 16.2531
R38142 vss.n5585 vss.n4690 16.2531
R38143 vss.n4690 vss.n4687 16.2531
R38144 vss.n5600 vss.n4687 16.2531
R38145 vss.n5607 vss.n5600 16.2531
R38146 vss.n5607 vss.n5606 16.2531
R38147 vss.n5579 vss.n4707 16.2531
R38148 vss.n5579 vss.n5578 16.2531
R38149 vss.n5578 vss.n4708 16.2531
R38150 vss.n4711 vss.n4708 16.2531
R38151 vss.n4724 vss.n4711 16.2531
R38152 vss.n4725 vss.n4724 16.2531
R38153 vss.n5543 vss.n5542 16.2531
R38154 vss.n5542 vss.n4733 16.2531
R38155 vss.n4733 vss.n4730 16.2531
R38156 vss.n5557 vss.n4730 16.2531
R38157 vss.n5564 vss.n5557 16.2531
R38158 vss.n5564 vss.n5563 16.2531
R38159 vss.n5536 vss.n4750 16.2531
R38160 vss.n5536 vss.n5535 16.2531
R38161 vss.n5535 vss.n4751 16.2531
R38162 vss.n4754 vss.n4751 16.2531
R38163 vss.n4767 vss.n4754 16.2531
R38164 vss.n4768 vss.n4767 16.2531
R38165 vss.n5500 vss.n5499 16.2531
R38166 vss.n5499 vss.n4776 16.2531
R38167 vss.n4776 vss.n4773 16.2531
R38168 vss.n5514 vss.n4773 16.2531
R38169 vss.n5521 vss.n5514 16.2531
R38170 vss.n5521 vss.n5520 16.2531
R38171 vss.n5493 vss.n4793 16.2531
R38172 vss.n5493 vss.n5492 16.2531
R38173 vss.n5492 vss.n4794 16.2531
R38174 vss.n4797 vss.n4794 16.2531
R38175 vss.n4810 vss.n4797 16.2531
R38176 vss.n4811 vss.n4810 16.2531
R38177 vss.n5457 vss.n5456 16.2531
R38178 vss.n5456 vss.n4819 16.2531
R38179 vss.n4819 vss.n4816 16.2531
R38180 vss.n5471 vss.n4816 16.2531
R38181 vss.n5478 vss.n5471 16.2531
R38182 vss.n5478 vss.n5477 16.2531
R38183 vss.n5450 vss.n4836 16.2531
R38184 vss.n5450 vss.n5449 16.2531
R38185 vss.n5449 vss.n4837 16.2531
R38186 vss.n4840 vss.n4837 16.2531
R38187 vss.n4853 vss.n4840 16.2531
R38188 vss.n4854 vss.n4853 16.2531
R38189 vss.n5414 vss.n5413 16.2531
R38190 vss.n5413 vss.n4862 16.2531
R38191 vss.n4862 vss.n4859 16.2531
R38192 vss.n5428 vss.n4859 16.2531
R38193 vss.n5435 vss.n5428 16.2531
R38194 vss.n5435 vss.n5434 16.2531
R38195 vss.n5407 vss.n4879 16.2531
R38196 vss.n5407 vss.n5406 16.2531
R38197 vss.n5406 vss.n5331 16.2531
R38198 vss.n5334 vss.n5331 16.2531
R38199 vss.n5347 vss.n5334 16.2531
R38200 vss.n5348 vss.n5347 16.2531
R38201 vss.n5379 vss.n5378 16.2531
R38202 vss.n5380 vss.n5379 16.2531
R38203 vss.n5380 vss.n5356 16.2531
R38204 vss.n5384 vss.n5356 16.2531
R38205 vss.n5392 vss.n5384 16.2531
R38206 vss.n5392 vss.n5391 16.2531
R38207 vss.n9825 vss.n9824 16.2531
R38208 vss.n9824 vss.n2873 16.2531
R38209 vss.n9843 vss.n2873 16.2531
R38210 vss.n9843 vss.n9842 16.2531
R38211 vss.n9842 vss.n2874 16.2531
R38212 vss.n9838 vss.n2874 16.2531
R38213 vss.n2949 vss.n2948 16.2531
R38214 vss.n2972 vss.n2949 16.2531
R38215 vss.n2972 vss.n2971 16.2531
R38216 vss.n2971 vss.n2968 16.2531
R38217 vss.n2968 vss.n2952 16.2531
R38218 vss.n2964 vss.n2952 16.2531
R38219 vss.n2902 vss.n2901 16.2531
R38220 vss.n2926 vss.n2902 16.2531
R38221 vss.n2926 vss.n2925 16.2531
R38222 vss.n2925 vss.n2921 16.2531
R38223 vss.n2921 vss.n2905 16.2531
R38224 vss.n2917 vss.n2905 16.2531
R38225 vss.n4945 vss.n4944 16.2531
R38226 vss.n4944 vss.n4924 16.2531
R38227 vss.n4963 vss.n4924 16.2531
R38228 vss.n4963 vss.n4962 16.2531
R38229 vss.n4962 vss.n4925 16.2531
R38230 vss.n4958 vss.n4925 16.2531
R38231 vss.n5147 vss.n5146 16.2531
R38232 vss.n5146 vss.n5126 16.2531
R38233 vss.n5165 vss.n5126 16.2531
R38234 vss.n5165 vss.n5164 16.2531
R38235 vss.n5164 vss.n5127 16.2531
R38236 vss.n5160 vss.n5127 16.2531
R38237 vss.n3128 vss.n3127 16.2531
R38238 vss.n3127 vss.n3106 16.2531
R38239 vss.n3146 vss.n3106 16.2531
R38240 vss.n3146 vss.n3145 16.2531
R38241 vss.n3145 vss.n3107 16.2531
R38242 vss.n3141 vss.n3107 16.2531
R38243 vss.n4479 vss.n4478 16.2531
R38244 vss.n4478 vss.n4462 16.2531
R38245 vss.n4502 vss.n4462 16.2531
R38246 vss.n4502 vss.n4501 16.2531
R38247 vss.n4501 vss.n4463 16.2531
R38248 vss.n4493 vss.n4463 16.2531
R38249 vss.n4387 vss.n4386 16.2531
R38250 vss.n4386 vss.n4370 16.2531
R38251 vss.n4410 vss.n4370 16.2531
R38252 vss.n4410 vss.n4409 16.2531
R38253 vss.n4409 vss.n4371 16.2531
R38254 vss.n4401 vss.n4371 16.2531
R38255 vss.n4339 vss.n4338 16.2531
R38256 vss.n4338 vss.n4322 16.2531
R38257 vss.n4362 vss.n4322 16.2531
R38258 vss.n4362 vss.n4361 16.2531
R38259 vss.n4361 vss.n4323 16.2531
R38260 vss.n4353 vss.n4323 16.2531
R38261 vss.n3739 vss.n3738 16.2531
R38262 vss.n3738 vss.n3722 16.2531
R38263 vss.n3762 vss.n3722 16.2531
R38264 vss.n3762 vss.n3761 16.2531
R38265 vss.n3761 vss.n3723 16.2531
R38266 vss.n3753 vss.n3723 16.2531
R38267 vss.n4041 vss.n4040 16.2531
R38268 vss.n4040 vss.n4024 16.2531
R38269 vss.n4064 vss.n4024 16.2531
R38270 vss.n4064 vss.n4063 16.2531
R38271 vss.n4063 vss.n4025 16.2531
R38272 vss.n4055 vss.n4025 16.2531
R38273 vss.n3694 vss.n3693 16.2531
R38274 vss.n3693 vss.n3677 16.2531
R38275 vss.n3717 vss.n3677 16.2531
R38276 vss.n3717 vss.n3716 16.2531
R38277 vss.n3716 vss.n3678 16.2531
R38278 vss.n3708 vss.n3678 16.2531
R38279 vss.n4095 vss.n4094 16.2531
R38280 vss.n4094 vss.n4078 16.2531
R38281 vss.n4118 vss.n4078 16.2531
R38282 vss.n4118 vss.n4117 16.2531
R38283 vss.n4117 vss.n4079 16.2531
R38284 vss.n4109 vss.n4079 16.2531
R38285 vss.n3519 vss.n3518 16.2531
R38286 vss.n3518 vss.n3502 16.2531
R38287 vss.n3542 vss.n3502 16.2531
R38288 vss.n3542 vss.n3541 16.2531
R38289 vss.n3541 vss.n3503 16.2531
R38290 vss.n3533 vss.n3503 16.2531
R38291 vss.n3474 vss.n3473 16.2531
R38292 vss.n3473 vss.n3457 16.2531
R38293 vss.n3497 vss.n3457 16.2531
R38294 vss.n3497 vss.n3496 16.2531
R38295 vss.n3496 vss.n3458 16.2531
R38296 vss.n3488 vss.n3458 16.2531
R38297 vss.n5762 vss.n5761 16.2531
R38298 vss.n5761 vss.n5745 16.2531
R38299 vss.n5785 vss.n5745 16.2531
R38300 vss.n5785 vss.n5784 16.2531
R38301 vss.n5784 vss.n5746 16.2531
R38302 vss.n5776 vss.n5746 16.2531
R38303 vss.n4515 vss.n4446 16.2531
R38304 vss.n4515 vss.n4449 16.2531
R38305 vss.n4508 vss.n4449 16.2531
R38306 vss.n4529 vss.n4508 16.2531
R38307 vss.n4529 vss.n4528 16.2531
R38308 vss.n4528 vss.n4527 16.2531
R38309 vss.n4537 vss.n4435 16.2531
R38310 vss.n4545 vss.n4435 16.2531
R38311 vss.n4546 vss.n4545 16.2531
R38312 vss.n4548 vss.n4546 16.2531
R38313 vss.n4548 vss.n4547 16.2531
R38314 vss.n4547 vss.n4425 16.2531
R38315 vss.n4569 vss.n4568 16.2531
R38316 vss.n4568 vss.n4414 16.2531
R38317 vss.n4609 vss.n4414 16.2531
R38318 vss.n4609 vss.n4608 16.2531
R38319 vss.n4608 vss.n4415 16.2531
R38320 vss.n4600 vss.n4415 16.2531
R38321 vss.n4573 vss.n4572 16.2531
R38322 vss.n4573 vss.n3645 16.2531
R38323 vss.n4617 vss.n3645 16.2531
R38324 vss.n4619 vss.n4617 16.2531
R38325 vss.n4619 vss.n4618 16.2531
R38326 vss.n4618 vss.n3633 16.2531
R38327 vss.n3783 vss.n3782 16.2531
R38328 vss.n3782 vss.n3764 16.2531
R38329 vss.n4206 vss.n3764 16.2531
R38330 vss.n4206 vss.n4205 16.2531
R38331 vss.n4205 vss.n3765 16.2531
R38332 vss.n4197 vss.n3765 16.2531
R38333 vss.n3796 vss.n3786 16.2531
R38334 vss.n4175 vss.n3796 16.2531
R38335 vss.n4175 vss.n4174 16.2531
R38336 vss.n4174 vss.n3799 16.2531
R38337 vss.n3815 vss.n3799 16.2531
R38338 vss.n3815 vss.n3814 16.2531
R38339 vss.n3839 vss.n3838 16.2531
R38340 vss.n3838 vss.n3804 16.2531
R38341 vss.n4171 vss.n3804 16.2531
R38342 vss.n4171 vss.n4170 16.2531
R38343 vss.n4170 vss.n3805 16.2531
R38344 vss.n4162 vss.n3805 16.2531
R38345 vss.n3852 vss.n3842 16.2531
R38346 vss.n4140 vss.n3852 16.2531
R38347 vss.n4140 vss.n4139 16.2531
R38348 vss.n4139 vss.n4138 16.2531
R38349 vss.n4138 vss.n3856 16.2531
R38350 vss.n3862 vss.n3856 16.2531
R38351 vss.n3937 vss.n3884 16.2531
R38352 vss.n3945 vss.n3884 16.2531
R38353 vss.n4124 vss.n3945 16.2531
R38354 vss.n4126 vss.n4124 16.2531
R38355 vss.n4126 vss.n4125 16.2531
R38356 vss.n4125 vss.n3872 16.2531
R38357 vss.n3904 vss.n3894 16.2531
R38358 vss.n3927 vss.n3904 16.2531
R38359 vss.n3927 vss.n3926 16.2531
R38360 vss.n3926 vss.n3925 16.2531
R38361 vss.n3925 vss.n3907 16.2531
R38362 vss.n3913 vss.n3907 16.2531
R38363 vss.n3562 vss.n3561 16.2531
R38364 vss.n3561 vss.n3545 16.2531
R38365 vss.n5838 vss.n3545 16.2531
R38366 vss.n5838 vss.n5837 16.2531
R38367 vss.n5837 vss.n3546 16.2531
R38368 vss.n5829 vss.n3546 16.2531
R38369 vss.n3575 vss.n3565 16.2531
R38370 vss.n5807 vss.n3575 16.2531
R38371 vss.n5807 vss.n5806 16.2531
R38372 vss.n5806 vss.n5805 16.2531
R38373 vss.n5805 vss.n3580 16.2531
R38374 vss.n3616 vss.n3580 16.2531
R38375 vss.n5665 vss.n5662 16.2531
R38376 vss.n5665 vss.n3598 16.2531
R38377 vss.n5791 vss.n3598 16.2531
R38378 vss.n5793 vss.n5791 16.2531
R38379 vss.n5793 vss.n5792 16.2531
R38380 vss.n5792 vss.n3586 16.2531
R38381 vss.n5658 vss.n5657 16.2531
R38382 vss.n5657 vss.n3604 16.2531
R38383 vss.n5738 vss.n3604 16.2531
R38384 vss.n5738 vss.n5737 16.2531
R38385 vss.n5737 vss.n3605 16.2531
R38386 vss.n5647 vss.n3605 16.2531
R38387 vss.n5714 vss.n5706 16.2531
R38388 vss.n5722 vss.n5706 16.2531
R38389 vss.n5723 vss.n5722 16.2531
R38390 vss.n5725 vss.n5723 16.2531
R38391 vss.n5725 vss.n5724 16.2531
R38392 vss.n5724 vss.n5694 16.2531
R38393 vss.n9966 vss.n9965 16.2531
R38394 vss.n9965 vss.n2632 16.2531
R38395 vss.n9989 vss.n2632 16.2531
R38396 vss.n9989 vss.n9988 16.2531
R38397 vss.n9988 vss.n2633 16.2531
R38398 vss.n9980 vss.n2633 16.2531
R38399 vss.n2663 vss.n2654 16.2531
R38400 vss.n2671 vss.n2654 16.2531
R38401 vss.n2674 vss.n2671 16.2531
R38402 vss.n2676 vss.n2674 16.2531
R38403 vss.n2676 vss.n2675 16.2531
R38404 vss.n2675 vss.n2642 16.2531
R38405 vss.n3399 vss.n3398 16.2531
R38406 vss.n3398 vss.n3382 16.2531
R38407 vss.n3422 vss.n3382 16.2531
R38408 vss.n3422 vss.n3421 16.2531
R38409 vss.n3421 vss.n3383 16.2531
R38410 vss.n3413 vss.n3383 16.2531
R38411 vss.n3996 vss.n3995 16.2531
R38412 vss.n3995 vss.n3979 16.2531
R38413 vss.n4019 vss.n3979 16.2531
R38414 vss.n4019 vss.n4018 16.2531
R38415 vss.n4018 vss.n3980 16.2531
R38416 vss.n4010 vss.n3980 16.2531
R38417 vss.n4263 vss.n4262 16.2531
R38418 vss.n4262 vss.n4246 16.2531
R38419 vss.n4286 vss.n4246 16.2531
R38420 vss.n4286 vss.n4285 16.2531
R38421 vss.n4285 vss.n4247 16.2531
R38422 vss.n4277 vss.n4247 16.2531
R38423 vss.n5906 vss.n5905 16.2531
R38424 vss.n5905 vss.n5890 16.2531
R38425 vss.n5930 vss.n5890 16.2531
R38426 vss.n5930 vss.n5929 16.2531
R38427 vss.n5929 vss.n5891 16.2531
R38428 vss.n5920 vss.n5891 16.2531
R38429 vss.n14069 vss.n14068 16.2531
R38430 vss.n14068 vss.n476 16.2531
R38431 vss.n14087 vss.n476 16.2531
R38432 vss.n14087 vss.n14086 16.2531
R38433 vss.n14086 vss.n477 16.2531
R38434 vss.n14082 vss.n477 16.2531
R38435 vss.n10124 vss.n10123 16.2531
R38436 vss.n10123 vss.n10103 16.2531
R38437 vss.n10142 vss.n10103 16.2531
R38438 vss.n10142 vss.n10141 16.2531
R38439 vss.n10141 vss.n10104 16.2531
R38440 vss.n10137 vss.n10104 16.2531
R38441 vss.n12882 vss.n12881 16.2531
R38442 vss.n12881 vss.n12861 16.2531
R38443 vss.n12900 vss.n12861 16.2531
R38444 vss.n12900 vss.n12899 16.2531
R38445 vss.n12899 vss.n12862 16.2531
R38446 vss.n12895 vss.n12862 16.2531
R38447 vss.n10165 vss.n10164 16.2531
R38448 vss.n10164 vss.n10144 16.2531
R38449 vss.n10183 vss.n10144 16.2531
R38450 vss.n10183 vss.n10182 16.2531
R38451 vss.n10182 vss.n10145 16.2531
R38452 vss.n10178 vss.n10145 16.2531
R38453 vss.n12431 vss.n12430 16.2531
R38454 vss.n12430 vss.n12410 16.2531
R38455 vss.n12449 vss.n12410 16.2531
R38456 vss.n12449 vss.n12448 16.2531
R38457 vss.n12448 vss.n12411 16.2531
R38458 vss.n12444 vss.n12411 16.2531
R38459 vss.n11760 vss.n11759 16.2531
R38460 vss.n11759 vss.n11739 16.2531
R38461 vss.n11778 vss.n11739 16.2531
R38462 vss.n11778 vss.n11777 16.2531
R38463 vss.n11777 vss.n11740 16.2531
R38464 vss.n11773 vss.n11740 16.2531
R38465 vss.n12476 vss.n12475 16.2531
R38466 vss.n12475 vss.n12455 16.2531
R38467 vss.n12494 vss.n12455 16.2531
R38468 vss.n12494 vss.n12493 16.2531
R38469 vss.n12493 vss.n12456 16.2531
R38470 vss.n12489 vss.n12456 16.2531
R38471 vss.n2319 vss.n2318 16.2531
R38472 vss.n2342 vss.n2319 16.2531
R38473 vss.n2342 vss.n2341 16.2531
R38474 vss.n2341 vss.n2338 16.2531
R38475 vss.n2338 vss.n2322 16.2531
R38476 vss.n2334 vss.n2322 16.2531
R38477 vss.n12301 vss.n12300 16.2531
R38478 vss.n12300 vss.n12280 16.2531
R38479 vss.n12319 vss.n12280 16.2531
R38480 vss.n12319 vss.n12318 16.2531
R38481 vss.n12318 vss.n12281 16.2531
R38482 vss.n12314 vss.n12281 16.2531
R38483 vss.n12346 vss.n12345 16.2531
R38484 vss.n12345 vss.n12325 16.2531
R38485 vss.n12364 vss.n12325 16.2531
R38486 vss.n12364 vss.n12363 16.2531
R38487 vss.n12363 vss.n12326 16.2531
R38488 vss.n12359 vss.n12326 16.2531
R38489 vss.n10242 vss.n10241 16.2531
R38490 vss.n10241 vss.n10221 16.2531
R38491 vss.n10260 vss.n10221 16.2531
R38492 vss.n10260 vss.n10259 16.2531
R38493 vss.n10259 vss.n10222 16.2531
R38494 vss.n10255 vss.n10222 16.2531
R38495 vss.n2422 vss.n2421 16.2531
R38496 vss.n2421 vss.n2401 16.2531
R38497 vss.n2440 vss.n2401 16.2531
R38498 vss.n2440 vss.n2439 16.2531
R38499 vss.n2439 vss.n2402 16.2531
R38500 vss.n2435 vss.n2402 16.2531
R38501 vss.n2379 vss.n2378 16.2531
R38502 vss.n12967 vss.n2379 16.2531
R38503 vss.n12967 vss.n12966 16.2531
R38504 vss.n12966 vss.n2398 16.2531
R38505 vss.n2398 vss.n2382 16.2531
R38506 vss.n2394 vss.n2382 16.2531
R38507 vss.n10034 vss.n10033 16.2531
R38508 vss.n10033 vss.n10018 16.2531
R38509 vss.n12951 vss.n10018 16.2531
R38510 vss.n12951 vss.n12950 16.2531
R38511 vss.n12950 vss.n10019 16.2531
R38512 vss.n10056 vss.n10019 16.2531
R38513 vss.n13088 vss.n2099 16.2531
R38514 vss.n13088 vss.n13087 16.2531
R38515 vss.n13087 vss.n2100 16.2531
R38516 vss.n2103 vss.n2100 16.2531
R38517 vss.n2116 vss.n2103 16.2531
R38518 vss.n2117 vss.n2116 16.2531
R38519 vss.n12927 vss.n12926 16.2531
R38520 vss.n12928 vss.n12927 16.2531
R38521 vss.n12928 vss.n10067 16.2531
R38522 vss.n12936 vss.n10067 16.2531
R38523 vss.n12937 vss.n12936 16.2531
R38524 vss.n12938 vss.n12937 16.2531
R38525 vss.n2502 vss.n2501 16.2531
R38526 vss.n2501 vss.n2480 16.2531
R38527 vss.n2520 vss.n2480 16.2531
R38528 vss.n2520 vss.n2519 16.2531
R38529 vss.n2519 vss.n2481 16.2531
R38530 vss.n2515 vss.n2481 16.2531
R38531 vss.n13073 vss.n13072 16.2531
R38532 vss.n13072 vss.n13071 16.2531
R38533 vss.n13071 vss.n2124 16.2531
R38534 vss.n2139 vss.n2124 16.2531
R38535 vss.n13061 vss.n2139 16.2531
R38536 vss.n13061 vss.n13060 16.2531
R38537 vss.n12105 vss.n12104 16.2531
R38538 vss.n12106 vss.n12105 16.2531
R38539 vss.n12106 vss.n11836 16.2531
R38540 vss.n12116 vss.n11836 16.2531
R38541 vss.n12117 vss.n12116 16.2531
R38542 vss.n12118 vss.n12117 16.2531
R38543 vss.n11820 vss.n11819 16.2531
R38544 vss.n12145 vss.n11820 16.2531
R38545 vss.n12145 vss.n12144 16.2531
R38546 vss.n12144 vss.n12137 16.2531
R38547 vss.n12137 vss.n11823 16.2531
R38548 vss.n12133 vss.n11823 16.2531
R38549 vss.n12158 vss.n12157 16.2531
R38550 vss.n12159 vss.n12158 16.2531
R38551 vss.n12159 vss.n11792 16.2531
R38552 vss.n12169 vss.n11792 16.2531
R38553 vss.n12170 vss.n12169 16.2531
R38554 vss.n12171 vss.n12170 16.2531
R38555 vss.n12256 vss.n12255 16.2531
R38556 vss.n12256 vss.n11781 16.2531
R38557 vss.n12275 vss.n11781 16.2531
R38558 vss.n12275 vss.n12274 16.2531
R38559 vss.n12274 vss.n11782 16.2531
R38560 vss.n12270 vss.n11782 16.2531
R38561 vss.n12202 vss.n12201 16.2531
R38562 vss.n12243 vss.n12202 16.2531
R38563 vss.n12243 vss.n12242 16.2531
R38564 vss.n12242 vss.n12239 16.2531
R38565 vss.n12239 vss.n12205 16.2531
R38566 vss.n12207 vss.n12205 16.2531
R38567 vss.n11732 vss.n11731 16.2531
R38568 vss.n12541 vss.n11732 16.2531
R38569 vss.n12541 vss.n12540 16.2531
R38570 vss.n12540 vss.n11735 16.2531
R38571 vss.n12222 vss.n11735 16.2531
R38572 vss.n12223 vss.n12222 16.2531
R38573 vss.n12554 vss.n12553 16.2531
R38574 vss.n12555 vss.n12554 16.2531
R38575 vss.n12555 vss.n11705 16.2531
R38576 vss.n12565 vss.n11705 16.2531
R38577 vss.n12566 vss.n12565 16.2531
R38578 vss.n12567 vss.n12566 16.2531
R38579 vss.n12583 vss.n12582 16.2531
R38580 vss.n12582 vss.n12581 16.2531
R38581 vss.n12581 vss.n11628 16.2531
R38582 vss.n12577 vss.n11628 16.2531
R38583 vss.n12577 vss.n12576 16.2531
R38584 vss.n12576 vss.n12575 16.2531
R38585 vss.n11653 vss.n11652 16.2531
R38586 vss.n11678 vss.n11653 16.2531
R38587 vss.n11678 vss.n11677 16.2531
R38588 vss.n11677 vss.n11674 16.2531
R38589 vss.n11674 vss.n11656 16.2531
R38590 vss.n11658 vss.n11656 16.2531
R38591 vss.n12836 vss.n12835 16.2531
R38592 vss.n12836 vss.n10304 16.2531
R38593 vss.n12855 vss.n10304 16.2531
R38594 vss.n12855 vss.n12854 16.2531
R38595 vss.n12854 vss.n10305 16.2531
R38596 vss.n12850 vss.n10305 16.2531
R38597 vss.n12784 vss.n12783 16.2531
R38598 vss.n12823 vss.n12784 16.2531
R38599 vss.n12823 vss.n12822 16.2531
R38600 vss.n12822 vss.n12821 16.2531
R38601 vss.n12821 vss.n12787 16.2531
R38602 vss.n12789 vss.n12787 16.2531
R38603 vss.n10097 vss.n10096 16.2531
R38604 vss.n12914 vss.n10097 16.2531
R38605 vss.n12914 vss.n12913 16.2531
R38606 vss.n12913 vss.n10100 16.2531
R38607 vss.n12804 vss.n10100 16.2531
R38608 vss.n12805 vss.n12804 16.2531
R38609 vss.n11880 vss.n11872 16.2531
R38610 vss.n11888 vss.n11872 16.2531
R38611 vss.n12076 vss.n11888 16.2531
R38612 vss.n12078 vss.n12076 16.2531
R38613 vss.n12078 vss.n12077 16.2531
R38614 vss.n12077 vss.n11860 16.2531
R38615 vss.n10479 vss.n10478 16.2531
R38616 vss.n10478 vss.n10462 16.2531
R38617 vss.n10501 vss.n10462 16.2531
R38618 vss.n10501 vss.n10500 16.2531
R38619 vss.n10500 vss.n10463 16.2531
R38620 vss.n10492 vss.n10463 16.2531
R38621 vss.n10700 vss.n10699 16.2531
R38622 vss.n10699 vss.n10683 16.2531
R38623 vss.n10722 vss.n10683 16.2531
R38624 vss.n10722 vss.n10721 16.2531
R38625 vss.n10721 vss.n10684 16.2531
R38626 vss.n10713 vss.n10684 16.2531
R38627 vss.n11014 vss.n11013 16.2531
R38628 vss.n11013 vss.n10997 16.2531
R38629 vss.n11036 vss.n10997 16.2531
R38630 vss.n11036 vss.n11035 16.2531
R38631 vss.n11035 vss.n10998 16.2531
R38632 vss.n11027 vss.n10998 16.2531
R38633 vss.n11122 vss.n11121 16.2531
R38634 vss.n11121 vss.n11106 16.2531
R38635 vss.n11145 vss.n11106 16.2531
R38636 vss.n11145 vss.n11144 16.2531
R38637 vss.n11144 vss.n11107 16.2531
R38638 vss.n11135 vss.n11107 16.2531
R38639 vss.n11153 vss.n11152 15.2779
R38640 vss.n11152 vss.n11151 15.2779
R38641 vss.n11104 vss.n11103 15.2779
R38642 vss.n11103 vss.n11102 15.2779
R38643 vss.n11102 vss.n11101 15.2779
R38644 vss.n11172 vss.n11171 15.2779
R38645 vss.n11171 vss.n11043 15.2779
R38646 vss.n11356 vss.n11355 15.2779
R38647 vss.n11355 vss.n11354 15.2779
R38648 vss.n11354 vss.n11353 15.2779
R38649 vss.n11234 vss.n11233 15.2779
R38650 vss.n11233 vss.n11232 15.2779
R38651 vss.n11230 vss.n11229 15.2779
R38652 vss.n11229 vss.n11228 15.2779
R38653 vss.n11228 vss.n11227 15.2779
R38654 vss.n11295 vss.n11294 15.2779
R38655 vss.n11294 vss.n11293 15.2779
R38656 vss.n11291 vss.n11290 15.2779
R38657 vss.n11290 vss.n11289 15.2779
R38658 vss.n11289 vss.n11288 15.2779
R38659 vss.n14765 vss.n104 15.2779
R38660 vss.n14765 vss.n14764 15.2779
R38661 vss.n14764 vss.n14763 15.2779
R38662 vss.n393 vss.n392 15.2779
R38663 vss.n392 vss.n391 15.2779
R38664 vss.n391 vss.n381 15.2779
R38665 vss.n270 vss.n269 15.2779
R38666 vss.n269 vss.n268 15.2779
R38667 vss.n268 vss.n258 15.2779
R38668 vss.n14427 vss.n14426 15.2779
R38669 vss.n14426 vss.n14425 15.2779
R38670 vss.n14425 vss.n14415 15.2779
R38671 vss.n211 vss.n210 15.2779
R38672 vss.n210 vss.n209 15.2779
R38673 vss.n209 vss.n199 15.2779
R38674 vss.n14622 vss.n14621 15.2779
R38675 vss.n14621 vss.n14620 15.2779
R38676 vss.n14620 vss.n14610 15.2779
R38677 vss.n134 vss.n133 15.2779
R38678 vss.n133 vss.n132 15.2779
R38679 vss.n132 vss.n122 15.2779
R38680 vss.n376 vss.n375 15.2779
R38681 vss.n377 vss.n376 15.2779
R38682 vss.n378 vss.n377 15.2779
R38683 vss.n7377 vss.n7376 15.2779
R38684 vss.n7376 vss.n7375 15.2779
R38685 vss.n7375 vss.n7374 15.2779
R38686 vss.n7828 vss.n7826 15.2779
R38687 vss.n7828 vss.n7827 15.2779
R38688 vss.n7827 vss.n7812 15.2779
R38689 vss.n7641 vss.n7639 15.2779
R38690 vss.n7641 vss.n7640 15.2779
R38691 vss.n7640 vss.n7625 15.2779
R38692 vss.n7452 vss.n7450 15.2779
R38693 vss.n7452 vss.n7451 15.2779
R38694 vss.n7451 vss.n7436 15.2779
R38695 vss.n8983 vss.n8982 15.2779
R38696 vss.n8982 vss.n8981 15.2779
R38697 vss.n8981 vss.n8980 15.2779
R38698 vss.n7606 vss.n7604 15.2779
R38699 vss.n7606 vss.n7605 15.2779
R38700 vss.n7605 vss.n7590 15.2779
R38701 vss.n7749 vss.n7747 15.2779
R38702 vss.n7749 vss.n7748 15.2779
R38703 vss.n7748 vss.n7733 15.2779
R38704 vss.n7970 vss.n7968 15.2779
R38705 vss.n7970 vss.n7969 15.2779
R38706 vss.n7969 vss.n7954 15.2779
R38707 vss.n3241 vss.n3236 15.2779
R38708 vss.n3237 vss.n3236 15.2779
R38709 vss.n3237 vss.n3227 15.2779
R38710 vss.n3084 vss.n3079 15.2779
R38711 vss.n3080 vss.n3079 15.2779
R38712 vss.n3080 vss.n3070 15.2779
R38713 vss.n5058 vss.n5053 15.2779
R38714 vss.n5054 vss.n5053 15.2779
R38715 vss.n5054 vss.n5044 15.2779
R38716 vss.n2850 vss.n2845 15.2779
R38717 vss.n2846 vss.n2845 15.2779
R38718 vss.n2846 vss.n2836 15.2779
R38719 vss.n9851 vss.n2827 15.2779
R38720 vss.n9854 vss.n9851 15.2779
R38721 vss.n9854 vss.n9853 15.2779
R38722 vss.n4981 vss.n4976 15.2779
R38723 vss.n4977 vss.n4976 15.2779
R38724 vss.n4977 vss.n4967 15.2779
R38725 vss.n5183 vss.n5178 15.2779
R38726 vss.n5179 vss.n5178 15.2779
R38727 vss.n5179 vss.n5169 15.2779
R38728 vss.n3164 vss.n3159 15.2779
R38729 vss.n3160 vss.n3159 15.2779
R38730 vss.n3160 vss.n3150 15.2779
R38731 vss.n10200 vss.n10195 15.2779
R38732 vss.n10196 vss.n10195 15.2779
R38733 vss.n10196 vss.n10186 15.2779
R38734 vss.n10218 vss.n10187 15.2779
R38735 vss.n10214 vss.n10187 15.2779
R38736 vss.n12511 vss.n12506 15.2779
R38737 vss.n12507 vss.n12506 15.2779
R38738 vss.n12507 vss.n12497 15.2779
R38739 vss.n12529 vss.n12498 15.2779
R38740 vss.n12525 vss.n12498 15.2779
R38741 vss.n2219 vss.n2214 15.2779
R38742 vss.n2215 vss.n2214 15.2779
R38743 vss.n2215 vss.n2205 15.2779
R38744 vss.n2237 vss.n2206 15.2779
R38745 vss.n2233 vss.n2206 15.2779
R38746 vss.n12382 vss.n12377 15.2779
R38747 vss.n12378 vss.n12377 15.2779
R38748 vss.n12378 vss.n12368 15.2779
R38749 vss.n12400 vss.n12369 15.2779
R38750 vss.n12396 vss.n12369 15.2779
R38751 vss.n10278 vss.n10273 15.2779
R38752 vss.n10274 vss.n10273 15.2779
R38753 vss.n10274 vss.n10264 15.2779
R38754 vss.n10296 vss.n10265 15.2779
R38755 vss.n10292 vss.n10265 15.2779
R38756 vss.n2458 vss.n2453 15.2779
R38757 vss.n2454 vss.n2453 15.2779
R38758 vss.n2454 vss.n2444 15.2779
R38759 vss.n2476 vss.n2445 15.2779
R38760 vss.n2472 vss.n2445 15.2779
R38761 vss.n2537 vss.n2532 15.2779
R38762 vss.n2533 vss.n2532 15.2779
R38763 vss.n2533 vss.n2523 15.2779
R38764 vss.n2555 vss.n2524 15.2779
R38765 vss.n2551 vss.n2524 15.2779
R38766 vss.n13029 vss.n13025 15.2779
R38767 vss.n13041 vss.n13025 15.2779
R38768 vss.n13041 vss.n13040 15.2779
R38769 vss.n13046 vss.n13045 15.2779
R38770 vss.n13048 vss.n13046 15.2779
R38771 vss.n11325 vss.n11324 15.2779
R38772 vss.n11324 vss.n11323 15.2779
R38773 vss.n11309 vss.n11308 15.2779
R38774 vss.n11310 vss.n11309 15.2779
R38775 vss.n11311 vss.n11310 15.2779
R38776 vss.n11264 vss.n11263 15.2779
R38777 vss.n11263 vss.n11262 15.2779
R38778 vss.n11248 vss.n11247 15.2779
R38779 vss.n11249 vss.n11248 15.2779
R38780 vss.n11250 vss.n11249 15.2779
R38781 vss.n11203 vss.n11202 15.2779
R38782 vss.n11202 vss.n11201 15.2779
R38783 vss.n11199 vss.n11198 15.2779
R38784 vss.n11198 vss.n11197 15.2779
R38785 vss.n11197 vss.n11196 15.2779
R38786 vss.n12669 vss.n12668 15.2779
R38787 vss.n12668 vss.n12667 15.2779
R38788 vss.n11342 vss.n10459 15.2779
R38789 vss.n11347 vss.n11342 15.2779
R38790 vss.n11347 vss.n11346 15.2779
R38791 vss.n11151 vss.n11150 14.9682
R38792 vss.n11357 vss.n11043 14.9682
R38793 vss.n11232 vss.n11231 14.9682
R38794 vss.n11293 vss.n11292 14.9682
R38795 vss.n14762 vss.n121 14.9682
R38796 vss.n411 vss.n410 14.9682
R38797 vss.n288 vss.n287 14.9682
R38798 vss.n14445 vss.n14444 14.9682
R38799 vss.n229 vss.n228 14.9682
R38800 vss.n14640 vss.n14639 14.9682
R38801 vss.n152 vss.n151 14.9682
R38802 vss.n380 vss.n379 14.9682
R38803 vss.n7373 vss.n7372 14.9682
R38804 vss.n7846 vss.n7845 14.9682
R38805 vss.n7659 vss.n7658 14.9682
R38806 vss.n7470 vss.n7469 14.9682
R38807 vss.n8979 vss.n7435 14.9682
R38808 vss.n7624 vss.n7623 14.9682
R38809 vss.n7767 vss.n7766 14.9682
R38810 vss.n7988 vss.n7987 14.9682
R38811 vss.n3260 vss.n3259 14.9682
R38812 vss.n3103 vss.n3102 14.9682
R38813 vss.n5077 vss.n5076 14.9682
R38814 vss.n2869 vss.n2868 14.9682
R38815 vss.n9860 vss.n9849 14.9682
R38816 vss.n5000 vss.n4999 14.9682
R38817 vss.n5202 vss.n5201 14.9682
R38818 vss.n3183 vss.n3182 14.9682
R38819 vss.n10219 vss.n10218 14.9682
R38820 vss.n12530 vss.n12529 14.9682
R38821 vss.n2238 vss.n2237 14.9682
R38822 vss.n12401 vss.n12400 14.9682
R38823 vss.n10297 vss.n10296 14.9682
R38824 vss.n2477 vss.n2476 14.9682
R38825 vss.n2556 vss.n2555 14.9682
R38826 vss.n13045 vss.n13023 14.9682
R38827 vss.n11323 vss.n10460 14.9682
R38828 vss.n11262 vss.n10681 14.9682
R38829 vss.n11201 vss.n11200 14.9682
R38830 vss.n12667 vss.n12666 14.9682
R38831 vss.n120 vss.n109 13.5231
R38832 vss.n121 vss.n120 13.5231
R38833 vss.n409 vss.n382 13.5231
R38834 vss.n410 vss.n409 13.5231
R38835 vss.n286 vss.n259 13.5231
R38836 vss.n287 vss.n286 13.5231
R38837 vss.n14443 vss.n14416 13.5231
R38838 vss.n14444 vss.n14443 13.5231
R38839 vss.n227 vss.n200 13.5231
R38840 vss.n228 vss.n227 13.5231
R38841 vss.n14638 vss.n14611 13.5231
R38842 vss.n14639 vss.n14638 13.5231
R38843 vss.n150 vss.n123 13.5231
R38844 vss.n151 vss.n150 13.5231
R38845 vss.n69 vss.n66 13.5231
R38846 vss.n379 vss.n69 13.5231
R38847 vss.n14048 vss.n14035 13.5231
R38848 vss.n508 vss.n507 13.5231
R38849 vss.n511 vss.n507 13.5231
R38850 vss.n14034 vss.n511 13.5231
R38851 vss.n14049 vss.n14034 13.5231
R38852 vss.n14049 vss.n14048 13.5231
R38853 vss.n1594 vss.n1593 13.5231
R38854 vss.n1581 vss.n1580 13.5231
R38855 vss.n1581 vss.n1572 13.5231
R38856 vss.n1605 vss.n1572 13.5231
R38857 vss.n1605 vss.n1573 13.5231
R38858 vss.n1594 vss.n1573 13.5231
R38859 vss.n1299 vss.n1298 13.5231
R38860 vss.n1286 vss.n1285 13.5231
R38861 vss.n1286 vss.n1277 13.5231
R38862 vss.n1310 vss.n1277 13.5231
R38863 vss.n1310 vss.n1278 13.5231
R38864 vss.n1299 vss.n1278 13.5231
R38865 vss.n1038 vss.n1037 13.5231
R38866 vss.n1025 vss.n1024 13.5231
R38867 vss.n1025 vss.n1016 13.5231
R38868 vss.n1049 vss.n1016 13.5231
R38869 vss.n1049 vss.n1017 13.5231
R38870 vss.n1038 vss.n1017 13.5231
R38871 vss.n1431 vss.n1430 13.5231
R38872 vss.n1418 vss.n1417 13.5231
R38873 vss.n1418 vss.n1409 13.5231
R38874 vss.n1442 vss.n1409 13.5231
R38875 vss.n1442 vss.n1410 13.5231
R38876 vss.n1431 vss.n1410 13.5231
R38877 vss.n1511 vss.n1510 13.5231
R38878 vss.n1498 vss.n1497 13.5231
R38879 vss.n1498 vss.n1489 13.5231
R38880 vss.n1522 vss.n1489 13.5231
R38881 vss.n1522 vss.n1490 13.5231
R38882 vss.n1511 vss.n1490 13.5231
R38883 vss.n953 vss.n952 13.5231
R38884 vss.n967 vss.n966 13.5231
R38885 vss.n966 vss.n965 13.5231
R38886 vss.n965 vss.n964 13.5231
R38887 vss.n964 vss.n938 13.5231
R38888 vss.n953 vss.n938 13.5231
R38889 vss.n1005 vss.n1004 13.5231
R38890 vss.n13207 vss.n13206 13.5231
R38891 vss.n13206 vss.n13205 13.5231
R38892 vss.n13205 vss.n13204 13.5231
R38893 vss.n13204 vss.n990 13.5231
R38894 vss.n1005 vss.n990 13.5231
R38895 vss.n7362 vss.n7346 13.5231
R38896 vss.n7372 vss.n7346 13.5231
R38897 vss.n7844 vss.n7813 13.5231
R38898 vss.n7845 vss.n7844 13.5231
R38899 vss.n7657 vss.n7626 13.5231
R38900 vss.n7658 vss.n7657 13.5231
R38901 vss.n7468 vss.n7437 13.5231
R38902 vss.n7469 vss.n7468 13.5231
R38903 vss.n7434 vss.n7411 13.5231
R38904 vss.n7435 vss.n7434 13.5231
R38905 vss.n7622 vss.n7591 13.5231
R38906 vss.n7623 vss.n7622 13.5231
R38907 vss.n7765 vss.n7734 13.5231
R38908 vss.n7766 vss.n7765 13.5231
R38909 vss.n7986 vss.n7955 13.5231
R38910 vss.n7987 vss.n7986 13.5231
R38911 vss.n6248 vss.n6232 13.5231
R38912 vss.n6255 vss.n6254 13.5231
R38913 vss.n6254 vss.n6253 13.5231
R38914 vss.n6253 vss.n6007 13.5231
R38915 vss.n6249 vss.n6007 13.5231
R38916 vss.n6249 vss.n6248 13.5231
R38917 vss.n6617 vss.n6603 13.5231
R38918 vss.n6609 vss.n6608 13.5231
R38919 vss.n6608 vss.n6596 13.5231
R38920 vss.n6628 vss.n6596 13.5231
R38921 vss.n6628 vss.n6597 13.5231
R38922 vss.n6603 vss.n6597 13.5231
R38923 vss.n6390 vss.n6376 13.5231
R38924 vss.n6382 vss.n6381 13.5231
R38925 vss.n6381 vss.n6369 13.5231
R38926 vss.n6401 vss.n6369 13.5231
R38927 vss.n6401 vss.n6370 13.5231
R38928 vss.n6376 vss.n6370 13.5231
R38929 vss.n9277 vss.n9261 13.5231
R38930 vss.n9284 vss.n9283 13.5231
R38931 vss.n9283 vss.n9282 13.5231
R38932 vss.n9282 vss.n9257 13.5231
R38933 vss.n9278 vss.n9257 13.5231
R38934 vss.n9278 vss.n9277 13.5231
R38935 vss.n6926 vss.n6912 13.5231
R38936 vss.n6918 vss.n6917 13.5231
R38937 vss.n6917 vss.n6905 13.5231
R38938 vss.n6937 vss.n6905 13.5231
R38939 vss.n6937 vss.n6906 13.5231
R38940 vss.n6912 vss.n6906 13.5231
R38941 vss.n7115 vss.n7101 13.5231
R38942 vss.n7107 vss.n7106 13.5231
R38943 vss.n7106 vss.n7094 13.5231
R38944 vss.n7126 vss.n7094 13.5231
R38945 vss.n7126 vss.n7095 13.5231
R38946 vss.n7101 vss.n7095 13.5231
R38947 vss.n6286 vss.n6270 13.5231
R38948 vss.n6293 vss.n6292 13.5231
R38949 vss.n6292 vss.n6291 13.5231
R38950 vss.n6291 vss.n6266 13.5231
R38951 vss.n6287 vss.n6266 13.5231
R38952 vss.n6287 vss.n6286 13.5231
R38953 vss.n9299 vss.n9298 13.5231
R38954 vss.n9314 vss.n9313 13.5231
R38955 vss.n9313 vss.n6214 13.5231
R38956 vss.n9319 vss.n6214 13.5231
R38957 vss.n9319 vss.n6215 13.5231
R38958 vss.n9299 vss.n6215 13.5231
R38959 vss.n3320 vss.n3319 13.5231
R38960 vss.n3329 vss.n3328 13.5231
R38961 vss.n3329 vss.n3308 13.5231
R38962 vss.n5888 vss.n3308 13.5231
R38963 vss.n5888 vss.n3309 13.5231
R38964 vss.n3319 vss.n3309 13.5231
R38965 vss.n3255 vss.n3228 13.5231
R38966 vss.n3259 vss.n3228 13.5231
R38967 vss.n3098 vss.n3071 13.5231
R38968 vss.n3102 vss.n3071 13.5231
R38969 vss.n5072 vss.n5045 13.5231
R38970 vss.n5076 vss.n5045 13.5231
R38971 vss.n2864 vss.n2837 13.5231
R38972 vss.n2868 vss.n2837 13.5231
R38973 vss.n9861 vss.n2835 13.5231
R38974 vss.n9861 vss.n9860 13.5231
R38975 vss.n4995 vss.n4968 13.5231
R38976 vss.n4999 vss.n4968 13.5231
R38977 vss.n5197 vss.n5170 13.5231
R38978 vss.n5201 vss.n5170 13.5231
R38979 vss.n3178 vss.n3151 13.5231
R38980 vss.n3182 vss.n3151 13.5231
R38981 vss.n4297 vss.n4296 13.5231
R38982 vss.n4308 vss.n4307 13.5231
R38983 vss.n4308 vss.n4291 13.5231
R38984 vss.n4320 vss.n4291 13.5231
R38985 vss.n4320 vss.n4292 13.5231
R38986 vss.n4297 vss.n4292 13.5231
R38987 vss.n3652 vss.n3651 13.5231
R38988 vss.n3663 vss.n3662 13.5231
R38989 vss.n3663 vss.n3646 13.5231
R38990 vss.n3675 vss.n3646 13.5231
R38991 vss.n3675 vss.n3647 13.5231
R38992 vss.n3652 vss.n3647 13.5231
R38993 vss.n3432 vss.n3431 13.5231
R38994 vss.n3443 vss.n3442 13.5231
R38995 vss.n3443 vss.n3426 13.5231
R38996 vss.n3455 vss.n3426 13.5231
R38997 vss.n3455 vss.n3427 13.5231
R38998 vss.n3432 vss.n3427 13.5231
R38999 vss.n5870 vss.n5869 13.5231
R39000 vss.n9997 vss.n9996 13.5231
R39001 vss.n9996 vss.n9995 13.5231
R39002 vss.n9995 vss.n9994 13.5231
R39003 vss.n9994 vss.n2628 13.5231
R39004 vss.n5870 vss.n2628 13.5231
R39005 vss.n3369 vss.n3368 13.5231
R39006 vss.n5851 vss.n3363 13.5231
R39007 vss.n5851 vss.n5850 13.5231
R39008 vss.n5850 vss.n5849 13.5231
R39009 vss.n5849 vss.n3364 13.5231
R39010 vss.n3369 vss.n3364 13.5231
R39011 vss.n3954 vss.n3953 13.5231
R39012 vss.n3965 vss.n3964 13.5231
R39013 vss.n3965 vss.n3948 13.5231
R39014 vss.n3977 vss.n3948 13.5231
R39015 vss.n3977 vss.n3949 13.5231
R39016 vss.n3954 vss.n3949 13.5231
R39017 vss.n4221 vss.n4220 13.5231
R39018 vss.n4232 vss.n4231 13.5231
R39019 vss.n4232 vss.n4215 13.5231
R39020 vss.n4244 vss.n4215 13.5231
R39021 vss.n4244 vss.n4216 13.5231
R39022 vss.n4221 vss.n4216 13.5231
R39023 vss.n10000 vss.n9999 12.1759
R39024 vss.t1197 vss.n3269 8.39745
R39025 vss.t973 vss.n442 8.39745
R39026 vss.n13155 vss 7.1255
R39027 vss.n13150 vss.n13149 7.05642
R39028 vss.n13152 vss.n13151 6.93142
R39029 vss.n13154 vss.n13153 6.93142
R39030 vss.n14093 vss.n14092 5.17978
R39031 vss.n9634 vss.n9633 5.17978
R39032 vss.n9732 vss.n9731 5.17978
R39033 vss.n12960 vss.n10014 5.17978
R39034 vss.n13151 vss.n13150 5.10905
R39035 vss.n13153 vss.n13152 5.10905
R39036 vss.n13155 vss.n13154 5.10905
R39037 vss vss.n9682 4.95527
R39038 vss.n9730 vss 4.83932
R39039 vss.n14091 vss 4.83932
R39040 vss vss.n10010 4.7579
R39041 vss vss.n9628 4.7579
R39042 vss.n9632 vss 4.64195
R39043 vss.n14092 vss 4.35741
R39044 vss.n9633 vss 4.35741
R39045 vss.n9731 vss 4.35741
R39046 vss vss.n10014 4.35741
R39047 vss.n6220 vss.n5970 3.88057
R39048 vss.n10014 vss.n10013 3.55067
R39049 vss.n13653 vss.n13649 2.88866
R39050 vss.n13758 vss.n13754 2.88866
R39051 vss.n13863 vss.n13859 2.88866
R39052 vss.n1906 vss.n1201 2.88866
R39053 vss.n1802 vss.n1697 2.88866
R39054 vss.n13290 vss.n13289 2.88866
R39055 vss.n9247 vss.n6489 2.88866
R39056 vss.n7084 vss.n6717 2.88866
R39057 vss.n9145 vss.n6546 2.88866
R39058 vss.n5739 vss.n3602 2.88866
R39059 vss.n5839 vss.n3543 2.88866
R39060 vss.n4173 vss.n4172 2.88866
R39061 vss.n4610 vss.n4412 2.88866
R39062 vss.n12953 vss.n12952 2.88866
R39063 vss.n12075 vss.n12074 2.88866
R39064 vss.n12610 vss.n10590 2.88866
R39065 vss.n11539 vss.n10811 2.88866
R39066 vss.n12740 vss.n12739 2.88866
R39067 vss.n14145 vss.n14142 2.88866
R39068 vss.n13991 vss.n13990 2.88866
R39069 vss.n8477 vss.n8474 2.88866
R39070 vss.n8379 vss.n8376 2.88866
R39071 vss.n8258 vss.n7906 2.88866
R39072 vss.n9641 vss.n6004 2.88866
R39073 vss.n9540 vss.n9539 2.88866
R39074 vss.n5330 vss.n5327 2.88866
R39075 vss.n5269 vss.n5268 2.88866
R39076 vss.n5210 vss.n5209 2.88866
R39077 vss.n9740 vss.n9739 2.88866
R39078 vss.n12143 vss.n12140 2.88866
R39079 vss.n12539 vss.n11736 2.88866
R39080 vss.n12856 vss.n10302 2.88866
R39081 vss.n14092 vss.n14091 2.43143
R39082 vss.n9633 vss.n9632 2.43143
R39083 vss.n9731 vss.n9730 2.43143
R39084 vss.n14139 vss.n14138 1.89112
R39085 vss.n9638 vss.n9637 1.89112
R39086 vss.n9736 vss.n9735 1.89112
R39087 vss.n12957 vss.n12956 1.89112
R39088 vss.n13203 vss 1.87386
R39089 vss vss.n9364 1.87386
R39090 vss.n9993 vss 1.87386
R39091 vss.n12665 vss 1.87386
R39092 vss.n14034 vss.n14033 1.52776
R39093 vss.n1649 vss.n1605 1.52776
R39094 vss.n1357 vss.n1310 1.52776
R39095 vss.n1094 vss.n1049 1.52776
R39096 vss.n1487 vss.n1442 1.52776
R39097 vss.n1570 vss.n1522 1.52776
R39098 vss.n964 vss.n515 1.52776
R39099 vss.n13204 vss.n13203 1.52776
R39100 vss.n9582 vss.n6007 1.52776
R39101 vss.n7093 vss.n6628 1.52776
R39102 vss.n6446 vss.n6401 1.52776
R39103 vss.n9257 vss.n9256 1.52776
R39104 vss.n6983 vss.n6937 1.52776
R39105 vss.n7174 vss.n7126 1.52776
R39106 vss.n6266 vss.n6054 1.52776
R39107 vss.n9364 vss.n9319 1.52776
R39108 vss.n5934 vss.n5888 1.52776
R39109 vss.n4365 vss.n4320 1.52776
R39110 vss.n3720 vss.n3675 1.52776
R39111 vss.n3500 vss.n3455 1.52776
R39112 vss.n9994 vss.n9993 1.52776
R39113 vss.n5849 vss.n5848 1.52776
R39114 vss.n4073 vss.n3977 1.52776
R39115 vss.n4290 vss.n4244 1.52776
R39116 vss.n9874 vss.n2783 1.44407
R39117 vss.n11401 vss.n11042 1.44293
R39118 vss.n10995 vss.n10769 1.44293
R39119 vss.n11549 vss.n10548 1.44293
R39120 vss.n12665 vss.n12620 1.44293
R39121 vss.n14093 vss.n412 1.44293
R39122 vss.n14369 vss.n289 1.44293
R39123 vss.n14252 vss.n289 1.44293
R39124 vss.n14252 vss.n14251 1.44293
R39125 vss.n14446 vss.n14369 1.44293
R39126 vss.n14564 vss.n230 1.44293
R39127 vss.n14447 vss.n230 1.44293
R39128 vss.n14641 vss.n14564 1.44293
R39129 vss.n14759 vss.n153 1.44293
R39130 vss.n14642 vss.n153 1.44293
R39131 vss.n14642 vss.n14641 1.44293
R39132 vss.n14251 vss.n14250 1.44293
R39133 vss.n14250 vss.n412 1.44293
R39134 vss.n1649 vss.n1571 1.44293
R39135 vss.n1408 vss.n1357 1.44293
R39136 vss.n1984 vss.n1094 1.44293
R39137 vss.n1356 vss.n1094 1.44293
R39138 vss.n1357 vss.n1356 1.44293
R39139 vss.n1487 vss.n1408 1.44293
R39140 vss.n1650 vss.n1649 1.44293
R39141 vss.n1571 vss.n1570 1.44293
R39142 vss.n1570 vss.n1569 1.44293
R39143 vss.n1569 vss.n515 1.44293
R39144 vss.n14032 vss.n515 1.44293
R39145 vss.n14033 vss.n14032 1.44293
R39146 vss.n13203 vss.n1984 1.44293
R39147 vss.n9634 vss.n6006 1.44293
R39148 vss.n8250 vss.n7847 1.44293
R39149 vss.n8741 vss.n7660 1.44293
R39150 vss.n8860 vss.n7471 1.44293
R39151 vss.n8978 vss.n8977 1.44293
R39152 vss.n8977 vss.n7471 1.44293
R39153 vss.n8860 vss.n8859 1.44293
R39154 vss.n8859 vss.n8858 1.44293
R39155 vss.n8858 vss.n7660 1.44293
R39156 vss.n8740 vss.n8739 1.44293
R39157 vss.n8739 vss.n7847 1.44293
R39158 vss.n8250 vss.n8249 1.44293
R39159 vss.n8249 vss.n8248 1.44293
R39160 vss.n8248 vss.n6006 1.44293
R39161 vss.n7175 vss.n7093 1.44293
R39162 vss.n6984 vss.n6446 1.44293
R39163 vss.n9256 vss.n6213 1.44293
R39164 vss.n9256 vss.n9255 1.44293
R39165 vss.n9255 vss.n6446 1.44293
R39166 vss.n6984 vss.n6983 1.44293
R39167 vss.n7093 vss.n7092 1.44293
R39168 vss.n7175 vss.n7174 1.44293
R39169 vss.n7174 vss.n7173 1.44293
R39170 vss.n7173 vss.n6054 1.44293
R39171 vss.n9581 vss.n6054 1.44293
R39172 vss.n9582 vss.n9581 1.44293
R39173 vss.n9364 vss.n6213 1.44293
R39174 vss.n9732 vss.n3261 1.44293
R39175 vss.n9790 vss.n3104 1.44293
R39176 vss.n5260 vss.n5078 1.44293
R39177 vss.n5319 vss.n2870 1.44293
R39178 vss.n9848 vss.n9847 1.44293
R39179 vss.n9847 vss.n2870 1.44293
R39180 vss.n5319 vss.n5318 1.44293
R39181 vss.n5318 vss.n5317 1.44293
R39182 vss.n5317 vss.n5078 1.44293
R39183 vss.n5259 vss.n5258 1.44293
R39184 vss.n5258 vss.n3104 1.44293
R39185 vss.n9790 vss.n9789 1.44293
R39186 vss.n9789 vss.n9788 1.44293
R39187 vss.n9788 vss.n3261 1.44293
R39188 vss.n4365 vss.n3307 1.44293
R39189 vss.n4214 vss.n3720 1.44293
R39190 vss.n4074 vss.n3500 1.44293
R39191 vss.n9993 vss.n2630 1.44293
R39192 vss.n5848 vss.n2630 1.44293
R39193 vss.n5848 vss.n5847 1.44293
R39194 vss.n5847 vss.n3500 1.44293
R39195 vss.n4074 vss.n4073 1.44293
R39196 vss.n4072 vss.n3720 1.44293
R39197 vss.n4290 vss.n4214 1.44293
R39198 vss.n4366 vss.n4290 1.44293
R39199 vss.n4366 vss.n4365 1.44293
R39200 vss.n5934 vss.n3307 1.44293
R39201 vss.n12906 vss.n12905 1.44293
R39202 vss.n12531 vss.n12453 1.44293
R39203 vss.n12323 vss.n2239 1.44293
R39204 vss.n12402 vss.n12323 1.44293
R39205 vss.n12532 vss.n12402 1.44293
R39206 vss.n12532 vss.n12531 1.44293
R39207 vss.n12904 vss.n10298 1.44293
R39208 vss.n12905 vss.n12904 1.44293
R39209 vss.n12906 vss.n2478 1.44293
R39210 vss.n12962 vss.n2478 1.44293
R39211 vss.n12962 vss.n12961 1.44293
R39212 vss.n12961 vss.n12960 1.44293
R39213 vss.n13022 vss.n13021 1.44293
R39214 vss.n13021 vss.n2239 1.44293
R39215 vss.n12620 vss.n12619 1.44293
R39216 vss.n12619 vss.n12618 1.44293
R39217 vss.n12618 vss.n10548 1.44293
R39218 vss.n11549 vss.n11548 1.44293
R39219 vss.n11547 vss.n10769 1.44293
R39220 vss.n11040 vss.n10995 1.44293
R39221 vss.n11402 vss.n11040 1.44293
R39222 vss.n11402 vss.n11401 1.44293
R39223 vss.n11149 vss.n11042 1.44293
R39224 vss.n14761 vss.n14759 1.44293
R39225 vss.n14255 vss.n316 1.19376
R39226 vss.n14366 vss.n290 1.19376
R39227 vss.n14450 vss.n257 1.19376
R39228 vss.n14561 vss.n231 1.19376
R39229 vss.n14645 vss.n198 1.19376
R39230 vss.n14756 vss.n154 1.19376
R39231 vss.n14247 vss.n413 1.19376
R39232 vss.n1910 vss.n1200 1.19376
R39233 vss.n1405 vss.n1404 1.19376
R39234 vss.n1806 vss.n1694 1.19376
R39235 vss.n13236 vss.n13235 1.19376
R39236 vss.n13954 vss.n13953 1.19376
R39237 vss.n14029 vss.n14028 1.19376
R39238 vss.n1981 vss.n1980 1.19376
R39239 vss.n13200 vss.n13158 1.19376
R39240 vss.n8974 vss.n7472 1.19376
R39241 vss.n8863 vss.n7544 1.19376
R39242 vss.n8855 vss.n7661 1.19376
R39243 vss.n8744 vss.n7687 1.19376
R39244 vss.n8736 vss.n7848 1.19376
R39245 vss.n8254 vss.n8253 1.19376
R39246 vss.n8245 vss.n7991 1.19376
R39247 vss.n9252 vss.n9251 1.19376
R39248 vss.n7030 vss.n7029 1.19376
R39249 vss.n7089 vss.n7088 1.19376
R39250 vss.n7221 vss.n7220 1.19376
R39251 vss.n9503 vss.n9502 1.19376
R39252 vss.n9578 vss.n9577 1.19376
R39253 vss.n9193 vss.n9192 1.19376
R39254 vss.n9367 vss.n2028 1.19376
R39255 vss.n9844 vss.n2871 1.19376
R39256 vss.n5323 vss.n5322 1.19376
R39257 vss.n5314 vss.n5272 1.19376
R39258 vss.n5264 vss.n5263 1.19376
R39259 vss.n5255 vss.n5213 1.19376
R39260 vss.n9793 vss.n3026 1.19376
R39261 vss.n9785 vss.n9743 1.19376
R39262 vss.n9990 vss.n2029 1.19376
R39263 vss.n5787 vss.n5786 1.19376
R39264 vss.n5844 vss.n5843 1.19376
R39265 vss.n4120 vss.n4119 1.19376
R39266 vss.n4069 vss.n4068 1.19376
R39267 vss.n4211 vss.n4210 1.19376
R39268 vss.n4614 vss.n4411 1.19376
R39269 vss.n4504 vss.n4503 1.19376
R39270 vss.n12320 vss.n12278 1.19376
R39271 vss.n12536 vss.n12535 1.19376
R39272 vss.n12450 vss.n12408 1.19376
R39273 vss.n12901 vss.n12859 1.19376
R39274 vss.n12910 vss.n12909 1.19376
R39275 vss.n12965 vss.n2399 1.19376
R39276 vss.n13018 vss.n2240 1.19376
R39277 vss.n11968 vss.n11967 1.19376
R39278 vss.n12615 vss.n12614 1.19376
R39279 vss.n11594 vss.n11593 1.19376
R39280 vss.n11544 vss.n11543 1.19376
R39281 vss.n10992 vss.n10991 1.19376
R39282 vss.n11449 vss.n11446 1.19376
R39283 vss.n12697 vss.n12696 1.19376
R39284 vss.n13149 vss.n13148 1.19376
R39285 vss.n9730 vss.n9729 1.11974
R39286 vss.n9632 vss.n9631 1.11974
R39287 vss.n14091 vss.n14090 1.11974
R39288 vss.n14033 vss 1.0778
R39289 vss vss.n1487 1.0778
R39290 vss vss.n9582 1.0778
R39291 vss.n6983 vss 1.0778
R39292 vss.n4073 vss 1.0778
R39293 vss vss.n5934 1.0778
R39294 vss.n11548 vss 1.0778
R39295 vss.n11149 vss 1.0778
R39296 vss.n13055 vss.n2159 1.05976
R39297 vss vss.n14446 1.04491
R39298 vss vss.n8740 1.04491
R39299 vss vss.n5259 1.04491
R39300 vss vss.n10298 1.04491
R39301 vss.n13022 vss 1.02517
R39302 vss.n8978 vss 1.02517
R39303 vss.n9848 vss 1.02517
R39304 vss.n14761 vss 1.02517
R39305 vss.n1404 vss 0.887013
R39306 vss.n13236 vss 0.887013
R39307 vss.n14028 vss 0.887013
R39308 vss.n1980 vss 0.887013
R39309 vss.n7030 vss 0.887013
R39310 vss.n7221 vss 0.887013
R39311 vss.n9577 vss 0.887013
R39312 vss.n9193 vss 0.887013
R39313 vss.n5787 vss 0.887013
R39314 vss.n4120 vss 0.887013
R39315 vss.n4210 vss 0.887013
R39316 vss.n4504 vss 0.887013
R39317 vss.n11968 vss 0.887013
R39318 vss.n11594 vss 0.887013
R39319 vss.n10991 vss 0.887013
R39320 vss.n12697 vss 0.887013
R39321 vss.n12614 vss 0.854118
R39322 vss.n11543 vss 0.854118
R39323 vss vss.n11449 0.854118
R39324 vss vss.n290 0.854118
R39325 vss vss.n231 0.854118
R39326 vss vss.n154 0.854118
R39327 vss vss.n413 0.854118
R39328 vss vss.n1806 0.854118
R39329 vss vss.n1910 0.854118
R39330 vss vss.n13954 0.854118
R39331 vss vss.n7472 0.854118
R39332 vss vss.n7661 0.854118
R39333 vss vss.n7848 0.854118
R39334 vss.n7991 vss 0.854118
R39335 vss.n7088 vss 0.854118
R39336 vss.n9251 vss 0.854118
R39337 vss vss.n9503 0.854118
R39338 vss vss.n2871 0.854118
R39339 vss.n5272 vss 0.854118
R39340 vss.n5213 vss 0.854118
R39341 vss.n9743 vss 0.854118
R39342 vss.n5843 vss 0.854118
R39343 vss.n4068 vss 0.854118
R39344 vss vss.n4614 0.854118
R39345 vss vss.n2240 0.854118
R39346 vss vss.n12536 0.854118
R39347 vss.n12859 vss 0.854118
R39348 vss vss.n2399 0.854118
R39349 vss vss.n198 0.821224
R39350 vss vss.n257 0.821224
R39351 vss vss.n316 0.821224
R39352 vss.n8254 vss 0.821224
R39353 vss vss.n7687 0.821224
R39354 vss vss.n7544 0.821224
R39355 vss vss.n3026 0.821224
R39356 vss.n5264 vss 0.821224
R39357 vss.n5323 vss 0.821224
R39358 vss vss.n12910 0.821224
R39359 vss.n12408 vss 0.821224
R39360 vss.n12278 vss 0.821224
R39361 vss.n13549 vss.n413 0.697868
R39362 vss.n13650 vss.n316 0.697868
R39363 vss.n13702 vss.n290 0.697868
R39364 vss.n13755 vss.n257 0.697868
R39365 vss.n13807 vss.n231 0.697868
R39366 vss.n13860 vss.n198 0.697868
R39367 vss.n13318 vss.n154 0.697868
R39368 vss.n1910 vss.n1909 0.697868
R39369 vss.n1404 vss.n1403 0.697868
R39370 vss.n1806 vss.n1805 0.697868
R39371 vss.n13237 vss.n13236 0.697868
R39372 vss.n13954 vss.n593 0.697868
R39373 vss.n14028 vss.n14027 0.697868
R39374 vss.n13158 vss.n13157 0.697868
R39375 vss.n1980 vss.n1979 0.697868
R39376 vss.n8057 vss.n7991 0.697868
R39377 vss.n7871 vss.n7848 0.697868
R39378 vss.n8402 vss.n7661 0.697868
R39379 vss.n8500 vss.n7472 0.697868
R39380 vss.n8471 vss.n7544 0.697868
R39381 vss.n8373 vss.n7687 0.697868
R39382 vss.n8255 vss.n8254 0.697868
R39383 vss.n9251 vss.n9250 0.697868
R39384 vss.n7031 vss.n7030 0.697868
R39385 vss.n7088 vss.n7087 0.697868
R39386 vss.n7222 vss.n7221 0.697868
R39387 vss.n9503 vss.n6133 0.697868
R39388 vss.n9577 vss.n9576 0.697868
R39389 vss.n6543 vss.n2028 0.697868
R39390 vss.n9194 vss.n9193 0.697868
R39391 vss.n9743 vss.n3262 0.697868
R39392 vss.n5213 vss.n5205 0.697868
R39393 vss.n5272 vss.n5081 0.697868
R39394 vss.n5353 vss.n2871 0.697868
R39395 vss.n5324 vss.n5323 0.697868
R39396 vss.n5265 vss.n5264 0.697868
R39397 vss.n5206 vss.n3026 0.697868
R39398 vss.n3599 vss.n2029 0.697868
R39399 vss.n5788 vss.n5787 0.697868
R39400 vss.n5843 vss.n5842 0.697868
R39401 vss.n4121 vss.n4120 0.697868
R39402 vss.n4068 vss.n4067 0.697868
R39403 vss.n4210 vss.n4209 0.697868
R39404 vss.n4614 vss.n4613 0.697868
R39405 vss.n4505 vss.n4504 0.697868
R39406 vss.n12859 vss.n10299 0.697868
R39407 vss.n12536 vss.n11737 0.697868
R39408 vss.n12278 vss.n11779 0.697868
R39409 vss.n12408 vss.n12405 0.697868
R39410 vss.n12910 vss.n10101 0.697868
R39411 vss.n10064 vss.n2399 0.697868
R39412 vss.n11833 vss.n2240 0.697868
R39413 vss.n13149 vss.n2030 0.697868
R39414 vss.n11969 vss.n11968 0.697868
R39415 vss.n12614 vss.n12613 0.697868
R39416 vss.n11595 vss.n11594 0.697868
R39417 vss.n11543 vss.n11542 0.697868
R39418 vss.n10991 vss.n10990 0.697868
R39419 vss.n11449 vss.n11448 0.697868
R39420 vss.n12698 vss.n12697 0.697868
R39421 vss.n643 vss 0.672375
R39422 vss.n1091 vss 0.672375
R39423 vss.n1484 vss 0.672375
R39424 vss.n1565 vss 0.672375
R39425 vss.n6051 vss 0.672375
R39426 vss.n6366 vss 0.672375
R39427 vss.n6980 vss 0.672375
R39428 vss.n7169 vss 0.672375
R39429 vss.n3423 vss 0.672375
R39430 vss.n4020 vss 0.672375
R39431 vss.n4287 vss 0.672375
R39432 vss.n5931 vss 0.672375
R39433 vss.n10502 vss 0.672375
R39434 vss.n10723 vss 0.672375
R39435 vss.n11037 vss 0.672375
R39436 vss.n11146 vss 0.672375
R39437 vss.n14412 vss 0.606586
R39438 vss.n14607 vss 0.606586
R39439 vss.n359 vss 0.606586
R39440 vss.n7587 vss 0.606586
R39441 vss.n7730 vss 0.606586
R39442 vss.n7951 vss 0.606586
R39443 vss.n4964 vss 0.606586
R39444 vss.n5166 vss 0.606586
R39445 vss.n3147 vss 0.606586
R39446 vss.n12365 vss 0.606586
R39447 vss.n10261 vss 0.606586
R39448 vss.n2441 vss 0.606586
R39449 vss.n7497 vss 0.588493
R39450 vss.n2924 vss 0.588493
R39451 vss.n2265 vss 0.588493
R39452 vss vss.n14793 0.588493
R39453 vss.n11401 vss 0.431421
R39454 vss.n10769 vss 0.431421
R39455 vss.n10548 vss 0.431421
R39456 vss.n14033 vss 0.431421
R39457 vss.n1649 vss 0.431421
R39458 vss.n1357 vss 0.431421
R39459 vss.n1094 vss 0.431421
R39460 vss.n1356 vss 0.431421
R39461 vss.n1408 vss 0.431421
R39462 vss.n1487 vss 0.431421
R39463 vss vss.n1650 0.431421
R39464 vss.n1571 vss 0.431421
R39465 vss.n1570 vss 0.431421
R39466 vss.n1569 vss 0.431421
R39467 vss vss.n515 0.431421
R39468 vss.n14032 vss 0.431421
R39469 vss.n1984 vss 0.431421
R39470 vss.n13203 vss 0.431421
R39471 vss.n9582 vss 0.431421
R39472 vss.n7093 vss 0.431421
R39473 vss.n6446 vss 0.431421
R39474 vss.n9256 vss 0.431421
R39475 vss.n9255 vss 0.431421
R39476 vss vss.n6984 0.431421
R39477 vss.n6983 vss 0.431421
R39478 vss.n7092 vss 0.431421
R39479 vss vss.n7175 0.431421
R39480 vss.n7174 vss 0.431421
R39481 vss.n7173 vss 0.431421
R39482 vss vss.n6054 0.431421
R39483 vss.n9581 vss 0.431421
R39484 vss vss.n6213 0.431421
R39485 vss.n9364 vss 0.431421
R39486 vss.n4365 vss 0.431421
R39487 vss.n3720 vss 0.431421
R39488 vss.n3500 vss 0.431421
R39489 vss.n9993 vss 0.431421
R39490 vss vss.n2630 0.431421
R39491 vss.n5848 vss 0.431421
R39492 vss.n5847 vss 0.431421
R39493 vss vss.n4074 0.431421
R39494 vss.n4073 vss 0.431421
R39495 vss.n4072 vss 0.431421
R39496 vss.n4214 vss 0.431421
R39497 vss.n4290 vss 0.431421
R39498 vss vss.n4366 0.431421
R39499 vss vss.n3307 0.431421
R39500 vss.n5934 vss 0.431421
R39501 vss.n12620 vss 0.431421
R39502 vss.n12619 vss 0.431421
R39503 vss.n12618 vss 0.431421
R39504 vss vss.n11549 0.431421
R39505 vss.n11548 vss 0.431421
R39506 vss.n11547 vss 0.431421
R39507 vss.n10995 vss 0.431421
R39508 vss.n11040 vss 0.431421
R39509 vss vss.n11402 0.431421
R39510 vss.n11042 vss 0.431421
R39511 vss.n11149 vss 0.431421
R39512 vss.n12665 vss 0.431421
R39513 vss vss.n412 0.398526
R39514 vss vss.n289 0.398526
R39515 vss vss.n14252 0.398526
R39516 vss.n14369 vss 0.398526
R39517 vss.n14446 vss 0.398526
R39518 vss vss.n230 0.398526
R39519 vss.n14447 vss 0.398526
R39520 vss vss.n14447 0.398526
R39521 vss.n14564 vss 0.398526
R39522 vss.n14641 vss 0.398526
R39523 vss vss.n153 0.398526
R39524 vss vss.n14642 0.398526
R39525 vss.n14759 vss 0.398526
R39526 vss.n14251 vss 0.398526
R39527 vss.n14250 vss 0.398526
R39528 vss vss.n14093 0.398526
R39529 vss vss.n6006 0.398526
R39530 vss.n7847 vss 0.398526
R39531 vss vss.n7660 0.398526
R39532 vss vss.n7471 0.398526
R39533 vss.n8978 vss 0.398526
R39534 vss.n8977 vss 0.398526
R39535 vss vss.n8860 0.398526
R39536 vss.n8859 vss 0.398526
R39537 vss.n8858 vss 0.398526
R39538 vss vss.n8741 0.398526
R39539 vss.n8741 vss 0.398526
R39540 vss.n8740 vss 0.398526
R39541 vss.n8739 vss 0.398526
R39542 vss vss.n8250 0.398526
R39543 vss.n8249 vss 0.398526
R39544 vss.n8248 vss 0.398526
R39545 vss vss.n9634 0.398526
R39546 vss.n3261 vss 0.398526
R39547 vss.n3104 vss 0.398526
R39548 vss.n5078 vss 0.398526
R39549 vss vss.n2870 0.398526
R39550 vss.n9848 vss 0.398526
R39551 vss.n9847 vss 0.398526
R39552 vss vss.n5319 0.398526
R39553 vss.n5318 vss 0.398526
R39554 vss.n5317 vss 0.398526
R39555 vss vss.n5260 0.398526
R39556 vss.n5260 vss 0.398526
R39557 vss.n5259 vss 0.398526
R39558 vss.n5258 vss 0.398526
R39559 vss vss.n9790 0.398526
R39560 vss.n9789 vss 0.398526
R39561 vss.n9788 vss 0.398526
R39562 vss vss.n9732 0.398526
R39563 vss.n12905 vss 0.398526
R39564 vss.n12531 vss 0.398526
R39565 vss vss.n2239 0.398526
R39566 vss.n12323 vss 0.398526
R39567 vss.n12402 vss 0.398526
R39568 vss vss.n12532 0.398526
R39569 vss.n12453 vss 0.398526
R39570 vss.n12453 vss 0.398526
R39571 vss.n10298 vss 0.398526
R39572 vss.n12904 vss 0.398526
R39573 vss vss.n12906 0.398526
R39574 vss.n2478 vss 0.398526
R39575 vss vss.n12962 0.398526
R39576 vss.n12961 vss 0.398526
R39577 vss.n12960 vss 0.398526
R39578 vss.n13022 vss 0.398526
R39579 vss.n13021 vss 0.398526
R39580 vss.n14761 vss 0.398526
R39581 vss.n1650 vss 0.365632
R39582 vss.n7092 vss 0.365632
R39583 vss vss.n4072 0.365632
R39584 vss vss.n11547 0.365632
R39585 vss.n11400 vss.n11399 0.317934
R39586 vss.n10768 vss.n10767 0.317934
R39587 vss.n10547 vss.n10546 0.317934
R39588 vss.n11971 vss.n11970 0.317934
R39589 vss.n12014 vss.n12013 0.317934
R39590 vss.n11597 vss.n11596 0.317934
R39591 vss.n10844 vss.n10843 0.317934
R39592 vss.n10989 vss.n10988 0.317934
R39593 vss.n11451 vss.n11450 0.317934
R39594 vss.n12700 vss.n12699 0.317934
R39595 vss.n1978 vss.n1977 0.317934
R39596 vss.n14182 vss.n14181 0.317934
R39597 vss.n13551 vss.n13550 0.317934
R39598 vss.n13370 vss.n13369 0.317934
R39599 vss.n13450 vss.n13449 0.317934
R39600 vss.n13530 vss.n13529 0.317934
R39601 vss.n14301 vss.n14300 0.317934
R39602 vss.n14254 vss.n14253 0.317934
R39603 vss.n13652 vss.n13651 0.317934
R39604 vss.n13648 vss.n13647 0.317934
R39605 vss.n13704 vss.n13703 0.317934
R39606 vss.n14368 vss.n14367 0.317934
R39607 vss.n14414 vss.n14413 0.317934
R39608 vss.n14496 vss.n14495 0.317934
R39609 vss.n14449 vss.n14448 0.317934
R39610 vss.n13757 vss.n13756 0.317934
R39611 vss.n13753 vss.n13752 0.317934
R39612 vss.n13809 vss.n13808 0.317934
R39613 vss.n14563 vss.n14562 0.317934
R39614 vss.n14609 vss.n14608 0.317934
R39615 vss.n14691 vss.n14690 0.317934
R39616 vss.n14644 vss.n14643 0.317934
R39617 vss.n13862 vss.n13861 0.317934
R39618 vss.n13858 vss.n13857 0.317934
R39619 vss.n14758 vss.n14757 0.317934
R39620 vss.n13320 vss.n13319 0.317934
R39621 vss.n361 vss.n360 0.317934
R39622 vss.n14249 vss.n14248 0.317934
R39623 vss.n14144 vss.n14143 0.317934
R39624 vss.n14141 vss.n14140 0.317934
R39625 vss.n14095 vss.n14094 0.317934
R39626 vss.n642 vss.n641 0.317934
R39627 vss.n13239 vss.n13238 0.317934
R39628 vss.n1808 vss.n1807 0.317934
R39629 vss.n1648 vss.n1647 0.317934
R39630 vss.n1402 vss.n1401 0.317934
R39631 vss.n1912 vss.n1911 0.317934
R39632 vss.n1353 vss.n1352 0.317934
R39633 vss.n1093 vss.n1092 0.317934
R39634 vss.n1355 vss.n1354 0.317934
R39635 vss.n1908 vss.n1907 0.317934
R39636 vss.n1400 vss.n1399 0.317934
R39637 vss.n1407 vss.n1406 0.317934
R39638 vss.n1486 vss.n1485 0.317934
R39639 vss.n1652 vss.n1651 0.317934
R39640 vss.n1804 vss.n1803 0.317934
R39641 vss.n1696 vss.n1695 0.317934
R39642 vss.n1488 vss.n793 0.317934
R39643 vss.n1567 vss.n1566 0.317934
R39644 vss.n554 vss.n553 0.317934
R39645 vss.n592 vss.n555 0.317934
R39646 vss.n13956 vss.n13955 0.317934
R39647 vss.n1568 vss.n594 0.317934
R39648 vss.n891 vss.n890 0.317934
R39649 vss.n14031 vss.n14030 0.317934
R39650 vss.n14026 vss.n14025 0.317934
R39651 vss.n13156 vss.n706 0.317934
R39652 vss.n1136 vss.n705 0.317934
R39653 vss.n1983 vss.n1982 0.317934
R39654 vss.n2027 vss.n2026 0.317934
R39655 vss.n13202 vss.n13201 0.317934
R39656 vss.n9196 vss.n9195 0.317934
R39657 vss.n8059 vss.n8058 0.317934
R39658 vss.n8180 vss.n8179 0.317934
R39659 vss.n7811 vss.n7810 0.317934
R39660 vss.n8790 vss.n8789 0.317934
R39661 vss.n7908 vss.n7907 0.317934
R39662 vss.n7873 vss.n7872 0.317934
R39663 vss.n8329 vss.n8328 0.317934
R39664 vss.n8404 vss.n8403 0.317934
R39665 vss.n8427 vss.n8426 0.317934
R39666 vss.n8502 vss.n8501 0.317934
R39667 vss.n8909 vss.n8908 0.317934
R39668 vss.n7496 vss.n7495 0.317934
R39669 vss.n8976 vss.n8975 0.317934
R39670 vss.n8476 vss.n8475 0.317934
R39671 vss.n8473 vss.n8472 0.317934
R39672 vss.n8862 vss.n8861 0.317934
R39673 vss.n7589 vss.n7588 0.317934
R39674 vss.n8857 vss.n8856 0.317934
R39675 vss.n8378 vss.n8377 0.317934
R39676 vss.n8375 vss.n8374 0.317934
R39677 vss.n8743 vss.n8742 0.317934
R39678 vss.n7732 vss.n7731 0.317934
R39679 vss.n8738 vss.n8737 0.317934
R39680 vss.n7905 vss.n7904 0.317934
R39681 vss.n8257 vss.n8256 0.317934
R39682 vss.n8252 vss.n8251 0.317934
R39683 vss.n7953 vss.n7952 0.317934
R39684 vss.n8247 vss.n8246 0.317934
R39685 vss.n7990 vss.n7989 0.317934
R39686 vss.n9640 vss.n9639 0.317934
R39687 vss.n9636 vss.n9635 0.317934
R39688 vss.n6053 vss.n6052 0.317934
R39689 vss.n7224 vss.n7223 0.317934
R39690 vss.n7050 vss.n7049 0.317934
R39691 vss.n6672 vss.n6671 0.317934
R39692 vss.n7033 vss.n7032 0.317934
R39693 vss.n9213 vss.n9212 0.317934
R39694 vss.n6445 vss.n6444 0.317934
R39695 vss.n6368 vss.n6367 0.317934
R39696 vss.n9254 vss.n9253 0.317934
R39697 vss.n9249 vss.n9248 0.317934
R39698 vss.n6904 vss.n6903 0.317934
R39699 vss.n6986 vss.n6985 0.317934
R39700 vss.n6982 vss.n6981 0.317934
R39701 vss.n7091 vss.n7090 0.317934
R39702 vss.n7086 vss.n7085 0.317934
R39703 vss.n6716 vss.n6715 0.317934
R39704 vss.n7177 vss.n7176 0.317934
R39705 vss.n7171 vss.n7170 0.317934
R39706 vss.n6094 vss.n6093 0.317934
R39707 vss.n6132 vss.n6095 0.317934
R39708 vss.n9505 vss.n9504 0.317934
R39709 vss.n7172 vss.n6134 0.317934
R39710 vss.n9429 vss.n9428 0.317934
R39711 vss.n9580 vss.n9579 0.317934
R39712 vss.n9575 vss.n9574 0.317934
R39713 vss.n6545 vss.n6544 0.317934
R39714 vss.n9147 vss.n9146 0.317934
R39715 vss.n9149 vss.n9148 0.317934
R39716 vss.n9363 vss.n9362 0.317934
R39717 vss.n9366 vss.n9365 0.317934
R39718 vss.n3226 vss.n3225 0.317934
R39719 vss.n3069 vss.n3068 0.317934
R39720 vss.n5043 vss.n5042 0.317934
R39721 vss.n4642 vss.n4641 0.317934
R39722 vss.n4633 vss.n4632 0.317934
R39723 vss.n5204 vss.n5203 0.317934
R39724 vss.n5083 vss.n5082 0.317934
R39725 vss.n5080 vss.n5079 0.317934
R39726 vss.n4881 vss.n4880 0.317934
R39727 vss.n5355 vss.n5354 0.317934
R39728 vss.n2970 vss.n2969 0.317934
R39729 vss.n2923 vss.n2922 0.317934
R39730 vss.n9846 vss.n9845 0.317934
R39731 vss.n5329 vss.n5328 0.317934
R39732 vss.n5326 vss.n5325 0.317934
R39733 vss.n5321 vss.n5320 0.317934
R39734 vss.n4966 vss.n4965 0.317934
R39735 vss.n5316 vss.n5315 0.317934
R39736 vss.n5271 vss.n5270 0.317934
R39737 vss.n5267 vss.n5266 0.317934
R39738 vss.n5262 vss.n5261 0.317934
R39739 vss.n5168 vss.n5167 0.317934
R39740 vss.n5257 vss.n5256 0.317934
R39741 vss.n5212 vss.n5211 0.317934
R39742 vss.n5208 vss.n5207 0.317934
R39743 vss.n9792 vss.n9791 0.317934
R39744 vss.n3149 vss.n3148 0.317934
R39745 vss.n9787 vss.n9786 0.317934
R39746 vss.n9742 vss.n9741 0.317934
R39747 vss.n9738 vss.n9737 0.317934
R39748 vss.n9734 vss.n9733 0.317934
R39749 vss.n4364 vss.n4363 0.317934
R39750 vss.n3719 vss.n3718 0.317934
R39751 vss.n3499 vss.n3498 0.317934
R39752 vss.n5790 vss.n5789 0.317934
R39753 vss.n3579 vss.n3578 0.317934
R39754 vss.n4123 vss.n4122 0.317934
R39755 vss.n4065 vss.n3855 0.317934
R39756 vss.n4208 vss.n4207 0.317934
R39757 vss.n4616 vss.n4615 0.317934
R39758 vss.n4507 vss.n4506 0.317934
R39759 vss.n2673 vss.n2672 0.317934
R39760 vss.n9992 vss.n9991 0.317934
R39761 vss.n3601 vss.n3600 0.317934
R39762 vss.n5741 vss.n5740 0.317934
R39763 vss.n5743 vss.n5742 0.317934
R39764 vss.n3425 vss.n3424 0.317934
R39765 vss.n5846 vss.n5845 0.317934
R39766 vss.n5841 vss.n5840 0.317934
R39767 vss.n3947 vss.n3946 0.317934
R39768 vss.n4076 vss.n4075 0.317934
R39769 vss.n4022 vss.n4021 0.317934
R39770 vss.n4071 vss.n4070 0.317934
R39771 vss.n4066 vss.n3802 0.317934
R39772 vss.n3801 vss.n3800 0.317934
R39773 vss.n4213 vss.n4212 0.317934
R39774 vss.n4289 vss.n4288 0.317934
R39775 vss.n4368 vss.n4367 0.317934
R39776 vss.n4612 vss.n4611 0.317934
R39777 vss.n4458 vss.n4457 0.317934
R39778 vss.n4460 vss.n4459 0.317934
R39779 vss.n5933 vss.n5932 0.317934
R39780 vss.n10012 vss.n10011 0.317934
R39781 vss.n5935 vss.n2557 0.317934
R39782 vss.n9684 vss.n9683 0.317934
R39783 vss.n9583 vss.n5936 0.317934
R39784 vss.n9630 vss.n9629 0.317934
R39785 vss.n9585 vss.n9584 0.317934
R39786 vss.n14089 vss.n14088 0.317934
R39787 vss.n12912 vss.n12911 0.317934
R39788 vss.n11676 vss.n11675 0.317934
R39789 vss.n10185 vss.n10184 0.317934
R39790 vss.n12407 vss.n12406 0.317934
R39791 vss.n12241 vss.n12240 0.317934
R39792 vss.n12496 vss.n12495 0.317934
R39793 vss.n2340 vss.n2339 0.317934
R39794 vss.n12277 vss.n12276 0.317934
R39795 vss.n12142 vss.n12141 0.317934
R39796 vss.n12139 vss.n12138 0.317934
R39797 vss.n12322 vss.n12321 0.317934
R39798 vss.n12367 vss.n12366 0.317934
R39799 vss.n12534 vss.n12533 0.317934
R39800 vss.n12538 vss.n12537 0.317934
R39801 vss.n12404 vss.n12403 0.317934
R39802 vss.n12452 vss.n12451 0.317934
R39803 vss.n10263 vss.n10262 0.317934
R39804 vss.n12903 vss.n12902 0.317934
R39805 vss.n12858 vss.n12857 0.317934
R39806 vss.n10301 vss.n10300 0.317934
R39807 vss.n12908 vss.n12907 0.317934
R39808 vss.n2443 vss.n2442 0.317934
R39809 vss.n12955 vss.n12954 0.317934
R39810 vss.n10016 vss.n10015 0.317934
R39811 vss.n10066 vss.n10065 0.317934
R39812 vss.n12964 vss.n12963 0.317934
R39813 vss.n2522 vss.n2521 0.317934
R39814 vss.n12959 vss.n12958 0.317934
R39815 vss.n2264 vss.n2263 0.317934
R39816 vss.n13020 vss.n13019 0.317934
R39817 vss.n11835 vss.n11834 0.317934
R39818 vss.n11890 vss.n11889 0.317934
R39819 vss.n11923 vss.n11891 0.317934
R39820 vss.n11925 vss.n11924 0.317934
R39821 vss.n10504 vss.n10503 0.317934
R39822 vss.n12617 vss.n12616 0.317934
R39823 vss.n12612 vss.n12611 0.317934
R39824 vss.n10680 vss.n10679 0.317934
R39825 vss.n11551 vss.n11550 0.317934
R39826 vss.n10725 vss.n10724 0.317934
R39827 vss.n11546 vss.n11545 0.317934
R39828 vss.n11541 vss.n11540 0.317934
R39829 vss.n10975 vss.n10974 0.317934
R39830 vss.n10994 vss.n10993 0.317934
R39831 vss.n11039 vss.n11038 0.317934
R39832 vss.n11404 vss.n11403 0.317934
R39833 vss.n11447 vss.n10339 0.317934
R39834 vss.n10372 vss.n10340 0.317934
R39835 vss.n11041 vss.n10373 0.317934
R39836 vss.n11148 vss.n11147 0.317934
R39837 vss.n12663 vss.n12662 0.317934
R39838 vss.n12664 vss.n2031 0.317934
R39839 vss.n14760 vss.n0 0.317934
R39840 vss.n11150 vss.n11104 0.310177
R39841 vss.n11357 vss.n11356 0.310177
R39842 vss.n11231 vss.n11230 0.310177
R39843 vss.n11292 vss.n11291 0.310177
R39844 vss.n14763 vss.n14762 0.310177
R39845 vss.n411 vss.n381 0.310177
R39846 vss.n288 vss.n258 0.310177
R39847 vss.n14445 vss.n14415 0.310177
R39848 vss.n229 vss.n199 0.310177
R39849 vss.n14640 vss.n14610 0.310177
R39850 vss.n152 vss.n122 0.310177
R39851 vss.n380 vss.n378 0.310177
R39852 vss.n7374 vss.n7373 0.310177
R39853 vss.n7846 vss.n7812 0.310177
R39854 vss.n7659 vss.n7625 0.310177
R39855 vss.n7470 vss.n7436 0.310177
R39856 vss.n8980 vss.n8979 0.310177
R39857 vss.n7624 vss.n7590 0.310177
R39858 vss.n7767 vss.n7733 0.310177
R39859 vss.n7988 vss.n7954 0.310177
R39860 vss.n3260 vss.n3227 0.310177
R39861 vss.n3103 vss.n3070 0.310177
R39862 vss.n5077 vss.n5044 0.310177
R39863 vss.n2869 vss.n2836 0.310177
R39864 vss.n9853 vss.n9849 0.310177
R39865 vss.n5000 vss.n4967 0.310177
R39866 vss.n5202 vss.n5169 0.310177
R39867 vss.n3183 vss.n3150 0.310177
R39868 vss.n10219 vss.n10186 0.310177
R39869 vss.n12530 vss.n12497 0.310177
R39870 vss.n2238 vss.n2205 0.310177
R39871 vss.n12401 vss.n12368 0.310177
R39872 vss.n10297 vss.n10264 0.310177
R39873 vss.n2477 vss.n2444 0.310177
R39874 vss.n2556 vss.n2523 0.310177
R39875 vss.n13040 vss.n13023 0.310177
R39876 vss.n11308 vss.n10460 0.310177
R39877 vss.n11247 vss.n10681 0.310177
R39878 vss.n11200 vss.n11199 0.310177
R39879 vss.n12666 vss.n10459 0.310177
R39880 vss.n11399 vss.n11398 0.271061
R39881 vss.n10767 vss.n10766 0.271061
R39882 vss.n10546 vss.n10545 0.271061
R39883 vss.n11972 vss.n11971 0.271061
R39884 vss.n12015 vss.n12014 0.271061
R39885 vss.n11598 vss.n11597 0.271061
R39886 vss.n10848 vss.n10844 0.271061
R39887 vss.n10988 vss.n10987 0.271061
R39888 vss.n11452 vss.n11451 0.271061
R39889 vss.n12701 vss.n12700 0.271061
R39890 vss.n1977 vss.n1976 0.271061
R39891 vss.n14183 vss.n14182 0.271061
R39892 vss.n13552 vss.n13551 0.271061
R39893 vss.n13371 vss.n13370 0.271061
R39894 vss.n13451 vss.n13450 0.271061
R39895 vss.n13531 vss.n13530 0.271061
R39896 vss.n14302 vss.n14301 0.271061
R39897 vss.n13705 vss.n13704 0.271061
R39898 vss.n14497 vss.n14496 0.271061
R39899 vss.n13810 vss.n13809 0.271061
R39900 vss.n14692 vss.n14691 0.271061
R39901 vss.n13912 vss.n13320 0.271061
R39902 vss.n13240 vss.n13239 0.271061
R39903 vss.n1809 vss.n1808 0.271061
R39904 vss.n1647 vss.n1646 0.271061
R39905 vss.n1401 vss.n1245 0.271061
R39906 vss.n1913 vss.n1912 0.271061
R39907 vss.n1352 vss.n1351 0.271061
R39908 vss.n13957 vss.n13956 0.271061
R39909 vss.n892 vss.n891 0.271061
R39910 vss.n14025 vss.n14024 0.271061
R39911 vss.n2026 vss.n2025 0.271061
R39912 vss.n9197 vss.n9196 0.271061
R39913 vss.n8060 vss.n8059 0.271061
R39914 vss.n8181 vss.n8180 0.271061
R39915 vss.n7810 vss.n7809 0.271061
R39916 vss.n8791 vss.n8790 0.271061
R39917 vss.n7907 vss.n7272 0.271061
R39918 vss.n7874 vss.n7873 0.271061
R39919 vss.n8330 vss.n8329 0.271061
R39920 vss.n8405 vss.n8404 0.271061
R39921 vss.n8428 vss.n8427 0.271061
R39922 vss.n8503 vss.n8502 0.271061
R39923 vss.n8910 vss.n8909 0.271061
R39924 vss.n7225 vss.n7224 0.271061
R39925 vss.n7051 vss.n7050 0.271061
R39926 vss.n6671 vss.n6670 0.271061
R39927 vss.n7034 vss.n7033 0.271061
R39928 vss.n9214 vss.n9213 0.271061
R39929 vss.n6444 vss.n6443 0.271061
R39930 vss.n9506 vss.n9505 0.271061
R39931 vss.n9430 vss.n9429 0.271061
R39932 vss.n9574 vss.n9573 0.271061
R39933 vss.n9362 vss.n9361 0.271061
R39934 vss.n3225 vss.n3224 0.271061
R39935 vss.n3068 vss.n3067 0.271061
R39936 vss.n5042 vss.n5041 0.271061
R39937 vss.n4643 vss.n4642 0.271061
R39938 vss.n4634 vss.n4633 0.271061
R39939 vss.n5203 vss.n4730 0.271061
R39940 vss.n5082 vss.n4751 0.271061
R39941 vss.n5079 vss.n4816 0.271061
R39942 vss.n4880 vss.n4837 0.271061
R39943 vss.n5356 vss.n5355 0.271061
R39944 vss.n2971 vss.n2970 0.271061
R39945 vss.n4363 vss.n4362 0.271061
R39946 vss.n3718 vss.n3717 0.271061
R39947 vss.n3498 vss.n3497 0.271061
R39948 vss.n5791 vss.n5790 0.271061
R39949 vss.n5806 vss.n3579 0.271061
R39950 vss.n4124 vss.n4123 0.271061
R39951 vss.n4139 vss.n3855 0.271061
R39952 vss.n4207 vss.n4206 0.271061
R39953 vss.n4617 vss.n4616 0.271061
R39954 vss.n4508 vss.n4507 0.271061
R39955 vss.n2674 vss.n2673 0.271061
R39956 vss.n12913 vss.n12912 0.271061
R39957 vss.n11677 vss.n11676 0.271061
R39958 vss.n10184 vss.n10183 0.271061
R39959 vss.n12406 vss.n11628 0.271061
R39960 vss.n12242 vss.n12241 0.271061
R39961 vss.n12495 vss.n12494 0.271061
R39962 vss.n2341 vss.n2340 0.271061
R39963 vss.n12276 vss.n12275 0.271061
R39964 vss.n10067 vss.n10066 0.271061
R39965 vss.n2521 vss.n2520 0.271061
R39966 vss.n11836 vss.n11835 0.271061
R39967 vss.n12662 vss.n12661 0.271061
R39968 vss.n14255 vss.n14254 0.271059
R39969 vss.n13653 vss.n13652 0.271059
R39970 vss.n13649 vss.n13648 0.271059
R39971 vss.n14367 vss.n14366 0.271059
R39972 vss.n14413 vss.n14412 0.271059
R39973 vss.n14450 vss.n14449 0.271059
R39974 vss.n13758 vss.n13757 0.271059
R39975 vss.n13754 vss.n13753 0.271059
R39976 vss.n14562 vss.n14561 0.271059
R39977 vss.n14608 vss.n14607 0.271059
R39978 vss.n14645 vss.n14644 0.271059
R39979 vss.n13863 vss.n13862 0.271059
R39980 vss.n13859 vss.n13858 0.271059
R39981 vss.n14757 vss.n14756 0.271059
R39982 vss.n360 vss.n359 0.271059
R39983 vss.n14248 vss.n14247 0.271059
R39984 vss.n14145 vss.n14144 0.271059
R39985 vss.n14142 vss.n14141 0.271059
R39986 vss.n14138 vss.n14095 0.271059
R39987 vss.n643 vss.n642 0.271059
R39988 vss.n1092 vss.n1091 0.271059
R39989 vss.n1354 vss.n1200 0.271059
R39990 vss.n1907 vss.n1906 0.271059
R39991 vss.n1399 vss.n1201 0.271059
R39992 vss.n1406 vss.n1405 0.271059
R39993 vss.n1485 vss.n1484 0.271059
R39994 vss.n1694 vss.n1652 0.271059
R39995 vss.n1803 vss.n1802 0.271059
R39996 vss.n1697 vss.n1696 0.271059
R39997 vss.n13235 vss.n793 0.271059
R39998 vss.n1566 vss.n1565 0.271059
R39999 vss.n13991 vss.n554 0.271059
R40000 vss.n13990 vss.n555 0.271059
R40001 vss.n13953 vss.n594 0.271059
R40002 vss.n14030 vss.n14029 0.271059
R40003 vss.n13289 vss.n706 0.271059
R40004 vss.n13290 vss.n705 0.271059
R40005 vss.n1982 vss.n1981 0.271059
R40006 vss.n13201 vss.n13200 0.271059
R40007 vss.n7497 vss.n7496 0.271059
R40008 vss.n8975 vss.n8974 0.271059
R40009 vss.n8477 vss.n8476 0.271059
R40010 vss.n8474 vss.n8473 0.271059
R40011 vss.n8863 vss.n8862 0.271059
R40012 vss.n7588 vss.n7587 0.271059
R40013 vss.n8856 vss.n8855 0.271059
R40014 vss.n8379 vss.n8378 0.271059
R40015 vss.n8376 vss.n8375 0.271059
R40016 vss.n8744 vss.n8743 0.271059
R40017 vss.n7731 vss.n7730 0.271059
R40018 vss.n8737 vss.n8736 0.271059
R40019 vss.n7906 vss.n7905 0.271059
R40020 vss.n8258 vss.n8257 0.271059
R40021 vss.n8253 vss.n8252 0.271059
R40022 vss.n7952 vss.n7951 0.271059
R40023 vss.n8246 vss.n8245 0.271059
R40024 vss.n7989 vss.n6004 0.271059
R40025 vss.n9641 vss.n9640 0.271059
R40026 vss.n9637 vss.n9636 0.271059
R40027 vss.n6052 vss.n6051 0.271059
R40028 vss.n6367 vss.n6366 0.271059
R40029 vss.n9253 vss.n9252 0.271059
R40030 vss.n9248 vss.n9247 0.271059
R40031 vss.n6903 vss.n6489 0.271059
R40032 vss.n7029 vss.n6986 0.271059
R40033 vss.n6981 vss.n6980 0.271059
R40034 vss.n7090 vss.n7089 0.271059
R40035 vss.n7085 vss.n7084 0.271059
R40036 vss.n6717 vss.n6716 0.271059
R40037 vss.n7220 vss.n7177 0.271059
R40038 vss.n7170 vss.n7169 0.271059
R40039 vss.n9540 vss.n6094 0.271059
R40040 vss.n9539 vss.n6095 0.271059
R40041 vss.n9502 vss.n6134 0.271059
R40042 vss.n9579 vss.n9578 0.271059
R40043 vss.n6546 vss.n6545 0.271059
R40044 vss.n9146 vss.n9145 0.271059
R40045 vss.n9192 vss.n9149 0.271059
R40046 vss.n9367 vss.n9366 0.271059
R40047 vss.n2924 vss.n2923 0.271059
R40048 vss.n9845 vss.n9844 0.271059
R40049 vss.n5330 vss.n5329 0.271059
R40050 vss.n5327 vss.n5326 0.271059
R40051 vss.n5322 vss.n5321 0.271059
R40052 vss.n4965 vss.n4964 0.271059
R40053 vss.n5315 vss.n5314 0.271059
R40054 vss.n5270 vss.n5269 0.271059
R40055 vss.n5268 vss.n5267 0.271059
R40056 vss.n5263 vss.n5262 0.271059
R40057 vss.n5167 vss.n5166 0.271059
R40058 vss.n5256 vss.n5255 0.271059
R40059 vss.n5211 vss.n5210 0.271059
R40060 vss.n5209 vss.n5208 0.271059
R40061 vss.n9793 vss.n9792 0.271059
R40062 vss.n3148 vss.n3147 0.271059
R40063 vss.n9786 vss.n9785 0.271059
R40064 vss.n9741 vss.n9740 0.271059
R40065 vss.n9739 vss.n9738 0.271059
R40066 vss.n9735 vss.n9734 0.271059
R40067 vss.n9991 vss.n9990 0.271059
R40068 vss.n3602 vss.n3601 0.271059
R40069 vss.n5740 vss.n5739 0.271059
R40070 vss.n5786 vss.n5743 0.271059
R40071 vss.n3424 vss.n3423 0.271059
R40072 vss.n5845 vss.n5844 0.271059
R40073 vss.n5840 vss.n5839 0.271059
R40074 vss.n3946 vss.n3543 0.271059
R40075 vss.n4119 vss.n4076 0.271059
R40076 vss.n4021 vss.n4020 0.271059
R40077 vss.n4070 vss.n4069 0.271059
R40078 vss.n4172 vss.n3802 0.271059
R40079 vss.n4173 vss.n3801 0.271059
R40080 vss.n4212 vss.n4211 0.271059
R40081 vss.n4288 vss.n4287 0.271059
R40082 vss.n4411 vss.n4368 0.271059
R40083 vss.n4611 vss.n4610 0.271059
R40084 vss.n4457 vss.n4412 0.271059
R40085 vss.n4503 vss.n4460 0.271059
R40086 vss.n5932 vss.n5931 0.271059
R40087 vss.n10013 vss.n10012 0.271059
R40088 vss.n10010 vss.n2557 0.271059
R40089 vss.n9729 vss.n9684 0.271059
R40090 vss.n9682 vss.n5936 0.271059
R40091 vss.n9631 vss.n9630 0.271059
R40092 vss.n9628 vss.n9585 0.271059
R40093 vss.n14090 vss.n14089 0.271059
R40094 vss.n12143 vss.n12142 0.271059
R40095 vss.n12140 vss.n12139 0.271059
R40096 vss.n12321 vss.n12320 0.271059
R40097 vss.n12366 vss.n12365 0.271059
R40098 vss.n12535 vss.n12534 0.271059
R40099 vss.n12539 vss.n12538 0.271059
R40100 vss.n12403 vss.n11736 0.271059
R40101 vss.n12451 vss.n12450 0.271059
R40102 vss.n10262 vss.n10261 0.271059
R40103 vss.n12902 vss.n12901 0.271059
R40104 vss.n12857 vss.n12856 0.271059
R40105 vss.n10302 vss.n10301 0.271059
R40106 vss.n12909 vss.n12908 0.271059
R40107 vss.n2442 vss.n2441 0.271059
R40108 vss.n12954 vss.n12953 0.271059
R40109 vss.n12952 vss.n10016 0.271059
R40110 vss.n12965 vss.n12964 0.271059
R40111 vss.n12958 vss.n12957 0.271059
R40112 vss.n2265 vss.n2264 0.271059
R40113 vss.n13019 vss.n13018 0.271059
R40114 vss.n12075 vss.n11890 0.271059
R40115 vss.n12074 vss.n11891 0.271059
R40116 vss.n11967 vss.n11925 0.271059
R40117 vss.n10503 vss.n10502 0.271059
R40118 vss.n12616 vss.n12615 0.271059
R40119 vss.n12611 vss.n12610 0.271059
R40120 vss.n10679 vss.n10590 0.271059
R40121 vss.n11593 vss.n11551 0.271059
R40122 vss.n10724 vss.n10723 0.271059
R40123 vss.n11545 vss.n11544 0.271059
R40124 vss.n11540 vss.n11539 0.271059
R40125 vss.n10974 vss.n10811 0.271059
R40126 vss.n10993 vss.n10992 0.271059
R40127 vss.n11038 vss.n11037 0.271059
R40128 vss.n11446 vss.n11404 0.271059
R40129 vss.n12740 vss.n10339 0.271059
R40130 vss.n12739 vss.n10340 0.271059
R40131 vss.n12696 vss.n10373 0.271059
R40132 vss.n11147 vss.n11146 0.271059
R40133 vss.n13148 vss.n2031 0.271059
R40134 vss.n14793 vss.n0 0.271059
R40135 vss.n13150 vss 0.194579
R40136 vss.n13154 vss 0.194579
R40137 vss.n13152 vss 0.194579
R40138 vss.n114 vss.n97 0.1305
R40139 vss.n14772 vss.n97 0.1305
R40140 vss.n111 vss.n98 0.1305
R40141 vss.n14772 vss.n98 0.1305
R40142 vss.n103 vss.n99 0.1305
R40143 vss.n14772 vss.n99 0.1305
R40144 vss.n14771 vss.n14770 0.1305
R40145 vss.n14772 vss.n14771 0.1305
R40146 vss.n109 vss.n37 0.1305
R40147 vss.n14782 vss.n37 0.1305
R40148 vss.n121 vss.n36 0.1305
R40149 vss.n14782 vss.n36 0.1305
R40150 vss.n14764 vss.n35 0.1305
R40151 vss.n14782 vss.n35 0.1305
R40152 vss.n104 vss.n34 0.1305
R40153 vss.n14782 vss.n34 0.1305
R40154 vss.n144 vss.n93 0.1305
R40155 vss.n14772 vss.n93 0.1305
R40156 vss.n141 vss.n94 0.1305
R40157 vss.n14772 vss.n94 0.1305
R40158 vss.n139 vss.n95 0.1305
R40159 vss.n14772 vss.n95 0.1305
R40160 vss.n137 vss.n96 0.1305
R40161 vss.n14772 vss.n96 0.1305
R40162 vss.n123 vss.n41 0.1305
R40163 vss.n14782 vss.n41 0.1305
R40164 vss.n151 vss.n40 0.1305
R40165 vss.n14782 vss.n40 0.1305
R40166 vss.n132 vss.n39 0.1305
R40167 vss.n14782 vss.n39 0.1305
R40168 vss.n134 vss.n38 0.1305
R40169 vss.n14782 vss.n38 0.1305
R40170 vss.n14632 vss.n89 0.1305
R40171 vss.n14772 vss.n89 0.1305
R40172 vss.n14629 vss.n90 0.1305
R40173 vss.n14772 vss.n90 0.1305
R40174 vss.n14627 vss.n91 0.1305
R40175 vss.n14772 vss.n91 0.1305
R40176 vss.n14625 vss.n92 0.1305
R40177 vss.n14772 vss.n92 0.1305
R40178 vss.n14611 vss.n45 0.1305
R40179 vss.n14782 vss.n45 0.1305
R40180 vss.n14639 vss.n44 0.1305
R40181 vss.n14782 vss.n44 0.1305
R40182 vss.n14620 vss.n43 0.1305
R40183 vss.n14782 vss.n43 0.1305
R40184 vss.n14622 vss.n42 0.1305
R40185 vss.n14782 vss.n42 0.1305
R40186 vss.n221 vss.n85 0.1305
R40187 vss.n14772 vss.n85 0.1305
R40188 vss.n218 vss.n86 0.1305
R40189 vss.n14772 vss.n86 0.1305
R40190 vss.n216 vss.n87 0.1305
R40191 vss.n14772 vss.n87 0.1305
R40192 vss.n214 vss.n88 0.1305
R40193 vss.n14772 vss.n88 0.1305
R40194 vss.n200 vss.n49 0.1305
R40195 vss.n14782 vss.n49 0.1305
R40196 vss.n228 vss.n48 0.1305
R40197 vss.n14782 vss.n48 0.1305
R40198 vss.n209 vss.n47 0.1305
R40199 vss.n14782 vss.n47 0.1305
R40200 vss.n211 vss.n46 0.1305
R40201 vss.n14782 vss.n46 0.1305
R40202 vss.n14437 vss.n81 0.1305
R40203 vss.n14772 vss.n81 0.1305
R40204 vss.n14434 vss.n82 0.1305
R40205 vss.n14772 vss.n82 0.1305
R40206 vss.n14432 vss.n83 0.1305
R40207 vss.n14772 vss.n83 0.1305
R40208 vss.n14430 vss.n84 0.1305
R40209 vss.n14772 vss.n84 0.1305
R40210 vss.n14416 vss.n53 0.1305
R40211 vss.n14782 vss.n53 0.1305
R40212 vss.n14444 vss.n52 0.1305
R40213 vss.n14782 vss.n52 0.1305
R40214 vss.n14425 vss.n51 0.1305
R40215 vss.n14782 vss.n51 0.1305
R40216 vss.n14427 vss.n50 0.1305
R40217 vss.n14782 vss.n50 0.1305
R40218 vss.n280 vss.n77 0.1305
R40219 vss.n14772 vss.n77 0.1305
R40220 vss.n277 vss.n78 0.1305
R40221 vss.n14772 vss.n78 0.1305
R40222 vss.n275 vss.n79 0.1305
R40223 vss.n14772 vss.n79 0.1305
R40224 vss.n273 vss.n80 0.1305
R40225 vss.n14772 vss.n80 0.1305
R40226 vss.n259 vss.n57 0.1305
R40227 vss.n14782 vss.n57 0.1305
R40228 vss.n287 vss.n56 0.1305
R40229 vss.n14782 vss.n56 0.1305
R40230 vss.n268 vss.n55 0.1305
R40231 vss.n14782 vss.n55 0.1305
R40232 vss.n270 vss.n54 0.1305
R40233 vss.n14782 vss.n54 0.1305
R40234 vss.n403 vss.n71 0.1305
R40235 vss.n14772 vss.n71 0.1305
R40236 vss.n400 vss.n72 0.1305
R40237 vss.n14772 vss.n72 0.1305
R40238 vss.n398 vss.n73 0.1305
R40239 vss.n14772 vss.n73 0.1305
R40240 vss.n396 vss.n74 0.1305
R40241 vss.n14772 vss.n74 0.1305
R40242 vss.n382 vss.n64 0.1305
R40243 vss.n14782 vss.n64 0.1305
R40244 vss.n410 vss.n63 0.1305
R40245 vss.n14782 vss.n63 0.1305
R40246 vss.n391 vss.n62 0.1305
R40247 vss.n14782 vss.n62 0.1305
R40248 vss.n393 vss.n61 0.1305
R40249 vss.n14782 vss.n61 0.1305
R40250 vss.n14781 vss.n66 0.1305
R40251 vss.n14782 vss.n14781 0.1305
R40252 vss.n14778 vss.n67 0.1305
R40253 vss.n14772 vss.n67 0.1305
R40254 vss.n14773 vss.n68 0.1305
R40255 vss.n14773 vss.n14772 0.1305
R40256 vss.n371 vss.n75 0.1305
R40257 vss.n14772 vss.n75 0.1305
R40258 vss.n373 vss.n76 0.1305
R40259 vss.n14772 vss.n76 0.1305
R40260 vss.n14782 vss.n60 0.1305
R40261 vss.n379 vss.n60 0.1305
R40262 vss.n14782 vss.n59 0.1305
R40263 vss.n377 vss.n59 0.1305
R40264 vss.n14782 vss.n58 0.1305
R40265 vss.n375 vss.n58 0.1305
R40266 vss.n9298 vss.n9294 0.1305
R40267 vss.n9294 vss.n6220 0.1305
R40268 vss.n9289 vss.n6215 0.1305
R40269 vss.n9289 vss.n6220 0.1305
R40270 vss.n9304 vss.n6214 0.1305
R40271 vss.n9304 vss.n6220 0.1305
R40272 vss.n9314 vss.n9306 0.1305
R40273 vss.n9306 vss.n6220 0.1305
R40274 vss.n9307 vss.n9303 0.1305
R40275 vss.n9303 vss.n6219 0.1305
R40276 vss.n9310 vss.n9309 0.1305
R40277 vss.n9309 vss.n6219 0.1305
R40278 vss.n9292 vss.n9291 0.1305
R40279 vss.n9291 vss.n6219 0.1305
R40280 vss.n9296 vss.n9295 0.1305
R40281 vss.n9295 vss.n6219 0.1305
R40282 vss.n9261 vss.n9260 0.1305
R40283 vss.n9260 vss.n6220 0.1305
R40284 vss.n9279 vss.n9278 0.1305
R40285 vss.n9279 vss.n6220 0.1305
R40286 vss.n9282 vss.n9281 0.1305
R40287 vss.n9281 vss.n6220 0.1305
R40288 vss.n9284 vss.n6321 0.1305
R40289 vss.n6321 vss.n6220 0.1305
R40290 vss.n6322 vss.n6320 0.1305
R40291 vss.n6320 vss.n6219 0.1305
R40292 vss.n9269 vss.n9268 0.1305
R40293 vss.n9269 vss.n6219 0.1305
R40294 vss.n9271 vss.n9262 0.1305
R40295 vss.n9271 vss.n6219 0.1305
R40296 vss.n9274 vss.n9273 0.1305
R40297 vss.n9273 vss.n6219 0.1305
R40298 vss.n6390 vss.n6389 0.1305
R40299 vss.n6389 vss.n6220 0.1305
R40300 vss.n6387 vss.n6370 0.1305
R40301 vss.n6387 vss.n6220 0.1305
R40302 vss.n6385 vss.n6369 0.1305
R40303 vss.n6385 vss.n6220 0.1305
R40304 vss.n6383 vss.n6382 0.1305
R40305 vss.n6383 vss.n6220 0.1305
R40306 vss.n6378 vss.n6377 0.1305
R40307 vss.n6377 vss.n6219 0.1305
R40308 vss.n6398 vss.n6397 0.1305
R40309 vss.n6397 vss.n6219 0.1305
R40310 vss.n6395 vss.n6371 0.1305
R40311 vss.n6395 vss.n6219 0.1305
R40312 vss.n6393 vss.n6392 0.1305
R40313 vss.n6393 vss.n6219 0.1305
R40314 vss.n6926 vss.n6925 0.1305
R40315 vss.n6925 vss.n6220 0.1305
R40316 vss.n6923 vss.n6906 0.1305
R40317 vss.n6923 vss.n6220 0.1305
R40318 vss.n6921 vss.n6905 0.1305
R40319 vss.n6921 vss.n6220 0.1305
R40320 vss.n6919 vss.n6918 0.1305
R40321 vss.n6919 vss.n6220 0.1305
R40322 vss.n6914 vss.n6913 0.1305
R40323 vss.n6913 vss.n6219 0.1305
R40324 vss.n6934 vss.n6933 0.1305
R40325 vss.n6933 vss.n6219 0.1305
R40326 vss.n6931 vss.n6907 0.1305
R40327 vss.n6931 vss.n6219 0.1305
R40328 vss.n6929 vss.n6928 0.1305
R40329 vss.n6929 vss.n6219 0.1305
R40330 vss.n6617 vss.n6616 0.1305
R40331 vss.n6616 vss.n6220 0.1305
R40332 vss.n6614 vss.n6597 0.1305
R40333 vss.n6614 vss.n6220 0.1305
R40334 vss.n6612 vss.n6596 0.1305
R40335 vss.n6612 vss.n6220 0.1305
R40336 vss.n6610 vss.n6609 0.1305
R40337 vss.n6610 vss.n6220 0.1305
R40338 vss.n6605 vss.n6604 0.1305
R40339 vss.n6604 vss.n6219 0.1305
R40340 vss.n6625 vss.n6624 0.1305
R40341 vss.n6624 vss.n6219 0.1305
R40342 vss.n6622 vss.n6598 0.1305
R40343 vss.n6622 vss.n6219 0.1305
R40344 vss.n6620 vss.n6619 0.1305
R40345 vss.n6620 vss.n6219 0.1305
R40346 vss.n7115 vss.n7114 0.1305
R40347 vss.n7114 vss.n6220 0.1305
R40348 vss.n7112 vss.n7095 0.1305
R40349 vss.n7112 vss.n6220 0.1305
R40350 vss.n7110 vss.n7094 0.1305
R40351 vss.n7110 vss.n6220 0.1305
R40352 vss.n7108 vss.n7107 0.1305
R40353 vss.n7108 vss.n6220 0.1305
R40354 vss.n7103 vss.n7102 0.1305
R40355 vss.n7102 vss.n6219 0.1305
R40356 vss.n7123 vss.n7122 0.1305
R40357 vss.n7122 vss.n6219 0.1305
R40358 vss.n7120 vss.n7096 0.1305
R40359 vss.n7120 vss.n6219 0.1305
R40360 vss.n7118 vss.n7117 0.1305
R40361 vss.n7118 vss.n6219 0.1305
R40362 vss.n6270 vss.n6269 0.1305
R40363 vss.n6269 vss.n6220 0.1305
R40364 vss.n6288 vss.n6287 0.1305
R40365 vss.n6288 vss.n6220 0.1305
R40366 vss.n6291 vss.n6290 0.1305
R40367 vss.n6290 vss.n6220 0.1305
R40368 vss.n6293 vss.n6263 0.1305
R40369 vss.n6263 vss.n6220 0.1305
R40370 vss.n6264 vss.n6262 0.1305
R40371 vss.n6262 vss.n6219 0.1305
R40372 vss.n6278 vss.n6277 0.1305
R40373 vss.n6278 vss.n6219 0.1305
R40374 vss.n6280 vss.n6271 0.1305
R40375 vss.n6280 vss.n6219 0.1305
R40376 vss.n6283 vss.n6282 0.1305
R40377 vss.n6282 vss.n6219 0.1305
R40378 vss.n6232 vss.n6231 0.1305
R40379 vss.n6231 vss.n6220 0.1305
R40380 vss.n6250 vss.n6249 0.1305
R40381 vss.n6250 vss.n6220 0.1305
R40382 vss.n6253 vss.n6252 0.1305
R40383 vss.n6252 vss.n6220 0.1305
R40384 vss.n6255 vss.n6226 0.1305
R40385 vss.n6226 vss.n6220 0.1305
R40386 vss.n6227 vss.n6225 0.1305
R40387 vss.n6225 vss.n6219 0.1305
R40388 vss.n6240 vss.n6239 0.1305
R40389 vss.n6240 vss.n6219 0.1305
R40390 vss.n6242 vss.n6233 0.1305
R40391 vss.n6242 vss.n6219 0.1305
R40392 vss.n6245 vss.n6244 0.1305
R40393 vss.n6244 vss.n6219 0.1305
R40394 vss.n3253 vss.n3252 0.1305
R40395 vss.n3252 vss.n2793 0.1305
R40396 vss.n3250 vss.n3249 0.1305
R40397 vss.n3250 vss.n2793 0.1305
R40398 vss.n3247 vss.n3246 0.1305
R40399 vss.n3246 vss.n2793 0.1305
R40400 vss.n3244 vss.n3243 0.1305
R40401 vss.n3244 vss.n2793 0.1305
R40402 vss.n3256 vss.n3255 0.1305
R40403 vss.n3256 vss.n2783 0.1305
R40404 vss.n3259 vss.n3258 0.1305
R40405 vss.n3258 vss.n2783 0.1305
R40406 vss.n3238 vss.n3237 0.1305
R40407 vss.n3238 vss.n2783 0.1305
R40408 vss.n3241 vss.n3240 0.1305
R40409 vss.n3240 vss.n2783 0.1305
R40410 vss.n3176 vss.n3175 0.1305
R40411 vss.n3175 vss.n2793 0.1305
R40412 vss.n3173 vss.n3172 0.1305
R40413 vss.n3173 vss.n2793 0.1305
R40414 vss.n3170 vss.n3169 0.1305
R40415 vss.n3169 vss.n2793 0.1305
R40416 vss.n3167 vss.n3166 0.1305
R40417 vss.n3167 vss.n2793 0.1305
R40418 vss.n3179 vss.n3178 0.1305
R40419 vss.n3179 vss.n2783 0.1305
R40420 vss.n3182 vss.n3181 0.1305
R40421 vss.n3181 vss.n2783 0.1305
R40422 vss.n3161 vss.n3160 0.1305
R40423 vss.n3161 vss.n2783 0.1305
R40424 vss.n3164 vss.n3163 0.1305
R40425 vss.n3163 vss.n2783 0.1305
R40426 vss.n3096 vss.n3095 0.1305
R40427 vss.n3095 vss.n2793 0.1305
R40428 vss.n3093 vss.n3092 0.1305
R40429 vss.n3093 vss.n2793 0.1305
R40430 vss.n3090 vss.n3089 0.1305
R40431 vss.n3089 vss.n2793 0.1305
R40432 vss.n3087 vss.n3086 0.1305
R40433 vss.n3087 vss.n2793 0.1305
R40434 vss.n3099 vss.n3098 0.1305
R40435 vss.n3099 vss.n2783 0.1305
R40436 vss.n3102 vss.n3101 0.1305
R40437 vss.n3101 vss.n2783 0.1305
R40438 vss.n3081 vss.n3080 0.1305
R40439 vss.n3081 vss.n2783 0.1305
R40440 vss.n3084 vss.n3083 0.1305
R40441 vss.n3083 vss.n2783 0.1305
R40442 vss.n5195 vss.n5194 0.1305
R40443 vss.n5194 vss.n2793 0.1305
R40444 vss.n5192 vss.n5191 0.1305
R40445 vss.n5192 vss.n2793 0.1305
R40446 vss.n5189 vss.n5188 0.1305
R40447 vss.n5188 vss.n2793 0.1305
R40448 vss.n5186 vss.n5185 0.1305
R40449 vss.n5186 vss.n2793 0.1305
R40450 vss.n5198 vss.n5197 0.1305
R40451 vss.n5198 vss.n2783 0.1305
R40452 vss.n5201 vss.n5200 0.1305
R40453 vss.n5200 vss.n2783 0.1305
R40454 vss.n5180 vss.n5179 0.1305
R40455 vss.n5180 vss.n2783 0.1305
R40456 vss.n5183 vss.n5182 0.1305
R40457 vss.n5182 vss.n2783 0.1305
R40458 vss.n5070 vss.n5069 0.1305
R40459 vss.n5069 vss.n2793 0.1305
R40460 vss.n5067 vss.n5066 0.1305
R40461 vss.n5067 vss.n2793 0.1305
R40462 vss.n5064 vss.n5063 0.1305
R40463 vss.n5063 vss.n2793 0.1305
R40464 vss.n5061 vss.n5060 0.1305
R40465 vss.n5061 vss.n2793 0.1305
R40466 vss.n5073 vss.n5072 0.1305
R40467 vss.n5073 vss.n2783 0.1305
R40468 vss.n5076 vss.n5075 0.1305
R40469 vss.n5075 vss.n2783 0.1305
R40470 vss.n5055 vss.n5054 0.1305
R40471 vss.n5055 vss.n2783 0.1305
R40472 vss.n5058 vss.n5057 0.1305
R40473 vss.n5057 vss.n2783 0.1305
R40474 vss.n4993 vss.n4992 0.1305
R40475 vss.n4992 vss.n2793 0.1305
R40476 vss.n4990 vss.n4989 0.1305
R40477 vss.n4990 vss.n2793 0.1305
R40478 vss.n4987 vss.n4986 0.1305
R40479 vss.n4986 vss.n2793 0.1305
R40480 vss.n4984 vss.n4983 0.1305
R40481 vss.n4984 vss.n2793 0.1305
R40482 vss.n4996 vss.n4995 0.1305
R40483 vss.n4996 vss.n2783 0.1305
R40484 vss.n4999 vss.n4998 0.1305
R40485 vss.n4998 vss.n2783 0.1305
R40486 vss.n4978 vss.n4977 0.1305
R40487 vss.n4978 vss.n2783 0.1305
R40488 vss.n4981 vss.n4980 0.1305
R40489 vss.n4980 vss.n2783 0.1305
R40490 vss.n2862 vss.n2861 0.1305
R40491 vss.n2861 vss.n2793 0.1305
R40492 vss.n2859 vss.n2858 0.1305
R40493 vss.n2859 vss.n2793 0.1305
R40494 vss.n2856 vss.n2855 0.1305
R40495 vss.n2855 vss.n2793 0.1305
R40496 vss.n2853 vss.n2852 0.1305
R40497 vss.n2853 vss.n2793 0.1305
R40498 vss.n2865 vss.n2864 0.1305
R40499 vss.n2865 vss.n2783 0.1305
R40500 vss.n2868 vss.n2867 0.1305
R40501 vss.n2867 vss.n2783 0.1305
R40502 vss.n2847 vss.n2846 0.1305
R40503 vss.n2847 vss.n2783 0.1305
R40504 vss.n2850 vss.n2849 0.1305
R40505 vss.n2849 vss.n2783 0.1305
R40506 vss.n2833 vss.n2832 0.1305
R40507 vss.n2832 vss.n2793 0.1305
R40508 vss.n9865 vss.n9864 0.1305
R40509 vss.n9865 vss.n2793 0.1305
R40510 vss.n9868 vss.n9867 0.1305
R40511 vss.n9867 vss.n2793 0.1305
R40512 vss.n9870 vss.n2826 0.1305
R40513 vss.n2826 vss.n2793 0.1305
R40514 vss.n9857 vss.n2835 0.1305
R40515 vss.n9857 vss.n2783 0.1305
R40516 vss.n9860 vss.n9859 0.1305
R40517 vss.n9859 vss.n2783 0.1305
R40518 vss.n9855 vss.n9854 0.1305
R40519 vss.n9855 vss.n2783 0.1305
R40520 vss.n2827 vss.n2825 0.1305
R40521 vss.n2825 vss.n2783 0.1305
R40522 vss.n1004 vss.n925 0.1305
R40523 vss.n13209 vss.n925 0.1305
R40524 vss.n990 vss.n984 0.1305
R40525 vss.n13209 vss.n984 0.1305
R40526 vss.n13205 vss.n985 0.1305
R40527 vss.n13209 vss.n985 0.1305
R40528 vss.n13208 vss.n13207 0.1305
R40529 vss.n13209 vss.n13208 0.1305
R40530 vss.n995 vss.n994 0.1305
R40531 vss.n994 vss.n497 0.1305
R40532 vss.n998 vss.n997 0.1305
R40533 vss.n998 vss.n497 0.1305
R40534 vss.n1011 vss.n1010 0.1305
R40535 vss.n1011 vss.n497 0.1305
R40536 vss.n1001 vss.n1000 0.1305
R40537 vss.n1001 vss.n497 0.1305
R40538 vss.n1037 vss.n926 0.1305
R40539 vss.n13209 vss.n926 0.1305
R40540 vss.n1017 vss.n981 0.1305
R40541 vss.n13209 vss.n981 0.1305
R40542 vss.n1016 vss.n982 0.1305
R40543 vss.n13209 vss.n982 0.1305
R40544 vss.n1024 vss.n983 0.1305
R40545 vss.n13209 vss.n983 0.1305
R40546 vss.n1021 vss.n1020 0.1305
R40547 vss.n1021 vss.n497 0.1305
R40548 vss.n1031 vss.n1030 0.1305
R40549 vss.n1031 vss.n497 0.1305
R40550 vss.n1044 vss.n1043 0.1305
R40551 vss.n1044 vss.n497 0.1305
R40552 vss.n1034 vss.n1033 0.1305
R40553 vss.n1034 vss.n497 0.1305
R40554 vss.n1298 vss.n927 0.1305
R40555 vss.n13209 vss.n927 0.1305
R40556 vss.n1278 vss.n978 0.1305
R40557 vss.n13209 vss.n978 0.1305
R40558 vss.n1277 vss.n979 0.1305
R40559 vss.n13209 vss.n979 0.1305
R40560 vss.n1285 vss.n980 0.1305
R40561 vss.n13209 vss.n980 0.1305
R40562 vss.n1282 vss.n1281 0.1305
R40563 vss.n1282 vss.n497 0.1305
R40564 vss.n1292 vss.n1291 0.1305
R40565 vss.n1292 vss.n497 0.1305
R40566 vss.n1305 vss.n1304 0.1305
R40567 vss.n1305 vss.n497 0.1305
R40568 vss.n1295 vss.n1294 0.1305
R40569 vss.n1295 vss.n497 0.1305
R40570 vss.n1430 vss.n928 0.1305
R40571 vss.n13209 vss.n928 0.1305
R40572 vss.n1410 vss.n975 0.1305
R40573 vss.n13209 vss.n975 0.1305
R40574 vss.n1409 vss.n976 0.1305
R40575 vss.n13209 vss.n976 0.1305
R40576 vss.n1417 vss.n977 0.1305
R40577 vss.n13209 vss.n977 0.1305
R40578 vss.n1414 vss.n1413 0.1305
R40579 vss.n1414 vss.n497 0.1305
R40580 vss.n1424 vss.n1423 0.1305
R40581 vss.n1424 vss.n497 0.1305
R40582 vss.n1437 vss.n1436 0.1305
R40583 vss.n1437 vss.n497 0.1305
R40584 vss.n1427 vss.n1426 0.1305
R40585 vss.n1427 vss.n497 0.1305
R40586 vss.n1593 vss.n929 0.1305
R40587 vss.n13209 vss.n929 0.1305
R40588 vss.n1573 vss.n972 0.1305
R40589 vss.n13209 vss.n972 0.1305
R40590 vss.n1572 vss.n973 0.1305
R40591 vss.n13209 vss.n973 0.1305
R40592 vss.n1580 vss.n974 0.1305
R40593 vss.n13209 vss.n974 0.1305
R40594 vss.n1577 vss.n1576 0.1305
R40595 vss.n1577 vss.n497 0.1305
R40596 vss.n1587 vss.n1586 0.1305
R40597 vss.n1587 vss.n497 0.1305
R40598 vss.n1600 vss.n1599 0.1305
R40599 vss.n1600 vss.n497 0.1305
R40600 vss.n1590 vss.n1589 0.1305
R40601 vss.n1590 vss.n497 0.1305
R40602 vss.n1510 vss.n930 0.1305
R40603 vss.n13209 vss.n930 0.1305
R40604 vss.n1490 vss.n969 0.1305
R40605 vss.n13209 vss.n969 0.1305
R40606 vss.n1489 vss.n970 0.1305
R40607 vss.n13209 vss.n970 0.1305
R40608 vss.n1497 vss.n971 0.1305
R40609 vss.n13209 vss.n971 0.1305
R40610 vss.n1494 vss.n1493 0.1305
R40611 vss.n1494 vss.n497 0.1305
R40612 vss.n1504 vss.n1503 0.1305
R40613 vss.n1504 vss.n497 0.1305
R40614 vss.n1517 vss.n1516 0.1305
R40615 vss.n1517 vss.n497 0.1305
R40616 vss.n1507 vss.n1506 0.1305
R40617 vss.n1507 vss.n497 0.1305
R40618 vss.n952 vss.n931 0.1305
R40619 vss.n13209 vss.n931 0.1305
R40620 vss.n938 vss.n932 0.1305
R40621 vss.n13209 vss.n932 0.1305
R40622 vss.n965 vss.n933 0.1305
R40623 vss.n13209 vss.n933 0.1305
R40624 vss.n968 vss.n967 0.1305
R40625 vss.n13209 vss.n968 0.1305
R40626 vss.n943 vss.n942 0.1305
R40627 vss.n942 vss.n497 0.1305
R40628 vss.n946 vss.n945 0.1305
R40629 vss.n946 vss.n497 0.1305
R40630 vss.n959 vss.n958 0.1305
R40631 vss.n959 vss.n497 0.1305
R40632 vss.n949 vss.n948 0.1305
R40633 vss.n949 vss.n497 0.1305
R40634 vss.n7358 vss.n7357 0.1305
R40635 vss.n7358 vss.n496 0.1305
R40636 vss.n7355 vss.n7354 0.1305
R40637 vss.n7354 vss.n496 0.1305
R40638 vss.n7375 vss.n7340 0.1305
R40639 vss.n8985 vss.n7340 0.1305
R40640 vss.n7378 vss.n7377 0.1305
R40641 vss.n8985 vss.n7378 0.1305
R40642 vss.n7982 vss.n7981 0.1305
R40643 vss.n7982 vss.n496 0.1305
R40644 vss.n7978 vss.n7977 0.1305
R40645 vss.n7978 vss.n496 0.1305
R40646 vss.n7975 vss.n7974 0.1305
R40647 vss.n7974 vss.n496 0.1305
R40648 vss.n7965 vss.n7963 0.1305
R40649 vss.n7963 vss.n496 0.1305
R40650 vss.n7955 vss.n7379 0.1305
R40651 vss.n8985 vss.n7379 0.1305
R40652 vss.n7987 vss.n7380 0.1305
R40653 vss.n8985 vss.n7380 0.1305
R40654 vss.n7969 vss.n7381 0.1305
R40655 vss.n8985 vss.n7381 0.1305
R40656 vss.n7968 vss.n7382 0.1305
R40657 vss.n8985 vss.n7382 0.1305
R40658 vss.n7840 vss.n7839 0.1305
R40659 vss.n7840 vss.n496 0.1305
R40660 vss.n7836 vss.n7835 0.1305
R40661 vss.n7836 vss.n496 0.1305
R40662 vss.n7833 vss.n7832 0.1305
R40663 vss.n7832 vss.n496 0.1305
R40664 vss.n7823 vss.n7821 0.1305
R40665 vss.n7821 vss.n496 0.1305
R40666 vss.n7813 vss.n7383 0.1305
R40667 vss.n8985 vss.n7383 0.1305
R40668 vss.n7845 vss.n7384 0.1305
R40669 vss.n8985 vss.n7384 0.1305
R40670 vss.n7827 vss.n7385 0.1305
R40671 vss.n8985 vss.n7385 0.1305
R40672 vss.n7826 vss.n7386 0.1305
R40673 vss.n8985 vss.n7386 0.1305
R40674 vss.n7761 vss.n7760 0.1305
R40675 vss.n7761 vss.n496 0.1305
R40676 vss.n7757 vss.n7756 0.1305
R40677 vss.n7757 vss.n496 0.1305
R40678 vss.n7754 vss.n7753 0.1305
R40679 vss.n7753 vss.n496 0.1305
R40680 vss.n7744 vss.n7742 0.1305
R40681 vss.n7742 vss.n496 0.1305
R40682 vss.n7734 vss.n7387 0.1305
R40683 vss.n8985 vss.n7387 0.1305
R40684 vss.n7766 vss.n7388 0.1305
R40685 vss.n8985 vss.n7388 0.1305
R40686 vss.n7748 vss.n7389 0.1305
R40687 vss.n8985 vss.n7389 0.1305
R40688 vss.n7747 vss.n7390 0.1305
R40689 vss.n8985 vss.n7390 0.1305
R40690 vss.n7653 vss.n7652 0.1305
R40691 vss.n7653 vss.n496 0.1305
R40692 vss.n7649 vss.n7648 0.1305
R40693 vss.n7649 vss.n496 0.1305
R40694 vss.n7646 vss.n7645 0.1305
R40695 vss.n7645 vss.n496 0.1305
R40696 vss.n7636 vss.n7634 0.1305
R40697 vss.n7634 vss.n496 0.1305
R40698 vss.n7626 vss.n7391 0.1305
R40699 vss.n8985 vss.n7391 0.1305
R40700 vss.n7658 vss.n7392 0.1305
R40701 vss.n8985 vss.n7392 0.1305
R40702 vss.n7640 vss.n7393 0.1305
R40703 vss.n8985 vss.n7393 0.1305
R40704 vss.n7639 vss.n7394 0.1305
R40705 vss.n8985 vss.n7394 0.1305
R40706 vss.n7618 vss.n7617 0.1305
R40707 vss.n7618 vss.n496 0.1305
R40708 vss.n7614 vss.n7613 0.1305
R40709 vss.n7614 vss.n496 0.1305
R40710 vss.n7611 vss.n7610 0.1305
R40711 vss.n7610 vss.n496 0.1305
R40712 vss.n7601 vss.n7599 0.1305
R40713 vss.n7599 vss.n496 0.1305
R40714 vss.n7591 vss.n7395 0.1305
R40715 vss.n8985 vss.n7395 0.1305
R40716 vss.n7623 vss.n7396 0.1305
R40717 vss.n8985 vss.n7396 0.1305
R40718 vss.n7605 vss.n7397 0.1305
R40719 vss.n8985 vss.n7397 0.1305
R40720 vss.n7604 vss.n7398 0.1305
R40721 vss.n8985 vss.n7398 0.1305
R40722 vss.n7464 vss.n7463 0.1305
R40723 vss.n7464 vss.n496 0.1305
R40724 vss.n7460 vss.n7459 0.1305
R40725 vss.n7460 vss.n496 0.1305
R40726 vss.n7457 vss.n7456 0.1305
R40727 vss.n7456 vss.n496 0.1305
R40728 vss.n7447 vss.n7445 0.1305
R40729 vss.n7445 vss.n496 0.1305
R40730 vss.n7437 vss.n7399 0.1305
R40731 vss.n8985 vss.n7399 0.1305
R40732 vss.n7469 vss.n7400 0.1305
R40733 vss.n8985 vss.n7400 0.1305
R40734 vss.n7451 vss.n7401 0.1305
R40735 vss.n8985 vss.n7401 0.1305
R40736 vss.n7450 vss.n7402 0.1305
R40737 vss.n8985 vss.n7402 0.1305
R40738 vss.n7430 vss.n7429 0.1305
R40739 vss.n7430 vss.n496 0.1305
R40740 vss.n7426 vss.n7425 0.1305
R40741 vss.n7426 vss.n496 0.1305
R40742 vss.n7423 vss.n7422 0.1305
R40743 vss.n7422 vss.n496 0.1305
R40744 vss.n7419 vss.n7418 0.1305
R40745 vss.n7419 vss.n496 0.1305
R40746 vss.n7411 vss.n7403 0.1305
R40747 vss.n8985 vss.n7403 0.1305
R40748 vss.n7435 vss.n7404 0.1305
R40749 vss.n8985 vss.n7404 0.1305
R40750 vss.n8981 vss.n7405 0.1305
R40751 vss.n8985 vss.n7405 0.1305
R40752 vss.n8984 vss.n8983 0.1305
R40753 vss.n8985 vss.n8984 0.1305
R40754 vss.n14035 vss.n513 0.1305
R40755 vss.n14051 vss.n513 0.1305
R40756 vss.n14050 vss.n14049 0.1305
R40757 vss.n14051 vss.n14050 0.1305
R40758 vss.n14052 vss.n511 0.1305
R40759 vss.n14052 vss.n14051 0.1305
R40760 vss.n509 vss.n508 0.1305
R40761 vss.n14051 vss.n509 0.1305
R40762 vss.n14058 vss.n14057 0.1305
R40763 vss.n14059 vss.n14058 0.1305
R40764 vss.n506 vss.n502 0.1305
R40765 vss.n14059 vss.n502 0.1305
R40766 vss.n14040 vss.n501 0.1305
R40767 vss.n14059 vss.n501 0.1305
R40768 vss.n14043 vss.n500 0.1305
R40769 vss.n14059 vss.n500 0.1305
R40770 vss.n7366 vss.n7365 0.1305
R40771 vss.n7365 vss.n499 0.1305
R40772 vss.n7361 vss.n7360 0.1305
R40773 vss.n7360 vss.n499 0.1305
R40774 vss.n7362 vss.n7348 0.1305
R40775 vss.n7348 vss.n7332 0.1305
R40776 vss.n7372 vss.n7371 0.1305
R40777 vss.n7371 vss.n7332 0.1305
R40778 vss.n2549 vss.n2548 0.1305
R40779 vss.n2548 vss.n2171 0.1305
R40780 vss.n2546 vss.n2545 0.1305
R40781 vss.n2546 vss.n2171 0.1305
R40782 vss.n2543 vss.n2542 0.1305
R40783 vss.n2542 vss.n2171 0.1305
R40784 vss.n2540 vss.n2539 0.1305
R40785 vss.n2540 vss.n2171 0.1305
R40786 vss.n2552 vss.n2551 0.1305
R40787 vss.n2552 vss.n2159 0.1305
R40788 vss.n2555 vss.n2554 0.1305
R40789 vss.n2554 vss.n2159 0.1305
R40790 vss.n2534 vss.n2533 0.1305
R40791 vss.n2534 vss.n2159 0.1305
R40792 vss.n2537 vss.n2536 0.1305
R40793 vss.n2536 vss.n2159 0.1305
R40794 vss.n2470 vss.n2469 0.1305
R40795 vss.n2469 vss.n2171 0.1305
R40796 vss.n2467 vss.n2466 0.1305
R40797 vss.n2467 vss.n2171 0.1305
R40798 vss.n2464 vss.n2463 0.1305
R40799 vss.n2463 vss.n2171 0.1305
R40800 vss.n2461 vss.n2460 0.1305
R40801 vss.n2461 vss.n2171 0.1305
R40802 vss.n2473 vss.n2472 0.1305
R40803 vss.n2473 vss.n2159 0.1305
R40804 vss.n2476 vss.n2475 0.1305
R40805 vss.n2475 vss.n2159 0.1305
R40806 vss.n2455 vss.n2454 0.1305
R40807 vss.n2455 vss.n2159 0.1305
R40808 vss.n2458 vss.n2457 0.1305
R40809 vss.n2457 vss.n2159 0.1305
R40810 vss.n10212 vss.n10211 0.1305
R40811 vss.n10211 vss.n2171 0.1305
R40812 vss.n10209 vss.n10208 0.1305
R40813 vss.n10209 vss.n2171 0.1305
R40814 vss.n10206 vss.n10205 0.1305
R40815 vss.n10205 vss.n2171 0.1305
R40816 vss.n10203 vss.n10202 0.1305
R40817 vss.n10203 vss.n2171 0.1305
R40818 vss.n10215 vss.n10214 0.1305
R40819 vss.n10215 vss.n2159 0.1305
R40820 vss.n10218 vss.n10217 0.1305
R40821 vss.n10217 vss.n2159 0.1305
R40822 vss.n10197 vss.n10196 0.1305
R40823 vss.n10197 vss.n2159 0.1305
R40824 vss.n10200 vss.n10199 0.1305
R40825 vss.n10199 vss.n2159 0.1305
R40826 vss.n10290 vss.n10289 0.1305
R40827 vss.n10289 vss.n2171 0.1305
R40828 vss.n10287 vss.n10286 0.1305
R40829 vss.n10287 vss.n2171 0.1305
R40830 vss.n10284 vss.n10283 0.1305
R40831 vss.n10283 vss.n2171 0.1305
R40832 vss.n10281 vss.n10280 0.1305
R40833 vss.n10281 vss.n2171 0.1305
R40834 vss.n10293 vss.n10292 0.1305
R40835 vss.n10293 vss.n2159 0.1305
R40836 vss.n10296 vss.n10295 0.1305
R40837 vss.n10295 vss.n2159 0.1305
R40838 vss.n10275 vss.n10274 0.1305
R40839 vss.n10275 vss.n2159 0.1305
R40840 vss.n10278 vss.n10277 0.1305
R40841 vss.n10277 vss.n2159 0.1305
R40842 vss.n12523 vss.n12522 0.1305
R40843 vss.n12522 vss.n2171 0.1305
R40844 vss.n12520 vss.n12519 0.1305
R40845 vss.n12520 vss.n2171 0.1305
R40846 vss.n12517 vss.n12516 0.1305
R40847 vss.n12516 vss.n2171 0.1305
R40848 vss.n12514 vss.n12513 0.1305
R40849 vss.n12514 vss.n2171 0.1305
R40850 vss.n12526 vss.n12525 0.1305
R40851 vss.n12526 vss.n2159 0.1305
R40852 vss.n12529 vss.n12528 0.1305
R40853 vss.n12528 vss.n2159 0.1305
R40854 vss.n12508 vss.n12507 0.1305
R40855 vss.n12508 vss.n2159 0.1305
R40856 vss.n12511 vss.n12510 0.1305
R40857 vss.n12510 vss.n2159 0.1305
R40858 vss.n12394 vss.n12393 0.1305
R40859 vss.n12393 vss.n2171 0.1305
R40860 vss.n12391 vss.n12390 0.1305
R40861 vss.n12391 vss.n2171 0.1305
R40862 vss.n12388 vss.n12387 0.1305
R40863 vss.n12387 vss.n2171 0.1305
R40864 vss.n12385 vss.n12384 0.1305
R40865 vss.n12385 vss.n2171 0.1305
R40866 vss.n12397 vss.n12396 0.1305
R40867 vss.n12397 vss.n2159 0.1305
R40868 vss.n12400 vss.n12399 0.1305
R40869 vss.n12399 vss.n2159 0.1305
R40870 vss.n12379 vss.n12378 0.1305
R40871 vss.n12379 vss.n2159 0.1305
R40872 vss.n12382 vss.n12381 0.1305
R40873 vss.n12381 vss.n2159 0.1305
R40874 vss.n2231 vss.n2230 0.1305
R40875 vss.n2230 vss.n2171 0.1305
R40876 vss.n2228 vss.n2227 0.1305
R40877 vss.n2228 vss.n2171 0.1305
R40878 vss.n2225 vss.n2224 0.1305
R40879 vss.n2224 vss.n2171 0.1305
R40880 vss.n2222 vss.n2221 0.1305
R40881 vss.n2222 vss.n2171 0.1305
R40882 vss.n2234 vss.n2233 0.1305
R40883 vss.n2234 vss.n2159 0.1305
R40884 vss.n2237 vss.n2236 0.1305
R40885 vss.n2236 vss.n2159 0.1305
R40886 vss.n2216 vss.n2215 0.1305
R40887 vss.n2216 vss.n2159 0.1305
R40888 vss.n2219 vss.n2218 0.1305
R40889 vss.n2218 vss.n2159 0.1305
R40890 vss.n5869 vss.n2592 0.1305
R40891 vss.n9999 vss.n2592 0.1305
R40892 vss.n2628 vss.n2622 0.1305
R40893 vss.n9999 vss.n2622 0.1305
R40894 vss.n9995 vss.n2623 0.1305
R40895 vss.n9999 vss.n2623 0.1305
R40896 vss.n9998 vss.n9997 0.1305
R40897 vss.n9999 vss.n9998 0.1305
R40898 vss.n5881 vss.n5880 0.1305
R40899 vss.n5882 vss.n5881 0.1305
R40900 vss.n5878 vss.n5863 0.1305
R40901 vss.n5882 vss.n5863 0.1305
R40902 vss.n5876 vss.n5859 0.1305
R40903 vss.n5882 vss.n5859 0.1305
R40904 vss.n5866 vss.n5858 0.1305
R40905 vss.n5882 vss.n5858 0.1305
R40906 vss.n3368 vss.n2593 0.1305
R40907 vss.n9999 vss.n2593 0.1305
R40908 vss.n3364 vss.n2619 0.1305
R40909 vss.n9999 vss.n2619 0.1305
R40910 vss.n5850 vss.n2620 0.1305
R40911 vss.n9999 vss.n2620 0.1305
R40912 vss.n3363 vss.n2621 0.1305
R40913 vss.n9999 vss.n2621 0.1305
R40914 vss.n5857 vss.n5856 0.1305
R40915 vss.n5882 vss.n5857 0.1305
R40916 vss.n3362 vss.n3358 0.1305
R40917 vss.n5882 vss.n3358 0.1305
R40918 vss.n3375 vss.n3357 0.1305
R40919 vss.n5882 vss.n3357 0.1305
R40920 vss.n3365 vss.n3356 0.1305
R40921 vss.n5882 vss.n3356 0.1305
R40922 vss.n3431 vss.n2594 0.1305
R40923 vss.n9999 vss.n2594 0.1305
R40924 vss.n3427 vss.n2616 0.1305
R40925 vss.n9999 vss.n2616 0.1305
R40926 vss.n3426 vss.n2617 0.1305
R40927 vss.n9999 vss.n2617 0.1305
R40928 vss.n3442 vss.n2618 0.1305
R40929 vss.n9999 vss.n2618 0.1305
R40930 vss.n3439 vss.n3355 0.1305
R40931 vss.n5882 vss.n3355 0.1305
R40932 vss.n3449 vss.n3354 0.1305
R40933 vss.n5882 vss.n3354 0.1305
R40934 vss.n3438 vss.n3353 0.1305
R40935 vss.n5882 vss.n3353 0.1305
R40936 vss.n3428 vss.n3352 0.1305
R40937 vss.n5882 vss.n3352 0.1305
R40938 vss.n3953 vss.n2595 0.1305
R40939 vss.n9999 vss.n2595 0.1305
R40940 vss.n3949 vss.n2613 0.1305
R40941 vss.n9999 vss.n2613 0.1305
R40942 vss.n3948 vss.n2614 0.1305
R40943 vss.n9999 vss.n2614 0.1305
R40944 vss.n3964 vss.n2615 0.1305
R40945 vss.n9999 vss.n2615 0.1305
R40946 vss.n3961 vss.n3351 0.1305
R40947 vss.n5882 vss.n3351 0.1305
R40948 vss.n3971 vss.n3350 0.1305
R40949 vss.n5882 vss.n3350 0.1305
R40950 vss.n3960 vss.n3349 0.1305
R40951 vss.n5882 vss.n3349 0.1305
R40952 vss.n3950 vss.n3348 0.1305
R40953 vss.n5882 vss.n3348 0.1305
R40954 vss.n3651 vss.n2596 0.1305
R40955 vss.n9999 vss.n2596 0.1305
R40956 vss.n3647 vss.n2610 0.1305
R40957 vss.n9999 vss.n2610 0.1305
R40958 vss.n3646 vss.n2611 0.1305
R40959 vss.n9999 vss.n2611 0.1305
R40960 vss.n3662 vss.n2612 0.1305
R40961 vss.n9999 vss.n2612 0.1305
R40962 vss.n3659 vss.n3347 0.1305
R40963 vss.n5882 vss.n3347 0.1305
R40964 vss.n3669 vss.n3346 0.1305
R40965 vss.n5882 vss.n3346 0.1305
R40966 vss.n3658 vss.n3345 0.1305
R40967 vss.n5882 vss.n3345 0.1305
R40968 vss.n3648 vss.n3344 0.1305
R40969 vss.n5882 vss.n3344 0.1305
R40970 vss.n4220 vss.n2597 0.1305
R40971 vss.n9999 vss.n2597 0.1305
R40972 vss.n4216 vss.n2607 0.1305
R40973 vss.n9999 vss.n2607 0.1305
R40974 vss.n4215 vss.n2608 0.1305
R40975 vss.n9999 vss.n2608 0.1305
R40976 vss.n4231 vss.n2609 0.1305
R40977 vss.n9999 vss.n2609 0.1305
R40978 vss.n4228 vss.n3343 0.1305
R40979 vss.n5882 vss.n3343 0.1305
R40980 vss.n4238 vss.n3342 0.1305
R40981 vss.n5882 vss.n3342 0.1305
R40982 vss.n4227 vss.n3341 0.1305
R40983 vss.n5882 vss.n3341 0.1305
R40984 vss.n4217 vss.n3340 0.1305
R40985 vss.n5882 vss.n3340 0.1305
R40986 vss.n4296 vss.n2598 0.1305
R40987 vss.n9999 vss.n2598 0.1305
R40988 vss.n4292 vss.n2604 0.1305
R40989 vss.n9999 vss.n2604 0.1305
R40990 vss.n4291 vss.n2605 0.1305
R40991 vss.n9999 vss.n2605 0.1305
R40992 vss.n4307 vss.n2606 0.1305
R40993 vss.n9999 vss.n2606 0.1305
R40994 vss.n4304 vss.n3339 0.1305
R40995 vss.n5882 vss.n3339 0.1305
R40996 vss.n4314 vss.n3338 0.1305
R40997 vss.n5882 vss.n3338 0.1305
R40998 vss.n4303 vss.n3337 0.1305
R40999 vss.n5882 vss.n3337 0.1305
R41000 vss.n4293 vss.n3336 0.1305
R41001 vss.n5882 vss.n3336 0.1305
R41002 vss.n3320 vss.n2599 0.1305
R41003 vss.n9999 vss.n2599 0.1305
R41004 vss.n3309 vss.n2601 0.1305
R41005 vss.n9999 vss.n2601 0.1305
R41006 vss.n3308 vss.n2602 0.1305
R41007 vss.n9999 vss.n2602 0.1305
R41008 vss.n3328 vss.n2603 0.1305
R41009 vss.n9999 vss.n2603 0.1305
R41010 vss.n3335 vss.n3334 0.1305
R41011 vss.n5882 vss.n3335 0.1305
R41012 vss.n3327 vss.n3311 0.1305
R41013 vss.n5882 vss.n3311 0.1305
R41014 vss.n5883 vss.n3313 0.1305
R41015 vss.n5883 vss.n5882 0.1305
R41016 vss.n3323 vss.n3322 0.1305
R41017 vss.n5882 vss.n3323 0.1305
R41018 vss.n13051 vss.n13050 0.1305
R41019 vss.n13051 vss.n2171 0.1305
R41020 vss.n13037 vss.n2203 0.1305
R41021 vss.n2203 vss.n2171 0.1305
R41022 vss.n13036 vss.n13035 0.1305
R41023 vss.n13035 vss.n2171 0.1305
R41024 vss.n13032 vss.n13031 0.1305
R41025 vss.n13032 vss.n2171 0.1305
R41026 vss.n13048 vss.n13047 0.1305
R41027 vss.n13047 vss.n2159 0.1305
R41028 vss.n13045 vss.n13044 0.1305
R41029 vss.n13044 vss.n2159 0.1305
R41030 vss.n13042 vss.n13041 0.1305
R41031 vss.n13042 vss.n2159 0.1305
R41032 vss.n13029 vss.n13028 0.1305
R41033 vss.n13028 vss.n2159 0.1305
R41034 vss.n11311 vss.n10424 0.1305
R41035 vss.n12671 vss.n10424 0.1305
R41036 vss.n11309 vss.n10449 0.1305
R41037 vss.n12671 vss.n10449 0.1305
R41038 vss.n11323 vss.n10450 0.1305
R41039 vss.n12671 vss.n10450 0.1305
R41040 vss.n11325 vss.n10451 0.1305
R41041 vss.n12671 vss.n10451 0.1305
R41042 vss.n11302 vss.n11301 0.1305
R41043 vss.n11301 vss.n11048 0.1305
R41044 vss.n11320 vss.n11319 0.1305
R41045 vss.n11319 vss.n11048 0.1305
R41046 vss.n11317 vss.n11316 0.1305
R41047 vss.n11317 vss.n11048 0.1305
R41048 vss.n11314 vss.n11313 0.1305
R41049 vss.n11313 vss.n11048 0.1305
R41050 vss.n11288 vss.n10425 0.1305
R41051 vss.n12671 vss.n10425 0.1305
R41052 vss.n11290 vss.n10446 0.1305
R41053 vss.n12671 vss.n10446 0.1305
R41054 vss.n11293 vss.n10447 0.1305
R41055 vss.n12671 vss.n10447 0.1305
R41056 vss.n11295 vss.n10448 0.1305
R41057 vss.n12671 vss.n10448 0.1305
R41058 vss.n11271 vss.n11270 0.1305
R41059 vss.n11270 vss.n11048 0.1305
R41060 vss.n11280 vss.n11279 0.1305
R41061 vss.n11279 vss.n11048 0.1305
R41062 vss.n11283 vss.n11282 0.1305
R41063 vss.n11283 vss.n11048 0.1305
R41064 vss.n11286 vss.n11285 0.1305
R41065 vss.n11285 vss.n11048 0.1305
R41066 vss.n11250 vss.n10426 0.1305
R41067 vss.n12671 vss.n10426 0.1305
R41068 vss.n11248 vss.n10443 0.1305
R41069 vss.n12671 vss.n10443 0.1305
R41070 vss.n11262 vss.n10444 0.1305
R41071 vss.n12671 vss.n10444 0.1305
R41072 vss.n11264 vss.n10445 0.1305
R41073 vss.n12671 vss.n10445 0.1305
R41074 vss.n11241 vss.n11240 0.1305
R41075 vss.n11240 vss.n11048 0.1305
R41076 vss.n11259 vss.n11258 0.1305
R41077 vss.n11258 vss.n11048 0.1305
R41078 vss.n11256 vss.n11255 0.1305
R41079 vss.n11256 vss.n11048 0.1305
R41080 vss.n11253 vss.n11252 0.1305
R41081 vss.n11252 vss.n11048 0.1305
R41082 vss.n11227 vss.n10427 0.1305
R41083 vss.n12671 vss.n10427 0.1305
R41084 vss.n11229 vss.n10440 0.1305
R41085 vss.n12671 vss.n10440 0.1305
R41086 vss.n11232 vss.n10441 0.1305
R41087 vss.n12671 vss.n10441 0.1305
R41088 vss.n11234 vss.n10442 0.1305
R41089 vss.n12671 vss.n10442 0.1305
R41090 vss.n11210 vss.n11209 0.1305
R41091 vss.n11209 vss.n11048 0.1305
R41092 vss.n11219 vss.n11218 0.1305
R41093 vss.n11218 vss.n11048 0.1305
R41094 vss.n11222 vss.n11221 0.1305
R41095 vss.n11222 vss.n11048 0.1305
R41096 vss.n11225 vss.n11224 0.1305
R41097 vss.n11224 vss.n11048 0.1305
R41098 vss.n11196 vss.n10428 0.1305
R41099 vss.n12671 vss.n10428 0.1305
R41100 vss.n11198 vss.n10437 0.1305
R41101 vss.n12671 vss.n10437 0.1305
R41102 vss.n11201 vss.n10438 0.1305
R41103 vss.n12671 vss.n10438 0.1305
R41104 vss.n11203 vss.n10439 0.1305
R41105 vss.n12671 vss.n10439 0.1305
R41106 vss.n11179 vss.n11178 0.1305
R41107 vss.n11178 vss.n11048 0.1305
R41108 vss.n11188 vss.n11187 0.1305
R41109 vss.n11187 vss.n11048 0.1305
R41110 vss.n11191 vss.n11190 0.1305
R41111 vss.n11191 vss.n11048 0.1305
R41112 vss.n11194 vss.n11193 0.1305
R41113 vss.n11193 vss.n11048 0.1305
R41114 vss.n11353 vss.n10429 0.1305
R41115 vss.n12671 vss.n10429 0.1305
R41116 vss.n11355 vss.n10434 0.1305
R41117 vss.n12671 vss.n10434 0.1305
R41118 vss.n11043 vss.n10435 0.1305
R41119 vss.n12671 vss.n10435 0.1305
R41120 vss.n11172 vss.n10436 0.1305
R41121 vss.n12671 vss.n10436 0.1305
R41122 vss.n11159 vss.n11158 0.1305
R41123 vss.n11158 vss.n11048 0.1305
R41124 vss.n11168 vss.n11167 0.1305
R41125 vss.n11167 vss.n11048 0.1305
R41126 vss.n11165 vss.n11164 0.1305
R41127 vss.n11165 vss.n11048 0.1305
R41128 vss.n11047 vss.n11046 0.1305
R41129 vss.n11048 vss.n11047 0.1305
R41130 vss.n11101 vss.n10430 0.1305
R41131 vss.n12671 vss.n10430 0.1305
R41132 vss.n11103 vss.n10431 0.1305
R41133 vss.n12671 vss.n10431 0.1305
R41134 vss.n11151 vss.n10432 0.1305
R41135 vss.n12671 vss.n10432 0.1305
R41136 vss.n11153 vss.n10433 0.1305
R41137 vss.n12671 vss.n10433 0.1305
R41138 vss.n11084 vss.n11083 0.1305
R41139 vss.n11083 vss.n11048 0.1305
R41140 vss.n11093 vss.n11092 0.1305
R41141 vss.n11092 vss.n11048 0.1305
R41142 vss.n11096 vss.n11095 0.1305
R41143 vss.n11096 vss.n11048 0.1305
R41144 vss.n11099 vss.n11098 0.1305
R41145 vss.n11098 vss.n11048 0.1305
R41146 vss.n11334 vss.n11333 0.1305
R41147 vss.n11333 vss.n11048 0.1305
R41148 vss.n11337 vss.n11336 0.1305
R41149 vss.n11337 vss.n11048 0.1305
R41150 vss.n11340 vss.n11339 0.1305
R41151 vss.n11339 vss.n11048 0.1305
R41152 vss.n11344 vss.n11343 0.1305
R41153 vss.n11343 vss.n11048 0.1305
R41154 vss.n11346 vss.n10452 0.1305
R41155 vss.n12671 vss.n10452 0.1305
R41156 vss.n11342 vss.n10453 0.1305
R41157 vss.n12671 vss.n10453 0.1305
R41158 vss.n12667 vss.n10454 0.1305
R41159 vss.n12671 vss.n10454 0.1305
R41160 vss.n12670 vss.n12669 0.1305
R41161 vss.n12671 vss.n12670 0.1305
R41162 vss.n13158 vss.n13155 0.1255
R41163 vss.n13153 vss.n2028 0.1255
R41164 vss.n13151 vss.n2029 0.1255
R41165 vss.n14181 vss 0.0745132
R41166 vss.n13369 vss 0.0745132
R41167 vss.n13449 vss 0.0745132
R41168 vss.n13529 vss 0.0745132
R41169 vss.n14300 vss 0.0745132
R41170 vss.n14253 vss 0.0745132
R41171 vss.n13647 vss 0.0745132
R41172 vss vss.n14368 0.0745132
R41173 vss vss.n14414 0.0745132
R41174 vss.n14495 vss 0.0745132
R41175 vss.n14448 vss 0.0745132
R41176 vss.n13752 vss 0.0745132
R41177 vss vss.n14563 0.0745132
R41178 vss vss.n14609 0.0745132
R41179 vss.n14690 vss 0.0745132
R41180 vss.n14643 vss 0.0745132
R41181 vss.n13857 vss 0.0745132
R41182 vss vss.n14758 0.0745132
R41183 vss vss.n361 0.0745132
R41184 vss vss.n14249 0.0745132
R41185 vss.n14143 vss 0.0745132
R41186 vss.n14094 vss 0.0745132
R41187 vss.n8179 vss 0.0745132
R41188 vss vss.n7811 0.0745132
R41189 vss.n8789 vss 0.0745132
R41190 vss vss.n7908 0.0745132
R41191 vss.n8328 vss 0.0745132
R41192 vss.n8426 vss 0.0745132
R41193 vss.n8908 vss 0.0745132
R41194 vss.n7495 vss 0.0745132
R41195 vss vss.n8976 0.0745132
R41196 vss.n8475 vss 0.0745132
R41197 vss.n8861 vss 0.0745132
R41198 vss vss.n7589 0.0745132
R41199 vss vss.n8857 0.0745132
R41200 vss.n8377 vss 0.0745132
R41201 vss.n8742 vss 0.0745132
R41202 vss vss.n7732 0.0745132
R41203 vss vss.n8738 0.0745132
R41204 vss.n7904 vss 0.0745132
R41205 vss.n8251 vss 0.0745132
R41206 vss vss.n7953 0.0745132
R41207 vss vss.n8247 0.0745132
R41208 vss vss.n7990 0.0745132
R41209 vss.n9635 vss 0.0745132
R41210 vss vss.n3226 0.0745132
R41211 vss vss.n3069 0.0745132
R41212 vss vss.n5043 0.0745132
R41213 vss.n4632 vss 0.0745132
R41214 vss vss.n5083 0.0745132
R41215 vss vss.n4881 0.0745132
R41216 vss.n2969 vss 0.0745132
R41217 vss.n2922 vss 0.0745132
R41218 vss vss.n9846 0.0745132
R41219 vss.n5328 vss 0.0745132
R41220 vss.n5320 vss 0.0745132
R41221 vss vss.n4966 0.0745132
R41222 vss vss.n5316 0.0745132
R41223 vss vss.n5271 0.0745132
R41224 vss.n5261 vss 0.0745132
R41225 vss vss.n5168 0.0745132
R41226 vss vss.n5257 0.0745132
R41227 vss vss.n5212 0.0745132
R41228 vss.n9791 vss 0.0745132
R41229 vss vss.n3149 0.0745132
R41230 vss vss.n9787 0.0745132
R41231 vss vss.n9742 0.0745132
R41232 vss.n9733 vss 0.0745132
R41233 vss.n10011 vss 0.0745132
R41234 vss vss.n5935 0.0745132
R41235 vss.n9683 vss 0.0745132
R41236 vss vss.n9583 0.0745132
R41237 vss.n9629 vss 0.0745132
R41238 vss.n9584 vss 0.0745132
R41239 vss.n14088 vss 0.0745132
R41240 vss.n12911 vss 0.0745132
R41241 vss vss.n10185 0.0745132
R41242 vss vss.n12407 0.0745132
R41243 vss vss.n12496 0.0745132
R41244 vss.n2339 vss 0.0745132
R41245 vss vss.n12277 0.0745132
R41246 vss.n12141 vss 0.0745132
R41247 vss vss.n12322 0.0745132
R41248 vss vss.n12367 0.0745132
R41249 vss.n12533 vss 0.0745132
R41250 vss.n12537 vss 0.0745132
R41251 vss vss.n12452 0.0745132
R41252 vss vss.n10263 0.0745132
R41253 vss vss.n12903 0.0745132
R41254 vss vss.n12858 0.0745132
R41255 vss.n12907 vss 0.0745132
R41256 vss vss.n2443 0.0745132
R41257 vss.n10015 vss 0.0745132
R41258 vss.n12963 vss 0.0745132
R41259 vss vss.n2522 0.0745132
R41260 vss vss.n12959 0.0745132
R41261 vss.n2263 vss 0.0745132
R41262 vss vss.n13020 0.0745132
R41263 vss vss.n14760 0.0745132
R41264 vss.n2047 vss.n2046 0.0702092
R41265 vss.n2047 vss.t1439 0.0702092
R41266 vss.n10394 vss.t1344 0.0702092
R41267 vss.n10403 vss.t1460 0.0702092
R41268 vss.t1462 vss.n13144 0.0702092
R41269 vss.n13140 vss.t1439 0.0702092
R41270 vss.n13146 vss.n13145 0.0702092
R41271 vss.n13145 vss.t1462 0.0702092
R41272 vss.n10402 vss.n2033 0.0702092
R41273 vss.t1460 vss.n10402 0.0702092
R41274 vss.n10395 vss.n10393 0.0702092
R41275 vss.n10393 vss.t1344 0.0702092
R41276 vss.n10406 vss.n10394 0.0702092
R41277 vss.n10404 vss.n10403 0.0702092
R41278 vss.n13144 vss.n13143 0.0702092
R41279 vss.n13141 vss.n13140 0.0702092
R41280 vss.n12652 vss.n12651 0.0702092
R41281 vss.n12652 vss.t971 0.0702092
R41282 vss.t1374 vss.n12641 0.0702092
R41283 vss.n12645 vss.t121 0.0702092
R41284 vss.t123 vss.n12658 0.0702092
R41285 vss.n12654 vss.t971 0.0702092
R41286 vss.n12660 vss.n12659 0.0702092
R41287 vss.n12659 vss.t123 0.0702092
R41288 vss.n12644 vss.n12622 0.0702092
R41289 vss.t121 vss.n12644 0.0702092
R41290 vss.n12642 vss.n12638 0.0702092
R41291 vss.n12642 vss.t1374 0.0702092
R41292 vss.n12641 vss.n12640 0.0702092
R41293 vss.n12646 vss.n12645 0.0702092
R41294 vss.n12658 vss.n12657 0.0702092
R41295 vss.n12655 vss.n12654 0.0702092
R41296 vss.n12676 vss.n12675 0.0702092
R41297 vss.t574 vss.n12676 0.0702092
R41298 vss.n12681 vss.n12680 0.0702092
R41299 vss.n12680 vss.t1095 0.0702092
R41300 vss.n12683 vss.n10380 0.0702092
R41301 vss.t1094 vss.n10380 0.0702092
R41302 vss.n12689 vss.n12688 0.0702092
R41303 vss.n12689 vss.t1063 0.0702092
R41304 vss.n12686 vss.n12685 0.0702092
R41305 vss.n12685 vss.t1063 0.0702092
R41306 vss.n12694 vss.n12693 0.0702092
R41307 vss.n12693 vss.t1094 0.0702092
R41308 vss.n12679 vss.n10375 0.0702092
R41309 vss.t1095 vss.n12679 0.0702092
R41310 vss.n12677 vss.n10392 0.0702092
R41311 vss.n12677 vss.t574 0.0702092
R41312 vss.n11426 vss.n11425 0.0702092
R41313 vss.t207 vss.n11426 0.0702092
R41314 vss.n11431 vss.n11430 0.0702092
R41315 vss.n11430 vss.t102 0.0702092
R41316 vss.n11433 vss.n11411 0.0702092
R41317 vss.t101 vss.n11411 0.0702092
R41318 vss.n11439 vss.n11438 0.0702092
R41319 vss.n11439 vss.t1048 0.0702092
R41320 vss.n11436 vss.n11435 0.0702092
R41321 vss.n11435 vss.t1048 0.0702092
R41322 vss.n11444 vss.n11443 0.0702092
R41323 vss.n11443 vss.t101 0.0702092
R41324 vss.n11429 vss.n11406 0.0702092
R41325 vss.t102 vss.n11429 0.0702092
R41326 vss.n11427 vss.n11423 0.0702092
R41327 vss.n11427 vss.t207 0.0702092
R41328 vss.n11379 vss.n11378 0.0702092
R41329 vss.t19 vss.n11379 0.0702092
R41330 vss.n11384 vss.n11383 0.0702092
R41331 vss.n11383 vss.t420 0.0702092
R41332 vss.n11386 vss.n11364 0.0702092
R41333 vss.t422 vss.n11364 0.0702092
R41334 vss.n11392 vss.n11391 0.0702092
R41335 vss.n11392 vss.t1463 0.0702092
R41336 vss.n11389 vss.n11388 0.0702092
R41337 vss.n11388 vss.t1463 0.0702092
R41338 vss.n11397 vss.n11396 0.0702092
R41339 vss.n11396 vss.t422 0.0702092
R41340 vss.n11382 vss.n11359 0.0702092
R41341 vss.t420 vss.n11382 0.0702092
R41342 vss.n11380 vss.n11376 0.0702092
R41343 vss.n11380 vss.t19 0.0702092
R41344 vss.n10954 vss.n10953 0.0702092
R41345 vss.t1368 vss.n10954 0.0702092
R41346 vss.n10959 vss.n10958 0.0702092
R41347 vss.n10958 vss.t813 0.0702092
R41348 vss.n10961 vss.n10939 0.0702092
R41349 vss.t815 vss.n10939 0.0702092
R41350 vss.n10967 vss.n10966 0.0702092
R41351 vss.n10967 vss.t1311 0.0702092
R41352 vss.n10964 vss.n10963 0.0702092
R41353 vss.n10963 vss.t1311 0.0702092
R41354 vss.n10972 vss.n10971 0.0702092
R41355 vss.n10971 vss.t815 0.0702092
R41356 vss.n10957 vss.n10934 0.0702092
R41357 vss.t813 vss.n10957 0.0702092
R41358 vss.n10955 vss.n10951 0.0702092
R41359 vss.n10955 vss.t1368 0.0702092
R41360 vss.n10791 vss.n10790 0.0702092
R41361 vss.t21 vss.n10791 0.0702092
R41362 vss.n10796 vss.n10795 0.0702092
R41363 vss.n10795 vss.t168 0.0702092
R41364 vss.n10798 vss.n10776 0.0702092
R41365 vss.t170 vss.n10776 0.0702092
R41366 vss.n10804 vss.n10803 0.0702092
R41367 vss.n10804 vss.t276 0.0702092
R41368 vss.n10801 vss.n10800 0.0702092
R41369 vss.n10800 vss.t276 0.0702092
R41370 vss.n10809 vss.n10808 0.0702092
R41371 vss.n10808 vss.t170 0.0702092
R41372 vss.n10794 vss.n10771 0.0702092
R41373 vss.t168 vss.n10794 0.0702092
R41374 vss.n10792 vss.n10788 0.0702092
R41375 vss.n10792 vss.t21 0.0702092
R41376 vss.n10747 vss.n10746 0.0702092
R41377 vss.t576 vss.n10747 0.0702092
R41378 vss.n10752 vss.n10751 0.0702092
R41379 vss.n10751 vss.t319 0.0702092
R41380 vss.n10754 vss.n10732 0.0702092
R41381 vss.t321 vss.n10732 0.0702092
R41382 vss.n10760 vss.n10759 0.0702092
R41383 vss.n10760 vss.t81 0.0702092
R41384 vss.n10757 vss.n10756 0.0702092
R41385 vss.n10756 vss.t81 0.0702092
R41386 vss.n10765 vss.n10764 0.0702092
R41387 vss.n10764 vss.t321 0.0702092
R41388 vss.n10750 vss.n10727 0.0702092
R41389 vss.t319 vss.n10750 0.0702092
R41390 vss.n10748 vss.n10744 0.0702092
R41391 vss.n10748 vss.t576 0.0702092
R41392 vss.n11573 vss.n11572 0.0702092
R41393 vss.t1364 vss.n11573 0.0702092
R41394 vss.n11578 vss.n11577 0.0702092
R41395 vss.n11577 vss.t663 0.0702092
R41396 vss.n11580 vss.n11558 0.0702092
R41397 vss.t665 vss.n11558 0.0702092
R41398 vss.n11586 vss.n11585 0.0702092
R41399 vss.n11586 vss.t120 0.0702092
R41400 vss.n11583 vss.n11582 0.0702092
R41401 vss.n11582 vss.t120 0.0702092
R41402 vss.n11591 vss.n11590 0.0702092
R41403 vss.n11590 vss.t665 0.0702092
R41404 vss.n11576 vss.n11553 0.0702092
R41405 vss.t663 vss.n11576 0.0702092
R41406 vss.n11574 vss.n11570 0.0702092
R41407 vss.n11574 vss.t1364 0.0702092
R41408 vss.n10570 vss.n10569 0.0702092
R41409 vss.t201 vss.n10570 0.0702092
R41410 vss.n10575 vss.n10574 0.0702092
R41411 vss.n10574 vss.t1143 0.0702092
R41412 vss.n10577 vss.n10555 0.0702092
R41413 vss.t1142 vss.n10555 0.0702092
R41414 vss.n10583 vss.n10582 0.0702092
R41415 vss.n10583 vss.t1145 0.0702092
R41416 vss.n10580 vss.n10579 0.0702092
R41417 vss.n10579 vss.t1145 0.0702092
R41418 vss.n10588 vss.n10587 0.0702092
R41419 vss.n10587 vss.t1142 0.0702092
R41420 vss.n10573 vss.n10550 0.0702092
R41421 vss.t1143 vss.n10573 0.0702092
R41422 vss.n10571 vss.n10567 0.0702092
R41423 vss.n10571 vss.t201 0.0702092
R41424 vss.n10526 vss.n10525 0.0702092
R41425 vss.t11 vss.n10526 0.0702092
R41426 vss.n10531 vss.n10530 0.0702092
R41427 vss.n10530 vss.t1388 0.0702092
R41428 vss.n10533 vss.n10511 0.0702092
R41429 vss.t1390 vss.n10511 0.0702092
R41430 vss.n10539 vss.n10538 0.0702092
R41431 vss.n10539 vss.t104 0.0702092
R41432 vss.n10536 vss.n10535 0.0702092
R41433 vss.n10535 vss.t104 0.0702092
R41434 vss.n10544 vss.n10543 0.0702092
R41435 vss.n10543 vss.t1390 0.0702092
R41436 vss.n10529 vss.n10506 0.0702092
R41437 vss.t1388 vss.n10529 0.0702092
R41438 vss.n10527 vss.n10523 0.0702092
R41439 vss.n10527 vss.t11 0.0702092
R41440 vss.n11947 vss.n11946 0.0702092
R41441 vss.t1481 vss.n11947 0.0702092
R41442 vss.n11952 vss.n11951 0.0702092
R41443 vss.n11951 vss.t1068 0.0702092
R41444 vss.n11954 vss.n11932 0.0702092
R41445 vss.t1070 vss.n11932 0.0702092
R41446 vss.n11960 vss.n11959 0.0702092
R41447 vss.n11960 vss.t113 0.0702092
R41448 vss.n11957 vss.n11956 0.0702092
R41449 vss.n11956 vss.t113 0.0702092
R41450 vss.n11965 vss.n11964 0.0702092
R41451 vss.n11964 vss.t1070 0.0702092
R41452 vss.n11950 vss.n11927 0.0702092
R41453 vss.t1068 vss.n11950 0.0702092
R41454 vss.n11948 vss.n11944 0.0702092
R41455 vss.n11948 vss.t1481 0.0702092
R41456 vss.n12072 vss.n12071 0.0702092
R41457 vss.n12071 vss.t128 0.0702092
R41458 vss.n12064 vss.t176 0.0702092
R41459 vss.t126 vss.n12068 0.0702092
R41460 vss.n12091 vss.t128 0.0702092
R41461 vss.n12069 vss.n11893 0.0702092
R41462 vss.n12069 vss.t126 0.0702092
R41463 vss.n12063 vss.n12062 0.0702092
R41464 vss.t176 vss.n12063 0.0702092
R41465 vss.n12065 vss.n12064 0.0702092
R41466 vss.n12068 vss.n12067 0.0702092
R41467 vss.n12092 vss.n12091 0.0702092
R41468 vss.n11909 vss.n11908 0.0702092
R41469 vss.n11909 vss.t958 0.0702092
R41470 vss.n11911 vss.t958 0.0702092
R41471 vss.n11912 vss.n11911 0.0702092
R41472 vss.n12053 vss.t305 0.0702092
R41473 vss.n12051 vss.t304 0.0702092
R41474 vss.n12047 vss.t939 0.0702092
R41475 vss.n11980 vss.n11979 0.0702092
R41476 vss.n11980 vss.t939 0.0702092
R41477 vss.n11977 vss.n11976 0.0702092
R41478 vss.n11976 vss.t304 0.0702092
R41479 vss.n11974 vss.n11973 0.0702092
R41480 vss.n11974 vss.t305 0.0702092
R41481 vss.n12054 vss.n12053 0.0702092
R41482 vss.n12051 vss.n12050 0.0702092
R41483 vss.n12048 vss.n12047 0.0702092
R41484 vss.n12034 vss.n12033 0.0702092
R41485 vss.n12034 vss.t1191 0.0702092
R41486 vss.n12038 vss.t1191 0.0702092
R41487 vss.n12039 vss.n12038 0.0702092
R41488 vss.n12024 vss.t1471 0.0702092
R41489 vss.n12028 vss.t700 0.0702092
R41490 vss.n12030 vss.t702 0.0702092
R41491 vss.n12017 vss.n12016 0.0702092
R41492 vss.n12017 vss.t702 0.0702092
R41493 vss.n12020 vss.n12019 0.0702092
R41494 vss.n12019 vss.t700 0.0702092
R41495 vss.n12023 vss.n12022 0.0702092
R41496 vss.t1471 vss.n12023 0.0702092
R41497 vss.n12025 vss.n12024 0.0702092
R41498 vss.n12028 vss.n12027 0.0702092
R41499 vss.n12031 vss.n12030 0.0702092
R41500 vss.n11997 vss.n11996 0.0702092
R41501 vss.n11997 vss.t1046 0.0702092
R41502 vss.n11999 vss.t1046 0.0702092
R41503 vss.n12000 vss.n11999 0.0702092
R41504 vss.n12001 vss.t237 0.0702092
R41505 vss.t239 vss.n12606 0.0702092
R41506 vss.n12602 vss.t1161 0.0702092
R41507 vss.n10606 vss.n10605 0.0702092
R41508 vss.n10606 vss.t1161 0.0702092
R41509 vss.n12608 vss.n12607 0.0702092
R41510 vss.n12607 vss.t239 0.0702092
R41511 vss.n11991 vss.n10592 0.0702092
R41512 vss.n11991 vss.t237 0.0702092
R41513 vss.n12002 vss.n12001 0.0702092
R41514 vss.n12606 vss.n12605 0.0702092
R41515 vss.n12603 vss.n12602 0.0702092
R41516 vss.n10613 vss.n10612 0.0702092
R41517 vss.n10613 vss.t232 0.0702092
R41518 vss.n12593 vss.t232 0.0702092
R41519 vss.n12594 vss.n12593 0.0702092
R41520 vss.n10644 vss.t444 0.0702092
R41521 vss.n10664 vss.t869 0.0702092
R41522 vss.n10662 vss.t871 0.0702092
R41523 vss.n10657 vss.n10656 0.0702092
R41524 vss.n10656 vss.t871 0.0702092
R41525 vss.n10655 vss.n10654 0.0702092
R41526 vss.n10654 vss.t869 0.0702092
R41527 vss.n10645 vss.n10643 0.0702092
R41528 vss.n10643 vss.t444 0.0702092
R41529 vss.n10667 vss.n10644 0.0702092
R41530 vss.n10665 vss.n10664 0.0702092
R41531 vss.n10662 vss.n10610 0.0702092
R41532 vss.n10642 vss.n10641 0.0702092
R41533 vss.t841 vss.n10642 0.0702092
R41534 vss.n10672 vss.t841 0.0702092
R41535 vss.n10673 vss.n10672 0.0702092
R41536 vss.t1245 vss.n10676 0.0702092
R41537 vss.n11606 vss.t1247 0.0702092
R41538 vss.n10624 vss.t1248 0.0702092
R41539 vss.n10625 vss.n10623 0.0702092
R41540 vss.n10623 vss.t1248 0.0702092
R41541 vss.n11601 vss.n11600 0.0702092
R41542 vss.n11601 vss.t1247 0.0702092
R41543 vss.n10678 vss.n10677 0.0702092
R41544 vss.n10677 vss.t1245 0.0702092
R41545 vss.n10676 vss.n10675 0.0702092
R41546 vss.n11607 vss.n11606 0.0702092
R41547 vss.n11609 vss.n10624 0.0702092
R41548 vss.n10618 vss.n10616 0.0702092
R41549 vss.n10616 vss.t685 0.0702092
R41550 vss.n10617 vss.t685 0.0702092
R41551 vss.n11620 vss.n10617 0.0702092
R41552 vss.n10831 vss.t1393 0.0702092
R41553 vss.n10851 vss.t683 0.0702092
R41554 vss.n11617 vss.t682 0.0702092
R41555 vss.n10847 vss.n10846 0.0702092
R41556 vss.n10846 vss.t682 0.0702092
R41557 vss.n10850 vss.n10849 0.0702092
R41558 vss.t683 vss.n10850 0.0702092
R41559 vss.n10832 vss.n10830 0.0702092
R41560 vss.n10830 vss.t1393 0.0702092
R41561 vss.n10854 vss.n10831 0.0702092
R41562 vss.n10852 vss.n10851 0.0702092
R41563 vss.n11618 vss.n11617 0.0702092
R41564 vss.n10862 vss.n10829 0.0702092
R41565 vss.n10862 vss.t950 0.0702092
R41566 vss.t950 vss.n10861 0.0702092
R41567 vss.n10861 vss.n10860 0.0702092
R41568 vss.n10865 vss.t401 0.0702092
R41569 vss.t400 vss.n11535 0.0702092
R41570 vss.n11531 vss.t403 0.0702092
R41571 vss.n10872 vss.n10871 0.0702092
R41572 vss.n10872 vss.t403 0.0702092
R41573 vss.n11537 vss.n11536 0.0702092
R41574 vss.n11536 vss.t400 0.0702092
R41575 vss.n10864 vss.n10813 0.0702092
R41576 vss.t401 vss.n10864 0.0702092
R41577 vss.n10866 vss.n10865 0.0702092
R41578 vss.n11535 vss.n11534 0.0702092
R41579 vss.n11532 vss.n11531 0.0702092
R41580 vss.n11519 vss.n11518 0.0702092
R41581 vss.n11519 vss.t142 0.0702092
R41582 vss.n11522 vss.t142 0.0702092
R41583 vss.n11523 vss.n11522 0.0702092
R41584 vss.n11509 vss.t861 0.0702092
R41585 vss.n11513 vss.t376 0.0702092
R41586 vss.n11515 vss.t378 0.0702092
R41587 vss.n11502 vss.n11501 0.0702092
R41588 vss.n11502 vss.t378 0.0702092
R41589 vss.n11505 vss.n11504 0.0702092
R41590 vss.n11504 vss.t376 0.0702092
R41591 vss.n11508 vss.n11507 0.0702092
R41592 vss.t861 vss.n11508 0.0702092
R41593 vss.n11510 vss.n11509 0.0702092
R41594 vss.n11513 vss.n11512 0.0702092
R41595 vss.n11516 vss.n11515 0.0702092
R41596 vss.n10888 vss.n10887 0.0702092
R41597 vss.n10888 vss.t993 0.0702092
R41598 vss.n10890 vss.t993 0.0702092
R41599 vss.n10891 vss.n10890 0.0702092
R41600 vss.n11488 vss.t693 0.0702092
R41601 vss.n11486 vss.t692 0.0702092
R41602 vss.n11482 vss.t711 0.0702092
R41603 vss.n10978 vss.n10898 0.0702092
R41604 vss.n10898 vss.t711 0.0702092
R41605 vss.n10986 vss.n10985 0.0702092
R41606 vss.n10985 vss.t692 0.0702092
R41607 vss.n10980 vss.n10977 0.0702092
R41608 vss.n10980 vss.t693 0.0702092
R41609 vss.n11489 vss.n11488 0.0702092
R41610 vss.n11486 vss.n11485 0.0702092
R41611 vss.n11483 vss.n11482 0.0702092
R41612 vss.n11471 vss.n11470 0.0702092
R41613 vss.n11471 vss.t1459 0.0702092
R41614 vss.n11473 vss.t1459 0.0702092
R41615 vss.n11474 vss.n11473 0.0702092
R41616 vss.n11461 vss.t593 0.0702092
R41617 vss.n11465 vss.t1099 0.0702092
R41618 vss.n11467 vss.t1098 0.0702092
R41619 vss.n11454 vss.n11453 0.0702092
R41620 vss.n11454 vss.t1098 0.0702092
R41621 vss.n11457 vss.n11456 0.0702092
R41622 vss.n11456 vss.t1099 0.0702092
R41623 vss.n11460 vss.n11459 0.0702092
R41624 vss.t593 vss.n11460 0.0702092
R41625 vss.n11462 vss.n11461 0.0702092
R41626 vss.n11465 vss.n11464 0.0702092
R41627 vss.n11468 vss.n11467 0.0702092
R41628 vss.n10917 vss.n10916 0.0702092
R41629 vss.n10917 vss.t954 0.0702092
R41630 vss.n10919 vss.t954 0.0702092
R41631 vss.n10920 vss.n10919 0.0702092
R41632 vss.n10921 vss.t976 0.0702092
R41633 vss.n12749 vss.t978 0.0702092
R41634 vss.n10331 vss.t317 0.0702092
R41635 vss.n10332 vss.n10330 0.0702092
R41636 vss.n10330 vss.t317 0.0702092
R41637 vss.n12744 vss.n12743 0.0702092
R41638 vss.n12744 vss.t978 0.0702092
R41639 vss.n10911 vss.n10338 0.0702092
R41640 vss.n10911 vss.t976 0.0702092
R41641 vss.n10922 vss.n10921 0.0702092
R41642 vss.n12750 vss.n12749 0.0702092
R41643 vss.n12752 vss.n10331 0.0702092
R41644 vss.n10325 vss.n10323 0.0702092
R41645 vss.n10323 vss.t1147 0.0702092
R41646 vss.n10324 vss.t1147 0.0702092
R41647 vss.n12763 vss.n10324 0.0702092
R41648 vss.n12729 vss.t655 0.0702092
R41649 vss.t1216 vss.n12733 0.0702092
R41650 vss.n12760 vss.t1218 0.0702092
R41651 vss.n12737 vss.n12736 0.0702092
R41652 vss.n12736 vss.t1218 0.0702092
R41653 vss.n12734 vss.n10342 0.0702092
R41654 vss.n12734 vss.t1216 0.0702092
R41655 vss.n12728 vss.n12727 0.0702092
R41656 vss.t655 vss.n12728 0.0702092
R41657 vss.n12730 vss.n12729 0.0702092
R41658 vss.n12733 vss.n12732 0.0702092
R41659 vss.n12761 vss.n12760 0.0702092
R41660 vss.n10358 vss.n10357 0.0702092
R41661 vss.n10358 vss.t1001 0.0702092
R41662 vss.n10360 vss.t1001 0.0702092
R41663 vss.n10361 vss.n10360 0.0702092
R41664 vss.n12718 vss.t1250 0.0702092
R41665 vss.n12716 vss.t1252 0.0702092
R41666 vss.n12712 vss.t1172 0.0702092
R41667 vss.n12709 vss.n12708 0.0702092
R41668 vss.n12709 vss.t1172 0.0702092
R41669 vss.n12706 vss.n12705 0.0702092
R41670 vss.n12705 vss.t1252 0.0702092
R41671 vss.n12703 vss.n12702 0.0702092
R41672 vss.n12703 vss.t1250 0.0702092
R41673 vss.n12719 vss.n12718 0.0702092
R41674 vss.n12716 vss.n12715 0.0702092
R41675 vss.n12713 vss.n12712 0.0702092
R41676 vss.n2300 vss.n2260 0.0702092
R41677 vss.n2260 vss.t1241 0.0702092
R41678 vss.n2287 vss.n2286 0.0702092
R41679 vss.n2286 vss.t1511 0.0702092
R41680 vss.n2281 vss.n2279 0.0702092
R41681 vss.t185 vss.n2279 0.0702092
R41682 vss.n2298 vss.n2297 0.0702092
R41683 vss.n2297 vss.t187 0.0702092
R41684 vss.n2261 vss.n2259 0.0702092
R41685 vss.n2259 vss.t1241 0.0702092
R41686 vss.n2296 vss.n2295 0.0702092
R41687 vss.t187 vss.n2296 0.0702092
R41688 vss.n2293 vss.n2292 0.0702092
R41689 vss.n2292 vss.t185 0.0702092
R41690 vss.n2284 vss.n2283 0.0702092
R41691 vss.n2284 vss.t1511 0.0702092
R41692 vss.n12998 vss.n2258 0.0702092
R41693 vss.n12998 vss.t926 0.0702092
R41694 vss.n13009 vss.n13008 0.0702092
R41695 vss.t500 vss.n13009 0.0702092
R41696 vss.n13016 vss.n13015 0.0702092
R41697 vss.n13015 vss.t642 0.0702092
R41698 vss.n13000 vss.n2242 0.0702092
R41699 vss.t644 vss.n13000 0.0702092
R41700 vss.n12997 vss.n12996 0.0702092
R41701 vss.t926 vss.n12997 0.0702092
R41702 vss.n13002 vss.n13001 0.0702092
R41703 vss.n13001 vss.t644 0.0702092
R41704 vss.n13014 vss.n13013 0.0702092
R41705 vss.t642 vss.n13014 0.0702092
R41706 vss.n13011 vss.n13010 0.0702092
R41707 vss.n13010 vss.t500 0.0702092
R41708 vss.n13919 vss.n13918 0.0702092
R41709 vss.t434 vss.n13919 0.0702092
R41710 vss.n13916 vss.n13915 0.0702092
R41711 vss.n13915 vss.t249 0.0702092
R41712 vss.n13903 vss.n13902 0.0702092
R41713 vss.n13902 vss.t250 0.0702092
R41714 vss.t434 vss.n13304 0.0702092
R41715 vss.t249 vss.n13914 0.0702092
R41716 vss.n13910 vss.t250 0.0702092
R41717 vss.n13911 vss.n13910 0.0702092
R41718 vss.n13914 vss.n13913 0.0702092
R41719 vss.n13314 vss.n13304 0.0702092
R41720 vss.n13908 vss.n13323 0.0702092
R41721 vss.n13908 vss.t914 0.0702092
R41722 vss.n13907 vss.n13906 0.0702092
R41723 vss.t914 vss.n13907 0.0702092
R41724 vss.n13882 vss.n13881 0.0702092
R41725 vss.n13881 vss.t681 0.0702092
R41726 vss.n13886 vss.n13885 0.0702092
R41727 vss.n13886 vss.t679 0.0702092
R41728 vss.n13328 vss.n13326 0.0702092
R41729 vss.n13326 vss.t820 0.0702092
R41730 vss.t681 vss.n13880 0.0702092
R41731 vss.n13891 vss.t679 0.0702092
R41732 vss.n13327 vss.t820 0.0702092
R41733 vss.n13894 vss.n13327 0.0702092
R41734 vss.n13892 vss.n13891 0.0702092
R41735 vss.n13880 vss.n13879 0.0702092
R41736 vss.n13877 vss.n13876 0.0702092
R41737 vss.n13876 vss.t268 0.0702092
R41738 vss.n13875 vss.n13874 0.0702092
R41739 vss.t268 vss.n13875 0.0702092
R41740 vss.n13871 vss.n13870 0.0702092
R41741 vss.t1454 vss.n13871 0.0702092
R41742 vss.n13868 vss.n13867 0.0702092
R41743 vss.n13867 vss.t806 0.0702092
R41744 vss.n13848 vss.n13847 0.0702092
R41745 vss.n13847 vss.t807 0.0702092
R41746 vss.t1454 vss.n13346 0.0702092
R41747 vss.t806 vss.n13866 0.0702092
R41748 vss.n13855 vss.t807 0.0702092
R41749 vss.n13856 vss.n13855 0.0702092
R41750 vss.n13866 vss.n13865 0.0702092
R41751 vss.n13356 vss.n13346 0.0702092
R41752 vss.n13853 vss.n13362 0.0702092
R41753 vss.n13853 vss.t1024 0.0702092
R41754 vss.n13852 vss.n13851 0.0702092
R41755 vss.t1024 vss.n13852 0.0702092
R41756 vss.n13828 vss.n13827 0.0702092
R41757 vss.n13827 vss.t1415 0.0702092
R41758 vss.n13832 vss.n13831 0.0702092
R41759 vss.n13832 vss.t1413 0.0702092
R41760 vss.n13367 vss.n13365 0.0702092
R41761 vss.n13365 vss.t111 0.0702092
R41762 vss.t1415 vss.n13826 0.0702092
R41763 vss.n13837 vss.t1413 0.0702092
R41764 vss.n13366 vss.t111 0.0702092
R41765 vss.n13840 vss.n13366 0.0702092
R41766 vss.n13838 vss.n13837 0.0702092
R41767 vss.n13826 vss.n13825 0.0702092
R41768 vss.n13823 vss.n13822 0.0702092
R41769 vss.n13822 vss.t722 0.0702092
R41770 vss.n13821 vss.n13820 0.0702092
R41771 vss.t722 vss.n13821 0.0702092
R41772 vss.n13817 vss.n13816 0.0702092
R41773 vss.t730 vss.n13817 0.0702092
R41774 vss.n13814 vss.n13813 0.0702092
R41775 vss.n13813 vss.t715 0.0702092
R41776 vss.n13798 vss.n13797 0.0702092
R41777 vss.n13797 vss.t716 0.0702092
R41778 vss.t730 vss.n13387 0.0702092
R41779 vss.t715 vss.n13812 0.0702092
R41780 vss.n13805 vss.t716 0.0702092
R41781 vss.n13806 vss.n13805 0.0702092
R41782 vss.n13812 vss.n13811 0.0702092
R41783 vss.n13397 vss.n13387 0.0702092
R41784 vss.n13803 vss.n13403 0.0702092
R41785 vss.n13803 vss.t47 0.0702092
R41786 vss.n13802 vss.n13801 0.0702092
R41787 vss.t47 vss.n13802 0.0702092
R41788 vss.n13777 vss.n13776 0.0702092
R41789 vss.n13776 vss.t307 0.0702092
R41790 vss.n13781 vss.n13780 0.0702092
R41791 vss.n13781 vss.t308 0.0702092
R41792 vss.n13408 vss.n13406 0.0702092
R41793 vss.n13406 vss.t795 0.0702092
R41794 vss.t307 vss.n13775 0.0702092
R41795 vss.n13786 vss.t308 0.0702092
R41796 vss.n13407 vss.t795 0.0702092
R41797 vss.n13789 vss.n13407 0.0702092
R41798 vss.n13787 vss.n13786 0.0702092
R41799 vss.n13775 vss.n13774 0.0702092
R41800 vss.n13772 vss.n13771 0.0702092
R41801 vss.n13771 vss.t516 0.0702092
R41802 vss.n13770 vss.n13769 0.0702092
R41803 vss.t516 vss.n13770 0.0702092
R41804 vss.n13766 vss.n13765 0.0702092
R41805 vss.t1470 vss.n13766 0.0702092
R41806 vss.n13763 vss.n13762 0.0702092
R41807 vss.n13762 vss.t1416 0.0702092
R41808 vss.n13743 vss.n13742 0.0702092
R41809 vss.n13742 vss.t1417 0.0702092
R41810 vss.t1470 vss.n13426 0.0702092
R41811 vss.t1416 vss.n13761 0.0702092
R41812 vss.n13750 vss.t1417 0.0702092
R41813 vss.n13751 vss.n13750 0.0702092
R41814 vss.n13761 vss.n13760 0.0702092
R41815 vss.n13436 vss.n13426 0.0702092
R41816 vss.n13748 vss.n13442 0.0702092
R41817 vss.n13748 vss.t1026 0.0702092
R41818 vss.n13747 vss.n13746 0.0702092
R41819 vss.t1026 vss.n13747 0.0702092
R41820 vss.n13723 vss.n13722 0.0702092
R41821 vss.n13722 vss.t1432 0.0702092
R41822 vss.n13727 vss.n13726 0.0702092
R41823 vss.n13727 vss.t1433 0.0702092
R41824 vss.n13447 vss.n13445 0.0702092
R41825 vss.n13445 vss.t1391 0.0702092
R41826 vss.t1432 vss.n13721 0.0702092
R41827 vss.n13732 vss.t1433 0.0702092
R41828 vss.n13446 vss.t1391 0.0702092
R41829 vss.n13735 vss.n13446 0.0702092
R41830 vss.n13733 vss.n13732 0.0702092
R41831 vss.n13721 vss.n13720 0.0702092
R41832 vss.n13718 vss.n13717 0.0702092
R41833 vss.n13717 vss.t687 0.0702092
R41834 vss.n13716 vss.n13715 0.0702092
R41835 vss.t687 vss.n13716 0.0702092
R41836 vss.n13712 vss.n13711 0.0702092
R41837 vss.t1386 vss.n13712 0.0702092
R41838 vss.n13709 vss.n13708 0.0702092
R41839 vss.n13708 vss.t1288 0.0702092
R41840 vss.n13693 vss.n13692 0.0702092
R41841 vss.n13692 vss.t1289 0.0702092
R41842 vss.t1386 vss.n13467 0.0702092
R41843 vss.t1288 vss.n13707 0.0702092
R41844 vss.n13700 vss.t1289 0.0702092
R41845 vss.n13701 vss.n13700 0.0702092
R41846 vss.n13707 vss.n13706 0.0702092
R41847 vss.n13477 vss.n13467 0.0702092
R41848 vss.n13698 vss.n13483 0.0702092
R41849 vss.n13698 vss.t991 0.0702092
R41850 vss.n13697 vss.n13696 0.0702092
R41851 vss.t991 vss.n13697 0.0702092
R41852 vss.n13672 vss.n13671 0.0702092
R41853 vss.n13671 vss.t271 0.0702092
R41854 vss.n13676 vss.n13675 0.0702092
R41855 vss.n13676 vss.t269 0.0702092
R41856 vss.n13488 vss.n13486 0.0702092
R41857 vss.n13486 vss.t826 0.0702092
R41858 vss.t271 vss.n13670 0.0702092
R41859 vss.n13681 vss.t269 0.0702092
R41860 vss.n13487 vss.t826 0.0702092
R41861 vss.n13684 vss.n13487 0.0702092
R41862 vss.n13682 vss.n13681 0.0702092
R41863 vss.n13670 vss.n13669 0.0702092
R41864 vss.n13667 vss.n13666 0.0702092
R41865 vss.n13666 vss.t1128 0.0702092
R41866 vss.n13665 vss.n13664 0.0702092
R41867 vss.t1128 vss.n13665 0.0702092
R41868 vss.n13661 vss.n13660 0.0702092
R41869 vss.t261 vss.n13661 0.0702092
R41870 vss.n13658 vss.n13657 0.0702092
R41871 vss.n13657 vss.t630 0.0702092
R41872 vss.n13638 vss.n13637 0.0702092
R41873 vss.n13637 vss.t631 0.0702092
R41874 vss.t261 vss.n13506 0.0702092
R41875 vss.t630 vss.n13656 0.0702092
R41876 vss.n13645 vss.t631 0.0702092
R41877 vss.n13646 vss.n13645 0.0702092
R41878 vss.n13656 vss.n13655 0.0702092
R41879 vss.n13516 vss.n13506 0.0702092
R41880 vss.n13643 vss.n13522 0.0702092
R41881 vss.n13643 vss.t1040 0.0702092
R41882 vss.n13642 vss.n13641 0.0702092
R41883 vss.t1040 vss.n13642 0.0702092
R41884 vss.n13618 vss.n13617 0.0702092
R41885 vss.n13617 vss.t1383 0.0702092
R41886 vss.n13622 vss.n13621 0.0702092
R41887 vss.n13622 vss.t1384 0.0702092
R41888 vss.n13527 vss.n13525 0.0702092
R41889 vss.n13525 vss.t107 0.0702092
R41890 vss.t1383 vss.n13616 0.0702092
R41891 vss.n13627 vss.t1384 0.0702092
R41892 vss.n13526 vss.t107 0.0702092
R41893 vss.n13630 vss.n13526 0.0702092
R41894 vss.n13628 vss.n13627 0.0702092
R41895 vss.n13616 vss.n13615 0.0702092
R41896 vss.n13613 vss.n13612 0.0702092
R41897 vss.n13612 vss.t988 0.0702092
R41898 vss.n13611 vss.n13610 0.0702092
R41899 vss.t988 vss.n13611 0.0702092
R41900 vss.n13605 vss.n13546 0.0702092
R41901 vss.n13546 vss.t770 0.0702092
R41902 vss.n13585 vss.n13565 0.0702092
R41903 vss.t1262 vss.n13565 0.0702092
R41904 vss.n13603 vss.n13602 0.0702092
R41905 vss.n13602 vss.t1264 0.0702092
R41906 vss.n13547 vss.n13545 0.0702092
R41907 vss.n13545 vss.t770 0.0702092
R41908 vss.n13601 vss.n13600 0.0702092
R41909 vss.t1264 vss.n13601 0.0702092
R41910 vss.n13598 vss.n13597 0.0702092
R41911 vss.n13597 vss.t1262 0.0702092
R41912 vss.n14148 vss.n14147 0.0702092
R41913 vss.t1272 vss.n14148 0.0702092
R41914 vss.n13579 vss.n13567 0.0702092
R41915 vss.n13567 vss.t816 0.0702092
R41916 vss.n13572 vss.n474 0.0702092
R41917 vss.t1273 vss.n13572 0.0702092
R41918 vss.n14150 vss.n14149 0.0702092
R41919 vss.n14149 vss.t1272 0.0702092
R41920 vss.n13574 vss.n13573 0.0702092
R41921 vss.t1273 vss.n13574 0.0702092
R41922 vss.n13568 vss.n13566 0.0702092
R41923 vss.n13566 vss.t816 0.0702092
R41924 vss.n13592 vss.n13591 0.0702092
R41925 vss.n13591 vss.t1018 0.0702092
R41926 vss.n13590 vss.n13589 0.0702092
R41927 vss.t1018 vss.n13590 0.0702092
R41928 vss.n14736 vss.n172 0.0702092
R41929 vss.n14736 vss.t1192 0.0702092
R41930 vss.n14747 vss.n14746 0.0702092
R41931 vss.t613 vss.n14747 0.0702092
R41932 vss.n14754 vss.n14753 0.0702092
R41933 vss.n14753 vss.t1112 0.0702092
R41934 vss.n14738 vss.n156 0.0702092
R41935 vss.t1111 vss.n14738 0.0702092
R41936 vss.n14735 vss.n14734 0.0702092
R41937 vss.t1192 vss.n14735 0.0702092
R41938 vss.n14740 vss.n14739 0.0702092
R41939 vss.n14739 vss.t1111 0.0702092
R41940 vss.n14752 vss.n14751 0.0702092
R41941 vss.t1112 vss.n14752 0.0702092
R41942 vss.n14749 vss.n14748 0.0702092
R41943 vss.n14748 vss.t613 0.0702092
R41944 vss.n14680 vss.n195 0.0702092
R41945 vss.n195 vss.t430 0.0702092
R41946 vss.n14667 vss.n14666 0.0702092
R41947 vss.n14666 vss.t1497 0.0702092
R41948 vss.n14661 vss.n14659 0.0702092
R41949 vss.t1050 vss.n14659 0.0702092
R41950 vss.n14678 vss.n14677 0.0702092
R41951 vss.n14677 vss.t1052 0.0702092
R41952 vss.n196 vss.n194 0.0702092
R41953 vss.n194 vss.t430 0.0702092
R41954 vss.n14676 vss.n14675 0.0702092
R41955 vss.t1052 vss.n14676 0.0702092
R41956 vss.n14673 vss.n14672 0.0702092
R41957 vss.n14672 vss.t1050 0.0702092
R41958 vss.n14664 vss.n14663 0.0702092
R41959 vss.n14664 vss.t1497 0.0702092
R41960 vss.n14541 vss.n249 0.0702092
R41961 vss.n14541 vss.t1168 0.0702092
R41962 vss.n14552 vss.n14551 0.0702092
R41963 vss.t1324 vss.n14552 0.0702092
R41964 vss.n14559 vss.n14558 0.0702092
R41965 vss.n14558 vss.t362 0.0702092
R41966 vss.n14543 vss.n233 0.0702092
R41967 vss.t364 vss.n14543 0.0702092
R41968 vss.n14540 vss.n14539 0.0702092
R41969 vss.t1168 vss.n14540 0.0702092
R41970 vss.n14545 vss.n14544 0.0702092
R41971 vss.n14544 vss.t364 0.0702092
R41972 vss.n14557 vss.n14556 0.0702092
R41973 vss.t362 vss.n14557 0.0702092
R41974 vss.n14554 vss.n14553 0.0702092
R41975 vss.n14553 vss.t1324 0.0702092
R41976 vss.n14485 vss.n254 0.0702092
R41977 vss.n254 vss.t1285 0.0702092
R41978 vss.n14472 vss.n14471 0.0702092
R41979 vss.n14471 vss.t381 0.0702092
R41980 vss.n14466 vss.n14464 0.0702092
R41981 vss.t834 vss.n14464 0.0702092
R41982 vss.n14483 vss.n14482 0.0702092
R41983 vss.n14482 vss.t833 0.0702092
R41984 vss.n255 vss.n253 0.0702092
R41985 vss.n253 vss.t1285 0.0702092
R41986 vss.n14481 vss.n14480 0.0702092
R41987 vss.t833 vss.n14481 0.0702092
R41988 vss.n14478 vss.n14477 0.0702092
R41989 vss.n14477 vss.t834 0.0702092
R41990 vss.n14469 vss.n14468 0.0702092
R41991 vss.n14469 vss.t381 0.0702092
R41992 vss.n14346 vss.n308 0.0702092
R41993 vss.n14346 vss.t1049 0.0702092
R41994 vss.n14357 vss.n14356 0.0702092
R41995 vss.t1350 vss.n14357 0.0702092
R41996 vss.n14364 vss.n14363 0.0702092
R41997 vss.n14363 vss.t1102 0.0702092
R41998 vss.n14348 vss.n292 0.0702092
R41999 vss.t1101 vss.n14348 0.0702092
R42000 vss.n14345 vss.n14344 0.0702092
R42001 vss.t1049 vss.n14345 0.0702092
R42002 vss.n14350 vss.n14349 0.0702092
R42003 vss.n14349 vss.t1101 0.0702092
R42004 vss.n14362 vss.n14361 0.0702092
R42005 vss.t1102 vss.n14362 0.0702092
R42006 vss.n14359 vss.n14358 0.0702092
R42007 vss.n14358 vss.t1350 0.0702092
R42008 vss.n14290 vss.n313 0.0702092
R42009 vss.n313 vss.t300 0.0702092
R42010 vss.n14277 vss.n14276 0.0702092
R42011 vss.n14276 vss.t502 0.0702092
R42012 vss.n14271 vss.n14269 0.0702092
R42013 vss.t156 vss.n14269 0.0702092
R42014 vss.n14288 vss.n14287 0.0702092
R42015 vss.n14287 vss.t158 0.0702092
R42016 vss.n314 vss.n312 0.0702092
R42017 vss.n312 vss.t300 0.0702092
R42018 vss.n14286 vss.n14285 0.0702092
R42019 vss.t158 vss.n14286 0.0702092
R42020 vss.n14283 vss.n14282 0.0702092
R42021 vss.n14282 vss.t156 0.0702092
R42022 vss.n14274 vss.n14273 0.0702092
R42023 vss.n14274 vss.t502 0.0702092
R42024 vss.n14227 vss.n431 0.0702092
R42025 vss.n14227 vss.t429 0.0702092
R42026 vss.n14238 vss.n14237 0.0702092
R42027 vss.t1332 vss.n14238 0.0702092
R42028 vss.n14245 vss.n14244 0.0702092
R42029 vss.n14244 vss.t1189 0.0702092
R42030 vss.n14229 vss.n415 0.0702092
R42031 vss.t1188 vss.n14229 0.0702092
R42032 vss.n14226 vss.n14225 0.0702092
R42033 vss.t429 vss.n14226 0.0702092
R42034 vss.n14231 vss.n14230 0.0702092
R42035 vss.n14230 vss.t1188 0.0702092
R42036 vss.n14243 vss.n14242 0.0702092
R42037 vss.t1189 vss.n14243 0.0702092
R42038 vss.n14240 vss.n14239 0.0702092
R42039 vss.n14239 vss.t1332 0.0702092
R42040 vss.n14118 vss.n14113 0.0702092
R42041 vss.n14118 vss.t718 0.0702092
R42042 vss.n14129 vss.n14128 0.0702092
R42043 vss.t393 vss.n14129 0.0702092
R42044 vss.n14136 vss.n14135 0.0702092
R42045 vss.n14135 vss.t1225 0.0702092
R42046 vss.n14120 vss.n14097 0.0702092
R42047 vss.t1224 vss.n14120 0.0702092
R42048 vss.n14117 vss.n14116 0.0702092
R42049 vss.t718 vss.n14117 0.0702092
R42050 vss.n14122 vss.n14121 0.0702092
R42051 vss.n14121 vss.t1224 0.0702092
R42052 vss.n14134 vss.n14133 0.0702092
R42053 vss.t1225 vss.n14134 0.0702092
R42054 vss.n14131 vss.n14130 0.0702092
R42055 vss.n14130 vss.t393 0.0702092
R42056 vss.n14217 vss.n14178 0.0702092
R42057 vss.n14178 vss.t1524 0.0702092
R42058 vss.n14204 vss.n14203 0.0702092
R42059 vss.n14203 vss.t1316 0.0702092
R42060 vss.n14198 vss.n14196 0.0702092
R42061 vss.t1522 vss.n14196 0.0702092
R42062 vss.n14215 vss.n14214 0.0702092
R42063 vss.n14214 vss.t1521 0.0702092
R42064 vss.n14179 vss.n14177 0.0702092
R42065 vss.n14177 vss.t1524 0.0702092
R42066 vss.n14213 vss.n14212 0.0702092
R42067 vss.t1521 vss.n14213 0.0702092
R42068 vss.n14210 vss.n14209 0.0702092
R42069 vss.n14209 vss.t1522 0.0702092
R42070 vss.n14201 vss.n14200 0.0702092
R42071 vss.n14201 vss.t1316 0.0702092
R42072 vss.n339 vss.n334 0.0702092
R42073 vss.n339 vss.t88 0.0702092
R42074 vss.n350 vss.n349 0.0702092
R42075 vss.t1352 vss.n350 0.0702092
R42076 vss.n357 vss.n356 0.0702092
R42077 vss.n356 vss.t1404 0.0702092
R42078 vss.n341 vss.n318 0.0702092
R42079 vss.t1403 vss.n341 0.0702092
R42080 vss.n338 vss.n337 0.0702092
R42081 vss.t88 vss.n338 0.0702092
R42082 vss.n343 vss.n342 0.0702092
R42083 vss.n342 vss.t1403 0.0702092
R42084 vss.n355 vss.n354 0.0702092
R42085 vss.t1404 vss.n355 0.0702092
R42086 vss.n352 vss.n351 0.0702092
R42087 vss.n351 vss.t1352 0.0702092
R42088 vss.n14336 vss.n14297 0.0702092
R42089 vss.n14297 vss.t368 0.0702092
R42090 vss.n14323 vss.n14322 0.0702092
R42091 vss.n14322 vss.t1477 0.0702092
R42092 vss.n14317 vss.n14315 0.0702092
R42093 vss.t754 vss.n14315 0.0702092
R42094 vss.n14334 vss.n14333 0.0702092
R42095 vss.n14333 vss.t753 0.0702092
R42096 vss.n14298 vss.n14296 0.0702092
R42097 vss.n14296 vss.t368 0.0702092
R42098 vss.n14332 vss.n14331 0.0702092
R42099 vss.t753 vss.n14332 0.0702092
R42100 vss.n14329 vss.n14328 0.0702092
R42101 vss.n14328 vss.t754 0.0702092
R42102 vss.n14320 vss.n14319 0.0702092
R42103 vss.n14320 vss.t1477 0.0702092
R42104 vss.n14392 vss.n14387 0.0702092
R42105 vss.n14392 vss.t1312 0.0702092
R42106 vss.n14403 vss.n14402 0.0702092
R42107 vss.t466 vss.n14403 0.0702092
R42108 vss.n14410 vss.n14409 0.0702092
R42109 vss.n14409 vss.t1208 0.0702092
R42110 vss.n14394 vss.n14371 0.0702092
R42111 vss.t1207 vss.n14394 0.0702092
R42112 vss.n14391 vss.n14390 0.0702092
R42113 vss.t1312 vss.n14391 0.0702092
R42114 vss.n14396 vss.n14395 0.0702092
R42115 vss.n14395 vss.t1207 0.0702092
R42116 vss.n14408 vss.n14407 0.0702092
R42117 vss.t1208 vss.n14408 0.0702092
R42118 vss.n14405 vss.n14404 0.0702092
R42119 vss.n14404 vss.t466 0.0702092
R42120 vss.n14531 vss.n14492 0.0702092
R42121 vss.n14492 vss.t1053 0.0702092
R42122 vss.n14518 vss.n14517 0.0702092
R42123 vss.n14517 vss.t1077 0.0702092
R42124 vss.n14512 vss.n14510 0.0702092
R42125 vss.t266 vss.n14510 0.0702092
R42126 vss.n14529 vss.n14528 0.0702092
R42127 vss.n14528 vss.t265 0.0702092
R42128 vss.n14493 vss.n14491 0.0702092
R42129 vss.n14491 vss.t1053 0.0702092
R42130 vss.n14527 vss.n14526 0.0702092
R42131 vss.t265 vss.n14527 0.0702092
R42132 vss.n14524 vss.n14523 0.0702092
R42133 vss.n14523 vss.t266 0.0702092
R42134 vss.n14515 vss.n14514 0.0702092
R42135 vss.n14515 vss.t1077 0.0702092
R42136 vss.n14587 vss.n14582 0.0702092
R42137 vss.n14587 vss.t984 0.0702092
R42138 vss.n14598 vss.n14597 0.0702092
R42139 vss.t1336 vss.n14598 0.0702092
R42140 vss.n14605 vss.n14604 0.0702092
R42141 vss.n14604 vss.t74 0.0702092
R42142 vss.n14589 vss.n14566 0.0702092
R42143 vss.t73 vss.n14589 0.0702092
R42144 vss.n14586 vss.n14585 0.0702092
R42145 vss.t984 vss.n14586 0.0702092
R42146 vss.n14591 vss.n14590 0.0702092
R42147 vss.n14590 vss.t73 0.0702092
R42148 vss.n14603 vss.n14602 0.0702092
R42149 vss.t74 vss.n14603 0.0702092
R42150 vss.n14600 vss.n14599 0.0702092
R42151 vss.n14599 vss.t1336 0.0702092
R42152 vss.n14726 vss.n14687 0.0702092
R42153 vss.n14687 vss.t562 0.0702092
R42154 vss.n14713 vss.n14712 0.0702092
R42155 vss.n14712 vss.t474 0.0702092
R42156 vss.n14707 vss.n14705 0.0702092
R42157 vss.t346 vss.n14705 0.0702092
R42158 vss.n14724 vss.n14723 0.0702092
R42159 vss.n14723 vss.t345 0.0702092
R42160 vss.n14688 vss.n14686 0.0702092
R42161 vss.n14686 vss.t562 0.0702092
R42162 vss.n14722 vss.n14721 0.0702092
R42163 vss.t345 vss.n14722 0.0702092
R42164 vss.n14719 vss.n14718 0.0702092
R42165 vss.n14718 vss.t346 0.0702092
R42166 vss.n14710 vss.n14709 0.0702092
R42167 vss.n14710 vss.t474 0.0702092
R42168 vss.n186 vss.n174 0.0702092
R42169 vss.n174 vss.t853 0.0702092
R42170 vss.n17 vss.n16 0.0702092
R42171 vss.t1081 vss.n17 0.0702092
R42172 vss.n14791 vss.n14790 0.0702092
R42173 vss.n14790 vss.t1109 0.0702092
R42174 vss.n179 vss.n2 0.0702092
R42175 vss.t1108 vss.n179 0.0702092
R42176 vss.n175 vss.n173 0.0702092
R42177 vss.n173 vss.t853 0.0702092
R42178 vss.n181 vss.n180 0.0702092
R42179 vss.t1108 vss.n181 0.0702092
R42180 vss.n14789 vss.n14788 0.0702092
R42181 vss.t1109 vss.n14789 0.0702092
R42182 vss.n14786 vss.n14785 0.0702092
R42183 vss.n14785 vss.t1081 0.0702092
R42184 vss.n14010 vss.n14009 0.0702092
R42185 vss.n14009 vss.t294 0.0702092
R42186 vss.n14012 vss.n523 0.0702092
R42187 vss.t296 vss.n523 0.0702092
R42188 vss.n14018 vss.n14017 0.0702092
R42189 vss.n14018 vss.t512 0.0702092
R42190 vss.n14015 vss.n14014 0.0702092
R42191 vss.n14014 vss.t512 0.0702092
R42192 vss.n14023 vss.n14022 0.0702092
R42193 vss.n14022 vss.t296 0.0702092
R42194 vss.n14008 vss.n518 0.0702092
R42195 vss.t294 vss.n14008 0.0702092
R42196 vss.n14006 vss.n535 0.0702092
R42197 vss.t999 vss.n14005 0.0702092
R42198 vss.n14006 vss.t999 0.0702092
R42199 vss.n14005 vss.n14004 0.0702092
R42200 vss.n13998 vss.n538 0.0702092
R42201 vss.n538 vss.t653 0.0702092
R42202 vss.n13996 vss.n13995 0.0702092
R42203 vss.n13995 vss.t673 0.0702092
R42204 vss.n673 vss.n672 0.0702092
R42205 vss.n672 vss.t675 0.0702092
R42206 vss.n671 vss.n552 0.0702092
R42207 vss.t675 vss.n671 0.0702092
R42208 vss.n13994 vss.n13993 0.0702092
R42209 vss.t673 vss.n13994 0.0702092
R42210 vss.n539 vss.n537 0.0702092
R42211 vss.n537 vss.t653 0.0702092
R42212 vss.n662 vss.n660 0.0702092
R42213 vss.n661 vss.t1279 0.0702092
R42214 vss.n660 vss.t1279 0.0702092
R42215 vss.n675 vss.n661 0.0702092
R42216 vss.n13975 vss.n13974 0.0702092
R42217 vss.n13974 vss.t301 0.0702092
R42218 vss.n13977 vss.n562 0.0702092
R42219 vss.t303 vss.n562 0.0702092
R42220 vss.n13983 vss.n13982 0.0702092
R42221 vss.n13983 vss.t553 0.0702092
R42222 vss.n13980 vss.n13979 0.0702092
R42223 vss.n13979 vss.t553 0.0702092
R42224 vss.n13988 vss.n13987 0.0702092
R42225 vss.n13987 vss.t303 0.0702092
R42226 vss.n13973 vss.n557 0.0702092
R42227 vss.t301 vss.n13973 0.0702092
R42228 vss.n13971 vss.n574 0.0702092
R42229 vss.t952 vss.n13970 0.0702092
R42230 vss.n13971 vss.t952 0.0702092
R42231 vss.n13970 vss.n13969 0.0702092
R42232 vss.n13963 vss.n577 0.0702092
R42233 vss.n577 vss.t109 0.0702092
R42234 vss.n13961 vss.n13960 0.0702092
R42235 vss.n13960 vss.t767 0.0702092
R42236 vss.n772 vss.n771 0.0702092
R42237 vss.n771 vss.t769 0.0702092
R42238 vss.n770 vss.n591 0.0702092
R42239 vss.t769 vss.n770 0.0702092
R42240 vss.n13959 vss.n13958 0.0702092
R42241 vss.t767 vss.n13959 0.0702092
R42242 vss.n578 vss.n576 0.0702092
R42243 vss.n576 vss.t109 0.0702092
R42244 vss.n777 vss.n765 0.0702092
R42245 vss.t1148 vss.n763 0.0702092
R42246 vss.t1148 vss.n777 0.0702092
R42247 vss.n774 vss.n763 0.0702092
R42248 vss.n13244 vss.n13243 0.0702092
R42249 vss.n13243 vss.t527 0.0702092
R42250 vss.n781 vss.n760 0.0702092
R42251 vss.t529 vss.n760 0.0702092
R42252 vss.n787 vss.n786 0.0702092
R42253 vss.n787 vss.t125 0.0702092
R42254 vss.n784 vss.n783 0.0702092
R42255 vss.n783 vss.t125 0.0702092
R42256 vss.n792 vss.n791 0.0702092
R42257 vss.n791 vss.t529 0.0702092
R42258 vss.n13242 vss.n13241 0.0702092
R42259 vss.t527 vss.n13242 0.0702092
R42260 vss.n745 vss.n743 0.0702092
R42261 vss.n744 vss.t890 0.0702092
R42262 vss.n743 vss.t890 0.0702092
R42263 vss.n13246 vss.n744 0.0702092
R42264 vss.n1732 vss.n1731 0.0702092
R42265 vss.n1731 vss.t657 0.0702092
R42266 vss.n1735 vss.n1734 0.0702092
R42267 vss.t908 vss.n1735 0.0702092
R42268 vss.n1743 vss.n1742 0.0702092
R42269 vss.n1742 vss.t907 0.0702092
R42270 vss.n1741 vss.n1740 0.0702092
R42271 vss.t907 vss.n1741 0.0702092
R42272 vss.n1737 vss.n1736 0.0702092
R42273 vss.n1736 vss.t908 0.0702092
R42274 vss.n1730 vss.n1729 0.0702092
R42275 vss.t657 vss.n1730 0.0702092
R42276 vss.n1748 vss.n1709 0.0702092
R42277 vss.t545 vss.n1707 0.0702092
R42278 vss.t545 vss.n1748 0.0702092
R42279 vss.n1745 vss.n1707 0.0702092
R42280 vss.n1787 vss.n1786 0.0702092
R42281 vss.n1786 vss.t289 0.0702092
R42282 vss.n1789 vss.n1704 0.0702092
R42283 vss.t291 vss.n1704 0.0702092
R42284 vss.n1795 vss.n1794 0.0702092
R42285 vss.n1795 vss.t982 0.0702092
R42286 vss.n1792 vss.n1791 0.0702092
R42287 vss.n1791 vss.t982 0.0702092
R42288 vss.n1800 vss.n1799 0.0702092
R42289 vss.n1799 vss.t291 0.0702092
R42290 vss.n1785 vss.n1699 0.0702092
R42291 vss.t289 vss.n1785 0.0702092
R42292 vss.n1783 vss.n1761 0.0702092
R42293 vss.t1022 vss.n1782 0.0702092
R42294 vss.n1783 vss.t1022 0.0702092
R42295 vss.n1782 vss.n1781 0.0702092
R42296 vss.n1775 vss.n1763 0.0702092
R42297 vss.n1763 vss.t1159 0.0702092
R42298 vss.n1773 vss.n1772 0.0702092
R42299 vss.n1772 vss.t417 0.0702092
R42300 vss.n1814 vss.n1813 0.0702092
R42301 vss.n1813 vss.t419 0.0702092
R42302 vss.n1812 vss.n1811 0.0702092
R42303 vss.t419 vss.n1812 0.0702092
R42304 vss.n1771 vss.n1276 0.0702092
R42305 vss.t417 vss.n1771 0.0702092
R42306 vss.n1764 vss.n1762 0.0702092
R42307 vss.n1762 vss.t1159 0.0702092
R42308 vss.n1819 vss.n1266 0.0702092
R42309 vss.t1067 vss.n1264 0.0702092
R42310 vss.t1067 vss.n1819 0.0702092
R42311 vss.n1816 vss.n1264 0.0702092
R42312 vss.n1257 vss.n1239 0.0702092
R42313 vss.t279 vss.n1239 0.0702092
R42314 vss.n1259 vss.n1242 0.0702092
R42315 vss.t278 vss.n1242 0.0702092
R42316 vss.n1262 vss.n1261 0.0702092
R42317 vss.t281 vss.n1262 0.0702092
R42318 vss.n1823 vss.n1822 0.0702092
R42319 vss.n1822 vss.t281 0.0702092
R42320 vss.n1826 vss.n1825 0.0702092
R42321 vss.t278 vss.n1826 0.0702092
R42322 vss.n1828 vss.n1237 0.0702092
R42323 vss.n1828 vss.t279 0.0702092
R42324 vss.n1830 vss.n1234 0.0702092
R42325 vss.t997 vss.n1232 0.0702092
R42326 vss.t997 vss.n1830 0.0702092
R42327 vss.n1255 vss.n1232 0.0702092
R42328 vss.n1836 vss.n1835 0.0702092
R42329 vss.n1835 vss.t174 0.0702092
R42330 vss.n1839 vss.n1838 0.0702092
R42331 vss.t1455 vss.n1839 0.0702092
R42332 vss.n1847 vss.n1846 0.0702092
R42333 vss.n1846 vss.t1457 0.0702092
R42334 vss.n1845 vss.n1844 0.0702092
R42335 vss.t1457 vss.n1845 0.0702092
R42336 vss.n1841 vss.n1840 0.0702092
R42337 vss.n1840 vss.t1455 0.0702092
R42338 vss.n1834 vss.n1833 0.0702092
R42339 vss.t174 vss.n1834 0.0702092
R42340 vss.n1852 vss.n1213 0.0702092
R42341 vss.t315 vss.n1211 0.0702092
R42342 vss.t315 vss.n1852 0.0702092
R42343 vss.n1849 vss.n1211 0.0702092
R42344 vss.n1891 vss.n1890 0.0702092
R42345 vss.n1890 vss.t1276 0.0702092
R42346 vss.n1893 vss.n1208 0.0702092
R42347 vss.t1278 vss.n1208 0.0702092
R42348 vss.n1899 vss.n1898 0.0702092
R42349 vss.n1899 vss.t669 0.0702092
R42350 vss.n1896 vss.n1895 0.0702092
R42351 vss.n1895 vss.t669 0.0702092
R42352 vss.n1904 vss.n1903 0.0702092
R42353 vss.n1903 vss.t1278 0.0702092
R42354 vss.n1889 vss.n1203 0.0702092
R42355 vss.t1276 vss.n1889 0.0702092
R42356 vss.n1887 vss.n1865 0.0702092
R42357 vss.t847 vss.n1886 0.0702092
R42358 vss.n1887 vss.t847 0.0702092
R42359 vss.n1886 vss.n1885 0.0702092
R42360 vss.n1879 vss.n1867 0.0702092
R42361 vss.n1867 vss.t599 0.0702092
R42362 vss.n1877 vss.n1876 0.0702092
R42363 vss.n1876 vss.t150 0.0702092
R42364 vss.n1918 vss.n1917 0.0702092
R42365 vss.n1917 vss.t152 0.0702092
R42366 vss.n1916 vss.n1915 0.0702092
R42367 vss.t152 vss.n1916 0.0702092
R42368 vss.n1875 vss.n1158 0.0702092
R42369 vss.t150 vss.n1875 0.0702092
R42370 vss.n1868 vss.n1866 0.0702092
R42371 vss.n1866 vss.t599 0.0702092
R42372 vss.n1923 vss.n1148 0.0702092
R42373 vss.t1397 vss.n1146 0.0702092
R42374 vss.t1397 vss.n1923 0.0702092
R42375 vss.n1920 vss.n1146 0.0702092
R42376 vss.n1962 vss.n1961 0.0702092
R42377 vss.n1961 vss.t365 0.0702092
R42378 vss.n1964 vss.n1143 0.0702092
R42379 vss.t367 vss.n1143 0.0702092
R42380 vss.n1970 vss.n1969 0.0702092
R42381 vss.n1970 vss.t62 0.0702092
R42382 vss.n1967 vss.n1966 0.0702092
R42383 vss.n1966 vss.t62 0.0702092
R42384 vss.n1975 vss.n1974 0.0702092
R42385 vss.n1974 vss.t367 0.0702092
R42386 vss.n1960 vss.n1138 0.0702092
R42387 vss.t365 vss.n1960 0.0702092
R42388 vss.n1958 vss.n1936 0.0702092
R42389 vss.t886 vss.n1957 0.0702092
R42390 vss.n1958 vss.t886 0.0702092
R42391 vss.n1957 vss.n1956 0.0702092
R42392 vss.n1950 vss.n1938 0.0702092
R42393 vss.n1938 vss.t824 0.0702092
R42394 vss.n1948 vss.n1947 0.0702092
R42395 vss.n1947 vss.t114 0.0702092
R42396 vss.n13296 vss.n13295 0.0702092
R42397 vss.n13295 vss.t116 0.0702092
R42398 vss.n13294 vss.n13293 0.0702092
R42399 vss.t116 vss.n13294 0.0702092
R42400 vss.n1946 vss.n704 0.0702092
R42401 vss.t114 vss.n1946 0.0702092
R42402 vss.n1939 vss.n1937 0.0702092
R42403 vss.n1937 vss.t824 0.0702092
R42404 vss.n692 vss.n690 0.0702092
R42405 vss.n691 vss.t1412 0.0702092
R42406 vss.n690 vss.t1412 0.0702092
R42407 vss.n13298 vss.n691 0.0702092
R42408 vss.n13269 vss.n13268 0.0702092
R42409 vss.t876 vss.n13269 0.0702092
R42410 vss.n13274 vss.n13273 0.0702092
R42411 vss.n13273 vss.t780 0.0702092
R42412 vss.n13276 vss.n713 0.0702092
R42413 vss.t782 vss.n713 0.0702092
R42414 vss.n13282 vss.n13281 0.0702092
R42415 vss.n13282 vss.t645 0.0702092
R42416 vss.n13279 vss.n13278 0.0702092
R42417 vss.n13278 vss.t645 0.0702092
R42418 vss.n13287 vss.n13286 0.0702092
R42419 vss.n13286 vss.t782 0.0702092
R42420 vss.n13272 vss.n708 0.0702092
R42421 vss.t780 vss.n13272 0.0702092
R42422 vss.n13270 vss.n727 0.0702092
R42423 vss.n13270 vss.t876 0.0702092
R42424 vss.n13179 vss.n13178 0.0702092
R42425 vss.t1495 vss.n13179 0.0702092
R42426 vss.n13184 vss.n13183 0.0702092
R42427 vss.n13183 vss.t348 0.0702092
R42428 vss.n13186 vss.n13165 0.0702092
R42429 vss.t350 vss.n13165 0.0702092
R42430 vss.n13192 vss.n13191 0.0702092
R42431 vss.n13191 vss.t1097 0.0702092
R42432 vss.n13180 vss.n13176 0.0702092
R42433 vss.n13180 vss.t1495 0.0702092
R42434 vss.n13182 vss.n13160 0.0702092
R42435 vss.t348 vss.n13182 0.0702092
R42436 vss.n13198 vss.n13197 0.0702092
R42437 vss.n13197 vss.t350 0.0702092
R42438 vss.n13189 vss.n13188 0.0702092
R42439 vss.n13189 vss.t1097 0.0702092
R42440 vss.n1126 vss.n1125 0.0702092
R42441 vss.n1126 vss.t1299 0.0702092
R42442 vss.t578 vss.n1115 0.0702092
R42443 vss.n1119 vss.t323 0.0702092
R42444 vss.t325 vss.n1132 0.0702092
R42445 vss.n1128 vss.t1299 0.0702092
R42446 vss.n1134 vss.n1133 0.0702092
R42447 vss.n1133 vss.t325 0.0702092
R42448 vss.n1118 vss.n1096 0.0702092
R42449 vss.t323 vss.n1118 0.0702092
R42450 vss.n1116 vss.n1112 0.0702092
R42451 vss.n1116 vss.t578 0.0702092
R42452 vss.n1115 vss.n1114 0.0702092
R42453 vss.n1120 vss.n1119 0.0702092
R42454 vss.n1132 vss.n1131 0.0702092
R42455 vss.n1129 vss.n1128 0.0702092
R42456 vss.n1190 vss.n1189 0.0702092
R42457 vss.n1190 vss.t1146 0.0702092
R42458 vss.t13 vss.n1179 0.0702092
R42459 vss.n1183 vss.t542 0.0702092
R42460 vss.t544 vss.n1196 0.0702092
R42461 vss.n1192 vss.t1146 0.0702092
R42462 vss.n1198 vss.n1197 0.0702092
R42463 vss.n1197 vss.t544 0.0702092
R42464 vss.n1182 vss.n1160 0.0702092
R42465 vss.t542 vss.n1182 0.0702092
R42466 vss.n1180 vss.n1176 0.0702092
R42467 vss.n1180 vss.t13 0.0702092
R42468 vss.n1179 vss.n1178 0.0702092
R42469 vss.n1184 vss.n1183 0.0702092
R42470 vss.n1196 vss.n1195 0.0702092
R42471 vss.n1193 vss.n1192 0.0702092
R42472 vss.n1389 vss.n1388 0.0702092
R42473 vss.n1389 vss.t549 0.0702092
R42474 vss.t615 vss.n1378 0.0702092
R42475 vss.n1382 vss.t1407 0.0702092
R42476 vss.t1406 vss.n1395 0.0702092
R42477 vss.n1391 vss.t549 0.0702092
R42478 vss.n1397 vss.n1396 0.0702092
R42479 vss.n1396 vss.t1406 0.0702092
R42480 vss.n1381 vss.n1359 0.0702092
R42481 vss.t1407 vss.n1381 0.0702092
R42482 vss.n1379 vss.n1375 0.0702092
R42483 vss.n1379 vss.t615 0.0702092
R42484 vss.n1378 vss.n1377 0.0702092
R42485 vss.n1383 vss.n1382 0.0702092
R42486 vss.n1395 vss.n1394 0.0702092
R42487 vss.n1392 vss.n1391 0.0702092
R42488 vss.n1684 vss.n1683 0.0702092
R42489 vss.n1684 vss.t1270 0.0702092
R42490 vss.t1360 vss.n1673 0.0702092
R42491 vss.n1677 vss.t1531 0.0702092
R42492 vss.t1533 vss.n1690 0.0702092
R42493 vss.n1686 vss.t1270 0.0702092
R42494 vss.n1692 vss.n1691 0.0702092
R42495 vss.n1691 vss.t1533 0.0702092
R42496 vss.n1676 vss.n1654 0.0702092
R42497 vss.t1531 vss.n1676 0.0702092
R42498 vss.n1674 vss.n1670 0.0702092
R42499 vss.n1674 vss.t1360 0.0702092
R42500 vss.n1673 vss.n1672 0.0702092
R42501 vss.n1678 vss.n1677 0.0702092
R42502 vss.n1690 vss.n1689 0.0702092
R42503 vss.n1687 vss.n1686 0.0702092
R42504 vss.n13225 vss.n13224 0.0702092
R42505 vss.n13225 vss.t1177 0.0702092
R42506 vss.t506 vss.n13214 0.0702092
R42507 vss.n13218 vss.t1174 0.0702092
R42508 vss.t1176 vss.n13231 0.0702092
R42509 vss.n13227 vss.t1177 0.0702092
R42510 vss.n13233 vss.n13232 0.0702092
R42511 vss.n13232 vss.t1176 0.0702092
R42512 vss.n13217 vss.n795 0.0702092
R42513 vss.t1174 vss.n13217 0.0702092
R42514 vss.n13215 vss.n811 0.0702092
R42515 vss.n13215 vss.t506 0.0702092
R42516 vss.n13214 vss.n13213 0.0702092
R42517 vss.n13219 vss.n13218 0.0702092
R42518 vss.n13231 vss.n13230 0.0702092
R42519 vss.n13228 vss.n13227 0.0702092
R42520 vss.n610 vss.n609 0.0702092
R42521 vss.n610 vss.t222 0.0702092
R42522 vss.n818 vss.t17 0.0702092
R42523 vss.n827 vss.t358 0.0702092
R42524 vss.t360 vss.n13949 0.0702092
R42525 vss.n13945 vss.t222 0.0702092
R42526 vss.n13951 vss.n13950 0.0702092
R42527 vss.n13950 vss.t360 0.0702092
R42528 vss.n826 vss.n596 0.0702092
R42529 vss.t358 vss.n826 0.0702092
R42530 vss.n819 vss.n817 0.0702092
R42531 vss.n817 vss.t17 0.0702092
R42532 vss.n830 vss.n818 0.0702092
R42533 vss.n828 vss.n827 0.0702092
R42534 vss.n13949 vss.n13948 0.0702092
R42535 vss.n13946 vss.n13945 0.0702092
R42536 vss.n860 vss.n859 0.0702092
R42537 vss.n860 vss.t552 0.0702092
R42538 vss.n835 vss.t395 0.0702092
R42539 vss.n868 vss.t762 0.0702092
R42540 vss.n866 vss.t761 0.0702092
R42541 vss.n862 vss.t552 0.0702092
R42542 vss.n857 vss.n856 0.0702092
R42543 vss.n856 vss.t761 0.0702092
R42544 vss.n854 vss.n853 0.0702092
R42545 vss.n854 vss.t762 0.0702092
R42546 vss.n836 vss.n834 0.0702092
R42547 vss.n834 vss.t395 0.0702092
R42548 vss.n871 vss.n835 0.0702092
R42549 vss.n869 vss.n868 0.0702092
R42550 vss.n866 vss.n865 0.0702092
R42551 vss.n863 vss.n862 0.0702092
R42552 vss.n904 vss.n903 0.0702092
R42553 vss.n904 vss.t344 0.0702092
R42554 vss.n876 vss.t504 0.0702092
R42555 vss.n912 vss.t935 0.0702092
R42556 vss.n910 vss.t937 0.0702092
R42557 vss.n906 vss.t344 0.0702092
R42558 vss.n901 vss.n900 0.0702092
R42559 vss.n900 vss.t937 0.0702092
R42560 vss.n898 vss.n897 0.0702092
R42561 vss.n898 vss.t935 0.0702092
R42562 vss.n877 vss.n875 0.0702092
R42563 vss.n875 vss.t504 0.0702092
R42564 vss.n915 vss.n876 0.0702092
R42565 vss.n913 vss.n912 0.0702092
R42566 vss.n910 vss.n909 0.0702092
R42567 vss.n907 vss.n906 0.0702092
R42568 vss.n1554 vss.n1553 0.0702092
R42569 vss.n1554 vss.t983 0.0702092
R42570 vss.t397 vss.n1543 0.0702092
R42571 vss.n1547 vss.t1429 0.0702092
R42572 vss.t1431 vss.n1561 0.0702092
R42573 vss.n1557 vss.t983 0.0702092
R42574 vss.n1563 vss.n1562 0.0702092
R42575 vss.n1562 vss.t1431 0.0702092
R42576 vss.n1546 vss.n1524 0.0702092
R42577 vss.t1429 vss.n1546 0.0702092
R42578 vss.n1544 vss.n1540 0.0702092
R42579 vss.n1544 vss.t397 0.0702092
R42580 vss.n1543 vss.n1542 0.0702092
R42581 vss.n1548 vss.n1547 0.0702092
R42582 vss.n1561 vss.n1560 0.0702092
R42583 vss.n1558 vss.n1557 0.0702092
R42584 vss.n1637 vss.n1636 0.0702092
R42585 vss.n1637 vss.t166 0.0702092
R42586 vss.t621 vss.n1626 0.0702092
R42587 vss.n1630 vss.t583 0.0702092
R42588 vss.t582 vss.n1643 0.0702092
R42589 vss.n1639 vss.t166 0.0702092
R42590 vss.n1645 vss.n1644 0.0702092
R42591 vss.n1644 vss.t582 0.0702092
R42592 vss.n1629 vss.n1607 0.0702092
R42593 vss.t583 vss.n1629 0.0702092
R42594 vss.n1627 vss.n1623 0.0702092
R42595 vss.n1627 vss.t621 0.0702092
R42596 vss.n1626 vss.n1625 0.0702092
R42597 vss.n1631 vss.n1630 0.0702092
R42598 vss.n1643 vss.n1642 0.0702092
R42599 vss.n1640 vss.n1639 0.0702092
R42600 vss.n1474 vss.n1473 0.0702092
R42601 vss.n1474 vss.t1266 0.0702092
R42602 vss.t498 vss.n1463 0.0702092
R42603 vss.n1467 vss.t171 0.0702092
R42604 vss.t173 vss.n1480 0.0702092
R42605 vss.n1476 vss.t1266 0.0702092
R42606 vss.n1482 vss.n1481 0.0702092
R42607 vss.n1481 vss.t173 0.0702092
R42608 vss.n1466 vss.n1444 0.0702092
R42609 vss.t171 vss.n1466 0.0702092
R42610 vss.n1464 vss.n1460 0.0702092
R42611 vss.n1464 vss.t498 0.0702092
R42612 vss.n1463 vss.n1462 0.0702092
R42613 vss.n1468 vss.n1467 0.0702092
R42614 vss.n1480 vss.n1479 0.0702092
R42615 vss.n1477 vss.n1476 0.0702092
R42616 vss.n1342 vss.n1341 0.0702092
R42617 vss.n1342 vss.t541 0.0702092
R42618 vss.t1083 vss.n1331 0.0702092
R42619 vss.n1335 vss.t764 0.0702092
R42620 vss.t766 vss.n1348 0.0702092
R42621 vss.n1344 vss.t541 0.0702092
R42622 vss.n1350 vss.n1349 0.0702092
R42623 vss.n1349 vss.t766 0.0702092
R42624 vss.n1334 vss.n1312 0.0702092
R42625 vss.t764 vss.n1334 0.0702092
R42626 vss.n1332 vss.n1328 0.0702092
R42627 vss.n1332 vss.t1083 0.0702092
R42628 vss.n1331 vss.n1330 0.0702092
R42629 vss.n1336 vss.n1335 0.0702092
R42630 vss.n1348 vss.n1347 0.0702092
R42631 vss.n1345 vss.n1344 0.0702092
R42632 vss.n1081 vss.n1080 0.0702092
R42633 vss.n1081 vss.t1007 0.0702092
R42634 vss.t1372 vss.n1070 0.0702092
R42635 vss.n1074 vss.t923 0.0702092
R42636 vss.t925 vss.n1087 0.0702092
R42637 vss.n1083 vss.t1007 0.0702092
R42638 vss.n1089 vss.n1088 0.0702092
R42639 vss.n1088 vss.t925 0.0702092
R42640 vss.n1073 vss.n1051 0.0702092
R42641 vss.t923 vss.n1073 0.0702092
R42642 vss.n1071 vss.n1067 0.0702092
R42643 vss.n1071 vss.t1372 0.0702092
R42644 vss.n1070 vss.n1069 0.0702092
R42645 vss.n1075 vss.n1074 0.0702092
R42646 vss.n1087 vss.n1086 0.0702092
R42647 vss.n1084 vss.n1083 0.0702092
R42648 vss.n2016 vss.n2015 0.0702092
R42649 vss.n2016 vss.t1210 0.0702092
R42650 vss.t1320 vss.n2005 0.0702092
R42651 vss.n2009 vss.t521 0.0702092
R42652 vss.t523 vss.n2022 0.0702092
R42653 vss.n2018 vss.t1210 0.0702092
R42654 vss.n2024 vss.n2023 0.0702092
R42655 vss.n2023 vss.t523 0.0702092
R42656 vss.n2008 vss.n1986 0.0702092
R42657 vss.t521 vss.n2008 0.0702092
R42658 vss.n2006 vss.n2002 0.0702092
R42659 vss.n2006 vss.t1320 0.0702092
R42660 vss.n2005 vss.n2004 0.0702092
R42661 vss.n2010 vss.n2009 0.0702092
R42662 vss.n2022 vss.n2021 0.0702092
R42663 vss.n2019 vss.n2018 0.0702092
R42664 vss.n9608 vss.n9603 0.0702092
R42665 vss.n9608 vss.t244 0.0702092
R42666 vss.n9619 vss.n9618 0.0702092
R42667 vss.t1016 vss.n9619 0.0702092
R42668 vss.n9626 vss.n9625 0.0702092
R42669 vss.n9625 vss.t1140 0.0702092
R42670 vss.n9610 vss.n9587 0.0702092
R42671 vss.t1139 vss.n9610 0.0702092
R42672 vss.n9607 vss.n9606 0.0702092
R42673 vss.t244 vss.n9607 0.0702092
R42674 vss.n9612 vss.n9611 0.0702092
R42675 vss.n9611 vss.t1139 0.0702092
R42676 vss.n9624 vss.n9623 0.0702092
R42677 vss.t1140 vss.n9624 0.0702092
R42678 vss.n9621 vss.n9620 0.0702092
R42679 vss.n9620 vss.t1016 0.0702092
R42680 vss.n8050 vss.n8049 0.0702092
R42681 vss.t94 vss.n8050 0.0702092
R42682 vss.n8047 vss.n8046 0.0702092
R42683 vss.n8046 vss.t1528 0.0702092
R42684 vss.n8031 vss.n8030 0.0702092
R42685 vss.n8030 vss.t1529 0.0702092
R42686 vss.n8034 vss.n8033 0.0702092
R42687 vss.n8034 vss.t635 0.0702092
R42688 vss.t94 vss.n8013 0.0702092
R42689 vss.t1528 vss.n8045 0.0702092
R42690 vss.n8040 vss.t1529 0.0702092
R42691 vss.n8036 vss.t635 0.0702092
R42692 vss.n8037 vss.n8036 0.0702092
R42693 vss.n8040 vss.n8039 0.0702092
R42694 vss.n8045 vss.n8044 0.0702092
R42695 vss.n8042 vss.n8013 0.0702092
R42696 vss.n9665 vss.n5975 0.0702092
R42697 vss.n5975 vss.t1121 0.0702092
R42698 vss.n9652 vss.n9651 0.0702092
R42699 vss.n9651 vss.t41 0.0702092
R42700 vss.n5993 vss.n5991 0.0702092
R42701 vss.t736 vss.n5991 0.0702092
R42702 vss.n9663 vss.n9662 0.0702092
R42703 vss.n9662 vss.t735 0.0702092
R42704 vss.n5976 vss.n5974 0.0702092
R42705 vss.n5974 vss.t1121 0.0702092
R42706 vss.n9661 vss.n9660 0.0702092
R42707 vss.t735 vss.n9661 0.0702092
R42708 vss.n9658 vss.n9657 0.0702092
R42709 vss.n9657 vss.t736 0.0702092
R42710 vss.n5996 vss.n5995 0.0702092
R42711 vss.n5996 vss.t41 0.0702092
R42712 vss.n8148 vss.n8124 0.0702092
R42713 vss.n8124 vss.t1219 0.0702092
R42714 vss.n8146 vss.n8145 0.0702092
R42715 vss.n8145 vss.t691 0.0702092
R42716 vss.n8143 vss.n8128 0.0702092
R42717 vss.n8143 vss.t689 0.0702092
R42718 vss.n8137 vss.n8136 0.0702092
R42719 vss.n8136 vss.t1005 0.0702092
R42720 vss.n5999 vss.t1219 0.0702092
R42721 vss.n9644 vss.t691 0.0702092
R42722 vss.t689 vss.n8142 0.0702092
R42723 vss.n8140 vss.t1005 0.0702092
R42724 vss.n8140 vss.n8139 0.0702092
R42725 vss.n8142 vss.n6003 0.0702092
R42726 vss.n9644 vss.n9643 0.0702092
R42727 vss.n8149 vss.n5999 0.0702092
R42728 vss.n8155 vss.n8154 0.0702092
R42729 vss.t1061 vss.n8155 0.0702092
R42730 vss.n8156 vss.t1061 0.0702092
R42731 vss.n8157 vss.n8156 0.0702092
R42732 vss.n9032 vss.n9031 0.0702092
R42733 vss.n9031 vss.t719 0.0702092
R42734 vss.n9021 vss.n9020 0.0702092
R42735 vss.n9020 vss.t585 0.0702092
R42736 vss.n7287 vss.n7285 0.0702092
R42737 vss.t720 vss.n7285 0.0702092
R42738 vss.n9030 vss.n9029 0.0702092
R42739 vss.t719 vss.n9030 0.0702092
R42740 vss.n9027 vss.n9026 0.0702092
R42741 vss.n9026 vss.t720 0.0702092
R42742 vss.n7290 vss.n7289 0.0702092
R42743 vss.n7290 vss.t585 0.0702092
R42744 vss.n9012 vss.n9011 0.0702092
R42745 vss.n9011 vss.t946 0.0702092
R42746 vss.n7297 vss.n7296 0.0702092
R42747 vss.n7297 vss.t946 0.0702092
R42748 vss.n8261 vss.n7294 0.0702092
R42749 vss.n8261 vss.t773 0.0702092
R42750 vss.n8277 vss.n8276 0.0702092
R42751 vss.n8276 vss.t772 0.0702092
R42752 vss.n8279 vss.n7901 0.0702092
R42753 vss.n7901 vss.t703 0.0702092
R42754 vss.n7902 vss.n7900 0.0702092
R42755 vss.n7900 vss.t703 0.0702092
R42756 vss.n8275 vss.n8274 0.0702092
R42757 vss.t772 vss.n8275 0.0702092
R42758 vss.n8272 vss.n8271 0.0702092
R42759 vss.n8271 vss.t773 0.0702092
R42760 vss.n8287 vss.n8286 0.0702092
R42761 vss.n8286 vss.t1054 0.0702092
R42762 vss.n8285 vss.n8284 0.0702092
R42763 vss.t1054 vss.n8285 0.0702092
R42764 vss.n8300 vss.n7879 0.0702092
R42765 vss.n7879 vss.t65 0.0702092
R42766 vss.n8298 vss.n8297 0.0702092
R42767 vss.n8297 vss.t809 0.0702092
R42768 vss.n8290 vss.n8289 0.0702092
R42769 vss.t811 vss.n8290 0.0702092
R42770 vss.n8292 vss.n8291 0.0702092
R42771 vss.n8291 vss.t811 0.0702092
R42772 vss.n8296 vss.n8295 0.0702092
R42773 vss.t809 vss.n8296 0.0702092
R42774 vss.n7880 vss.n7878 0.0702092
R42775 vss.n7878 vss.t65 0.0702092
R42776 vss.n8706 vss.n7868 0.0702092
R42777 vss.n7868 vss.t912 0.0702092
R42778 vss.n7869 vss.n7867 0.0702092
R42779 vss.n7867 vss.t912 0.0702092
R42780 vss.n8704 vss.n8703 0.0702092
R42781 vss.n8703 vss.t95 0.0702092
R42782 vss.n8696 vss.n8695 0.0702092
R42783 vss.t97 vss.n8696 0.0702092
R42784 vss.n8693 vss.n8692 0.0702092
R42785 vss.n8692 vss.t80 0.0702092
R42786 vss.n8691 vss.n8690 0.0702092
R42787 vss.t80 vss.n8691 0.0702092
R42788 vss.n8698 vss.n8697 0.0702092
R42789 vss.n8697 vss.t97 0.0702092
R42790 vss.n8702 vss.n8701 0.0702092
R42791 vss.t95 vss.n8702 0.0702092
R42792 vss.n8327 vss.n8326 0.0702092
R42793 vss.n8326 vss.t272 0.0702092
R42794 vss.n8324 vss.n8323 0.0702092
R42795 vss.n8324 vss.t272 0.0702092
R42796 vss.n8348 vss.n8347 0.0702092
R42797 vss.t1153 vss.n8348 0.0702092
R42798 vss.n8680 vss.n8333 0.0702092
R42799 vss.n8680 vss.t1228 0.0702092
R42800 vss.n8683 vss.n8682 0.0702092
R42801 vss.n8682 vss.t1227 0.0702092
R42802 vss.n8340 vss.n8339 0.0702092
R42803 vss.n8339 vss.t1227 0.0702092
R42804 vss.n8679 vss.n8678 0.0702092
R42805 vss.t1228 vss.n8679 0.0702092
R42806 vss.n8676 vss.n8675 0.0702092
R42807 vss.n8675 vss.t1153 0.0702092
R42808 vss.n8668 vss.n8667 0.0702092
R42809 vss.n8667 vss.t1032 0.0702092
R42810 vss.n8665 vss.n8664 0.0702092
R42811 vss.n8665 vss.t1032 0.0702092
R42812 vss.n8662 vss.n8661 0.0702092
R42813 vss.n8661 vss.t667 0.0702092
R42814 vss.n8659 vss.n8355 0.0702092
R42815 vss.n8659 vss.t666 0.0702092
R42816 vss.n8649 vss.n8648 0.0702092
R42817 vss.t1088 vss.n8649 0.0702092
R42818 vss.n8651 vss.n8650 0.0702092
R42819 vss.n8650 vss.t1088 0.0702092
R42820 vss.n8658 vss.n8657 0.0702092
R42821 vss.t666 vss.n8658 0.0702092
R42822 vss.n8655 vss.n8654 0.0702092
R42823 vss.n8654 vss.t667 0.0702092
R42824 vss.n8372 vss.n8371 0.0702092
R42825 vss.n8371 vss.t1223 0.0702092
R42826 vss.n8369 vss.n8368 0.0702092
R42827 vss.n8369 vss.t1223 0.0702092
R42828 vss.n8398 vss.n8397 0.0702092
R42829 vss.t865 vss.n8398 0.0702092
R42830 vss.n8637 vss.n8383 0.0702092
R42831 vss.n8637 vss.t606 0.0702092
R42832 vss.n8640 vss.n8639 0.0702092
R42833 vss.n8639 vss.t608 0.0702092
R42834 vss.n8390 vss.n8389 0.0702092
R42835 vss.n8389 vss.t608 0.0702092
R42836 vss.n8636 vss.n8635 0.0702092
R42837 vss.t606 vss.n8636 0.0702092
R42838 vss.n8633 vss.n8632 0.0702092
R42839 vss.n8632 vss.t865 0.0702092
R42840 vss.n8625 vss.n8624 0.0702092
R42841 vss.n8624 vss.t956 0.0702092
R42842 vss.n8621 vss.n8620 0.0702092
R42843 vss.n8621 vss.t956 0.0702092
R42844 vss.n8618 vss.n8617 0.0702092
R42845 vss.n8617 vss.t148 0.0702092
R42846 vss.n8615 vss.n8408 0.0702092
R42847 vss.n8615 vss.t147 0.0702092
R42848 vss.n8605 vss.n8604 0.0702092
R42849 vss.t82 vss.n8605 0.0702092
R42850 vss.n8607 vss.n8606 0.0702092
R42851 vss.n8606 vss.t82 0.0702092
R42852 vss.n8614 vss.n8613 0.0702092
R42853 vss.t147 vss.n8614 0.0702092
R42854 vss.n8611 vss.n8610 0.0702092
R42855 vss.n8610 vss.t148 0.0702092
R42856 vss.n8425 vss.n8424 0.0702092
R42857 vss.n8424 vss.t1115 0.0702092
R42858 vss.n8422 vss.n8421 0.0702092
R42859 vss.n8422 vss.t1115 0.0702092
R42860 vss.n8446 vss.n8445 0.0702092
R42861 vss.t595 vss.n8446 0.0702092
R42862 vss.n8593 vss.n8431 0.0702092
R42863 vss.n8593 vss.t98 0.0702092
R42864 vss.n8596 vss.n8595 0.0702092
R42865 vss.n8595 vss.t100 0.0702092
R42866 vss.n8438 vss.n8437 0.0702092
R42867 vss.n8437 vss.t100 0.0702092
R42868 vss.n8592 vss.n8591 0.0702092
R42869 vss.t98 vss.n8592 0.0702092
R42870 vss.n8589 vss.n8588 0.0702092
R42871 vss.n8588 vss.t595 0.0702092
R42872 vss.n8581 vss.n8580 0.0702092
R42873 vss.n8580 vss.t1030 0.0702092
R42874 vss.n8578 vss.n8577 0.0702092
R42875 vss.n8578 vss.t1030 0.0702092
R42876 vss.n8575 vss.n8574 0.0702092
R42877 vss.n8574 vss.t944 0.0702092
R42878 vss.n8572 vss.n8453 0.0702092
R42879 vss.n8572 vss.t943 0.0702092
R42880 vss.n8562 vss.n8561 0.0702092
R42881 vss.t686 vss.n8562 0.0702092
R42882 vss.n8564 vss.n8563 0.0702092
R42883 vss.n8563 vss.t686 0.0702092
R42884 vss.n8571 vss.n8570 0.0702092
R42885 vss.t943 vss.n8571 0.0702092
R42886 vss.n8568 vss.n8567 0.0702092
R42887 vss.n8567 vss.t944 0.0702092
R42888 vss.n8470 vss.n8469 0.0702092
R42889 vss.n8469 vss.t424 0.0702092
R42890 vss.n8467 vss.n8466 0.0702092
R42891 vss.n8467 vss.t424 0.0702092
R42892 vss.n8496 vss.n8495 0.0702092
R42893 vss.t178 vss.n8496 0.0702092
R42894 vss.n8550 vss.n8481 0.0702092
R42895 vss.n8550 vss.t792 0.0702092
R42896 vss.n8553 vss.n8552 0.0702092
R42897 vss.n8552 vss.t794 0.0702092
R42898 vss.n8488 vss.n8487 0.0702092
R42899 vss.n8487 vss.t794 0.0702092
R42900 vss.n8549 vss.n8548 0.0702092
R42901 vss.t792 vss.n8549 0.0702092
R42902 vss.n8546 vss.n8545 0.0702092
R42903 vss.n8545 vss.t178 0.0702092
R42904 vss.n8523 vss.n8522 0.0702092
R42905 vss.t292 vss.n8523 0.0702092
R42906 vss.n8520 vss.n8519 0.0702092
R42907 vss.n8519 vss.t1105 0.0702092
R42908 vss.n8517 vss.n8516 0.0702092
R42909 vss.n8517 vss.t1106 0.0702092
R42910 vss.n8534 vss.n8533 0.0702092
R42911 vss.n8534 vss.t1028 0.0702092
R42912 vss.n8524 vss.t292 0.0702092
R42913 vss.n8528 vss.t1105 0.0702092
R42914 vss.n8530 vss.t1106 0.0702092
R42915 vss.n8537 vss.t1028 0.0702092
R42916 vss.n8538 vss.n8537 0.0702092
R42917 vss.n8531 vss.n8530 0.0702092
R42918 vss.n8528 vss.n8527 0.0702092
R42919 vss.n8525 vss.n8524 0.0702092
R42920 vss.n9559 vss.n9558 0.0702092
R42921 vss.n9558 vss.t1300 0.0702092
R42922 vss.n9561 vss.n6062 0.0702092
R42923 vss.t1302 vss.n6062 0.0702092
R42924 vss.n9567 vss.n9566 0.0702092
R42925 vss.n9567 vss.t1291 0.0702092
R42926 vss.n9564 vss.n9563 0.0702092
R42927 vss.n9563 vss.t1291 0.0702092
R42928 vss.n9572 vss.n9571 0.0702092
R42929 vss.n9571 vss.t1302 0.0702092
R42930 vss.n9557 vss.n6057 0.0702092
R42931 vss.t1300 vss.n9557 0.0702092
R42932 vss.n9555 vss.n6075 0.0702092
R42933 vss.t1042 vss.n9554 0.0702092
R42934 vss.n9555 vss.t1042 0.0702092
R42935 vss.n9554 vss.n9553 0.0702092
R42936 vss.n9547 vss.n6078 0.0702092
R42937 vss.n6078 vss.t822 0.0702092
R42938 vss.n9545 vss.n9544 0.0702092
R42939 vss.n9544 vss.t903 0.0702092
R42940 vss.n7261 vss.n7260 0.0702092
R42941 vss.n7260 vss.t905 0.0702092
R42942 vss.n7259 vss.n6092 0.0702092
R42943 vss.t905 vss.n7259 0.0702092
R42944 vss.n9543 vss.n9542 0.0702092
R42945 vss.t903 vss.n9543 0.0702092
R42946 vss.n6079 vss.n6077 0.0702092
R42947 vss.n6077 vss.t822 0.0702092
R42948 vss.n7250 vss.n7248 0.0702092
R42949 vss.n7249 vss.t839 0.0702092
R42950 vss.n7248 vss.t839 0.0702092
R42951 vss.n7263 vss.n7249 0.0702092
R42952 vss.n9524 vss.n9523 0.0702092
R42953 vss.n9523 vss.t258 0.0702092
R42954 vss.n9526 vss.n6102 0.0702092
R42955 vss.t260 vss.n6102 0.0702092
R42956 vss.n9532 vss.n9531 0.0702092
R42957 vss.n9532 vss.t892 0.0702092
R42958 vss.n9529 vss.n9528 0.0702092
R42959 vss.n9528 vss.t892 0.0702092
R42960 vss.n9537 vss.n9536 0.0702092
R42961 vss.n9536 vss.t260 0.0702092
R42962 vss.n9522 vss.n6097 0.0702092
R42963 vss.t258 vss.n9522 0.0702092
R42964 vss.n9520 vss.n6114 0.0702092
R42965 vss.t989 vss.n9519 0.0702092
R42966 vss.n9520 vss.t989 0.0702092
R42967 vss.n9519 vss.n9518 0.0702092
R42968 vss.n9512 vss.n6117 0.0702092
R42969 vss.n6117 vss.t105 0.0702092
R42970 vss.n9510 vss.n9509 0.0702092
R42971 vss.n9509 vss.t453 0.0702092
R42972 vss.n7242 vss.n7241 0.0702092
R42973 vss.n7241 vss.t452 0.0702092
R42974 vss.n7240 vss.n6131 0.0702092
R42975 vss.t452 vss.n7240 0.0702092
R42976 vss.n9508 vss.n9507 0.0702092
R42977 vss.t453 vss.n9508 0.0702092
R42978 vss.n6118 vss.n6116 0.0702092
R42979 vss.n6116 vss.t105 0.0702092
R42980 vss.n6577 vss.n6575 0.0702092
R42981 vss.n6576 vss.t910 0.0702092
R42982 vss.n6575 vss.t910 0.0702092
R42983 vss.n7244 vss.n6576 0.0702092
R42984 vss.n6759 vss.n6758 0.0702092
R42985 vss.t532 vss.n6759 0.0702092
R42986 vss.n7230 vss.n7229 0.0702092
R42987 vss.n7229 vss.t531 0.0702092
R42988 vss.n7232 vss.n6582 0.0702092
R42989 vss.n6582 vss.t1516 0.0702092
R42990 vss.n6583 vss.n6581 0.0702092
R42991 vss.n6581 vss.t1516 0.0702092
R42992 vss.n7228 vss.n7227 0.0702092
R42993 vss.t531 vss.n7228 0.0702092
R42994 vss.n6760 vss.n6595 0.0702092
R42995 vss.n6760 vss.t532 0.0702092
R42996 vss.n6762 vss.n6750 0.0702092
R42997 vss.t43 vss.n6748 0.0702092
R42998 vss.t43 vss.n6762 0.0702092
R42999 vss.n6756 vss.n6748 0.0702092
R43000 vss.n6768 vss.n6767 0.0702092
R43001 vss.n6767 vss.t446 0.0702092
R43002 vss.n6771 vss.n6770 0.0702092
R43003 vss.t246 vss.n6771 0.0702092
R43004 vss.n6779 vss.n6778 0.0702092
R43005 vss.n6778 vss.t245 0.0702092
R43006 vss.n6777 vss.n6776 0.0702092
R43007 vss.t245 vss.n6777 0.0702092
R43008 vss.n6773 vss.n6772 0.0702092
R43009 vss.n6772 vss.t246 0.0702092
R43010 vss.n6766 vss.n6765 0.0702092
R43011 vss.t446 vss.n6766 0.0702092
R43012 vss.n6784 vss.n6729 0.0702092
R43013 vss.t248 vss.n6727 0.0702092
R43014 vss.t248 vss.n6784 0.0702092
R43015 vss.n6781 vss.n6727 0.0702092
R43016 vss.n7069 vss.n7068 0.0702092
R43017 vss.n7068 vss.t327 0.0702092
R43018 vss.n7071 vss.n6724 0.0702092
R43019 vss.t326 vss.n6724 0.0702092
R43020 vss.n7077 vss.n7076 0.0702092
R43021 vss.n7077 vss.t646 0.0702092
R43022 vss.n7074 vss.n7073 0.0702092
R43023 vss.n7073 vss.t646 0.0702092
R43024 vss.n7082 vss.n7081 0.0702092
R43025 vss.n7081 vss.t326 0.0702092
R43026 vss.n7067 vss.n6719 0.0702092
R43027 vss.t327 vss.n7067 0.0702092
R43028 vss.n7065 vss.n6797 0.0702092
R43029 vss.t995 vss.n7064 0.0702092
R43030 vss.n7065 vss.t995 0.0702092
R43031 vss.n7064 vss.n7063 0.0702092
R43032 vss.n7057 vss.n6799 0.0702092
R43033 vss.n6799 vss.t1157 0.0702092
R43034 vss.n7055 vss.n7054 0.0702092
R43035 vss.n7054 vss.t555 0.0702092
R43036 vss.n6821 vss.n6815 0.0702092
R43037 vss.t554 vss.n6815 0.0702092
R43038 vss.n7048 vss.n7047 0.0702092
R43039 vss.n7047 vss.t554 0.0702092
R43040 vss.n7053 vss.n7052 0.0702092
R43041 vss.t555 vss.n7053 0.0702092
R43042 vss.n6800 vss.n6798 0.0702092
R43043 vss.n6798 vss.t1157 0.0702092
R43044 vss.n6826 vss.n6819 0.0702092
R43045 vss.t557 vss.n6818 0.0702092
R43046 vss.t557 vss.n6826 0.0702092
R43047 vss.n6823 vss.n6818 0.0702092
R43048 vss.n6900 vss.n6899 0.0702092
R43049 vss.t670 vss.n6900 0.0702092
R43050 vss.n7039 vss.n7038 0.0702092
R43051 vss.n7038 vss.t672 0.0702092
R43052 vss.n7041 vss.n6828 0.0702092
R43053 vss.n6828 vss.t33 0.0702092
R43054 vss.n6829 vss.n6827 0.0702092
R43055 vss.n6827 vss.t33 0.0702092
R43056 vss.n7037 vss.n7036 0.0702092
R43057 vss.t672 vss.n7037 0.0702092
R43058 vss.n6902 vss.n6901 0.0702092
R43059 vss.n6901 vss.t670 0.0702092
R43060 vss.n6895 vss.n6894 0.0702092
R43061 vss.n6896 vss.t918 0.0702092
R43062 vss.t918 vss.n6895 0.0702092
R43063 vss.n6897 vss.n6896 0.0702092
R43064 vss.n6889 vss.n6850 0.0702092
R43065 vss.n6850 vss.t797 0.0702092
R43066 vss.n6887 vss.n6886 0.0702092
R43067 vss.n6886 vss.t140 0.0702092
R43068 vss.n6872 vss.n6866 0.0702092
R43069 vss.t139 vss.n6866 0.0702092
R43070 vss.n6882 vss.n6881 0.0702092
R43071 vss.n6881 vss.t139 0.0702092
R43072 vss.n6885 vss.n6884 0.0702092
R43073 vss.t140 vss.n6885 0.0702092
R43074 vss.n6851 vss.n6849 0.0702092
R43075 vss.n6849 vss.t797 0.0702092
R43076 vss.n6877 vss.n6870 0.0702092
R43077 vss.t343 vss.n6869 0.0702092
R43078 vss.t343 vss.n6877 0.0702092
R43079 vss.n6874 vss.n6869 0.0702092
R43080 vss.n9232 vss.n9231 0.0702092
R43081 vss.n9231 vss.t255 0.0702092
R43082 vss.n9234 vss.n6496 0.0702092
R43083 vss.t254 vss.n6496 0.0702092
R43084 vss.n9240 vss.n9239 0.0702092
R43085 vss.n9240 vss.t1458 0.0702092
R43086 vss.n9237 vss.n9236 0.0702092
R43087 vss.n9236 vss.t1458 0.0702092
R43088 vss.n9245 vss.n9244 0.0702092
R43089 vss.n9244 vss.t254 0.0702092
R43090 vss.n9230 vss.n6491 0.0702092
R43091 vss.t255 vss.n9230 0.0702092
R43092 vss.n9228 vss.n6508 0.0702092
R43093 vss.t57 vss.n9227 0.0702092
R43094 vss.n9228 vss.t57 0.0702092
R43095 vss.n9227 vss.n9226 0.0702092
R43096 vss.n9220 vss.n6510 0.0702092
R43097 vss.n6510 vss.t589 0.0702092
R43098 vss.n9218 vss.n9217 0.0702092
R43099 vss.n9217 vss.t1410 0.0702092
R43100 vss.n6562 vss.n6526 0.0702092
R43101 vss.t1409 vss.n6526 0.0702092
R43102 vss.n9211 vss.n9210 0.0702092
R43103 vss.n9210 vss.t1409 0.0702092
R43104 vss.n9216 vss.n9215 0.0702092
R43105 vss.t1410 vss.n9216 0.0702092
R43106 vss.n6511 vss.n6509 0.0702092
R43107 vss.n6509 vss.t589 0.0702092
R43108 vss.n6560 vss.n6557 0.0702092
R43109 vss.n6559 vss.t285 0.0702092
R43110 vss.n6557 vss.t285 0.0702092
R43111 vss.n6564 vss.n6559 0.0702092
R43112 vss.n9077 vss.n9076 0.0702092
R43113 vss.t1204 vss.n9077 0.0702092
R43114 vss.n9202 vss.n9201 0.0702092
R43115 vss.n9201 vss.t1203 0.0702092
R43116 vss.n9204 vss.n6529 0.0702092
R43117 vss.n6529 vss.t1138 0.0702092
R43118 vss.n6530 vss.n6528 0.0702092
R43119 vss.n6528 vss.t1138 0.0702092
R43120 vss.n9200 vss.n9199 0.0702092
R43121 vss.t1203 vss.n9200 0.0702092
R43122 vss.n9078 vss.n6542 0.0702092
R43123 vss.n9078 vss.t1204 0.0702092
R43124 vss.n9080 vss.n9068 0.0702092
R43125 vss.t1034 vss.n9066 0.0702092
R43126 vss.t1034 vss.n9080 0.0702092
R43127 vss.n9074 vss.n9066 0.0702092
R43128 vss.n9085 vss.n9084 0.0702092
R43129 vss.t859 vss.n9085 0.0702092
R43130 vss.n9090 vss.n9089 0.0702092
R43131 vss.n9089 vss.t460 0.0702092
R43132 vss.n9092 vss.n6553 0.0702092
R43133 vss.t459 vss.n6553 0.0702092
R43134 vss.n9143 vss.n9142 0.0702092
R43135 vss.n9142 vss.t459 0.0702092
R43136 vss.n9088 vss.n6548 0.0702092
R43137 vss.t460 vss.n9088 0.0702092
R43138 vss.n9086 vss.n9064 0.0702092
R43139 vss.n9086 vss.t859 0.0702092
R43140 vss.n9097 vss.n9053 0.0702092
R43141 vss.t351 vss.n9052 0.0702092
R43142 vss.t351 vss.n9097 0.0702092
R43143 vss.n9094 vss.n9052 0.0702092
R43144 vss.n9123 vss.n9122 0.0702092
R43145 vss.n9122 vss.t888 0.0702092
R43146 vss.n9126 vss.n9125 0.0702092
R43147 vss.t1436 vss.n9126 0.0702092
R43148 vss.n9134 vss.n9133 0.0702092
R43149 vss.n9133 vss.t1435 0.0702092
R43150 vss.n9136 vss.n9099 0.0702092
R43151 vss.n9099 vss.t1179 0.0702092
R43152 vss.n9100 vss.n9098 0.0702092
R43153 vss.n9098 vss.t1179 0.0702092
R43154 vss.n9132 vss.n9131 0.0702092
R43155 vss.t1435 vss.n9132 0.0702092
R43156 vss.n9128 vss.n9127 0.0702092
R43157 vss.n9127 vss.t1436 0.0702092
R43158 vss.n9121 vss.n9120 0.0702092
R43159 vss.t888 vss.n9121 0.0702092
R43160 vss.n6187 vss.n6185 0.0702092
R43161 vss.n6185 vss.t1092 0.0702092
R43162 vss.n6206 vss.t1079 0.0702092
R43163 vss.t1090 vss.n6210 0.0702092
R43164 vss.n9376 vss.t1089 0.0702092
R43165 vss.n6186 vss.t1092 0.0702092
R43166 vss.n9371 vss.n9370 0.0702092
R43167 vss.n9371 vss.t1089 0.0702092
R43168 vss.n6212 vss.n6211 0.0702092
R43169 vss.n6211 vss.t1090 0.0702092
R43170 vss.n6205 vss.n6204 0.0702092
R43171 vss.t1079 vss.n6205 0.0702092
R43172 vss.n6207 vss.n6206 0.0702092
R43173 vss.n6210 vss.n6209 0.0702092
R43174 vss.n9377 vss.n9376 0.0702092
R43175 vss.n9379 vss.n6186 0.0702092
R43176 vss.n9182 vss.n9181 0.0702092
R43177 vss.n9182 vss.t899 0.0702092
R43178 vss.t472 vss.n9171 0.0702092
R43179 vss.n9175 vss.t897 0.0702092
R43180 vss.t896 vss.n9188 0.0702092
R43181 vss.n9184 vss.t899 0.0702092
R43182 vss.n9190 vss.n9189 0.0702092
R43183 vss.n9189 vss.t896 0.0702092
R43184 vss.n9174 vss.n9151 0.0702092
R43185 vss.t897 vss.n9174 0.0702092
R43186 vss.n9172 vss.n9167 0.0702092
R43187 vss.n9172 vss.t472 0.0702092
R43188 vss.n9171 vss.n9170 0.0702092
R43189 vss.n9176 vss.n9175 0.0702092
R43190 vss.n9188 vss.n9187 0.0702092
R43191 vss.n9185 vss.n9184 0.0702092
R43192 vss.n6479 vss.n6478 0.0702092
R43193 vss.n6479 vss.t771 0.0702092
R43194 vss.t1334 vss.n6468 0.0702092
R43195 vss.n6472 vss.t1465 0.0702092
R43196 vss.t1464 vss.n6485 0.0702092
R43197 vss.n6481 vss.t771 0.0702092
R43198 vss.n6487 vss.n6486 0.0702092
R43199 vss.n6486 vss.t1464 0.0702092
R43200 vss.n6471 vss.n6448 0.0702092
R43201 vss.t1465 vss.n6471 0.0702092
R43202 vss.n6469 vss.n6464 0.0702092
R43203 vss.n6469 vss.t1334 0.0702092
R43204 vss.n6468 vss.n6467 0.0702092
R43205 vss.n6473 vss.n6472 0.0702092
R43206 vss.n6485 vss.n6484 0.0702092
R43207 vss.n6482 vss.n6481 0.0702092
R43208 vss.n7019 vss.n7018 0.0702092
R43209 vss.n7019 vss.t87 0.0702092
R43210 vss.t1314 vss.n7008 0.0702092
R43211 vss.n7012 vss.t333 0.0702092
R43212 vss.t332 vss.n7025 0.0702092
R43213 vss.n7021 vss.t87 0.0702092
R43214 vss.n7027 vss.n7026 0.0702092
R43215 vss.n7026 vss.t332 0.0702092
R43216 vss.n7011 vss.n6988 0.0702092
R43217 vss.t333 vss.n7011 0.0702092
R43218 vss.n7009 vss.n7004 0.0702092
R43219 vss.n7009 vss.t1314 0.0702092
R43220 vss.n7008 vss.n7007 0.0702092
R43221 vss.n7013 vss.n7012 0.0702092
R43222 vss.n7025 vss.n7024 0.0702092
R43223 vss.n7022 vss.n7021 0.0702092
R43224 vss.n6705 vss.n6704 0.0702092
R43225 vss.n6705 vss.t1008 0.0702092
R43226 vss.t1370 vss.n6694 0.0702092
R43227 vss.n6698 vss.t985 0.0702092
R43228 vss.t987 vss.n6711 0.0702092
R43229 vss.n6707 vss.t1008 0.0702092
R43230 vss.n6713 vss.n6712 0.0702092
R43231 vss.n6712 vss.t987 0.0702092
R43232 vss.n6697 vss.n6674 0.0702092
R43233 vss.t985 vss.n6697 0.0702092
R43234 vss.n6695 vss.n6690 0.0702092
R43235 vss.n6695 vss.t1370 0.0702092
R43236 vss.n6694 vss.n6693 0.0702092
R43237 vss.n6699 vss.n6698 0.0702092
R43238 vss.n6711 vss.n6710 0.0702092
R43239 vss.n6708 vss.n6707 0.0702092
R43240 vss.n7210 vss.n7209 0.0702092
R43241 vss.n7210 vss.t314 0.0702092
R43242 vss.t213 vss.n7199 0.0702092
R43243 vss.n7203 vss.t85 0.0702092
R43244 vss.t84 vss.n7216 0.0702092
R43245 vss.n7212 vss.t314 0.0702092
R43246 vss.n7218 vss.n7217 0.0702092
R43247 vss.n7217 vss.t84 0.0702092
R43248 vss.n7202 vss.n7179 0.0702092
R43249 vss.t85 vss.n7202 0.0702092
R43250 vss.n7200 vss.n7195 0.0702092
R43251 vss.n7200 vss.t213 0.0702092
R43252 vss.n7199 vss.n7198 0.0702092
R43253 vss.n7204 vss.n7203 0.0702092
R43254 vss.n7216 vss.n7215 0.0702092
R43255 vss.n7213 vss.n7212 0.0702092
R43256 vss.n6167 vss.n6166 0.0702092
R43257 vss.n6167 vss.t1104 0.0702092
R43258 vss.t1340 vss.n6156 0.0702092
R43259 vss.n6160 vss.t1293 0.0702092
R43260 vss.t1292 vss.n9498 0.0702092
R43261 vss.n9494 vss.t1104 0.0702092
R43262 vss.n9500 vss.n9499 0.0702092
R43263 vss.n9499 vss.t1292 0.0702092
R43264 vss.n6159 vss.n6136 0.0702092
R43265 vss.t1293 vss.n6159 0.0702092
R43266 vss.n6157 vss.n6152 0.0702092
R43267 vss.n6157 vss.t1340 0.0702092
R43268 vss.n6156 vss.n6155 0.0702092
R43269 vss.n6161 vss.n6160 0.0702092
R43270 vss.n9498 vss.n9497 0.0702092
R43271 vss.n9495 vss.n9494 0.0702092
R43272 vss.n9447 vss.n9445 0.0702092
R43273 vss.n9445 vss.t1254 0.0702092
R43274 vss.n9466 vss.t510 0.0702092
R43275 vss.t230 vss.n9470 0.0702092
R43276 vss.n9480 vss.t229 0.0702092
R43277 vss.n9446 vss.t1254 0.0702092
R43278 vss.n9475 vss.n9474 0.0702092
R43279 vss.n9475 vss.t229 0.0702092
R43280 vss.n9471 vss.n9454 0.0702092
R43281 vss.n9471 vss.t230 0.0702092
R43282 vss.n9465 vss.n9464 0.0702092
R43283 vss.t510 vss.n9465 0.0702092
R43284 vss.n9467 vss.n9466 0.0702092
R43285 vss.n9470 vss.n9469 0.0702092
R43286 vss.n9481 vss.n9480 0.0702092
R43287 vss.n9483 vss.n9446 0.0702092
R43288 vss.n6040 vss.n6039 0.0702092
R43289 vss.n6040 vss.t1114 0.0702092
R43290 vss.t211 vss.n6029 0.0702092
R43291 vss.n6033 vss.t731 0.0702092
R43292 vss.t733 vss.n6047 0.0702092
R43293 vss.n6043 vss.t1114 0.0702092
R43294 vss.n6049 vss.n6048 0.0702092
R43295 vss.n6048 vss.t733 0.0702092
R43296 vss.n6032 vss.n6009 0.0702092
R43297 vss.t731 vss.n6032 0.0702092
R43298 vss.n6030 vss.n6025 0.0702092
R43299 vss.n6030 vss.t211 0.0702092
R43300 vss.n6029 vss.n6028 0.0702092
R43301 vss.n6034 vss.n6033 0.0702092
R43302 vss.n6047 vss.n6046 0.0702092
R43303 vss.n6044 vss.n6043 0.0702092
R43304 vss.n9402 vss.n9400 0.0702092
R43305 vss.n9400 vss.t153 0.0702092
R43306 vss.n9421 vss.t1487 0.0702092
R43307 vss.t941 vss.n9425 0.0702092
R43308 vss.n9438 vss.t940 0.0702092
R43309 vss.n9401 vss.t153 0.0702092
R43310 vss.n9433 vss.n9432 0.0702092
R43311 vss.n9433 vss.t940 0.0702092
R43312 vss.n9427 vss.n9426 0.0702092
R43313 vss.n9426 vss.t941 0.0702092
R43314 vss.n9420 vss.n9419 0.0702092
R43315 vss.t1487 vss.n9420 0.0702092
R43316 vss.n9422 vss.n9421 0.0702092
R43317 vss.n9425 vss.n9424 0.0702092
R43318 vss.n9439 vss.n9438 0.0702092
R43319 vss.n9441 vss.n9401 0.0702092
R43320 vss.n7159 vss.n7158 0.0702092
R43321 vss.n7159 vss.t1283 0.0702092
R43322 vss.t1501 vss.n7148 0.0702092
R43323 vss.n7152 vss.t1281 0.0702092
R43324 vss.t1280 vss.n7165 0.0702092
R43325 vss.n7161 vss.t1283 0.0702092
R43326 vss.n7167 vss.n7166 0.0702092
R43327 vss.n7166 vss.t1280 0.0702092
R43328 vss.n7151 vss.n7128 0.0702092
R43329 vss.t1281 vss.n7151 0.0702092
R43330 vss.n7149 vss.n7144 0.0702092
R43331 vss.n7149 vss.t1501 0.0702092
R43332 vss.n7148 vss.n7147 0.0702092
R43333 vss.n7153 vss.n7152 0.0702092
R43334 vss.n7165 vss.n7164 0.0702092
R43335 vss.n7162 vss.n7161 0.0702092
R43336 vss.n6661 vss.n6660 0.0702092
R43337 vss.n6661 vss.t1120 0.0702092
R43338 vss.t1330 vss.n6650 0.0702092
R43339 vss.n6654 vss.t1118 0.0702092
R43340 vss.t1117 vss.n6667 0.0702092
R43341 vss.n6663 vss.t1120 0.0702092
R43342 vss.n6669 vss.n6668 0.0702092
R43343 vss.n6668 vss.t1117 0.0702092
R43344 vss.n6653 vss.n6630 0.0702092
R43345 vss.t1118 vss.n6653 0.0702092
R43346 vss.n6651 vss.n6646 0.0702092
R43347 vss.n6651 vss.t1330 0.0702092
R43348 vss.n6650 vss.n6649 0.0702092
R43349 vss.n6655 vss.n6654 0.0702092
R43350 vss.n6667 vss.n6666 0.0702092
R43351 vss.n6664 vss.n6663 0.0702092
R43352 vss.n6970 vss.n6969 0.0702092
R43353 vss.n6970 vss.t550 0.0702092
R43354 vss.t482 vss.n6959 0.0702092
R43355 vss.n6963 vss.t547 0.0702092
R43356 vss.t546 vss.n6976 0.0702092
R43357 vss.n6972 vss.t550 0.0702092
R43358 vss.n6978 vss.n6977 0.0702092
R43359 vss.n6977 vss.t546 0.0702092
R43360 vss.n6962 vss.n6939 0.0702092
R43361 vss.t547 vss.n6962 0.0702092
R43362 vss.n6960 vss.n6955 0.0702092
R43363 vss.n6960 vss.t482 0.0702092
R43364 vss.n6959 vss.n6958 0.0702092
R43365 vss.n6964 vss.n6963 0.0702092
R43366 vss.n6976 vss.n6975 0.0702092
R43367 vss.n6973 vss.n6972 0.0702092
R43368 vss.n6434 vss.n6433 0.0702092
R43369 vss.n6434 vss.t1313 0.0702092
R43370 vss.t1491 vss.n6423 0.0702092
R43371 vss.n6427 vss.t900 0.0702092
R43372 vss.t902 vss.n6440 0.0702092
R43373 vss.n6436 vss.t1313 0.0702092
R43374 vss.n6442 vss.n6441 0.0702092
R43375 vss.n6441 vss.t902 0.0702092
R43376 vss.n6426 vss.n6403 0.0702092
R43377 vss.t900 vss.n6426 0.0702092
R43378 vss.n6424 vss.n6419 0.0702092
R43379 vss.n6424 vss.t1491 0.0702092
R43380 vss.n6423 vss.n6422 0.0702092
R43381 vss.n6428 vss.n6427 0.0702092
R43382 vss.n6440 vss.n6439 0.0702092
R43383 vss.n6437 vss.n6436 0.0702092
R43384 vss.n6356 vss.n6355 0.0702092
R43385 vss.n6356 vss.t1009 0.0702092
R43386 vss.t1356 vss.n6345 0.0702092
R43387 vss.n6349 vss.t189 0.0702092
R43388 vss.t188 vss.n6362 0.0702092
R43389 vss.n6358 vss.t1009 0.0702092
R43390 vss.n6364 vss.n6363 0.0702092
R43391 vss.n6363 vss.t188 0.0702092
R43392 vss.n6348 vss.n6325 0.0702092
R43393 vss.t189 vss.n6348 0.0702092
R43394 vss.n6346 vss.n6341 0.0702092
R43395 vss.n6346 vss.t1356 0.0702092
R43396 vss.n6345 vss.n6344 0.0702092
R43397 vss.n6350 vss.n6349 0.0702092
R43398 vss.n6362 vss.n6361 0.0702092
R43399 vss.n6359 vss.n6358 0.0702092
R43400 vss.n9352 vss.n9351 0.0702092
R43401 vss.n9352 vss.t1055 0.0702092
R43402 vss.t609 vss.n9341 0.0702092
R43403 vss.n9345 vss.t535 0.0702092
R43404 vss.t534 vss.n9358 0.0702092
R43405 vss.n9354 vss.t1055 0.0702092
R43406 vss.n9360 vss.n9359 0.0702092
R43407 vss.n9359 vss.t534 0.0702092
R43408 vss.n9344 vss.n9321 0.0702092
R43409 vss.t535 vss.n9344 0.0702092
R43410 vss.n9342 vss.n9337 0.0702092
R43411 vss.n9342 vss.t609 0.0702092
R43412 vss.n9341 vss.n9340 0.0702092
R43413 vss.n9346 vss.n9345 0.0702092
R43414 vss.n9358 vss.n9357 0.0702092
R43415 vss.n9355 vss.n9354 0.0702092
R43416 vss.n5958 vss.n5954 0.0702092
R43417 vss.n5958 vss.t1271 0.0702092
R43418 vss.n5969 vss.n5968 0.0702092
R43419 vss.t1214 vss.n5969 0.0702092
R43420 vss.n9680 vss.n9679 0.0702092
R43421 vss.n9679 vss.t564 0.0702092
R43422 vss.n5960 vss.n5938 0.0702092
R43423 vss.t563 vss.n5960 0.0702092
R43424 vss.n5957 vss.n5956 0.0702092
R43425 vss.t1271 vss.n5957 0.0702092
R43426 vss.n5962 vss.n5961 0.0702092
R43427 vss.n5961 vss.t563 0.0702092
R43428 vss.n9678 vss.n9677 0.0702092
R43429 vss.t564 vss.n9678 0.0702092
R43430 vss.n9675 vss.n9674 0.0702092
R43431 vss.n9674 vss.t1214 0.0702092
R43432 vss.n2579 vss.n2575 0.0702092
R43433 vss.n2579 vss.t1180 0.0702092
R43434 vss.n2590 vss.n2589 0.0702092
R43435 vss.t1014 vss.n2590 0.0702092
R43436 vss.n10008 vss.n10007 0.0702092
R43437 vss.n10007 vss.t1201 0.0702092
R43438 vss.n2581 vss.n2559 0.0702092
R43439 vss.t1200 vss.n2581 0.0702092
R43440 vss.n2578 vss.n2577 0.0702092
R43441 vss.t1180 vss.n2578 0.0702092
R43442 vss.n2583 vss.n2582 0.0702092
R43443 vss.n2582 vss.t1200 0.0702092
R43444 vss.n10006 vss.n10005 0.0702092
R43445 vss.t1201 vss.n10006 0.0702092
R43446 vss.n10003 vss.n10002 0.0702092
R43447 vss.n10002 vss.t1014 0.0702092
R43448 vss.n9762 vss.n9761 0.0702092
R43449 vss.n9761 vss.t641 0.0702092
R43450 vss.n9771 vss.n9770 0.0702092
R43451 vss.n9770 vss.t712 0.0702092
R43452 vss.n9774 vss.n9773 0.0702092
R43453 vss.n9774 vss.t713 0.0702092
R43454 vss.n9777 vss.n9776 0.0702092
R43455 vss.n9776 vss.t476 0.0702092
R43456 vss.n9767 vss.t641 0.0702092
R43457 vss.t712 vss.n9769 0.0702092
R43458 vss.n9782 vss.t713 0.0702092
R43459 vss.n9780 vss.t476 0.0702092
R43460 vss.n9780 vss.n9779 0.0702092
R43461 vss.n9783 vss.n9782 0.0702092
R43462 vss.n9769 vss.n9745 0.0702092
R43463 vss.n9767 vss.n9766 0.0702092
R43464 vss.n3202 vss.n3201 0.0702092
R43465 vss.n3201 vss.t451 0.0702092
R43466 vss.n3211 vss.n3210 0.0702092
R43467 vss.n3210 vss.t494 0.0702092
R43468 vss.n3214 vss.n3213 0.0702092
R43469 vss.n3214 vss.t492 0.0702092
R43470 vss.n3217 vss.n3216 0.0702092
R43471 vss.n3216 vss.t1358 0.0702092
R43472 vss.n3207 vss.t451 0.0702092
R43473 vss.t494 vss.n3209 0.0702092
R43474 vss.n3222 vss.t492 0.0702092
R43475 vss.n3220 vss.t1358 0.0702092
R43476 vss.n3220 vss.n3219 0.0702092
R43477 vss.n3223 vss.n3222 0.0702092
R43478 vss.n3209 vss.n3185 0.0702092
R43479 vss.n3207 vss.n3206 0.0702092
R43480 vss.n9801 vss.n9800 0.0702092
R43481 vss.t1056 vss.n9801 0.0702092
R43482 vss.n9798 vss.n9797 0.0702092
R43483 vss.n9797 vss.t968 0.0702092
R43484 vss.n3016 vss.n3015 0.0702092
R43485 vss.n3016 vss.t969 0.0702092
R43486 vss.n3019 vss.n3018 0.0702092
R43487 vss.n3018 vss.t625 0.0702092
R43488 vss.t1056 vss.n2995 0.0702092
R43489 vss.t968 vss.n9796 0.0702092
R43490 vss.n3024 vss.t969 0.0702092
R43491 vss.n3022 vss.t625 0.0702092
R43492 vss.n3022 vss.n3021 0.0702092
R43493 vss.n3025 vss.n3024 0.0702092
R43494 vss.n9796 vss.n9795 0.0702092
R43495 vss.n3005 vss.n2995 0.0702092
R43496 vss.n5232 vss.n5231 0.0702092
R43497 vss.n5231 vss.t399 0.0702092
R43498 vss.n5241 vss.n5240 0.0702092
R43499 vss.n5240 vss.t1185 0.0702092
R43500 vss.n5244 vss.n5243 0.0702092
R43501 vss.n5244 vss.t1186 0.0702092
R43502 vss.n5247 vss.n5246 0.0702092
R43503 vss.n5246 vss.t480 0.0702092
R43504 vss.n5237 vss.t399 0.0702092
R43505 vss.t1185 vss.n5239 0.0702092
R43506 vss.n5252 vss.t1186 0.0702092
R43507 vss.n5250 vss.t480 0.0702092
R43508 vss.n5250 vss.n5249 0.0702092
R43509 vss.n5253 vss.n5252 0.0702092
R43510 vss.n5239 vss.n5215 0.0702092
R43511 vss.n5237 vss.n5236 0.0702092
R43512 vss.n3045 vss.n3044 0.0702092
R43513 vss.n3044 vss.t517 0.0702092
R43514 vss.n3054 vss.n3053 0.0702092
R43515 vss.n3053 vss.t198 0.0702092
R43516 vss.n3057 vss.n3056 0.0702092
R43517 vss.n3057 vss.t199 0.0702092
R43518 vss.n3060 vss.n3059 0.0702092
R43519 vss.n3059 vss.t1366 0.0702092
R43520 vss.n3050 vss.t517 0.0702092
R43521 vss.t198 vss.n3052 0.0702092
R43522 vss.n3065 vss.t199 0.0702092
R43523 vss.n3063 vss.t1366 0.0702092
R43524 vss.n3063 vss.n3062 0.0702092
R43525 vss.n3066 vss.n3065 0.0702092
R43526 vss.n3052 vss.n3028 0.0702092
R43527 vss.n3050 vss.n3049 0.0702092
R43528 vss.n5102 vss.n5101 0.0702092
R43529 vss.n5101 vss.t441 0.0702092
R43530 vss.n5111 vss.n5110 0.0702092
R43531 vss.n5110 vss.t0 0.0702092
R43532 vss.n5114 vss.n5113 0.0702092
R43533 vss.n5114 vss.t1 0.0702092
R43534 vss.n5117 vss.n5116 0.0702092
R43535 vss.n5116 vss.t1485 0.0702092
R43536 vss.n5107 vss.t441 0.0702092
R43537 vss.t0 vss.n5109 0.0702092
R43538 vss.n5122 vss.t1 0.0702092
R43539 vss.n5120 vss.t1485 0.0702092
R43540 vss.n5120 vss.n5119 0.0702092
R43541 vss.n5123 vss.n5122 0.0702092
R43542 vss.n5109 vss.n5085 0.0702092
R43543 vss.n5107 vss.n5106 0.0702092
R43544 vss.n5291 vss.n5290 0.0702092
R43545 vss.n5290 vss.t707 0.0702092
R43546 vss.n5300 vss.n5299 0.0702092
R43547 vss.n5299 vss.t704 0.0702092
R43548 vss.n5303 vss.n5302 0.0702092
R43549 vss.n5303 vss.t705 0.0702092
R43550 vss.n5306 vss.n5305 0.0702092
R43551 vss.n5305 vss.t1348 0.0702092
R43552 vss.n5296 vss.t707 0.0702092
R43553 vss.t704 vss.n5298 0.0702092
R43554 vss.n5311 vss.t705 0.0702092
R43555 vss.n5309 vss.t1348 0.0702092
R43556 vss.n5309 vss.n5308 0.0702092
R43557 vss.n5312 vss.n5311 0.0702092
R43558 vss.n5298 vss.n5274 0.0702092
R43559 vss.n5296 vss.n5295 0.0702092
R43560 vss.n5019 vss.n5018 0.0702092
R43561 vss.n5018 vss.t637 0.0702092
R43562 vss.n5028 vss.n5027 0.0702092
R43563 vss.n5027 vss.t1162 0.0702092
R43564 vss.n5031 vss.n5030 0.0702092
R43565 vss.n5031 vss.t1163 0.0702092
R43566 vss.n5034 vss.n5033 0.0702092
R43567 vss.n5033 vss.t1380 0.0702092
R43568 vss.n5024 vss.t637 0.0702092
R43569 vss.t1162 vss.n5026 0.0702092
R43570 vss.n5039 vss.t1163 0.0702092
R43571 vss.n5037 vss.t1380 0.0702092
R43572 vss.n5037 vss.n5036 0.0702092
R43573 vss.n5040 vss.n5039 0.0702092
R43574 vss.n5026 vss.n5002 0.0702092
R43575 vss.n5024 vss.n5023 0.0702092
R43576 vss.n4900 vss.n4899 0.0702092
R43577 vss.n4899 vss.t436 0.0702092
R43578 vss.n4909 vss.n4908 0.0702092
R43579 vss.n4908 vss.t603 0.0702092
R43580 vss.n4912 vss.n4911 0.0702092
R43581 vss.n4912 vss.t604 0.0702092
R43582 vss.n4915 vss.n4914 0.0702092
R43583 vss.n4914 vss.t1085 0.0702092
R43584 vss.n4905 vss.t436 0.0702092
R43585 vss.t603 vss.n4907 0.0702092
R43586 vss.n4920 vss.t604 0.0702092
R43587 vss.n4918 vss.t1085 0.0702092
R43588 vss.n4918 vss.n4917 0.0702092
R43589 vss.n4921 vss.n4920 0.0702092
R43590 vss.n4907 vss.n4883 0.0702092
R43591 vss.n4905 vss.n4904 0.0702092
R43592 vss.n9924 vss.n9923 0.0702092
R43593 vss.n9923 vss.t777 0.0702092
R43594 vss.n9913 vss.n9912 0.0702092
R43595 vss.n9912 vss.t69 0.0702092
R43596 vss.n2728 vss.n2726 0.0702092
R43597 vss.t778 vss.n2726 0.0702092
R43598 vss.n9922 vss.n9921 0.0702092
R43599 vss.t777 vss.n9922 0.0702092
R43600 vss.n9919 vss.n9918 0.0702092
R43601 vss.n9918 vss.t778 0.0702092
R43602 vss.n2731 vss.n2730 0.0702092
R43603 vss.n2731 vss.t69 0.0702092
R43604 vss.n9904 vss.n9903 0.0702092
R43605 vss.n9903 vss.t1044 0.0702092
R43606 vss.n2738 vss.n2737 0.0702092
R43607 vss.n2738 vss.t1044 0.0702092
R43608 vss.n4645 vss.n2735 0.0702092
R43609 vss.n4645 vss.t28 0.0702092
R43610 vss.n4661 vss.n4660 0.0702092
R43611 vss.n4660 vss.t30 0.0702092
R43612 vss.n4663 vss.n4638 0.0702092
R43613 vss.n4638 vss.t31 0.0702092
R43614 vss.n4639 vss.n4637 0.0702092
R43615 vss.n4637 vss.t31 0.0702092
R43616 vss.n4659 vss.n4658 0.0702092
R43617 vss.t30 vss.n4659 0.0702092
R43618 vss.n4656 vss.n4655 0.0702092
R43619 vss.n4655 vss.t28 0.0702092
R43620 vss.n5628 vss.n4629 0.0702092
R43621 vss.n4629 vss.t752 0.0702092
R43622 vss.n4630 vss.n4628 0.0702092
R43623 vss.n4628 vss.t752 0.0702092
R43624 vss.n5615 vss.n5614 0.0702092
R43625 vss.n5614 vss.t587 0.0702092
R43626 vss.n4680 vss.n4678 0.0702092
R43627 vss.t750 vss.n4678 0.0702092
R43628 vss.n5626 vss.n5625 0.0702092
R43629 vss.n5625 vss.t749 0.0702092
R43630 vss.n5624 vss.n5623 0.0702092
R43631 vss.t749 vss.n5624 0.0702092
R43632 vss.n5621 vss.n5620 0.0702092
R43633 vss.n5620 vss.t750 0.0702092
R43634 vss.n4683 vss.n4682 0.0702092
R43635 vss.n4683 vss.t587 0.0702092
R43636 vss.n5606 vss.n5605 0.0702092
R43637 vss.n5605 vss.t787 0.0702092
R43638 vss.n5603 vss.n5602 0.0702092
R43639 vss.n5603 vss.t787 0.0702092
R43640 vss.n5600 vss.n5599 0.0702092
R43641 vss.n5599 vss.t1420 0.0702092
R43642 vss.n5597 vss.n4690 0.0702092
R43643 vss.n5597 vss.t1419 0.0702092
R43644 vss.n5587 vss.n5586 0.0702092
R43645 vss.t253 vss.n5587 0.0702092
R43646 vss.n5589 vss.n5588 0.0702092
R43647 vss.n5588 vss.t253 0.0702092
R43648 vss.n5596 vss.n5595 0.0702092
R43649 vss.t1419 vss.n5596 0.0702092
R43650 vss.n5593 vss.n5592 0.0702092
R43651 vss.n5592 vss.t1420 0.0702092
R43652 vss.n4707 vss.n4706 0.0702092
R43653 vss.n4706 vss.t699 0.0702092
R43654 vss.n4704 vss.n4703 0.0702092
R43655 vss.n4704 vss.t699 0.0702092
R43656 vss.n4726 vss.n4725 0.0702092
R43657 vss.t67 vss.n4726 0.0702092
R43658 vss.n5575 vss.n4711 0.0702092
R43659 vss.n5575 vss.t1233 0.0702092
R43660 vss.n5578 vss.n5577 0.0702092
R43661 vss.n5577 vss.t1232 0.0702092
R43662 vss.n4718 vss.n4717 0.0702092
R43663 vss.n4717 vss.t1232 0.0702092
R43664 vss.n5574 vss.n5573 0.0702092
R43665 vss.t1233 vss.n5574 0.0702092
R43666 vss.n5571 vss.n5570 0.0702092
R43667 vss.n5570 vss.t67 0.0702092
R43668 vss.n5563 vss.n5562 0.0702092
R43669 vss.n5562 vss.t845 0.0702092
R43670 vss.n5560 vss.n5559 0.0702092
R43671 vss.n5560 vss.t845 0.0702092
R43672 vss.n5557 vss.n5556 0.0702092
R43673 vss.n5556 vss.t659 0.0702092
R43674 vss.n5554 vss.n4733 0.0702092
R43675 vss.n5554 vss.t661 0.0702092
R43676 vss.n5544 vss.n5543 0.0702092
R43677 vss.t313 vss.n5544 0.0702092
R43678 vss.n5546 vss.n5545 0.0702092
R43679 vss.n5545 vss.t313 0.0702092
R43680 vss.n5553 vss.n5552 0.0702092
R43681 vss.t661 vss.n5553 0.0702092
R43682 vss.n5550 vss.n5549 0.0702092
R43683 vss.n5549 vss.t659 0.0702092
R43684 vss.n4750 vss.n4749 0.0702092
R43685 vss.n4749 vss.t938 0.0702092
R43686 vss.n4747 vss.n4746 0.0702092
R43687 vss.n4747 vss.t938 0.0702092
R43688 vss.n4769 vss.n4768 0.0702092
R43689 vss.t1155 vss.n4769 0.0702092
R43690 vss.n5532 vss.n4754 0.0702092
R43691 vss.n5532 vss.t804 0.0702092
R43692 vss.n5535 vss.n5534 0.0702092
R43693 vss.n5534 vss.t803 0.0702092
R43694 vss.n4761 vss.n4760 0.0702092
R43695 vss.n4760 vss.t803 0.0702092
R43696 vss.n5531 vss.n5530 0.0702092
R43697 vss.t804 vss.n5531 0.0702092
R43698 vss.n5528 vss.n5527 0.0702092
R43699 vss.n5527 vss.t1155 0.0702092
R43700 vss.n5520 vss.n5519 0.0702092
R43701 vss.n5519 vss.t966 0.0702092
R43702 vss.n5517 vss.n5516 0.0702092
R43703 vss.n5517 vss.t966 0.0702092
R43704 vss.n5514 vss.n5513 0.0702092
R43705 vss.n5513 vss.t1221 0.0702092
R43706 vss.n5511 vss.n4776 0.0702092
R43707 vss.n5511 vss.t1220 0.0702092
R43708 vss.n5501 vss.n5500 0.0702092
R43709 vss.t1286 vss.n5501 0.0702092
R43710 vss.n5503 vss.n5502 0.0702092
R43711 vss.n5502 vss.t1286 0.0702092
R43712 vss.n5510 vss.n5509 0.0702092
R43713 vss.t1220 vss.n5510 0.0702092
R43714 vss.n5507 vss.n5506 0.0702092
R43715 vss.n5506 vss.t1221 0.0702092
R43716 vss.n4793 vss.n4792 0.0702092
R43717 vss.n4792 vss.t812 0.0702092
R43718 vss.n4790 vss.n4789 0.0702092
R43719 vss.n4790 vss.t812 0.0702092
R43720 vss.n4812 vss.n4811 0.0702092
R43721 vss.t818 vss.n4812 0.0702092
R43722 vss.n5489 vss.n4797 0.0702092
R43723 vss.n5489 vss.t1537 0.0702092
R43724 vss.n5492 vss.n5491 0.0702092
R43725 vss.n5491 vss.t1539 0.0702092
R43726 vss.n4804 vss.n4803 0.0702092
R43727 vss.n4803 vss.t1539 0.0702092
R43728 vss.n5488 vss.n5487 0.0702092
R43729 vss.t1537 vss.n5488 0.0702092
R43730 vss.n5485 vss.n5484 0.0702092
R43731 vss.n5484 vss.t818 0.0702092
R43732 vss.n5477 vss.n5476 0.0702092
R43733 vss.n5476 vss.t878 0.0702092
R43734 vss.n5474 vss.n5473 0.0702092
R43735 vss.n5474 vss.t878 0.0702092
R43736 vss.n5471 vss.n5470 0.0702092
R43737 vss.n5470 vss.t337 0.0702092
R43738 vss.n5468 vss.n4819 0.0702092
R43739 vss.n5468 vss.t336 0.0702092
R43740 vss.n5458 vss.n5457 0.0702092
R43741 vss.t34 vss.n5458 0.0702092
R43742 vss.n5460 vss.n5459 0.0702092
R43743 vss.n5459 vss.t34 0.0702092
R43744 vss.n5467 vss.n5466 0.0702092
R43745 vss.t336 vss.n5467 0.0702092
R43746 vss.n5464 vss.n5463 0.0702092
R43747 vss.n5463 vss.t337 0.0702092
R43748 vss.n4836 vss.n4835 0.0702092
R43749 vss.n4835 vss.t1438 0.0702092
R43750 vss.n4833 vss.n4832 0.0702092
R43751 vss.n4833 vss.t1438 0.0702092
R43752 vss.n4855 vss.n4854 0.0702092
R43753 vss.t601 vss.n4855 0.0702092
R43754 vss.n5446 vss.n4840 0.0702092
R43755 vss.n5446 vss.t1526 0.0702092
R43756 vss.n5449 vss.n5448 0.0702092
R43757 vss.n5448 vss.t1525 0.0702092
R43758 vss.n4847 vss.n4846 0.0702092
R43759 vss.n4846 vss.t1525 0.0702092
R43760 vss.n5445 vss.n5444 0.0702092
R43761 vss.t1526 vss.n5445 0.0702092
R43762 vss.n5442 vss.n5441 0.0702092
R43763 vss.n5441 vss.t601 0.0702092
R43764 vss.n5434 vss.n5433 0.0702092
R43765 vss.n5433 vss.t964 0.0702092
R43766 vss.n5431 vss.n5430 0.0702092
R43767 vss.n5431 vss.t964 0.0702092
R43768 vss.n5428 vss.n5427 0.0702092
R43769 vss.n5427 vss.t1243 0.0702092
R43770 vss.n5425 vss.n4862 0.0702092
R43771 vss.n5425 vss.t1242 0.0702092
R43772 vss.n5415 vss.n5414 0.0702092
R43773 vss.t934 vss.n5415 0.0702092
R43774 vss.n5417 vss.n5416 0.0702092
R43775 vss.n5416 vss.t934 0.0702092
R43776 vss.n5424 vss.n5423 0.0702092
R43777 vss.t1242 vss.n5424 0.0702092
R43778 vss.n5421 vss.n5420 0.0702092
R43779 vss.n5420 vss.t1243 0.0702092
R43780 vss.n4879 vss.n4878 0.0702092
R43781 vss.n4878 vss.t1265 0.0702092
R43782 vss.n4876 vss.n4875 0.0702092
R43783 vss.n4876 vss.t1265 0.0702092
R43784 vss.n5349 vss.n5348 0.0702092
R43785 vss.t180 vss.n5349 0.0702092
R43786 vss.n5403 vss.n5334 0.0702092
R43787 vss.n5403 vss.t192 0.0702092
R43788 vss.n5406 vss.n5405 0.0702092
R43789 vss.n5405 vss.t191 0.0702092
R43790 vss.n5341 vss.n5340 0.0702092
R43791 vss.n5340 vss.t191 0.0702092
R43792 vss.n5402 vss.n5401 0.0702092
R43793 vss.t192 vss.n5402 0.0702092
R43794 vss.n5399 vss.n5398 0.0702092
R43795 vss.n5398 vss.t180 0.0702092
R43796 vss.n5376 vss.n5375 0.0702092
R43797 vss.t744 vss.n5376 0.0702092
R43798 vss.n5373 vss.n5372 0.0702092
R43799 vss.n5372 vss.t741 0.0702092
R43800 vss.n5370 vss.n5369 0.0702092
R43801 vss.n5370 vss.t742 0.0702092
R43802 vss.n5387 vss.n5386 0.0702092
R43803 vss.n5387 vss.t55 0.0702092
R43804 vss.n5377 vss.t744 0.0702092
R43805 vss.n5381 vss.t741 0.0702092
R43806 vss.n5383 vss.t742 0.0702092
R43807 vss.n5390 vss.t55 0.0702092
R43808 vss.n5391 vss.n5390 0.0702092
R43809 vss.n5384 vss.n5383 0.0702092
R43810 vss.n5381 vss.n5380 0.0702092
R43811 vss.n5378 vss.n5377 0.0702092
R43812 vss.n9821 vss.n9820 0.0702092
R43813 vss.n9820 vss.t154 0.0702092
R43814 vss.n9830 vss.n9829 0.0702092
R43815 vss.n9829 vss.t410 0.0702092
R43816 vss.n9833 vss.n9832 0.0702092
R43817 vss.n9833 vss.t408 0.0702092
R43818 vss.n9836 vss.n9835 0.0702092
R43819 vss.n9835 vss.t15 0.0702092
R43820 vss.n9826 vss.t154 0.0702092
R43821 vss.t410 vss.n9828 0.0702092
R43822 vss.n9841 vss.t408 0.0702092
R43823 vss.n9839 vss.t15 0.0702092
R43824 vss.n9839 vss.n9838 0.0702092
R43825 vss.n9842 vss.n9841 0.0702092
R43826 vss.n9828 vss.n2873 0.0702092
R43827 vss.n9826 vss.n9825 0.0702092
R43828 vss.n2978 vss.n2977 0.0702092
R43829 vss.t491 vss.n2978 0.0702092
R43830 vss.n2975 vss.n2974 0.0702092
R43831 vss.n2974 vss.t1425 0.0702092
R43832 vss.n2959 vss.n2958 0.0702092
R43833 vss.n2959 vss.t1423 0.0702092
R43834 vss.n2962 vss.n2961 0.0702092
R43835 vss.n2961 vss.t1318 0.0702092
R43836 vss.t491 vss.n2938 0.0702092
R43837 vss.t1425 vss.n2973 0.0702092
R43838 vss.n2967 vss.t1423 0.0702092
R43839 vss.n2965 vss.t1318 0.0702092
R43840 vss.n2965 vss.n2964 0.0702092
R43841 vss.n2968 vss.n2967 0.0702092
R43842 vss.n2973 vss.n2972 0.0702092
R43843 vss.n2948 vss.n2938 0.0702092
R43844 vss.n2932 vss.n2931 0.0702092
R43845 vss.t335 vss.n2932 0.0702092
R43846 vss.n2929 vss.n2928 0.0702092
R43847 vss.n2928 vss.t789 0.0702092
R43848 vss.n2912 vss.n2911 0.0702092
R43849 vss.n2912 vss.t790 0.0702092
R43850 vss.n2915 vss.n2914 0.0702092
R43851 vss.n2914 vss.t470 0.0702092
R43852 vss.t335 vss.n2891 0.0702092
R43853 vss.t789 vss.n2927 0.0702092
R43854 vss.n2920 vss.t790 0.0702092
R43855 vss.n2918 vss.t470 0.0702092
R43856 vss.n2918 vss.n2917 0.0702092
R43857 vss.n2921 vss.n2920 0.0702092
R43858 vss.n2927 vss.n2926 0.0702092
R43859 vss.n2901 vss.n2891 0.0702092
R43860 vss.n4941 vss.n4940 0.0702092
R43861 vss.n4940 vss.t832 0.0702092
R43862 vss.n4950 vss.n4949 0.0702092
R43863 vss.n4949 vss.t1237 0.0702092
R43864 vss.n4953 vss.n4952 0.0702092
R43865 vss.n4953 vss.t1235 0.0702092
R43866 vss.n4956 vss.n4955 0.0702092
R43867 vss.n4955 vss.t1509 0.0702092
R43868 vss.n4946 vss.t832 0.0702092
R43869 vss.t1237 vss.n4948 0.0702092
R43870 vss.n4961 vss.t1235 0.0702092
R43871 vss.n4959 vss.t1509 0.0702092
R43872 vss.n4959 vss.n4958 0.0702092
R43873 vss.n4962 vss.n4961 0.0702092
R43874 vss.n4948 vss.n4924 0.0702092
R43875 vss.n4946 vss.n4945 0.0702092
R43876 vss.n5143 vss.n5142 0.0702092
R43877 vss.n5142 vss.t146 0.0702092
R43878 vss.n5152 vss.n5151 0.0702092
R43879 vss.n5151 vss.t1307 0.0702092
R43880 vss.n5155 vss.n5154 0.0702092
R43881 vss.n5155 vss.t1308 0.0702092
R43882 vss.n5158 vss.n5157 0.0702092
R43883 vss.n5157 vss.t508 0.0702092
R43884 vss.n5148 vss.t146 0.0702092
R43885 vss.t1307 vss.n5150 0.0702092
R43886 vss.n5163 vss.t1308 0.0702092
R43887 vss.n5161 vss.t508 0.0702092
R43888 vss.n5161 vss.n5160 0.0702092
R43889 vss.n5164 vss.n5163 0.0702092
R43890 vss.n5150 vss.n5126 0.0702092
R43891 vss.n5148 vss.n5147 0.0702092
R43892 vss.n3124 vss.n3123 0.0702092
R43893 vss.n3123 vss.t240 0.0702092
R43894 vss.n3133 vss.n3132 0.0702092
R43895 vss.n3132 vss.t710 0.0702092
R43896 vss.n3136 vss.n3135 0.0702092
R43897 vss.n3136 vss.t708 0.0702092
R43898 vss.n3139 vss.n3138 0.0702092
R43899 vss.n3138 vss.t1342 0.0702092
R43900 vss.n3129 vss.t240 0.0702092
R43901 vss.t710 vss.n3131 0.0702092
R43902 vss.n3144 vss.t708 0.0702092
R43903 vss.n3142 vss.t1342 0.0702092
R43904 vss.n3142 vss.n3141 0.0702092
R43905 vss.n3145 vss.n3144 0.0702092
R43906 vss.n3131 vss.n3106 0.0702092
R43907 vss.n3129 vss.n3128 0.0702092
R43908 vss.n4483 vss.n4482 0.0702092
R43909 vss.t580 vss.n4483 0.0702092
R43910 vss.n4488 vss.n4487 0.0702092
R43911 vss.n4487 vss.t159 0.0702092
R43912 vss.n4490 vss.n4467 0.0702092
R43913 vss.t161 vss.n4467 0.0702092
R43914 vss.n4496 vss.n4495 0.0702092
R43915 vss.n4496 vss.t1206 0.0702092
R43916 vss.n4493 vss.n4492 0.0702092
R43917 vss.n4492 vss.t1206 0.0702092
R43918 vss.n4501 vss.n4500 0.0702092
R43919 vss.n4500 vss.t161 0.0702092
R43920 vss.n4486 vss.n4462 0.0702092
R43921 vss.t159 vss.n4486 0.0702092
R43922 vss.n4484 vss.n4479 0.0702092
R43923 vss.n4484 vss.t580 0.0702092
R43924 vss.n4391 vss.n4390 0.0702092
R43925 vss.t568 vss.n4391 0.0702092
R43926 vss.n4396 vss.n4395 0.0702092
R43927 vss.n4395 vss.t488 0.0702092
R43928 vss.n4398 vss.n4375 0.0702092
R43929 vss.t490 vss.n4375 0.0702092
R43930 vss.n4404 vss.n4403 0.0702092
R43931 vss.n4404 vss.t1062 0.0702092
R43932 vss.n4401 vss.n4400 0.0702092
R43933 vss.n4400 vss.t1062 0.0702092
R43934 vss.n4409 vss.n4408 0.0702092
R43935 vss.n4408 vss.t490 0.0702092
R43936 vss.n4394 vss.n4370 0.0702092
R43937 vss.t488 vss.n4394 0.0702092
R43938 vss.n4392 vss.n4387 0.0702092
R43939 vss.n4392 vss.t568 0.0702092
R43940 vss.n4343 vss.n4342 0.0702092
R43941 vss.t1503 vss.n4343 0.0702092
R43942 vss.n4348 vss.n4347 0.0702092
R43943 vss.n4347 vss.t1259 0.0702092
R43944 vss.n4350 vss.n4327 0.0702092
R43945 vss.t1261 vss.n4327 0.0702092
R43946 vss.n4356 vss.n4355 0.0702092
R43947 vss.n4356 vss.t975 0.0702092
R43948 vss.n4353 vss.n4352 0.0702092
R43949 vss.n4352 vss.t975 0.0702092
R43950 vss.n4361 vss.n4360 0.0702092
R43951 vss.n4360 vss.t1261 0.0702092
R43952 vss.n4346 vss.n4322 0.0702092
R43953 vss.t1259 vss.n4346 0.0702092
R43954 vss.n4344 vss.n4339 0.0702092
R43955 vss.n4344 vss.t1503 0.0702092
R43956 vss.n3743 vss.n3742 0.0702092
R43957 vss.t1071 vss.n3743 0.0702092
R43958 vss.n3748 vss.n3747 0.0702092
R43959 vss.n3747 vss.t1255 0.0702092
R43960 vss.n3750 vss.n3727 0.0702092
R43961 vss.t1257 vss.n3727 0.0702092
R43962 vss.n3756 vss.n3755 0.0702092
R43963 vss.n3756 vss.t1116 0.0702092
R43964 vss.n3753 vss.n3752 0.0702092
R43965 vss.n3752 vss.t1116 0.0702092
R43966 vss.n3761 vss.n3760 0.0702092
R43967 vss.n3760 vss.t1257 0.0702092
R43968 vss.n3746 vss.n3722 0.0702092
R43969 vss.t1255 vss.n3746 0.0702092
R43970 vss.n3744 vss.n3739 0.0702092
R43971 vss.n3744 vss.t1071 0.0702092
R43972 vss.n4045 vss.n4044 0.0702092
R43973 vss.t623 vss.n4045 0.0702092
R43974 vss.n4050 vss.n4049 0.0702092
R43975 vss.n4049 vss.t1126 0.0702092
R43976 vss.n4052 vss.n4029 0.0702092
R43977 vss.t1125 vss.n4029 0.0702092
R43978 vss.n4058 vss.n4057 0.0702092
R43979 vss.n4058 vss.t316 0.0702092
R43980 vss.n4055 vss.n4054 0.0702092
R43981 vss.n4054 vss.t316 0.0702092
R43982 vss.n4063 vss.n4062 0.0702092
R43983 vss.n4062 vss.t1125 0.0702092
R43984 vss.n4048 vss.n4024 0.0702092
R43985 vss.t1126 vss.n4048 0.0702092
R43986 vss.n4046 vss.n4041 0.0702092
R43987 vss.n4046 vss.t623 0.0702092
R43988 vss.n3698 vss.n3697 0.0702092
R43989 vss.t1493 vss.n3698 0.0702092
R43990 vss.n3703 vss.n3702 0.0702092
R43991 vss.n3702 vss.t1441 0.0702092
R43992 vss.n3705 vss.n3682 0.0702092
R43993 vss.t1440 vss.n3682 0.0702092
R43994 vss.n3711 vss.n3710 0.0702092
R43995 vss.n3711 vss.t1443 0.0702092
R43996 vss.n3708 vss.n3707 0.0702092
R43997 vss.n3707 vss.t1443 0.0702092
R43998 vss.n3716 vss.n3715 0.0702092
R43999 vss.n3715 vss.t1440 0.0702092
R44000 vss.n3701 vss.n3677 0.0702092
R44001 vss.t1441 vss.n3701 0.0702092
R44002 vss.n3699 vss.n3694 0.0702092
R44003 vss.n3699 vss.t1493 0.0702092
R44004 vss.n4099 vss.n4098 0.0702092
R44005 vss.t1483 vss.n4099 0.0702092
R44006 vss.n4104 vss.n4103 0.0702092
R44007 vss.n4103 vss.t352 0.0702092
R44008 vss.n4106 vss.n4083 0.0702092
R44009 vss.t354 vss.n4083 0.0702092
R44010 vss.n4112 vss.n4111 0.0702092
R44011 vss.n4112 vss.t197 0.0702092
R44012 vss.n4109 vss.n4108 0.0702092
R44013 vss.n4108 vss.t197 0.0702092
R44014 vss.n4117 vss.n4116 0.0702092
R44015 vss.n4116 vss.t354 0.0702092
R44016 vss.n4102 vss.n4078 0.0702092
R44017 vss.t352 vss.n4102 0.0702092
R44018 vss.n4100 vss.n4095 0.0702092
R44019 vss.n4100 vss.t1483 0.0702092
R44020 vss.n3523 vss.n3522 0.0702092
R44021 vss.t566 vss.n3523 0.0702092
R44022 vss.n3528 vss.n3527 0.0702092
R44023 vss.n3527 vss.t727 0.0702092
R44024 vss.n3530 vss.n3507 0.0702092
R44025 vss.t729 vss.n3507 0.0702092
R44026 vss.n3536 vss.n3535 0.0702092
R44027 vss.n3536 vss.t551 0.0702092
R44028 vss.n3533 vss.n3532 0.0702092
R44029 vss.n3532 vss.t551 0.0702092
R44030 vss.n3541 vss.n3540 0.0702092
R44031 vss.n3540 vss.t729 0.0702092
R44032 vss.n3526 vss.n3502 0.0702092
R44033 vss.t727 vss.n3526 0.0702092
R44034 vss.n3524 vss.n3519 0.0702092
R44035 vss.n3524 vss.t566 0.0702092
R44036 vss.n3478 vss.n3477 0.0702092
R44037 vss.t617 vss.n3478 0.0702092
R44038 vss.n3483 vss.n3482 0.0702092
R44039 vss.n3482 vss.t1212 0.0702092
R44040 vss.n3485 vss.n3462 0.0702092
R44041 vss.t1211 vss.n3462 0.0702092
R44042 vss.n3491 vss.n3490 0.0702092
R44043 vss.n3491 vss.t124 0.0702092
R44044 vss.n3488 vss.n3487 0.0702092
R44045 vss.n3487 vss.t124 0.0702092
R44046 vss.n3496 vss.n3495 0.0702092
R44047 vss.n3495 vss.t1211 0.0702092
R44048 vss.n3481 vss.n3457 0.0702092
R44049 vss.t1212 vss.n3481 0.0702092
R44050 vss.n3479 vss.n3474 0.0702092
R44051 vss.n3479 vss.t617 0.0702092
R44052 vss.n5766 vss.n5765 0.0702092
R44053 vss.t379 vss.n5766 0.0702092
R44054 vss.n5771 vss.n5770 0.0702092
R44055 vss.n5770 vss.t746 0.0702092
R44056 vss.n5773 vss.n5750 0.0702092
R44057 vss.t748 vss.n5750 0.0702092
R44058 vss.n5779 vss.n5778 0.0702092
R44059 vss.n5779 vss.t78 0.0702092
R44060 vss.n5776 vss.n5775 0.0702092
R44061 vss.n5775 vss.t78 0.0702092
R44062 vss.n5784 vss.n5783 0.0702092
R44063 vss.n5783 vss.t748 0.0702092
R44064 vss.n5769 vss.n5745 0.0702092
R44065 vss.t746 vss.n5769 0.0702092
R44066 vss.n5767 vss.n5762 0.0702092
R44067 vss.n5767 vss.t379 0.0702092
R44068 vss.n4520 vss.n4451 0.0702092
R44069 vss.t724 vss.n4451 0.0702092
R44070 vss.n4522 vss.n4454 0.0702092
R44071 vss.t726 vss.n4454 0.0702092
R44072 vss.n4525 vss.n4524 0.0702092
R44073 vss.t1178 vss.n4525 0.0702092
R44074 vss.n4527 vss.n4526 0.0702092
R44075 vss.n4526 vss.t1178 0.0702092
R44076 vss.n4530 vss.n4529 0.0702092
R44077 vss.t726 vss.n4530 0.0702092
R44078 vss.n4532 vss.n4449 0.0702092
R44079 vss.n4532 vss.t724 0.0702092
R44080 vss.n4534 vss.n4446 0.0702092
R44081 vss.t948 vss.n4444 0.0702092
R44082 vss.t948 vss.n4534 0.0702092
R44083 vss.n4518 vss.n4444 0.0702092
R44084 vss.n4540 vss.n4539 0.0702092
R44085 vss.n4539 vss.t442 0.0702092
R44086 vss.n4543 vss.n4542 0.0702092
R44087 vss.t456 vss.n4543 0.0702092
R44088 vss.n4551 vss.n4550 0.0702092
R44089 vss.n4550 vss.t458 0.0702092
R44090 vss.n4549 vss.n4548 0.0702092
R44091 vss.t458 vss.n4549 0.0702092
R44092 vss.n4545 vss.n4544 0.0702092
R44093 vss.n4544 vss.t456 0.0702092
R44094 vss.n4538 vss.n4537 0.0702092
R44095 vss.t442 vss.n4538 0.0702092
R44096 vss.n4556 vss.n4425 0.0702092
R44097 vss.t155 vss.n4423 0.0702092
R44098 vss.t155 vss.n4556 0.0702092
R44099 vss.n4553 vss.n4423 0.0702092
R44100 vss.n4595 vss.n4594 0.0702092
R44101 vss.n4594 vss.t695 0.0702092
R44102 vss.n4597 vss.n4419 0.0702092
R44103 vss.t697 vss.n4419 0.0702092
R44104 vss.n4603 vss.n4602 0.0702092
R44105 vss.n4603 vss.t698 0.0702092
R44106 vss.n4600 vss.n4599 0.0702092
R44107 vss.n4599 vss.t698 0.0702092
R44108 vss.n4608 vss.n4607 0.0702092
R44109 vss.n4607 vss.t697 0.0702092
R44110 vss.n4593 vss.n4414 0.0702092
R44111 vss.t695 vss.n4593 0.0702092
R44112 vss.n4591 vss.n4569 0.0702092
R44113 vss.t916 vss.n4590 0.0702092
R44114 vss.n4591 vss.t916 0.0702092
R44115 vss.n4590 vss.n4589 0.0702092
R44116 vss.n4583 vss.n4571 0.0702092
R44117 vss.n4571 vss.t597 0.0702092
R44118 vss.n4581 vss.n4580 0.0702092
R44119 vss.n4580 vss.t1267 0.0702092
R44120 vss.n4622 vss.n4621 0.0702092
R44121 vss.n4621 vss.t1269 0.0702092
R44122 vss.n4620 vss.n4619 0.0702092
R44123 vss.t1269 vss.n4620 0.0702092
R44124 vss.n4579 vss.n3645 0.0702092
R44125 vss.t1267 vss.n4579 0.0702092
R44126 vss.n4572 vss.n4570 0.0702092
R44127 vss.n4570 vss.t597 0.0702092
R44128 vss.n3633 vss.n3631 0.0702092
R44129 vss.n3632 vss.t465 0.0702092
R44130 vss.n3631 vss.t465 0.0702092
R44131 vss.n4624 vss.n3632 0.0702092
R44132 vss.n4192 vss.n4191 0.0702092
R44133 vss.n4191 vss.t234 0.0702092
R44134 vss.n4194 vss.n3769 0.0702092
R44135 vss.t233 vss.n3769 0.0702092
R44136 vss.n4200 vss.n4199 0.0702092
R44137 vss.n4200 vss.t89 0.0702092
R44138 vss.n4197 vss.n4196 0.0702092
R44139 vss.n4196 vss.t89 0.0702092
R44140 vss.n4205 vss.n4204 0.0702092
R44141 vss.n4204 vss.t233 0.0702092
R44142 vss.n4190 vss.n3764 0.0702092
R44143 vss.t234 vss.n4190 0.0702092
R44144 vss.n4188 vss.n3783 0.0702092
R44145 vss.t1036 vss.n4187 0.0702092
R44146 vss.n4188 vss.t1036 0.0702092
R44147 vss.n4187 vss.n4186 0.0702092
R44148 vss.n4180 vss.n3785 0.0702092
R44149 vss.n3785 vss.t867 0.0702092
R44150 vss.n4178 vss.n4177 0.0702092
R44151 vss.n4177 vss.t373 0.0702092
R44152 vss.n3821 vss.n3820 0.0702092
R44153 vss.n3820 vss.t375 0.0702092
R44154 vss.n3819 vss.n3799 0.0702092
R44155 vss.t375 vss.n3819 0.0702092
R44156 vss.n4176 vss.n4175 0.0702092
R44157 vss.t373 vss.n4176 0.0702092
R44158 vss.n3786 vss.n3784 0.0702092
R44159 vss.n3784 vss.t867 0.0702092
R44160 vss.n3826 vss.n3814 0.0702092
R44161 vss.t1284 vss.n3812 0.0702092
R44162 vss.t1284 vss.n3826 0.0702092
R44163 vss.n3823 vss.n3812 0.0702092
R44164 vss.n4157 vss.n4156 0.0702092
R44165 vss.n4156 vss.t525 0.0702092
R44166 vss.n4159 vss.n3809 0.0702092
R44167 vss.t524 vss.n3809 0.0702092
R44168 vss.n4165 vss.n4164 0.0702092
R44169 vss.n4165 vss.t1193 0.0702092
R44170 vss.n4162 vss.n4161 0.0702092
R44171 vss.n4161 vss.t1193 0.0702092
R44172 vss.n4170 vss.n4169 0.0702092
R44173 vss.n4169 vss.t524 0.0702092
R44174 vss.n4155 vss.n3804 0.0702092
R44175 vss.t525 vss.n4155 0.0702092
R44176 vss.n4153 vss.n3839 0.0702092
R44177 vss.t962 vss.n4152 0.0702092
R44178 vss.n4153 vss.t962 0.0702092
R44179 vss.n4152 vss.n4151 0.0702092
R44180 vss.n4145 vss.n3841 0.0702092
R44181 vss.n3841 vss.t1151 0.0702092
R44182 vss.n4143 vss.n4142 0.0702092
R44183 vss.n4142 vss.t426 0.0702092
R44184 vss.n3864 vss.n3858 0.0702092
R44185 vss.t428 vss.n3858 0.0702092
R44186 vss.n4138 vss.n4137 0.0702092
R44187 vss.n4137 vss.t428 0.0702092
R44188 vss.n4141 vss.n4140 0.0702092
R44189 vss.t426 vss.n4141 0.0702092
R44190 vss.n3842 vss.n3840 0.0702092
R44191 vss.n3840 vss.t1151 0.0702092
R44192 vss.n3869 vss.n3862 0.0702092
R44193 vss.t423 vss.n3861 0.0702092
R44194 vss.t423 vss.n3869 0.0702092
R44195 vss.n3866 vss.n3861 0.0702092
R44196 vss.n3943 vss.n3942 0.0702092
R44197 vss.t1194 vss.n3943 0.0702092
R44198 vss.n4129 vss.n4128 0.0702092
R44199 vss.n4128 vss.t1196 0.0702092
R44200 vss.n4131 vss.n3871 0.0702092
R44201 vss.n3871 vss.t1428 0.0702092
R44202 vss.n3872 vss.n3870 0.0702092
R44203 vss.n3870 vss.t1428 0.0702092
R44204 vss.n4127 vss.n4126 0.0702092
R44205 vss.t1196 vss.n4127 0.0702092
R44206 vss.n3945 vss.n3944 0.0702092
R44207 vss.n3944 vss.t1194 0.0702092
R44208 vss.n3938 vss.n3937 0.0702092
R44209 vss.n3939 vss.t849 0.0702092
R44210 vss.t849 vss.n3938 0.0702092
R44211 vss.n3940 vss.n3939 0.0702092
R44212 vss.n3932 vss.n3893 0.0702092
R44213 vss.n3893 vss.t448 0.0702092
R44214 vss.n3930 vss.n3929 0.0702092
R44215 vss.n3929 vss.t117 0.0702092
R44216 vss.n3915 vss.n3909 0.0702092
R44217 vss.t119 vss.n3909 0.0702092
R44218 vss.n3925 vss.n3924 0.0702092
R44219 vss.n3924 vss.t119 0.0702092
R44220 vss.n3928 vss.n3927 0.0702092
R44221 vss.t117 vss.n3928 0.0702092
R44222 vss.n3894 vss.n3892 0.0702092
R44223 vss.n3892 vss.t448 0.0702092
R44224 vss.n3920 vss.n3913 0.0702092
R44225 vss.t629 vss.n3912 0.0702092
R44226 vss.t629 vss.n3920 0.0702092
R44227 vss.n3917 vss.n3912 0.0702092
R44228 vss.n5824 vss.n5823 0.0702092
R44229 vss.n5823 vss.t329 0.0702092
R44230 vss.n5826 vss.n3550 0.0702092
R44231 vss.t331 vss.n3550 0.0702092
R44232 vss.n5832 vss.n5831 0.0702092
R44233 vss.n5832 vss.t1306 0.0702092
R44234 vss.n5829 vss.n5828 0.0702092
R44235 vss.n5828 vss.t1306 0.0702092
R44236 vss.n5837 vss.n5836 0.0702092
R44237 vss.n5836 vss.t331 0.0702092
R44238 vss.n5822 vss.n3545 0.0702092
R44239 vss.t329 vss.n5822 0.0702092
R44240 vss.n5820 vss.n3562 0.0702092
R44241 vss.t51 vss.n5819 0.0702092
R44242 vss.n5820 vss.t51 0.0702092
R44243 vss.n5819 vss.n5818 0.0702092
R44244 vss.n5812 vss.n3564 0.0702092
R44245 vss.n3564 vss.t1475 0.0702092
R44246 vss.n5810 vss.n5809 0.0702092
R44247 vss.n5809 vss.t738 0.0702092
R44248 vss.n3618 vss.n3582 0.0702092
R44249 vss.t740 vss.n3582 0.0702092
R44250 vss.n5805 vss.n5804 0.0702092
R44251 vss.n5804 vss.t740 0.0702092
R44252 vss.n5808 vss.n5807 0.0702092
R44253 vss.t738 vss.n5808 0.0702092
R44254 vss.n3565 vss.n3563 0.0702092
R44255 vss.n3563 vss.t1475 0.0702092
R44256 vss.n3616 vss.n3613 0.0702092
R44257 vss.n3615 vss.t1093 0.0702092
R44258 vss.n3613 vss.t1093 0.0702092
R44259 vss.n3620 vss.n3615 0.0702092
R44260 vss.n5671 vss.n5670 0.0702092
R44261 vss.t1136 vss.n5671 0.0702092
R44262 vss.n5796 vss.n5795 0.0702092
R44263 vss.n5795 vss.t1135 0.0702092
R44264 vss.n5798 vss.n3585 0.0702092
R44265 vss.n3585 vss.t906 0.0702092
R44266 vss.n3586 vss.n3584 0.0702092
R44267 vss.n3584 vss.t906 0.0702092
R44268 vss.n5794 vss.n5793 0.0702092
R44269 vss.t1135 vss.n5794 0.0702092
R44270 vss.n5672 vss.n3598 0.0702092
R44271 vss.n5672 vss.t1136 0.0702092
R44272 vss.n5674 vss.n5662 0.0702092
R44273 vss.t1003 vss.n5660 0.0702092
R44274 vss.t1003 vss.n5674 0.0702092
R44275 vss.n5668 vss.n5660 0.0702092
R44276 vss.n5679 vss.n5678 0.0702092
R44277 vss.t63 vss.n5679 0.0702092
R44278 vss.n5684 vss.n5683 0.0702092
R44279 vss.n5683 vss.t1513 0.0702092
R44280 vss.n5686 vss.n3609 0.0702092
R44281 vss.t1515 vss.n3609 0.0702092
R44282 vss.n5737 vss.n5736 0.0702092
R44283 vss.n5736 vss.t1515 0.0702092
R44284 vss.n5682 vss.n3604 0.0702092
R44285 vss.t1513 vss.n5682 0.0702092
R44286 vss.n5680 vss.n5658 0.0702092
R44287 vss.n5680 vss.t63 0.0702092
R44288 vss.n5691 vss.n5647 0.0702092
R44289 vss.t688 vss.n5646 0.0702092
R44290 vss.t688 vss.n5691 0.0702092
R44291 vss.n5688 vss.n5646 0.0702092
R44292 vss.n5717 vss.n5716 0.0702092
R44293 vss.n5716 vss.t884 0.0702092
R44294 vss.n5720 vss.n5719 0.0702092
R44295 vss.t513 vss.n5720 0.0702092
R44296 vss.n5728 vss.n5727 0.0702092
R44297 vss.n5727 vss.t515 0.0702092
R44298 vss.n5730 vss.n5693 0.0702092
R44299 vss.n5693 vss.t1427 0.0702092
R44300 vss.n5694 vss.n5692 0.0702092
R44301 vss.n5692 vss.t1427 0.0702092
R44302 vss.n5726 vss.n5725 0.0702092
R44303 vss.t515 vss.n5726 0.0702092
R44304 vss.n5722 vss.n5721 0.0702092
R44305 vss.n5721 vss.t513 0.0702092
R44306 vss.n5715 vss.n5714 0.0702092
R44307 vss.t884 vss.n5715 0.0702092
R44308 vss.n9970 vss.n9969 0.0702092
R44309 vss.t1322 vss.n9970 0.0702092
R44310 vss.n9975 vss.n9974 0.0702092
R44311 vss.n9974 vss.t518 0.0702092
R44312 vss.n9977 vss.n2637 0.0702092
R44313 vss.t520 vss.n2637 0.0702092
R44314 vss.n9983 vss.n9982 0.0702092
R44315 vss.n9983 vss.t277 0.0702092
R44316 vss.n9980 vss.n9979 0.0702092
R44317 vss.n9979 vss.t277 0.0702092
R44318 vss.n9988 vss.n9987 0.0702092
R44319 vss.n9987 vss.t520 0.0702092
R44320 vss.n9973 vss.n2632 0.0702092
R44321 vss.t518 vss.n9973 0.0702092
R44322 vss.n9971 vss.n9966 0.0702092
R44323 vss.n9971 vss.t1322 0.0702092
R44324 vss.n2666 vss.n2665 0.0702092
R44325 vss.n2665 vss.t1075 0.0702092
R44326 vss.n2669 vss.n2668 0.0702092
R44327 vss.t405 vss.n2669 0.0702092
R44328 vss.n2679 vss.n2678 0.0702092
R44329 vss.n2678 vss.t407 0.0702092
R44330 vss.n2681 vss.n2641 0.0702092
R44331 vss.n2641 vss.t450 0.0702092
R44332 vss.n2642 vss.n2640 0.0702092
R44333 vss.n2640 vss.t450 0.0702092
R44334 vss.n2677 vss.n2676 0.0702092
R44335 vss.t407 vss.n2677 0.0702092
R44336 vss.n2671 vss.n2670 0.0702092
R44337 vss.n2670 vss.t405 0.0702092
R44338 vss.n2664 vss.n2663 0.0702092
R44339 vss.t1075 vss.n2664 0.0702092
R44340 vss.n3403 vss.n3402 0.0702092
R44341 vss.t3 vss.n3403 0.0702092
R44342 vss.n3408 vss.n3407 0.0702092
R44343 vss.n3407 vss.t647 0.0702092
R44344 vss.n3410 vss.n3387 0.0702092
R44345 vss.t649 vss.n3387 0.0702092
R44346 vss.n3416 vss.n3415 0.0702092
R44347 vss.n3416 vss.t495 0.0702092
R44348 vss.n3413 vss.n3412 0.0702092
R44349 vss.n3412 vss.t495 0.0702092
R44350 vss.n3421 vss.n3420 0.0702092
R44351 vss.n3420 vss.t649 0.0702092
R44352 vss.n3406 vss.n3382 0.0702092
R44353 vss.t647 vss.n3406 0.0702092
R44354 vss.n3404 vss.n3399 0.0702092
R44355 vss.n3404 vss.t3 0.0702092
R44356 vss.n4000 vss.n3999 0.0702092
R44357 vss.t391 vss.n4000 0.0702092
R44358 vss.n4005 vss.n4004 0.0702092
R44359 vss.n4004 vss.t431 0.0702092
R44360 vss.n4007 vss.n3984 0.0702092
R44361 vss.t433 vss.n3984 0.0702092
R44362 vss.n4013 vss.n4012 0.0702092
R44363 vss.n4013 vss.t840 0.0702092
R44364 vss.n4010 vss.n4009 0.0702092
R44365 vss.n4009 vss.t840 0.0702092
R44366 vss.n4018 vss.n4017 0.0702092
R44367 vss.n4017 vss.t433 0.0702092
R44368 vss.n4003 vss.n3979 0.0702092
R44369 vss.t431 vss.n4003 0.0702092
R44370 vss.n4001 vss.n3996 0.0702092
R44371 vss.n4001 vss.t391 0.0702092
R44372 vss.n4267 vss.n4266 0.0702092
R44373 vss.t486 vss.n4267 0.0702092
R44374 vss.n4272 vss.n4271 0.0702092
R44375 vss.n4271 vss.t1452 0.0702092
R44376 vss.n4274 vss.n4251 0.0702092
R44377 vss.t1451 vss.n4251 0.0702092
R44378 vss.n4280 vss.n4279 0.0702092
R44379 vss.n4280 vss.t1253 0.0702092
R44380 vss.n4277 vss.n4276 0.0702092
R44381 vss.n4276 vss.t1253 0.0702092
R44382 vss.n4285 vss.n4284 0.0702092
R44383 vss.n4284 vss.t1451 0.0702092
R44384 vss.n4270 vss.n4246 0.0702092
R44385 vss.t1452 vss.n4270 0.0702092
R44386 vss.n4268 vss.n4263 0.0702092
R44387 vss.n4268 vss.t486 0.0702092
R44388 vss.n5921 vss.n5920 0.0702092
R44389 vss.n5921 vss.t236 0.0702092
R44390 vss.t478 vss.n5910 0.0702092
R44391 vss.n5914 vss.t1064 0.0702092
R44392 vss.t1066 vss.n5927 0.0702092
R44393 vss.n5923 vss.t236 0.0702092
R44394 vss.n5929 vss.n5928 0.0702092
R44395 vss.n5928 vss.t1066 0.0702092
R44396 vss.n5913 vss.n5890 0.0702092
R44397 vss.t1064 vss.n5913 0.0702092
R44398 vss.n5911 vss.n5906 0.0702092
R44399 vss.n5911 vss.t478 0.0702092
R44400 vss.n5910 vss.n5909 0.0702092
R44401 vss.n5915 vss.n5914 0.0702092
R44402 vss.n5927 vss.n5926 0.0702092
R44403 vss.n5924 vss.n5923 0.0702092
R44404 vss.n9926 vss.n2710 0.0702092
R44405 vss.n2710 vss.t339 0.0702092
R44406 vss.n2711 vss.n2709 0.0702092
R44407 vss.n2709 vss.t339 0.0702092
R44408 vss.n3286 vss.n3280 0.0702092
R44409 vss.n3286 vss.t1387 0.0702092
R44410 vss.n3298 vss.n3297 0.0702092
R44411 vss.t49 vss.n3298 0.0702092
R44412 vss.n3305 vss.n3304 0.0702092
R44413 vss.n3304 vss.t1197 0.0702092
R44414 vss.n3288 vss.n3264 0.0702092
R44415 vss.t1199 vss.n3288 0.0702092
R44416 vss.n3285 vss.n3284 0.0702092
R44417 vss.t1387 vss.n3285 0.0702092
R44418 vss.n3290 vss.n3289 0.0702092
R44419 vss.n3289 vss.t1199 0.0702092
R44420 vss.n3303 vss.n3302 0.0702092
R44421 vss.t1197 vss.n3303 0.0702092
R44422 vss.n3300 vss.n3299 0.0702092
R44423 vss.n3299 vss.t49 0.0702092
R44424 vss.n9708 vss.n9702 0.0702092
R44425 vss.n9708 vss.t1398 0.0702092
R44426 vss.n9719 vss.n9718 0.0702092
R44427 vss.t39 vss.n9719 0.0702092
R44428 vss.n9727 vss.n9726 0.0702092
R44429 vss.n9726 vss.t1445 0.0702092
R44430 vss.n9710 vss.n9686 0.0702092
R44431 vss.t1444 vss.n9710 0.0702092
R44432 vss.n9707 vss.n9706 0.0702092
R44433 vss.t1398 vss.n9707 0.0702092
R44434 vss.n9712 vss.n9711 0.0702092
R44435 vss.n9711 vss.t1444 0.0702092
R44436 vss.n9725 vss.n9724 0.0702092
R44437 vss.t1445 vss.n9725 0.0702092
R44438 vss.n9722 vss.n9721 0.0702092
R44439 vss.n9721 vss.t39 0.0702092
R44440 vss.n9892 vss.n2745 0.0702092
R44441 vss.n2745 vss.t322 0.0702092
R44442 vss.n9879 vss.n9878 0.0702092
R44443 vss.n9878 vss.t217 0.0702092
R44444 vss.n2763 vss.n2761 0.0702092
R44445 vss.t130 vss.n2761 0.0702092
R44446 vss.n9890 vss.n9889 0.0702092
R44447 vss.n9889 vss.t129 0.0702092
R44448 vss.n2746 vss.n2744 0.0702092
R44449 vss.n2744 vss.t322 0.0702092
R44450 vss.n9888 vss.n9887 0.0702092
R44451 vss.t129 vss.n9888 0.0702092
R44452 vss.n9885 vss.n9884 0.0702092
R44453 vss.n9884 vss.t130 0.0702092
R44454 vss.n2766 vss.n2765 0.0702092
R44455 vss.n2766 vss.t217 0.0702092
R44456 vss.n9034 vss.n7269 0.0702092
R44457 vss.n7269 vss.t1382 0.0702092
R44458 vss.n7270 vss.n7268 0.0702092
R44459 vss.n7268 vss.t1382 0.0702092
R44460 vss.n8083 vss.n8082 0.0702092
R44461 vss.n8082 vss.t537 0.0702092
R44462 vss.n8094 vss.n8093 0.0702092
R44463 vss.n8093 vss.t183 0.0702092
R44464 vss.n8086 vss.n8085 0.0702092
R44465 vss.t182 vss.n8086 0.0702092
R44466 vss.n8081 vss.n8080 0.0702092
R44467 vss.t537 vss.n8081 0.0702092
R44468 vss.n8088 vss.n8087 0.0702092
R44469 vss.n8087 vss.t182 0.0702092
R44470 vss.n8092 vss.n8091 0.0702092
R44471 vss.t183 vss.n8092 0.0702092
R44472 vss.n8096 vss.n8054 0.0702092
R44473 vss.n8054 vss.t960 0.0702092
R44474 vss.n8055 vss.n8053 0.0702092
R44475 vss.n8053 vss.t960 0.0702092
R44476 vss.n8170 vss.n8101 0.0702092
R44477 vss.n8101 vss.t863 0.0702092
R44478 vss.n8168 vss.n8167 0.0702092
R44479 vss.n8167 vss.t1059 0.0702092
R44480 vss.n8160 vss.n8159 0.0702092
R44481 vss.t1058 vss.n8160 0.0702092
R44482 vss.n8162 vss.n8161 0.0702092
R44483 vss.n8161 vss.t1058 0.0702092
R44484 vss.n8166 vss.n8165 0.0702092
R44485 vss.t1059 vss.n8166 0.0702092
R44486 vss.n8102 vss.n8100 0.0702092
R44487 vss.n8100 vss.t863 0.0702092
R44488 vss.n8954 vss.n7490 0.0702092
R44489 vss.n8954 vss.t1173 0.0702092
R44490 vss.n8965 vss.n8964 0.0702092
R44491 vss.t1505 vss.n8965 0.0702092
R44492 vss.n8972 vss.n8971 0.0702092
R44493 vss.n8971 vss.t262 0.0702092
R44494 vss.n8956 vss.n7474 0.0702092
R44495 vss.t264 vss.n8956 0.0702092
R44496 vss.n8953 vss.n8952 0.0702092
R44497 vss.t1173 vss.n8953 0.0702092
R44498 vss.n8958 vss.n8957 0.0702092
R44499 vss.n8957 vss.t264 0.0702092
R44500 vss.n8970 vss.n8969 0.0702092
R44501 vss.t262 vss.n8970 0.0702092
R44502 vss.n8967 vss.n8966 0.0702092
R44503 vss.n8966 vss.t1505 0.0702092
R44504 vss.n8898 vss.n7541 0.0702092
R44505 vss.n7541 vss.t1517 0.0702092
R44506 vss.n8885 vss.n8884 0.0702092
R44507 vss.n8884 vss.t572 0.0702092
R44508 vss.n8879 vss.n8877 0.0702092
R44509 vss.t195 vss.n8877 0.0702092
R44510 vss.n8896 vss.n8895 0.0702092
R44511 vss.n8895 vss.t194 0.0702092
R44512 vss.n7542 vss.n7540 0.0702092
R44513 vss.n7540 vss.t1517 0.0702092
R44514 vss.n8894 vss.n8893 0.0702092
R44515 vss.t194 vss.n8894 0.0702092
R44516 vss.n8891 vss.n8890 0.0702092
R44517 vss.n8890 vss.t195 0.0702092
R44518 vss.n8882 vss.n8881 0.0702092
R44519 vss.n8882 vss.t572 0.0702092
R44520 vss.n8835 vss.n7679 0.0702092
R44521 vss.n8835 vss.t786 0.0702092
R44522 vss.n8846 vss.n8845 0.0702092
R44523 vss.t1073 vss.n8846 0.0702092
R44524 vss.n8853 vss.n8852 0.0702092
R44525 vss.n8852 vss.t784 0.0702092
R44526 vss.n8837 vss.n7663 0.0702092
R44527 vss.t783 vss.n8837 0.0702092
R44528 vss.n8834 vss.n8833 0.0702092
R44529 vss.t786 vss.n8834 0.0702092
R44530 vss.n8839 vss.n8838 0.0702092
R44531 vss.n8838 vss.t783 0.0702092
R44532 vss.n8851 vss.n8850 0.0702092
R44533 vss.t784 vss.n8851 0.0702092
R44534 vss.n8848 vss.n8847 0.0702092
R44535 vss.n8847 vss.t1073 0.0702092
R44536 vss.n8779 vss.n7684 0.0702092
R44537 vss.n7684 vss.t1134 0.0702092
R44538 vss.n8766 vss.n8765 0.0702092
R44539 vss.n8765 vss.t1376 0.0702092
R44540 vss.n8760 vss.n8758 0.0702092
R44541 vss.t1535 vss.n8758 0.0702092
R44542 vss.n8777 vss.n8776 0.0702092
R44543 vss.n8776 vss.t1534 0.0702092
R44544 vss.n7685 vss.n7683 0.0702092
R44545 vss.n7683 vss.t1134 0.0702092
R44546 vss.n8775 vss.n8774 0.0702092
R44547 vss.t1534 vss.n8775 0.0702092
R44548 vss.n8772 vss.n8771 0.0702092
R44549 vss.n8771 vss.t1535 0.0702092
R44550 vss.n8763 vss.n8762 0.0702092
R44551 vss.n8763 vss.t1376 0.0702092
R44552 vss.n8716 vss.n7866 0.0702092
R44553 vss.n8716 vss.t1298 0.0702092
R44554 vss.n8727 vss.n8726 0.0702092
R44555 vss.t611 vss.n8727 0.0702092
R44556 vss.n8734 vss.n8733 0.0702092
R44557 vss.n8733 vss.t1296 0.0702092
R44558 vss.n8718 vss.n7850 0.0702092
R44559 vss.t1295 vss.n8718 0.0702092
R44560 vss.n8715 vss.n8714 0.0702092
R44561 vss.t1298 vss.n8715 0.0702092
R44562 vss.n8720 vss.n8719 0.0702092
R44563 vss.n8719 vss.t1295 0.0702092
R44564 vss.n8732 vss.n8731 0.0702092
R44565 vss.t1296 vss.n8732 0.0702092
R44566 vss.n8729 vss.n8728 0.0702092
R44567 vss.n8728 vss.t611 0.0702092
R44568 vss.n9003 vss.n7301 0.0702092
R44569 vss.n7301 vss.t561 0.0702092
R44570 vss.n8990 vss.n8989 0.0702092
R44571 vss.n8989 vss.t383 0.0702092
R44572 vss.n7319 vss.n7317 0.0702092
R44573 vss.t412 vss.n7317 0.0702092
R44574 vss.n9001 vss.n9000 0.0702092
R44575 vss.n9000 vss.t411 0.0702092
R44576 vss.n7302 vss.n7300 0.0702092
R44577 vss.n7300 vss.t561 0.0702092
R44578 vss.n8999 vss.n8998 0.0702092
R44579 vss.t411 vss.n8999 0.0702092
R44580 vss.n8996 vss.n8995 0.0702092
R44581 vss.n8995 vss.t412 0.0702092
R44582 vss.n7322 vss.n7321 0.0702092
R44583 vss.n7322 vss.t383 0.0702092
R44584 vss.n8225 vss.n8009 0.0702092
R44585 vss.n8225 vss.t440 0.0702092
R44586 vss.n8236 vss.n8235 0.0702092
R44587 vss.t1507 vss.n8236 0.0702092
R44588 vss.n8243 vss.n8242 0.0702092
R44589 vss.n8242 vss.t559 0.0702092
R44590 vss.n8227 vss.n7993 0.0702092
R44591 vss.t558 vss.n8227 0.0702092
R44592 vss.n8224 vss.n8223 0.0702092
R44593 vss.t440 vss.n8224 0.0702092
R44594 vss.n8229 vss.n8228 0.0702092
R44595 vss.n8228 vss.t558 0.0702092
R44596 vss.n8241 vss.n8240 0.0702092
R44597 vss.t559 vss.n8241 0.0702092
R44598 vss.n8238 vss.n8237 0.0702092
R44599 vss.n8237 vss.t1507 0.0702092
R44600 vss.n8215 vss.n8176 0.0702092
R44601 vss.n8176 vss.t756 0.0702092
R44602 vss.n8202 vss.n8201 0.0702092
R44603 vss.n8201 vss.t1346 0.0702092
R44604 vss.n8196 vss.n8194 0.0702092
R44605 vss.t371 vss.n8194 0.0702092
R44606 vss.n8213 vss.n8212 0.0702092
R44607 vss.n8212 vss.t370 0.0702092
R44608 vss.n8177 vss.n8175 0.0702092
R44609 vss.n8175 vss.t756 0.0702092
R44610 vss.n8211 vss.n8210 0.0702092
R44611 vss.t370 vss.n8211 0.0702092
R44612 vss.n8208 vss.n8207 0.0702092
R44613 vss.n8207 vss.t371 0.0702092
R44614 vss.n8199 vss.n8198 0.0702092
R44615 vss.n8199 vss.t1346 0.0702092
R44616 vss.n7931 vss.n7926 0.0702092
R44617 vss.n7931 vss.t241 0.0702092
R44618 vss.n7942 vss.n7941 0.0702092
R44619 vss.t484 vss.n7942 0.0702092
R44620 vss.n7949 vss.n7948 0.0702092
R44621 vss.n7948 vss.t651 0.0702092
R44622 vss.n7933 vss.n7910 0.0702092
R44623 vss.t650 vss.n7933 0.0702092
R44624 vss.n7930 vss.n7929 0.0702092
R44625 vss.t241 vss.n7930 0.0702092
R44626 vss.n7935 vss.n7934 0.0702092
R44627 vss.n7934 vss.t650 0.0702092
R44628 vss.n7947 vss.n7946 0.0702092
R44629 vss.t651 vss.n7947 0.0702092
R44630 vss.n7944 vss.n7943 0.0702092
R44631 vss.n7943 vss.t484 0.0702092
R44632 vss.n7790 vss.n7785 0.0702092
R44633 vss.n7790 vss.t165 0.0702092
R44634 vss.n7801 vss.n7800 0.0702092
R44635 vss.t496 vss.n7801 0.0702092
R44636 vss.n7808 vss.n7807 0.0702092
R44637 vss.n7807 vss.t163 0.0702092
R44638 vss.n7792 vss.n7769 0.0702092
R44639 vss.t162 vss.n7792 0.0702092
R44640 vss.n7789 vss.n7788 0.0702092
R44641 vss.t165 vss.n7789 0.0702092
R44642 vss.n7794 vss.n7793 0.0702092
R44643 vss.n7793 vss.t162 0.0702092
R44644 vss.n7806 vss.n7805 0.0702092
R44645 vss.t163 vss.n7806 0.0702092
R44646 vss.n7803 vss.n7802 0.0702092
R44647 vss.n7802 vss.t496 0.0702092
R44648 vss.n7710 vss.n7705 0.0702092
R44649 vss.n7710 vss.t425 0.0702092
R44650 vss.n7721 vss.n7720 0.0702092
R44651 vss.t5 vss.n7721 0.0702092
R44652 vss.n7728 vss.n7727 0.0702092
R44653 vss.n7727 vss.t223 0.0702092
R44654 vss.n7712 vss.n7689 0.0702092
R44655 vss.t225 vss.n7712 0.0702092
R44656 vss.n7709 vss.n7708 0.0702092
R44657 vss.t425 vss.n7709 0.0702092
R44658 vss.n7714 vss.n7713 0.0702092
R44659 vss.n7713 vss.t225 0.0702092
R44660 vss.n7726 vss.n7725 0.0702092
R44661 vss.t223 vss.n7726 0.0702092
R44662 vss.n7723 vss.n7722 0.0702092
R44663 vss.n7722 vss.t5 0.0702092
R44664 vss.n8825 vss.n8786 0.0702092
R44665 vss.n8786 vss.t1013 0.0702092
R44666 vss.n8812 vss.n8811 0.0702092
R44667 vss.n8811 vss.t205 0.0702092
R44668 vss.n8806 vss.n8804 0.0702092
R44669 vss.t1011 vss.n8804 0.0702092
R44670 vss.n8823 vss.n8822 0.0702092
R44671 vss.n8822 vss.t1010 0.0702092
R44672 vss.n8787 vss.n8785 0.0702092
R44673 vss.n8785 vss.t1013 0.0702092
R44674 vss.n8821 vss.n8820 0.0702092
R44675 vss.t1010 vss.n8821 0.0702092
R44676 vss.n8818 vss.n8817 0.0702092
R44677 vss.n8817 vss.t1011 0.0702092
R44678 vss.n8809 vss.n8808 0.0702092
R44679 vss.n8809 vss.t205 0.0702092
R44680 vss.n7567 vss.n7562 0.0702092
R44681 vss.n7567 vss.t1133 0.0702092
R44682 vss.n7578 vss.n7577 0.0702092
R44683 vss.t633 vss.n7578 0.0702092
R44684 vss.n7585 vss.n7584 0.0702092
R44685 vss.n7584 vss.t836 0.0702092
R44686 vss.n7569 vss.n7546 0.0702092
R44687 vss.t838 vss.n7569 0.0702092
R44688 vss.n7566 vss.n7565 0.0702092
R44689 vss.t1133 vss.n7566 0.0702092
R44690 vss.n7571 vss.n7570 0.0702092
R44691 vss.n7570 vss.t838 0.0702092
R44692 vss.n7583 vss.n7582 0.0702092
R44693 vss.t836 vss.n7583 0.0702092
R44694 vss.n7580 vss.n7579 0.0702092
R44695 vss.n7579 vss.t633 0.0702092
R44696 vss.n8944 vss.n8905 0.0702092
R44697 vss.n8905 vss.t361 0.0702092
R44698 vss.n8931 vss.n8930 0.0702092
R44699 vss.n8930 vss.t9 0.0702092
R44700 vss.n8925 vss.n8923 0.0702092
R44701 vss.t310 vss.n8923 0.0702092
R44702 vss.n8942 vss.n8941 0.0702092
R44703 vss.n8941 vss.t312 0.0702092
R44704 vss.n8906 vss.n8904 0.0702092
R44705 vss.n8904 vss.t361 0.0702092
R44706 vss.n8940 vss.n8939 0.0702092
R44707 vss.t312 vss.n8940 0.0702092
R44708 vss.n8937 vss.n8936 0.0702092
R44709 vss.n8936 vss.t310 0.0702092
R44710 vss.n8928 vss.n8927 0.0702092
R44711 vss.n8928 vss.t9 0.0702092
R44712 vss.n7532 vss.n7492 0.0702092
R44713 vss.n7492 vss.t662 0.0702092
R44714 vss.n7519 vss.n7518 0.0702092
R44715 vss.n7518 vss.t215 0.0702092
R44716 vss.n7513 vss.n7511 0.0702092
R44717 vss.t1468 vss.n7511 0.0702092
R44718 vss.n7530 vss.n7529 0.0702092
R44719 vss.n7529 vss.t1467 0.0702092
R44720 vss.n7493 vss.n7491 0.0702092
R44721 vss.n7491 vss.t662 0.0702092
R44722 vss.n7528 vss.n7527 0.0702092
R44723 vss.t1467 vss.n7528 0.0702092
R44724 vss.n7525 vss.n7524 0.0702092
R44725 vss.n7524 vss.t1468 0.0702092
R44726 vss.n7516 vss.n7515 0.0702092
R44727 vss.n7516 vss.t215 0.0702092
R44728 vss.n616 vss.n614 0.0702092
R44729 vss.n614 vss.t132 0.0702092
R44730 vss.n634 vss.t23 0.0702092
R44731 vss.t136 vss.n638 0.0702092
R44732 vss.n652 vss.t138 0.0702092
R44733 vss.n615 vss.t132 0.0702092
R44734 vss.n647 vss.n646 0.0702092
R44735 vss.n647 vss.t138 0.0702092
R44736 vss.n640 vss.n639 0.0702092
R44737 vss.n639 vss.t136 0.0702092
R44738 vss.n633 vss.n632 0.0702092
R44739 vss.t23 vss.n633 0.0702092
R44740 vss.n635 vss.n634 0.0702092
R44741 vss.n638 vss.n637 0.0702092
R44742 vss.n653 vss.n652 0.0702092
R44743 vss.n655 vss.n615 0.0702092
R44744 vss.n470 vss.n459 0.0702092
R44745 vss.t1275 vss.n459 0.0702092
R44746 vss.n14153 vss.n14152 0.0702092
R44747 vss.t1275 vss.n14153 0.0702092
R44748 vss.n14159 vss.n14158 0.0702092
R44749 vss.n14158 vss.t293 0.0702092
R44750 vss.n14172 vss.n435 0.0702092
R44751 vss.n435 vss.t880 0.0702092
R44752 vss.n14170 vss.n14169 0.0702092
R44753 vss.n14169 vss.t973 0.0702092
R44754 vss.n14162 vss.n14161 0.0702092
R44755 vss.t972 vss.n14162 0.0702092
R44756 vss.n14157 vss.n14156 0.0702092
R44757 vss.t293 vss.n14157 0.0702092
R44758 vss.n14164 vss.n14163 0.0702092
R44759 vss.n14163 vss.t972 0.0702092
R44760 vss.n14168 vss.n14167 0.0702092
R44761 vss.t973 vss.n14168 0.0702092
R44762 vss.n436 vss.n434 0.0702092
R44763 vss.n434 vss.t880 0.0702092
R44764 vss.n14065 vss.n14064 0.0702092
R44765 vss.n14064 vss.t734 0.0702092
R44766 vss.n14074 vss.n14073 0.0702092
R44767 vss.n14073 vss.t920 0.0702092
R44768 vss.n14077 vss.n14076 0.0702092
R44769 vss.n14077 vss.t921 0.0702092
R44770 vss.n14080 vss.n14079 0.0702092
R44771 vss.n14079 vss.t35 0.0702092
R44772 vss.n14070 vss.t734 0.0702092
R44773 vss.t920 vss.n14072 0.0702092
R44774 vss.n14085 vss.t921 0.0702092
R44775 vss.n14083 vss.t35 0.0702092
R44776 vss.n14083 vss.n14082 0.0702092
R44777 vss.n14086 vss.n14085 0.0702092
R44778 vss.n14072 vss.n476 0.0702092
R44779 vss.n14070 vss.n14069 0.0702092
R44780 vss.n10120 vss.n10119 0.0702092
R44781 vss.n10119 vss.t828 0.0702092
R44782 vss.n10129 vss.n10128 0.0702092
R44783 vss.n10128 vss.t1305 0.0702092
R44784 vss.n10132 vss.n10131 0.0702092
R44785 vss.n10132 vss.t1303 0.0702092
R44786 vss.n10135 vss.n10134 0.0702092
R44787 vss.n10134 vss.t468 0.0702092
R44788 vss.n10125 vss.t828 0.0702092
R44789 vss.t1305 vss.n10127 0.0702092
R44790 vss.n10140 vss.t1303 0.0702092
R44791 vss.n10138 vss.t468 0.0702092
R44792 vss.n10138 vss.n10137 0.0702092
R44793 vss.n10141 vss.n10140 0.0702092
R44794 vss.n10127 vss.n10103 0.0702092
R44795 vss.n10125 vss.n10124 0.0702092
R44796 vss.n12878 vss.n12877 0.0702092
R44797 vss.n12877 vss.t252 0.0702092
R44798 vss.n12887 vss.n12886 0.0702092
R44799 vss.n12886 vss.t288 0.0702092
R44800 vss.n12890 vss.n12889 0.0702092
R44801 vss.n12890 vss.t286 0.0702092
R44802 vss.n12893 vss.n12892 0.0702092
R44803 vss.n12892 vss.t1479 0.0702092
R44804 vss.n12883 vss.t252 0.0702092
R44805 vss.t288 vss.n12885 0.0702092
R44806 vss.n12898 vss.t286 0.0702092
R44807 vss.n12896 vss.t1479 0.0702092
R44808 vss.n12896 vss.n12895 0.0702092
R44809 vss.n12899 vss.n12898 0.0702092
R44810 vss.n12885 vss.n12861 0.0702092
R44811 vss.n12883 vss.n12882 0.0702092
R44812 vss.n10161 vss.n10160 0.0702092
R44813 vss.n10160 vss.t1230 0.0702092
R44814 vss.n10170 vss.n10169 0.0702092
R44815 vss.n10169 vss.t299 0.0702092
R44816 vss.n10173 vss.n10172 0.0702092
R44817 vss.n10173 vss.t297 0.0702092
R44818 vss.n10176 vss.n10175 0.0702092
R44819 vss.n10175 vss.t385 0.0702092
R44820 vss.n10166 vss.t1230 0.0702092
R44821 vss.t299 vss.n10168 0.0702092
R44822 vss.n10181 vss.t297 0.0702092
R44823 vss.n10179 vss.t385 0.0702092
R44824 vss.n10179 vss.n10178 0.0702092
R44825 vss.n10182 vss.n10181 0.0702092
R44826 vss.n10168 vss.n10144 0.0702092
R44827 vss.n10166 vss.n10165 0.0702092
R44828 vss.n12427 vss.n12426 0.0702092
R44829 vss.n12426 vss.t1450 0.0702092
R44830 vss.n12436 vss.n12435 0.0702092
R44831 vss.n12435 vss.t464 0.0702092
R44832 vss.n12439 vss.n12438 0.0702092
R44833 vss.n12439 vss.t462 0.0702092
R44834 vss.n12442 vss.n12441 0.0702092
R44835 vss.n12441 vss.t7 0.0702092
R44836 vss.n12432 vss.t1450 0.0702092
R44837 vss.t464 vss.n12434 0.0702092
R44838 vss.n12447 vss.t462 0.0702092
R44839 vss.n12445 vss.t7 0.0702092
R44840 vss.n12445 vss.n12444 0.0702092
R44841 vss.n12448 vss.n12447 0.0702092
R44842 vss.n12434 vss.n12410 0.0702092
R44843 vss.n12432 vss.n12431 0.0702092
R44844 vss.n11756 vss.n11755 0.0702092
R44845 vss.n11755 vss.t627 0.0702092
R44846 vss.n11765 vss.n11764 0.0702092
R44847 vss.n11764 vss.t228 0.0702092
R44848 vss.n11768 vss.n11767 0.0702092
R44849 vss.n11768 vss.t226 0.0702092
R44850 vss.n11771 vss.n11770 0.0702092
R44851 vss.n11770 vss.t209 0.0702092
R44852 vss.n11761 vss.t627 0.0702092
R44853 vss.t228 vss.n11763 0.0702092
R44854 vss.n11776 vss.t226 0.0702092
R44855 vss.n11774 vss.t209 0.0702092
R44856 vss.n11774 vss.n11773 0.0702092
R44857 vss.n11777 vss.n11776 0.0702092
R44858 vss.n11763 vss.n11739 0.0702092
R44859 vss.n11761 vss.n11760 0.0702092
R44860 vss.n12472 vss.n12471 0.0702092
R44861 vss.n12471 vss.t369 0.0702092
R44862 vss.n12481 vss.n12480 0.0702092
R44863 vss.n12480 vss.t221 0.0702092
R44864 vss.n12484 vss.n12483 0.0702092
R44865 vss.n12484 vss.t219 0.0702092
R44866 vss.n12487 vss.n12486 0.0702092
R44867 vss.n12486 vss.t1499 0.0702092
R44868 vss.n12477 vss.t369 0.0702092
R44869 vss.t221 vss.n12479 0.0702092
R44870 vss.n12492 vss.t219 0.0702092
R44871 vss.n12490 vss.t1499 0.0702092
R44872 vss.n12490 vss.n12489 0.0702092
R44873 vss.n12493 vss.n12492 0.0702092
R44874 vss.n12479 vss.n12455 0.0702092
R44875 vss.n12477 vss.n12476 0.0702092
R44876 vss.n2348 vss.n2347 0.0702092
R44877 vss.t1287 vss.n2348 0.0702092
R44878 vss.n2345 vss.n2344 0.0702092
R44879 vss.n2344 vss.t981 0.0702092
R44880 vss.n2329 vss.n2328 0.0702092
R44881 vss.n2329 vss.t979 0.0702092
R44882 vss.n2332 vss.n2331 0.0702092
R44883 vss.n2331 vss.t1362 0.0702092
R44884 vss.t1287 vss.n2308 0.0702092
R44885 vss.t981 vss.n2343 0.0702092
R44886 vss.n2337 vss.t979 0.0702092
R44887 vss.n2335 vss.t1362 0.0702092
R44888 vss.n2335 vss.n2334 0.0702092
R44889 vss.n2338 vss.n2337 0.0702092
R44890 vss.n2343 vss.n2342 0.0702092
R44891 vss.n2318 vss.n2308 0.0702092
R44892 vss.n12297 vss.n12296 0.0702092
R44893 vss.n12296 vss.t404 0.0702092
R44894 vss.n12306 vss.n12305 0.0702092
R44895 vss.n12305 vss.t1171 0.0702092
R44896 vss.n12309 vss.n12308 0.0702092
R44897 vss.n12309 vss.t1169 0.0702092
R44898 vss.n12312 vss.n12311 0.0702092
R44899 vss.n12311 vss.t1338 0.0702092
R44900 vss.n12302 vss.t404 0.0702092
R44901 vss.t1171 vss.n12304 0.0702092
R44902 vss.n12317 vss.t1169 0.0702092
R44903 vss.n12315 vss.t1338 0.0702092
R44904 vss.n12315 vss.n12314 0.0702092
R44905 vss.n12318 vss.n12317 0.0702092
R44906 vss.n12304 vss.n12280 0.0702092
R44907 vss.n12302 vss.n12301 0.0702092
R44908 vss.n12342 vss.n12341 0.0702092
R44909 vss.n12341 vss.t243 0.0702092
R44910 vss.n12351 vss.n12350 0.0702092
R44911 vss.n12350 vss.t933 0.0702092
R44912 vss.n12354 vss.n12353 0.0702092
R44913 vss.n12354 vss.t931 0.0702092
R44914 vss.n12357 vss.n12356 0.0702092
R44915 vss.n12356 vss.t1326 0.0702092
R44916 vss.n12347 vss.t243 0.0702092
R44917 vss.t933 vss.n12349 0.0702092
R44918 vss.n12362 vss.t931 0.0702092
R44919 vss.n12360 vss.t1326 0.0702092
R44920 vss.n12360 vss.n12359 0.0702092
R44921 vss.n12363 vss.n12362 0.0702092
R44922 vss.n12349 vss.n12325 0.0702092
R44923 vss.n12347 vss.n12346 0.0702092
R44924 vss.n10238 vss.n10237 0.0702092
R44925 vss.n10237 vss.t1399 0.0702092
R44926 vss.n10247 vss.n10246 0.0702092
R44927 vss.n10246 vss.t439 0.0702092
R44928 vss.n10250 vss.n10249 0.0702092
R44929 vss.n10250 vss.t437 0.0702092
R44930 vss.n10253 vss.n10252 0.0702092
R44931 vss.n10252 vss.t1354 0.0702092
R44932 vss.n10243 vss.t1399 0.0702092
R44933 vss.t439 vss.n10245 0.0702092
R44934 vss.n10258 vss.t437 0.0702092
R44935 vss.n10256 vss.t1354 0.0702092
R44936 vss.n10256 vss.n10255 0.0702092
R44937 vss.n10259 vss.n10258 0.0702092
R44938 vss.n10245 vss.n10221 0.0702092
R44939 vss.n10243 vss.n10242 0.0702092
R44940 vss.n2418 vss.n2417 0.0702092
R44941 vss.n2417 vss.t1422 0.0702092
R44942 vss.n2427 vss.n2426 0.0702092
R44943 vss.n2426 vss.t135 0.0702092
R44944 vss.n2430 vss.n2429 0.0702092
R44945 vss.n2430 vss.t133 0.0702092
R44946 vss.n2433 vss.n2432 0.0702092
R44947 vss.n2432 vss.t389 0.0702092
R44948 vss.n2423 vss.t1422 0.0702092
R44949 vss.t135 vss.n2425 0.0702092
R44950 vss.n2438 vss.t133 0.0702092
R44951 vss.n2436 vss.t389 0.0702092
R44952 vss.n2436 vss.n2435 0.0702092
R44953 vss.n2439 vss.n2438 0.0702092
R44954 vss.n2425 vss.n2401 0.0702092
R44955 vss.n2423 vss.n2422 0.0702092
R44956 vss.n12973 vss.n12972 0.0702092
R44957 vss.t1150 vss.n12973 0.0702092
R44958 vss.n12970 vss.n12969 0.0702092
R44959 vss.n12969 vss.t1165 0.0702092
R44960 vss.n2389 vss.n2388 0.0702092
R44961 vss.n2389 vss.t1166 0.0702092
R44962 vss.n2392 vss.n2391 0.0702092
R44963 vss.n2391 vss.t203 0.0702092
R44964 vss.t1150 vss.n2368 0.0702092
R44965 vss.t1165 vss.n12968 0.0702092
R44966 vss.n2397 vss.t1166 0.0702092
R44967 vss.n2395 vss.t203 0.0702092
R44968 vss.n2395 vss.n2394 0.0702092
R44969 vss.n2398 vss.n2397 0.0702092
R44970 vss.n12968 vss.n12967 0.0702092
R44971 vss.n2378 vss.n2368 0.0702092
R44972 vss.n10046 vss.n10034 0.0702092
R44973 vss.n10046 vss.t318 0.0702092
R44974 vss.n10045 vss.n10044 0.0702092
R44975 vss.t318 vss.n10045 0.0702092
R44976 vss.n10038 vss.n10036 0.0702092
R44977 vss.n10036 vss.t1087 0.0702092
R44978 vss.n10037 vss.t1087 0.0702092
R44979 vss.n10037 vss.n2099 0.0702092
R44980 vss.n2498 vss.n2497 0.0702092
R44981 vss.n2497 vss.t723 0.0702092
R44982 vss.n2507 vss.n2506 0.0702092
R44983 vss.n2506 vss.t61 0.0702092
R44984 vss.n2510 vss.n2509 0.0702092
R44985 vss.n2510 vss.t59 0.0702092
R44986 vss.n2513 vss.n2512 0.0702092
R44987 vss.n2512 vss.t570 0.0702092
R44988 vss.n2503 vss.t723 0.0702092
R44989 vss.t61 vss.n2505 0.0702092
R44990 vss.n2518 vss.t59 0.0702092
R44991 vss.n2516 vss.t570 0.0702092
R44992 vss.n2516 vss.n2515 0.0702092
R44993 vss.n2519 vss.n2518 0.0702092
R44994 vss.n2505 vss.n2480 0.0702092
R44995 vss.n2503 vss.n2502 0.0702092
R44996 vss.n13073 vss.n2121 0.0702092
R44997 vss.n2121 vss.t1149 0.0702092
R44998 vss.n13060 vss.n13059 0.0702092
R44999 vss.n13059 vss.t619 0.0702092
R45000 vss.n2139 vss.n2137 0.0702092
R45001 vss.t855 vss.n2137 0.0702092
R45002 vss.n13071 vss.n13070 0.0702092
R45003 vss.n13070 vss.t854 0.0702092
R45004 vss.n2122 vss.n2120 0.0702092
R45005 vss.n2120 vss.t1149 0.0702092
R45006 vss.n13069 vss.n13068 0.0702092
R45007 vss.t854 vss.n13069 0.0702092
R45008 vss.n13066 vss.n13065 0.0702092
R45009 vss.n13065 vss.t855 0.0702092
R45010 vss.n2142 vss.n2141 0.0702092
R45011 vss.n2142 vss.t619 0.0702092
R45012 vss.n12102 vss.n12101 0.0702092
R45013 vss.t435 vss.n12102 0.0702092
R45014 vss.n12109 vss.n12108 0.0702092
R45015 vss.n12108 vss.t540 0.0702092
R45016 vss.n12112 vss.n12111 0.0702092
R45017 vss.t538 vss.n12112 0.0702092
R45018 vss.n12103 vss.t435 0.0702092
R45019 vss.t540 vss.n12107 0.0702092
R45020 vss.n12115 vss.t538 0.0702092
R45021 vss.n12116 vss.n12115 0.0702092
R45022 vss.n12107 vss.n12106 0.0702092
R45023 vss.n12104 vss.n12103 0.0702092
R45024 vss.n12118 vss.n11827 0.0702092
R45025 vss.t1038 vss.n11827 0.0702092
R45026 vss.n12121 vss.n12120 0.0702092
R45027 vss.t1038 vss.n12121 0.0702092
R45028 vss.n12148 vss.n12147 0.0702092
R45029 vss.n12147 vss.t342 0.0702092
R45030 vss.n12128 vss.n12127 0.0702092
R45031 vss.n12128 vss.t340 0.0702092
R45032 vss.n12131 vss.n12130 0.0702092
R45033 vss.n12130 vss.t799 0.0702092
R45034 vss.t342 vss.n12146 0.0702092
R45035 vss.n12136 vss.t340 0.0702092
R45036 vss.n12134 vss.t799 0.0702092
R45037 vss.n12134 vss.n12133 0.0702092
R45038 vss.n12137 vss.n12136 0.0702092
R45039 vss.n12146 vss.n12145 0.0702092
R45040 vss.n11819 vss.n11808 0.0702092
R45041 vss.t1057 vss.n11808 0.0702092
R45042 vss.n12151 vss.n12150 0.0702092
R45043 vss.t1057 vss.n12151 0.0702092
R45044 vss.n12155 vss.n12154 0.0702092
R45045 vss.t745 vss.n12155 0.0702092
R45046 vss.n12162 vss.n12161 0.0702092
R45047 vss.n12161 vss.t1124 0.0702092
R45048 vss.n12165 vss.n12164 0.0702092
R45049 vss.t1122 vss.n12165 0.0702092
R45050 vss.n12156 vss.t745 0.0702092
R45051 vss.t1124 vss.n12160 0.0702092
R45052 vss.n12168 vss.t1122 0.0702092
R45053 vss.n12169 vss.n12168 0.0702092
R45054 vss.n12160 vss.n12159 0.0702092
R45055 vss.n12157 vss.n12156 0.0702092
R45056 vss.n12171 vss.n11787 0.0702092
R45057 vss.t872 vss.n11787 0.0702092
R45058 vss.n12174 vss.n12173 0.0702092
R45059 vss.t872 vss.n12174 0.0702092
R45060 vss.n12262 vss.n12261 0.0702092
R45061 vss.n12261 vss.t416 0.0702092
R45062 vss.n12265 vss.n12264 0.0702092
R45063 vss.n12265 vss.t414 0.0702092
R45064 vss.n12268 vss.n12267 0.0702092
R45065 vss.n12267 vss.t591 0.0702092
R45066 vss.t416 vss.n12260 0.0702092
R45067 vss.n12273 vss.t414 0.0702092
R45068 vss.n12271 vss.t591 0.0702092
R45069 vss.n12271 vss.n12270 0.0702092
R45070 vss.n12274 vss.n12273 0.0702092
R45071 vss.n12260 vss.n11781 0.0702092
R45072 vss.n12255 vss.n12186 0.0702092
R45073 vss.t1258 vss.n12186 0.0702092
R45074 vss.n12188 vss.n12187 0.0702092
R45075 vss.t1258 vss.n12188 0.0702092
R45076 vss.n12249 vss.n12248 0.0702092
R45077 vss.t455 vss.n12249 0.0702092
R45078 vss.n12246 vss.n12245 0.0702092
R45079 vss.n12245 vss.t93 0.0702092
R45080 vss.n12231 vss.n12230 0.0702092
R45081 vss.n12230 vss.t91 0.0702092
R45082 vss.t455 vss.n12191 0.0702092
R45083 vss.t93 vss.n12244 0.0702092
R45084 vss.n12238 vss.t91 0.0702092
R45085 vss.n12239 vss.n12238 0.0702092
R45086 vss.n12244 vss.n12243 0.0702092
R45087 vss.n12201 vss.n12191 0.0702092
R45088 vss.n12236 vss.n12207 0.0702092
R45089 vss.n12236 vss.t851 0.0702092
R45090 vss.n12235 vss.n12234 0.0702092
R45091 vss.t851 vss.n12235 0.0702092
R45092 vss.n12544 vss.n12543 0.0702092
R45093 vss.n12543 vss.t145 0.0702092
R45094 vss.n12218 vss.n12217 0.0702092
R45095 vss.t143 vss.n12218 0.0702092
R45096 vss.n12212 vss.n12210 0.0702092
R45097 vss.n12210 vss.t71 0.0702092
R45098 vss.t145 vss.n12542 0.0702092
R45099 vss.t143 vss.n12216 0.0702092
R45100 vss.n12211 vss.t71 0.0702092
R45101 vss.n12223 vss.n12211 0.0702092
R45102 vss.n12216 vss.n11735 0.0702092
R45103 vss.n12542 vss.n12541 0.0702092
R45104 vss.n11731 vss.n11720 0.0702092
R45105 vss.t1132 vss.n11720 0.0702092
R45106 vss.n12547 vss.n12546 0.0702092
R45107 vss.t1132 vss.n12547 0.0702092
R45108 vss.n12551 vss.n12550 0.0702092
R45109 vss.t1249 vss.n12551 0.0702092
R45110 vss.n12558 vss.n12557 0.0702092
R45111 vss.n12557 vss.t1402 0.0702092
R45112 vss.n12561 vss.n12560 0.0702092
R45113 vss.t1400 vss.n12561 0.0702092
R45114 vss.n12552 vss.t1249 0.0702092
R45115 vss.t1402 vss.n12556 0.0702092
R45116 vss.n12564 vss.t1400 0.0702092
R45117 vss.n12565 vss.n12564 0.0702092
R45118 vss.n12556 vss.n12555 0.0702092
R45119 vss.n12553 vss.n12552 0.0702092
R45120 vss.n12567 vss.n11700 0.0702092
R45121 vss.t874 vss.n11700 0.0702092
R45122 vss.n12570 vss.n12569 0.0702092
R45123 vss.t874 vss.n12570 0.0702092
R45124 vss.n11692 vss.n11691 0.0702092
R45125 vss.n11692 vss.t638 0.0702092
R45126 vss.n11695 vss.n11694 0.0702092
R45127 vss.n11694 vss.t639 0.0702092
R45128 vss.n11698 vss.n11697 0.0702092
R45129 vss.n11698 vss.t1395 0.0702092
R45130 vss.n12580 vss.t638 0.0702092
R45131 vss.n12578 vss.t639 0.0702092
R45132 vss.n12574 vss.t1395 0.0702092
R45133 vss.n12575 vss.n12574 0.0702092
R45134 vss.n12578 vss.n12577 0.0702092
R45135 vss.n12581 vss.n12580 0.0702092
R45136 vss.n12583 vss.n11625 0.0702092
R45137 vss.n11625 vss.t757 0.0702092
R45138 vss.n11626 vss.n11624 0.0702092
R45139 vss.n11624 vss.t757 0.0702092
R45140 vss.n11684 vss.n11683 0.0702092
R45141 vss.t1184 vss.n11684 0.0702092
R45142 vss.n11681 vss.n11680 0.0702092
R45143 vss.n11680 vss.t831 0.0702092
R45144 vss.n11666 vss.n11665 0.0702092
R45145 vss.n11665 vss.t829 0.0702092
R45146 vss.t1184 vss.n11642 0.0702092
R45147 vss.t831 vss.n11679 0.0702092
R45148 vss.n11673 vss.t829 0.0702092
R45149 vss.n11674 vss.n11673 0.0702092
R45150 vss.n11679 vss.n11678 0.0702092
R45151 vss.n11652 vss.n11642 0.0702092
R45152 vss.n11671 vss.n11658 0.0702092
R45153 vss.n11671 vss.t882 0.0702092
R45154 vss.n11670 vss.n11669 0.0702092
R45155 vss.t882 vss.n11670 0.0702092
R45156 vss.n12842 vss.n12841 0.0702092
R45157 vss.n12841 vss.t284 0.0702092
R45158 vss.n12845 vss.n12844 0.0702092
R45159 vss.n12845 vss.t282 0.0702092
R45160 vss.n12848 vss.n12847 0.0702092
R45161 vss.n12847 vss.t801 0.0702092
R45162 vss.t284 vss.n12840 0.0702092
R45163 vss.n12853 vss.t282 0.0702092
R45164 vss.n12851 vss.t801 0.0702092
R45165 vss.n12851 vss.n12850 0.0702092
R45166 vss.n12854 vss.n12853 0.0702092
R45167 vss.n12840 vss.n10304 0.0702092
R45168 vss.n12835 vss.n10318 0.0702092
R45169 vss.t32 vss.n10318 0.0702092
R45170 vss.n10320 vss.n10319 0.0702092
R45171 vss.t32 vss.n10320 0.0702092
R45172 vss.n12829 vss.n12828 0.0702092
R45173 vss.t1310 vss.n12829 0.0702092
R45174 vss.n12826 vss.n12825 0.0702092
R45175 vss.n12825 vss.t1240 0.0702092
R45176 vss.n12813 vss.n12812 0.0702092
R45177 vss.n12812 vss.t1238 0.0702092
R45178 vss.t1310 vss.n12773 0.0702092
R45179 vss.t1240 vss.n12824 0.0702092
R45180 vss.n12820 vss.t1238 0.0702092
R45181 vss.n12821 vss.n12820 0.0702092
R45182 vss.n12824 vss.n12823 0.0702092
R45183 vss.n12783 vss.n12773 0.0702092
R45184 vss.n12818 vss.n12789 0.0702092
R45185 vss.n12818 vss.t843 0.0702092
R45186 vss.n12817 vss.n12816 0.0702092
R45187 vss.t843 vss.n12817 0.0702092
R45188 vss.n12917 vss.n12916 0.0702092
R45189 vss.n12916 vss.t1447 0.0702092
R45190 vss.n12800 vss.n12799 0.0702092
R45191 vss.t1448 vss.n12800 0.0702092
R45192 vss.n12794 vss.n12792 0.0702092
R45193 vss.n12792 vss.t1473 0.0702092
R45194 vss.t1447 vss.n12915 0.0702092
R45195 vss.t1448 vss.n12798 0.0702092
R45196 vss.n12793 vss.t1473 0.0702092
R45197 vss.n12805 vss.n12793 0.0702092
R45198 vss.n12798 vss.n10100 0.0702092
R45199 vss.n12915 vss.n12914 0.0702092
R45200 vss.n10096 vss.n10085 0.0702092
R45201 vss.t1426 vss.n10085 0.0702092
R45202 vss.n12920 vss.n12919 0.0702092
R45203 vss.t1426 vss.n12920 0.0702092
R45204 vss.n12926 vss.n12925 0.0702092
R45205 vss.n12925 vss.t1231 0.0702092
R45206 vss.n12936 vss.n12935 0.0702092
R45207 vss.n12935 vss.t273 0.0702092
R45208 vss.n12929 vss.n12928 0.0702092
R45209 vss.t275 vss.n12929 0.0702092
R45210 vss.n12924 vss.n12923 0.0702092
R45211 vss.t1231 vss.n12924 0.0702092
R45212 vss.n12931 vss.n12930 0.0702092
R45213 vss.n12930 vss.t275 0.0702092
R45214 vss.n12934 vss.n12933 0.0702092
R45215 vss.t273 vss.n12934 0.0702092
R45216 vss.n10057 vss.n10056 0.0702092
R45217 vss.t857 vss.n10057 0.0702092
R45218 vss.n12950 vss.n12949 0.0702092
R45219 vss.n12949 vss.t1518 0.0702092
R45220 vss.n10048 vss.n10018 0.0702092
R45221 vss.t1520 vss.n10048 0.0702092
R45222 vss.n10050 vss.n10049 0.0702092
R45223 vss.n10049 vss.t1520 0.0702092
R45224 vss.n12948 vss.n12947 0.0702092
R45225 vss.t1518 vss.n12948 0.0702092
R45226 vss.n12945 vss.n12944 0.0702092
R45227 vss.n12944 vss.t857 0.0702092
R45228 vss.n12938 vss.n10059 0.0702092
R45229 vss.t45 vss.n10059 0.0702092
R45230 vss.n12941 vss.n12940 0.0702092
R45231 vss.t45 vss.n12941 0.0702092
R45232 vss.n2118 vss.n2117 0.0702092
R45233 vss.t53 vss.n2118 0.0702092
R45234 vss.n13084 vss.n2103 0.0702092
R45235 vss.n13084 vss.t676 0.0702092
R45236 vss.n13087 vss.n13086 0.0702092
R45237 vss.n13086 vss.t678 0.0702092
R45238 vss.n2110 vss.n2109 0.0702092
R45239 vss.n2109 vss.t678 0.0702092
R45240 vss.n13083 vss.n13082 0.0702092
R45241 vss.t676 vss.n13083 0.0702092
R45242 vss.n13080 vss.n13079 0.0702092
R45243 vss.n13079 vss.t53 0.0702092
R45244 vss.n13109 vss.n2074 0.0702092
R45245 vss.n2074 vss.t776 0.0702092
R45246 vss.n13096 vss.n13095 0.0702092
R45247 vss.n13095 vss.t37 0.0702092
R45248 vss.n2092 vss.n2090 0.0702092
R45249 vss.t1182 vss.n2090 0.0702092
R45250 vss.n13107 vss.n13106 0.0702092
R45251 vss.n13106 vss.t1181 0.0702092
R45252 vss.n2075 vss.n2073 0.0702092
R45253 vss.n2073 vss.t776 0.0702092
R45254 vss.n13105 vss.n13104 0.0702092
R45255 vss.t1181 vss.n13105 0.0702092
R45256 vss.n13102 vss.n13101 0.0702092
R45257 vss.n13101 vss.t1182 0.0702092
R45258 vss.n2095 vss.n2094 0.0702092
R45259 vss.n2095 vss.t37 0.0702092
R45260 vss.n11852 vss.t530 0.0702092
R45261 vss.n11853 vss.n11851 0.0702092
R45262 vss.n11851 vss.t530 0.0702092
R45263 vss.n12094 vss.n11852 0.0702092
R45264 vss.n11883 vss.n11882 0.0702092
R45265 vss.n11882 vss.t1020 0.0702092
R45266 vss.n11886 vss.n11885 0.0702092
R45267 vss.t893 vss.n11886 0.0702092
R45268 vss.n12081 vss.n12080 0.0702092
R45269 vss.n12080 vss.t895 0.0702092
R45270 vss.n12083 vss.n11859 0.0702092
R45271 vss.n11859 vss.t628 0.0702092
R45272 vss.n11860 vss.n11858 0.0702092
R45273 vss.n11858 vss.t628 0.0702092
R45274 vss.n12079 vss.n12078 0.0702092
R45275 vss.t895 vss.n12079 0.0702092
R45276 vss.n11888 vss.n11887 0.0702092
R45277 vss.n11887 vss.t893 0.0702092
R45278 vss.n11881 vss.n11880 0.0702092
R45279 vss.t1020 vss.n11881 0.0702092
R45280 vss.n10482 vss.n10481 0.0702092
R45281 vss.t387 vss.n10482 0.0702092
R45282 vss.n10487 vss.n10486 0.0702092
R45283 vss.n10486 vss.t758 0.0702092
R45284 vss.n10489 vss.n10467 0.0702092
R45285 vss.t760 vss.n10467 0.0702092
R45286 vss.n10495 vss.n10494 0.0702092
R45287 vss.n10495 vss.t775 0.0702092
R45288 vss.n10492 vss.n10491 0.0702092
R45289 vss.n10491 vss.t775 0.0702092
R45290 vss.n10500 vss.n10499 0.0702092
R45291 vss.n10499 vss.t760 0.0702092
R45292 vss.n10485 vss.n10462 0.0702092
R45293 vss.t758 vss.n10485 0.0702092
R45294 vss.n10483 vss.n10479 0.0702092
R45295 vss.n10483 vss.t387 0.0702092
R45296 vss.n10703 vss.n10702 0.0702092
R45297 vss.t1489 vss.n10703 0.0702092
R45298 vss.n10708 vss.n10707 0.0702092
R45299 vss.n10707 vss.t1129 0.0702092
R45300 vss.n10710 vss.n10688 0.0702092
R45301 vss.t1131 vss.n10688 0.0702092
R45302 vss.n10716 vss.n10715 0.0702092
R45303 vss.n10716 vss.t167 0.0702092
R45304 vss.n10713 vss.n10712 0.0702092
R45305 vss.n10712 vss.t167 0.0702092
R45306 vss.n10721 vss.n10720 0.0702092
R45307 vss.n10720 vss.t1131 0.0702092
R45308 vss.n10706 vss.n10683 0.0702092
R45309 vss.t1129 vss.n10706 0.0702092
R45310 vss.n10704 vss.n10700 0.0702092
R45311 vss.n10704 vss.t1489 0.0702092
R45312 vss.n11017 vss.n11016 0.0702092
R45313 vss.t1328 vss.n11017 0.0702092
R45314 vss.n11022 vss.n11021 0.0702092
R45315 vss.n11021 vss.t927 0.0702092
R45316 vss.n11024 vss.n11002 0.0702092
R45317 vss.t929 vss.n11002 0.0702092
R45318 vss.n11030 vss.n11029 0.0702092
R45319 vss.n11030 vss.t930 0.0702092
R45320 vss.n11027 vss.n11026 0.0702092
R45321 vss.n11026 vss.t930 0.0702092
R45322 vss.n11035 vss.n11034 0.0702092
R45323 vss.n11034 vss.t929 0.0702092
R45324 vss.n11020 vss.n10997 0.0702092
R45325 vss.t927 vss.n11020 0.0702092
R45326 vss.n11018 vss.n11014 0.0702092
R45327 vss.n11018 vss.t1328 0.0702092
R45328 vss.n11136 vss.n11135 0.0702092
R45329 vss.n11136 vss.t911 0.0702092
R45330 vss.t1378 vss.n11125 0.0702092
R45331 vss.n11129 vss.t355 0.0702092
R45332 vss.t357 vss.n11142 0.0702092
R45333 vss.n11138 vss.t911 0.0702092
R45334 vss.n11144 vss.n11143 0.0702092
R45335 vss.n11143 vss.t357 0.0702092
R45336 vss.n11128 vss.n11106 0.0702092
R45337 vss.t355 vss.n11128 0.0702092
R45338 vss.n11126 vss.n11122 0.0702092
R45339 vss.n11126 vss.t1378 0.0702092
R45340 vss.n11125 vss.n11124 0.0702092
R45341 vss.n11130 vss.n11129 0.0702092
R45342 vss.n11142 vss.n11141 0.0702092
R45343 vss.n11139 vss.n11138 0.0702092
R45344 vss.n2044 vss.n2043 0.0661418
R45345 vss.n2043 vss.n2038 0.0661418
R45346 vss.n2039 vss.n2032 0.0661418
R45347 vss.n2039 vss.n2037 0.0661418
R45348 vss.n10400 vss.n10397 0.0661418
R45349 vss.n10400 vss.n10399 0.0661418
R45350 vss.n10408 vss.n10407 0.0661418
R45351 vss.n10409 vss.n10408 0.0661418
R45352 vss.n13139 vss.n2045 0.0661418
R45353 vss.n13139 vss.n13138 0.0661418
R45354 vss.n12649 vss.n12648 0.0661418
R45355 vss.n12648 vss.n12627 0.0661418
R45356 vss.n12628 vss.n12621 0.0661418
R45357 vss.n12628 vss.n12626 0.0661418
R45358 vss.n12636 vss.n12634 0.0661418
R45359 vss.n12634 vss.n12633 0.0661418
R45360 vss.n12639 vss.n12635 0.0661418
R45361 vss.n12635 vss.n10410 0.0661418
R45362 vss.n12653 vss.n12650 0.0661418
R45363 vss.n12653 vss.n2049 0.0661418
R45364 vss.n10385 vss.n10374 0.0661418
R45365 vss.n10385 vss.n10379 0.0661418
R45366 vss.n10390 vss.n10388 0.0661418
R45367 vss.n10388 vss.n10387 0.0661418
R45368 vss.n12691 vss.n10381 0.0661418
R45369 vss.n12692 vss.n12691 0.0661418
R45370 vss.n12687 vss.n10382 0.0661418
R45371 vss.n10382 vss.n2068 0.0661418
R45372 vss.n12674 vss.n10389 0.0661418
R45373 vss.n12673 vss.n10389 0.0661418
R45374 vss.n11416 vss.n11405 0.0661418
R45375 vss.n11416 vss.n11410 0.0661418
R45376 vss.n11421 vss.n11419 0.0661418
R45377 vss.n11419 vss.n11418 0.0661418
R45378 vss.n11441 vss.n11412 0.0661418
R45379 vss.n11442 vss.n11441 0.0661418
R45380 vss.n11437 vss.n11413 0.0661418
R45381 vss.n11413 vss.n2065 0.0661418
R45382 vss.n11424 vss.n11420 0.0661418
R45383 vss.n11420 vss.n10411 0.0661418
R45384 vss.n11369 vss.n11358 0.0661418
R45385 vss.n11369 vss.n11363 0.0661418
R45386 vss.n11374 vss.n11372 0.0661418
R45387 vss.n11372 vss.n11371 0.0661418
R45388 vss.n11394 vss.n11365 0.0661418
R45389 vss.n11395 vss.n11394 0.0661418
R45390 vss.n11390 vss.n11366 0.0661418
R45391 vss.n11366 vss.n2067 0.0661418
R45392 vss.n11377 vss.n11373 0.0661418
R45393 vss.n11373 vss.n10412 0.0661418
R45394 vss.n10944 vss.n10933 0.0661418
R45395 vss.n10944 vss.n10938 0.0661418
R45396 vss.n10949 vss.n10947 0.0661418
R45397 vss.n10947 vss.n10946 0.0661418
R45398 vss.n10969 vss.n10940 0.0661418
R45399 vss.n10970 vss.n10969 0.0661418
R45400 vss.n10965 vss.n10941 0.0661418
R45401 vss.n10941 vss.n2062 0.0661418
R45402 vss.n10952 vss.n10948 0.0661418
R45403 vss.n10948 vss.n10413 0.0661418
R45404 vss.n10781 vss.n10770 0.0661418
R45405 vss.n10781 vss.n10775 0.0661418
R45406 vss.n10786 vss.n10784 0.0661418
R45407 vss.n10784 vss.n10783 0.0661418
R45408 vss.n10806 vss.n10777 0.0661418
R45409 vss.n10807 vss.n10806 0.0661418
R45410 vss.n10802 vss.n10778 0.0661418
R45411 vss.n10778 vss.n2059 0.0661418
R45412 vss.n10789 vss.n10785 0.0661418
R45413 vss.n10785 vss.n10414 0.0661418
R45414 vss.n10737 vss.n10726 0.0661418
R45415 vss.n10737 vss.n10731 0.0661418
R45416 vss.n10742 vss.n10740 0.0661418
R45417 vss.n10740 vss.n10739 0.0661418
R45418 vss.n10762 vss.n10733 0.0661418
R45419 vss.n10763 vss.n10762 0.0661418
R45420 vss.n10758 vss.n10734 0.0661418
R45421 vss.n10734 vss.n2061 0.0661418
R45422 vss.n10745 vss.n10741 0.0661418
R45423 vss.n10741 vss.n10415 0.0661418
R45424 vss.n11563 vss.n11552 0.0661418
R45425 vss.n11563 vss.n11557 0.0661418
R45426 vss.n11568 vss.n11566 0.0661418
R45427 vss.n11566 vss.n11565 0.0661418
R45428 vss.n11588 vss.n11559 0.0661418
R45429 vss.n11589 vss.n11588 0.0661418
R45430 vss.n11584 vss.n11560 0.0661418
R45431 vss.n11560 vss.n2056 0.0661418
R45432 vss.n11571 vss.n11567 0.0661418
R45433 vss.n11567 vss.n10416 0.0661418
R45434 vss.n10560 vss.n10549 0.0661418
R45435 vss.n10560 vss.n10554 0.0661418
R45436 vss.n10565 vss.n10563 0.0661418
R45437 vss.n10563 vss.n10562 0.0661418
R45438 vss.n10585 vss.n10556 0.0661418
R45439 vss.n10586 vss.n10585 0.0661418
R45440 vss.n10581 vss.n10557 0.0661418
R45441 vss.n10557 vss.n2053 0.0661418
R45442 vss.n10568 vss.n10564 0.0661418
R45443 vss.n10564 vss.n10417 0.0661418
R45444 vss.n10516 vss.n10505 0.0661418
R45445 vss.n10516 vss.n10510 0.0661418
R45446 vss.n10521 vss.n10519 0.0661418
R45447 vss.n10519 vss.n10518 0.0661418
R45448 vss.n10541 vss.n10512 0.0661418
R45449 vss.n10542 vss.n10541 0.0661418
R45450 vss.n10537 vss.n10513 0.0661418
R45451 vss.n10513 vss.n2055 0.0661418
R45452 vss.n10524 vss.n10520 0.0661418
R45453 vss.n10520 vss.n10418 0.0661418
R45454 vss.n11937 vss.n11926 0.0661418
R45455 vss.n11937 vss.n11931 0.0661418
R45456 vss.n11942 vss.n11940 0.0661418
R45457 vss.n11940 vss.n11939 0.0661418
R45458 vss.n11962 vss.n11933 0.0661418
R45459 vss.n11963 vss.n11962 0.0661418
R45460 vss.n11958 vss.n11934 0.0661418
R45461 vss.n11934 vss.n2050 0.0661418
R45462 vss.n11945 vss.n11941 0.0661418
R45463 vss.n11941 vss.n10419 0.0661418
R45464 vss.n12089 vss.n11854 0.0661418
R45465 vss.n12089 vss.n12088 0.0661418
R45466 vss.n11895 vss.n11892 0.0661418
R45467 vss.n11898 vss.n11895 0.0661418
R45468 vss.n11901 vss.n11900 0.0661418
R45469 vss.n11900 vss.n11897 0.0661418
R45470 vss.n11903 vss.n11902 0.0661418
R45471 vss.n12060 vss.n11903 0.0661418
R45472 vss.n11910 vss.n11907 0.0661418
R45473 vss.n11910 vss.n2051 0.0661418
R45474 vss.n11920 vss.n11917 0.0661418
R45475 vss.n11920 vss.n11919 0.0661418
R45476 vss.n11922 vss.n11914 0.0661418
R45477 vss.n11915 vss.n11914 0.0661418
R45478 vss.n12057 vss.n12056 0.0661418
R45479 vss.n12058 vss.n12057 0.0661418
R45480 vss.n12046 vss.n11918 0.0661418
R45481 vss.n12046 vss.n12045 0.0661418
R45482 vss.n12037 vss.n12032 0.0661418
R45483 vss.n12037 vss.n12036 0.0661418
R45484 vss.n12042 vss.n12041 0.0661418
R45485 vss.n12043 vss.n12042 0.0661418
R45486 vss.n12012 vss.n11985 0.0661418
R45487 vss.n11987 vss.n11985 0.0661418
R45488 vss.n12010 vss.n11988 0.0661418
R45489 vss.n12010 vss.n12009 0.0661418
R45490 vss.n11990 vss.n11989 0.0661418
R45491 vss.n12008 vss.n11990 0.0661418
R45492 vss.n11998 vss.n11995 0.0661418
R45493 vss.n11998 vss.n2054 0.0661418
R45494 vss.n10603 vss.n10602 0.0661418
R45495 vss.n10602 vss.n10597 0.0661418
R45496 vss.n10598 vss.n10591 0.0661418
R45497 vss.n10598 vss.n10596 0.0661418
R45498 vss.n12005 vss.n12004 0.0661418
R45499 vss.n12006 vss.n12005 0.0661418
R45500 vss.n12601 vss.n10604 0.0661418
R45501 vss.n12601 vss.n12600 0.0661418
R45502 vss.n12592 vss.n10611 0.0661418
R45503 vss.n12592 vss.n12591 0.0661418
R45504 vss.n12597 vss.n12596 0.0661418
R45505 vss.n12598 vss.n12597 0.0661418
R45506 vss.n10661 vss.n10659 0.0661418
R45507 vss.n10661 vss.n10660 0.0661418
R45508 vss.n10652 vss.n10646 0.0661418
R45509 vss.n10652 vss.n10651 0.0661418
R45510 vss.n10669 vss.n10668 0.0661418
R45511 vss.n10670 vss.n10669 0.0661418
R45512 vss.n10640 vss.n10639 0.0661418
R45513 vss.n10640 vss.n2057 0.0661418
R45514 vss.n11604 vss.n10626 0.0661418
R45515 vss.n11604 vss.n11603 0.0661418
R45516 vss.n10634 vss.n10630 0.0661418
R45517 vss.n10635 vss.n10634 0.0661418
R45518 vss.n10638 vss.n10637 0.0661418
R45519 vss.n10637 vss.n10633 0.0661418
R45520 vss.n11611 vss.n11610 0.0661418
R45521 vss.n11612 vss.n11611 0.0661418
R45522 vss.n11622 vss.n11621 0.0661418
R45523 vss.n11623 vss.n11622 0.0661418
R45524 vss.n11615 vss.n10619 0.0661418
R45525 vss.n11615 vss.n11614 0.0661418
R45526 vss.n10842 vss.n10841 0.0661418
R45527 vss.n10841 vss.n10836 0.0661418
R45528 vss.n10837 vss.n10833 0.0661418
R45529 vss.n10837 vss.n10835 0.0661418
R45530 vss.n10856 vss.n10855 0.0661418
R45531 vss.n10857 vss.n10856 0.0661418
R45532 vss.n10859 vss.n10826 0.0661418
R45533 vss.n10826 vss.n2060 0.0661418
R45534 vss.n10869 vss.n10868 0.0661418
R45535 vss.n10868 vss.n10818 0.0661418
R45536 vss.n10819 vss.n10812 0.0661418
R45537 vss.n10819 vss.n10817 0.0661418
R45538 vss.n10827 vss.n10825 0.0661418
R45539 vss.n10825 vss.n10824 0.0661418
R45540 vss.n11530 vss.n10870 0.0661418
R45541 vss.n11530 vss.n11529 0.0661418
R45542 vss.n11521 vss.n11517 0.0661418
R45543 vss.n11521 vss.n11520 0.0661418
R45544 vss.n11526 vss.n11525 0.0661418
R45545 vss.n11527 vss.n11526 0.0661418
R45546 vss.n11499 vss.n10877 0.0661418
R45547 vss.n10879 vss.n10877 0.0661418
R45548 vss.n11497 vss.n10880 0.0661418
R45549 vss.n11497 vss.n11496 0.0661418
R45550 vss.n10882 vss.n10881 0.0661418
R45551 vss.n11495 vss.n10882 0.0661418
R45552 vss.n10889 vss.n10886 0.0661418
R45553 vss.n10889 vss.n2063 0.0661418
R45554 vss.n10983 vss.n10896 0.0661418
R45555 vss.n10983 vss.n10982 0.0661418
R45556 vss.n10976 vss.n10893 0.0661418
R45557 vss.n10894 vss.n10893 0.0661418
R45558 vss.n11492 vss.n11491 0.0661418
R45559 vss.n11493 vss.n11492 0.0661418
R45560 vss.n11481 vss.n10897 0.0661418
R45561 vss.n11481 vss.n11480 0.0661418
R45562 vss.n11472 vss.n11469 0.0661418
R45563 vss.n11472 vss.n10322 0.0661418
R45564 vss.n11477 vss.n11476 0.0661418
R45565 vss.n11478 vss.n11477 0.0661418
R45566 vss.n10932 vss.n10903 0.0661418
R45567 vss.n10905 vss.n10903 0.0661418
R45568 vss.n10930 vss.n10906 0.0661418
R45569 vss.n10930 vss.n10929 0.0661418
R45570 vss.n10908 vss.n10907 0.0661418
R45571 vss.n10928 vss.n10908 0.0661418
R45572 vss.n10918 vss.n10915 0.0661418
R45573 vss.n10918 vss.n2066 0.0661418
R45574 vss.n12747 vss.n10333 0.0661418
R45575 vss.n12747 vss.n12746 0.0661418
R45576 vss.n10909 vss.n10337 0.0661418
R45577 vss.n10910 vss.n10909 0.0661418
R45578 vss.n10925 vss.n10924 0.0661418
R45579 vss.n10926 vss.n10925 0.0661418
R45580 vss.n12754 vss.n12753 0.0661418
R45581 vss.n12755 vss.n12754 0.0661418
R45582 vss.n12765 vss.n12764 0.0661418
R45583 vss.n12766 vss.n12765 0.0661418
R45584 vss.n12758 vss.n10326 0.0661418
R45585 vss.n12758 vss.n12757 0.0661418
R45586 vss.n10344 vss.n10341 0.0661418
R45587 vss.n10347 vss.n10344 0.0661418
R45588 vss.n10350 vss.n10349 0.0661418
R45589 vss.n10349 vss.n10346 0.0661418
R45590 vss.n10352 vss.n10351 0.0661418
R45591 vss.n12725 vss.n10352 0.0661418
R45592 vss.n10359 vss.n10356 0.0661418
R45593 vss.n10359 vss.n2069 0.0661418
R45594 vss.n10369 vss.n10366 0.0661418
R45595 vss.n10369 vss.n10368 0.0661418
R45596 vss.n10371 vss.n10363 0.0661418
R45597 vss.n10364 vss.n10363 0.0661418
R45598 vss.n12722 vss.n12721 0.0661418
R45599 vss.n12723 vss.n12722 0.0661418
R45600 vss.n12711 vss.n10367 0.0661418
R45601 vss.n12711 vss.n12710 0.0661418
R45602 vss.n2271 vss.n2262 0.0661418
R45603 vss.n2271 vss.n2269 0.0661418
R45604 vss.n2276 vss.n2275 0.0661418
R45605 vss.n2275 vss.n2270 0.0661418
R45606 vss.n2290 vss.n2289 0.0661418
R45607 vss.n2291 vss.n2290 0.0661418
R45608 vss.n2285 vss.n2282 0.0661418
R45609 vss.n2285 vss.n2143 0.0661418
R45610 vss.n2302 vss.n2301 0.0661418
R45611 vss.n2303 vss.n2302 0.0661418
R45612 vss.n2256 vss.n2254 0.0661418
R45613 vss.n2254 vss.n2253 0.0661418
R45614 vss.n2248 vss.n2241 0.0661418
R45615 vss.n2248 vss.n2246 0.0661418
R45616 vss.n13005 vss.n13004 0.0661418
R45617 vss.n13004 vss.n2247 0.0661418
R45618 vss.n13007 vss.n13006 0.0661418
R45619 vss.n13007 vss.n2144 0.0661418
R45620 vss.n12995 vss.n2255 0.0661418
R45621 vss.n12994 vss.n2255 0.0661418
R45622 vss.n13317 vss.n13316 0.0661418
R45623 vss.n13316 vss.n13310 0.0661418
R45624 vss.n13901 vss.n13322 0.0661418
R45625 vss.n13325 vss.n13322 0.0661418
R45626 vss.n13311 vss.n13307 0.0661418
R45627 vss.n13311 vss.n13303 0.0661418
R45628 vss.n13306 vss.n13302 0.0661418
R45629 vss.n13920 vss.n13302 0.0661418
R45630 vss.n13905 vss.n13324 0.0661418
R45631 vss.n13899 vss.n13324 0.0661418
R45632 vss.n13889 vss.n13329 0.0661418
R45633 vss.n13889 vss.n13888 0.0661418
R45634 vss.n13337 vss.n13333 0.0661418
R45635 vss.n13338 vss.n13337 0.0661418
R45636 vss.n13341 vss.n13340 0.0661418
R45637 vss.n13340 vss.n13336 0.0661418
R45638 vss.n13896 vss.n13895 0.0661418
R45639 vss.n13897 vss.n13896 0.0661418
R45640 vss.n13343 vss.n13342 0.0661418
R45641 vss.n13343 vss.n689 0.0661418
R45642 vss.n13359 vss.n13358 0.0661418
R45643 vss.n13358 vss.n13352 0.0661418
R45644 vss.n13846 vss.n13361 0.0661418
R45645 vss.n13364 vss.n13361 0.0661418
R45646 vss.n13353 vss.n13349 0.0661418
R45647 vss.n13353 vss.n13345 0.0661418
R45648 vss.n13348 vss.n13344 0.0661418
R45649 vss.n13872 vss.n13344 0.0661418
R45650 vss.n13850 vss.n13363 0.0661418
R45651 vss.n13363 vss.n192 0.0661418
R45652 vss.n13835 vss.n13368 0.0661418
R45653 vss.n13835 vss.n13834 0.0661418
R45654 vss.n13378 vss.n13374 0.0661418
R45655 vss.n13379 vss.n13378 0.0661418
R45656 vss.n13382 vss.n13381 0.0661418
R45657 vss.n13381 vss.n13377 0.0661418
R45658 vss.n13842 vss.n13841 0.0661418
R45659 vss.n13843 vss.n13842 0.0661418
R45660 vss.n13384 vss.n13383 0.0661418
R45661 vss.n13384 vss.n687 0.0661418
R45662 vss.n13400 vss.n13399 0.0661418
R45663 vss.n13399 vss.n13393 0.0661418
R45664 vss.n13796 vss.n13402 0.0661418
R45665 vss.n13405 vss.n13402 0.0661418
R45666 vss.n13394 vss.n13390 0.0661418
R45667 vss.n13394 vss.n13386 0.0661418
R45668 vss.n13389 vss.n13385 0.0661418
R45669 vss.n13818 vss.n13385 0.0661418
R45670 vss.n13800 vss.n13404 0.0661418
R45671 vss.n13794 vss.n13404 0.0661418
R45672 vss.n13784 vss.n13409 0.0661418
R45673 vss.n13784 vss.n13783 0.0661418
R45674 vss.n13417 vss.n13413 0.0661418
R45675 vss.n13418 vss.n13417 0.0661418
R45676 vss.n13421 vss.n13420 0.0661418
R45677 vss.n13420 vss.n13416 0.0661418
R45678 vss.n13791 vss.n13790 0.0661418
R45679 vss.n13792 vss.n13791 0.0661418
R45680 vss.n13423 vss.n13422 0.0661418
R45681 vss.n13423 vss.n685 0.0661418
R45682 vss.n13439 vss.n13438 0.0661418
R45683 vss.n13438 vss.n13432 0.0661418
R45684 vss.n13741 vss.n13441 0.0661418
R45685 vss.n13444 vss.n13441 0.0661418
R45686 vss.n13433 vss.n13429 0.0661418
R45687 vss.n13433 vss.n13425 0.0661418
R45688 vss.n13428 vss.n13424 0.0661418
R45689 vss.n13767 vss.n13424 0.0661418
R45690 vss.n13745 vss.n13443 0.0661418
R45691 vss.n13443 vss.n251 0.0661418
R45692 vss.n13730 vss.n13448 0.0661418
R45693 vss.n13730 vss.n13729 0.0661418
R45694 vss.n13458 vss.n13454 0.0661418
R45695 vss.n13459 vss.n13458 0.0661418
R45696 vss.n13462 vss.n13461 0.0661418
R45697 vss.n13461 vss.n13457 0.0661418
R45698 vss.n13737 vss.n13736 0.0661418
R45699 vss.n13738 vss.n13737 0.0661418
R45700 vss.n13464 vss.n13463 0.0661418
R45701 vss.n13464 vss.n683 0.0661418
R45702 vss.n13480 vss.n13479 0.0661418
R45703 vss.n13479 vss.n13473 0.0661418
R45704 vss.n13691 vss.n13482 0.0661418
R45705 vss.n13485 vss.n13482 0.0661418
R45706 vss.n13474 vss.n13470 0.0661418
R45707 vss.n13474 vss.n13466 0.0661418
R45708 vss.n13469 vss.n13465 0.0661418
R45709 vss.n13713 vss.n13465 0.0661418
R45710 vss.n13695 vss.n13484 0.0661418
R45711 vss.n13689 vss.n13484 0.0661418
R45712 vss.n13679 vss.n13489 0.0661418
R45713 vss.n13679 vss.n13678 0.0661418
R45714 vss.n13497 vss.n13493 0.0661418
R45715 vss.n13498 vss.n13497 0.0661418
R45716 vss.n13501 vss.n13500 0.0661418
R45717 vss.n13500 vss.n13496 0.0661418
R45718 vss.n13686 vss.n13685 0.0661418
R45719 vss.n13687 vss.n13686 0.0661418
R45720 vss.n13503 vss.n13502 0.0661418
R45721 vss.n13503 vss.n681 0.0661418
R45722 vss.n13519 vss.n13518 0.0661418
R45723 vss.n13518 vss.n13512 0.0661418
R45724 vss.n13636 vss.n13521 0.0661418
R45725 vss.n13524 vss.n13521 0.0661418
R45726 vss.n13513 vss.n13509 0.0661418
R45727 vss.n13513 vss.n13505 0.0661418
R45728 vss.n13508 vss.n13504 0.0661418
R45729 vss.n13662 vss.n13504 0.0661418
R45730 vss.n13640 vss.n13523 0.0661418
R45731 vss.n13523 vss.n310 0.0661418
R45732 vss.n13625 vss.n13528 0.0661418
R45733 vss.n13625 vss.n13624 0.0661418
R45734 vss.n13538 vss.n13534 0.0661418
R45735 vss.n13539 vss.n13538 0.0661418
R45736 vss.n13542 vss.n13541 0.0661418
R45737 vss.n13541 vss.n13537 0.0661418
R45738 vss.n13632 vss.n13631 0.0661418
R45739 vss.n13633 vss.n13632 0.0661418
R45740 vss.n13544 vss.n13543 0.0661418
R45741 vss.n13544 vss.n679 0.0661418
R45742 vss.n13557 vss.n13548 0.0661418
R45743 vss.n13557 vss.n13555 0.0661418
R45744 vss.n13562 vss.n13561 0.0661418
R45745 vss.n13561 vss.n13556 0.0661418
R45746 vss.n13595 vss.n13594 0.0661418
R45747 vss.n13596 vss.n13595 0.0661418
R45748 vss.n13607 vss.n13606 0.0661418
R45749 vss.n13608 vss.n13607 0.0661418
R45750 vss.n467 vss.n463 0.0661418
R45751 vss.n467 vss.n457 0.0661418
R45752 vss.n473 vss.n472 0.0661418
R45753 vss.n472 vss.n466 0.0661418
R45754 vss.n13577 vss.n13576 0.0661418
R45755 vss.n13576 vss.n13575 0.0661418
R45756 vss.n13581 vss.n13580 0.0661418
R45757 vss.n13582 vss.n13581 0.0661418
R45758 vss.n13587 vss.n13586 0.0661418
R45759 vss.n13588 vss.n13587 0.0661418
R45760 vss.n170 vss.n168 0.0661418
R45761 vss.n168 vss.n167 0.0661418
R45762 vss.n162 vss.n155 0.0661418
R45763 vss.n162 vss.n160 0.0661418
R45764 vss.n14743 vss.n14742 0.0661418
R45765 vss.n14742 vss.n161 0.0661418
R45766 vss.n14745 vss.n14744 0.0661418
R45767 vss.n14745 vss.n19 0.0661418
R45768 vss.n14733 vss.n169 0.0661418
R45769 vss.n14732 vss.n169 0.0661418
R45770 vss.n14651 vss.n197 0.0661418
R45771 vss.n14651 vss.n14649 0.0661418
R45772 vss.n14656 vss.n14655 0.0661418
R45773 vss.n14655 vss.n14650 0.0661418
R45774 vss.n14670 vss.n14669 0.0661418
R45775 vss.n14671 vss.n14670 0.0661418
R45776 vss.n14665 vss.n14662 0.0661418
R45777 vss.n14665 vss.n20 0.0661418
R45778 vss.n14682 vss.n14681 0.0661418
R45779 vss.n14683 vss.n14682 0.0661418
R45780 vss.n247 vss.n245 0.0661418
R45781 vss.n245 vss.n244 0.0661418
R45782 vss.n239 vss.n232 0.0661418
R45783 vss.n239 vss.n237 0.0661418
R45784 vss.n14548 vss.n14547 0.0661418
R45785 vss.n14547 vss.n238 0.0661418
R45786 vss.n14550 vss.n14549 0.0661418
R45787 vss.n14550 vss.n21 0.0661418
R45788 vss.n14538 vss.n246 0.0661418
R45789 vss.n14537 vss.n246 0.0661418
R45790 vss.n14456 vss.n256 0.0661418
R45791 vss.n14456 vss.n14454 0.0661418
R45792 vss.n14461 vss.n14460 0.0661418
R45793 vss.n14460 vss.n14455 0.0661418
R45794 vss.n14475 vss.n14474 0.0661418
R45795 vss.n14476 vss.n14475 0.0661418
R45796 vss.n14470 vss.n14467 0.0661418
R45797 vss.n14470 vss.n22 0.0661418
R45798 vss.n14487 vss.n14486 0.0661418
R45799 vss.n14488 vss.n14487 0.0661418
R45800 vss.n306 vss.n304 0.0661418
R45801 vss.n304 vss.n303 0.0661418
R45802 vss.n298 vss.n291 0.0661418
R45803 vss.n298 vss.n296 0.0661418
R45804 vss.n14353 vss.n14352 0.0661418
R45805 vss.n14352 vss.n297 0.0661418
R45806 vss.n14355 vss.n14354 0.0661418
R45807 vss.n14355 vss.n23 0.0661418
R45808 vss.n14343 vss.n305 0.0661418
R45809 vss.n14342 vss.n305 0.0661418
R45810 vss.n14261 vss.n315 0.0661418
R45811 vss.n14261 vss.n14259 0.0661418
R45812 vss.n14266 vss.n14265 0.0661418
R45813 vss.n14265 vss.n14260 0.0661418
R45814 vss.n14280 vss.n14279 0.0661418
R45815 vss.n14281 vss.n14280 0.0661418
R45816 vss.n14275 vss.n14272 0.0661418
R45817 vss.n14275 vss.n24 0.0661418
R45818 vss.n14292 vss.n14291 0.0661418
R45819 vss.n14293 vss.n14292 0.0661418
R45820 vss.n429 vss.n427 0.0661418
R45821 vss.n427 vss.n426 0.0661418
R45822 vss.n421 vss.n414 0.0661418
R45823 vss.n421 vss.n419 0.0661418
R45824 vss.n14234 vss.n14233 0.0661418
R45825 vss.n14233 vss.n420 0.0661418
R45826 vss.n14236 vss.n14235 0.0661418
R45827 vss.n14236 vss.n25 0.0661418
R45828 vss.n14224 vss.n428 0.0661418
R45829 vss.n14223 vss.n428 0.0661418
R45830 vss.n14111 vss.n14109 0.0661418
R45831 vss.n14109 vss.n14108 0.0661418
R45832 vss.n14103 vss.n14096 0.0661418
R45833 vss.n14103 vss.n14101 0.0661418
R45834 vss.n14125 vss.n14124 0.0661418
R45835 vss.n14124 vss.n14102 0.0661418
R45836 vss.n14127 vss.n14126 0.0661418
R45837 vss.n14127 vss.n26 0.0661418
R45838 vss.n14115 vss.n14110 0.0661418
R45839 vss.n14114 vss.n14110 0.0661418
R45840 vss.n14188 vss.n14180 0.0661418
R45841 vss.n14188 vss.n14186 0.0661418
R45842 vss.n14193 vss.n14192 0.0661418
R45843 vss.n14192 vss.n14187 0.0661418
R45844 vss.n14207 vss.n14206 0.0661418
R45845 vss.n14208 vss.n14207 0.0661418
R45846 vss.n14202 vss.n14199 0.0661418
R45847 vss.n14202 vss.n27 0.0661418
R45848 vss.n14219 vss.n14218 0.0661418
R45849 vss.n14220 vss.n14219 0.0661418
R45850 vss.n332 vss.n330 0.0661418
R45851 vss.n330 vss.n329 0.0661418
R45852 vss.n324 vss.n317 0.0661418
R45853 vss.n324 vss.n322 0.0661418
R45854 vss.n346 vss.n345 0.0661418
R45855 vss.n345 vss.n323 0.0661418
R45856 vss.n348 vss.n347 0.0661418
R45857 vss.n348 vss.n28 0.0661418
R45858 vss.n336 vss.n331 0.0661418
R45859 vss.n335 vss.n331 0.0661418
R45860 vss.n14307 vss.n14299 0.0661418
R45861 vss.n14307 vss.n14305 0.0661418
R45862 vss.n14312 vss.n14311 0.0661418
R45863 vss.n14311 vss.n14306 0.0661418
R45864 vss.n14326 vss.n14325 0.0661418
R45865 vss.n14327 vss.n14326 0.0661418
R45866 vss.n14321 vss.n14318 0.0661418
R45867 vss.n14321 vss.n29 0.0661418
R45868 vss.n14338 vss.n14337 0.0661418
R45869 vss.n14339 vss.n14338 0.0661418
R45870 vss.n14385 vss.n14383 0.0661418
R45871 vss.n14383 vss.n14382 0.0661418
R45872 vss.n14377 vss.n14370 0.0661418
R45873 vss.n14377 vss.n14375 0.0661418
R45874 vss.n14399 vss.n14398 0.0661418
R45875 vss.n14398 vss.n14376 0.0661418
R45876 vss.n14401 vss.n14400 0.0661418
R45877 vss.n14401 vss.n30 0.0661418
R45878 vss.n14389 vss.n14384 0.0661418
R45879 vss.n14388 vss.n14384 0.0661418
R45880 vss.n14502 vss.n14494 0.0661418
R45881 vss.n14502 vss.n14500 0.0661418
R45882 vss.n14507 vss.n14506 0.0661418
R45883 vss.n14506 vss.n14501 0.0661418
R45884 vss.n14521 vss.n14520 0.0661418
R45885 vss.n14522 vss.n14521 0.0661418
R45886 vss.n14516 vss.n14513 0.0661418
R45887 vss.n14516 vss.n31 0.0661418
R45888 vss.n14533 vss.n14532 0.0661418
R45889 vss.n14534 vss.n14533 0.0661418
R45890 vss.n14580 vss.n14578 0.0661418
R45891 vss.n14578 vss.n14577 0.0661418
R45892 vss.n14572 vss.n14565 0.0661418
R45893 vss.n14572 vss.n14570 0.0661418
R45894 vss.n14594 vss.n14593 0.0661418
R45895 vss.n14593 vss.n14571 0.0661418
R45896 vss.n14596 vss.n14595 0.0661418
R45897 vss.n14596 vss.n32 0.0661418
R45898 vss.n14584 vss.n14579 0.0661418
R45899 vss.n14583 vss.n14579 0.0661418
R45900 vss.n14697 vss.n14689 0.0661418
R45901 vss.n14697 vss.n14695 0.0661418
R45902 vss.n14702 vss.n14701 0.0661418
R45903 vss.n14701 vss.n14696 0.0661418
R45904 vss.n14716 vss.n14715 0.0661418
R45905 vss.n14717 vss.n14716 0.0661418
R45906 vss.n14711 vss.n14708 0.0661418
R45907 vss.n14711 vss.n33 0.0661418
R45908 vss.n14728 vss.n14727 0.0661418
R45909 vss.n14729 vss.n14728 0.0661418
R45910 vss.n184 vss.n183 0.0661418
R45911 vss.n183 vss.n182 0.0661418
R45912 vss.n8 vss.n1 0.0661418
R45913 vss.n8 vss.n6 0.0661418
R45914 vss.n13 vss.n12 0.0661418
R45915 vss.n12 vss.n7 0.0661418
R45916 vss.n15 vss.n14 0.0661418
R45917 vss.n14784 vss.n15 0.0661418
R45918 vss.n188 vss.n187 0.0661418
R45919 vss.n189 vss.n188 0.0661418
R45920 vss.n528 vss.n517 0.0661418
R45921 vss.n528 vss.n522 0.0661418
R45922 vss.n533 vss.n531 0.0661418
R45923 vss.n531 vss.n530 0.0661418
R45924 vss.n14020 vss.n524 0.0661418
R45925 vss.n14021 vss.n14020 0.0661418
R45926 vss.n14016 vss.n525 0.0661418
R45927 vss.n659 vss.n525 0.0661418
R45928 vss.n14003 vss.n532 0.0661418
R45929 vss.n536 vss.n532 0.0661418
R45930 vss.n551 vss.n550 0.0661418
R45931 vss.n550 vss.n545 0.0661418
R45932 vss.n546 vss.n540 0.0661418
R45933 vss.n546 vss.n544 0.0661418
R45934 vss.n669 vss.n664 0.0661418
R45935 vss.n669 vss.n668 0.0661418
R45936 vss.n14000 vss.n13999 0.0661418
R45937 vss.n14001 vss.n14000 0.0661418
R45938 vss.n677 vss.n676 0.0661418
R45939 vss.n678 vss.n677 0.0661418
R45940 vss.n567 vss.n556 0.0661418
R45941 vss.n567 vss.n561 0.0661418
R45942 vss.n572 vss.n570 0.0661418
R45943 vss.n570 vss.n569 0.0661418
R45944 vss.n13985 vss.n563 0.0661418
R45945 vss.n13986 vss.n13985 0.0661418
R45946 vss.n13981 vss.n564 0.0661418
R45947 vss.n666 vss.n564 0.0661418
R45948 vss.n13968 vss.n571 0.0661418
R45949 vss.n575 vss.n571 0.0661418
R45950 vss.n590 vss.n589 0.0661418
R45951 vss.n589 vss.n584 0.0661418
R45952 vss.n585 vss.n579 0.0661418
R45953 vss.n585 vss.n583 0.0661418
R45954 vss.n768 vss.n767 0.0661418
R45955 vss.n768 vss.n762 0.0661418
R45956 vss.n13965 vss.n13964 0.0661418
R45957 vss.n13966 vss.n13965 0.0661418
R45958 vss.n776 vss.n775 0.0661418
R45959 vss.n776 vss.n680 0.0661418
R45960 vss.n757 vss.n756 0.0661418
R45961 vss.n756 vss.n751 0.0661418
R45962 vss.n752 vss.n746 0.0661418
R45963 vss.n752 vss.n750 0.0661418
R45964 vss.n789 vss.n761 0.0661418
R45965 vss.n790 vss.n789 0.0661418
R45966 vss.n785 vss.n780 0.0661418
R45967 vss.n780 vss.n779 0.0661418
R45968 vss.n13248 vss.n13247 0.0661418
R45969 vss.n13249 vss.n13248 0.0661418
R45970 vss.n1718 vss.n1717 0.0661418
R45971 vss.n1717 vss.n1715 0.0661418
R45972 vss.n1724 vss.n1723 0.0661418
R45973 vss.n1723 vss.n1721 0.0661418
R45974 vss.n1713 vss.n1710 0.0661418
R45975 vss.n1713 vss.n1706 0.0661418
R45976 vss.n1726 vss.n1725 0.0661418
R45977 vss.n1728 vss.n1726 0.0661418
R45978 vss.n1747 vss.n1746 0.0661418
R45979 vss.n1747 vss.n682 0.0661418
R45980 vss.n1754 vss.n1698 0.0661418
R45981 vss.n1754 vss.n1703 0.0661418
R45982 vss.n1759 vss.n1757 0.0661418
R45983 vss.n1757 vss.n1756 0.0661418
R45984 vss.n1797 vss.n1705 0.0661418
R45985 vss.n1798 vss.n1797 0.0661418
R45986 vss.n1793 vss.n1751 0.0661418
R45987 vss.n1751 vss.n1750 0.0661418
R45988 vss.n1780 vss.n1758 0.0661418
R45989 vss.n1758 vss.n740 0.0661418
R45990 vss.n1275 vss.n1274 0.0661418
R45991 vss.n1274 vss.n1272 0.0661418
R45992 vss.n1769 vss.n1766 0.0661418
R45993 vss.n1769 vss.n1768 0.0661418
R45994 vss.n1270 vss.n1267 0.0661418
R45995 vss.n1270 vss.n1263 0.0661418
R45996 vss.n1777 vss.n1776 0.0661418
R45997 vss.n1778 vss.n1777 0.0661418
R45998 vss.n1818 vss.n1817 0.0661418
R45999 vss.n1818 vss.n684 0.0661418
R46000 vss.n1251 vss.n1240 0.0661418
R46001 vss.n1827 vss.n1240 0.0661418
R46002 vss.n1253 vss.n1235 0.0661418
R46003 vss.n1235 vss.n1231 0.0661418
R46004 vss.n1249 vss.n1246 0.0661418
R46005 vss.n1249 vss.n1243 0.0661418
R46006 vss.n1248 vss.n1247 0.0661418
R46007 vss.n1821 vss.n1248 0.0661418
R46008 vss.n1254 vss.n1233 0.0661418
R46009 vss.n1233 vss.n737 0.0661418
R46010 vss.n1222 vss.n1221 0.0661418
R46011 vss.n1221 vss.n1219 0.0661418
R46012 vss.n1228 vss.n1227 0.0661418
R46013 vss.n1227 vss.n1225 0.0661418
R46014 vss.n1217 vss.n1214 0.0661418
R46015 vss.n1217 vss.n1210 0.0661418
R46016 vss.n1230 vss.n1229 0.0661418
R46017 vss.n1832 vss.n1230 0.0661418
R46018 vss.n1851 vss.n1850 0.0661418
R46019 vss.n1851 vss.n686 0.0661418
R46020 vss.n1858 vss.n1202 0.0661418
R46021 vss.n1858 vss.n1207 0.0661418
R46022 vss.n1863 vss.n1861 0.0661418
R46023 vss.n1861 vss.n1860 0.0661418
R46024 vss.n1901 vss.n1209 0.0661418
R46025 vss.n1902 vss.n1901 0.0661418
R46026 vss.n1897 vss.n1855 0.0661418
R46027 vss.n1855 vss.n1854 0.0661418
R46028 vss.n1884 vss.n1862 0.0661418
R46029 vss.n1862 vss.n734 0.0661418
R46030 vss.n1157 vss.n1156 0.0661418
R46031 vss.n1156 vss.n1154 0.0661418
R46032 vss.n1873 vss.n1870 0.0661418
R46033 vss.n1873 vss.n1872 0.0661418
R46034 vss.n1152 vss.n1149 0.0661418
R46035 vss.n1152 vss.n1145 0.0661418
R46036 vss.n1881 vss.n1880 0.0661418
R46037 vss.n1882 vss.n1881 0.0661418
R46038 vss.n1922 vss.n1921 0.0661418
R46039 vss.n1922 vss.n688 0.0661418
R46040 vss.n1929 vss.n1137 0.0661418
R46041 vss.n1929 vss.n1142 0.0661418
R46042 vss.n1934 vss.n1932 0.0661418
R46043 vss.n1932 vss.n1931 0.0661418
R46044 vss.n1972 vss.n1144 0.0661418
R46045 vss.n1973 vss.n1972 0.0661418
R46046 vss.n1968 vss.n1926 0.0661418
R46047 vss.n1926 vss.n1925 0.0661418
R46048 vss.n1955 vss.n1933 0.0661418
R46049 vss.n1933 vss.n731 0.0661418
R46050 vss.n703 vss.n702 0.0661418
R46051 vss.n702 vss.n697 0.0661418
R46052 vss.n1944 vss.n1941 0.0661418
R46053 vss.n1944 vss.n1943 0.0661418
R46054 vss.n700 vss.n693 0.0661418
R46055 vss.n700 vss.n698 0.0661418
R46056 vss.n1952 vss.n1951 0.0661418
R46057 vss.n1953 vss.n1952 0.0661418
R46058 vss.n13300 vss.n13299 0.0661418
R46059 vss.n13301 vss.n13300 0.0661418
R46060 vss.n720 vss.n707 0.0661418
R46061 vss.n720 vss.n712 0.0661418
R46062 vss.n725 vss.n723 0.0661418
R46063 vss.n723 vss.n722 0.0661418
R46064 vss.n13284 vss.n714 0.0661418
R46065 vss.n13285 vss.n13284 0.0661418
R46066 vss.n13280 vss.n717 0.0661418
R46067 vss.n717 vss.n716 0.0661418
R46068 vss.n13267 vss.n724 0.0661418
R46069 vss.n13266 vss.n724 0.0661418
R46070 vss.n13195 vss.n13194 0.0661418
R46071 vss.n13196 vss.n13195 0.0661418
R46072 vss.n13169 vss.n13159 0.0661418
R46073 vss.n13169 vss.n13164 0.0661418
R46074 vss.n13174 vss.n13172 0.0661418
R46075 vss.n13172 vss.n13171 0.0661418
R46076 vss.n13190 vss.n13187 0.0661418
R46077 vss.n13190 vss.n728 0.0661418
R46078 vss.n13177 vss.n13173 0.0661418
R46079 vss.n13173 vss.n812 0.0661418
R46080 vss.n1123 vss.n1122 0.0661418
R46081 vss.n1122 vss.n1101 0.0661418
R46082 vss.n1102 vss.n1095 0.0661418
R46083 vss.n1102 vss.n1100 0.0661418
R46084 vss.n1110 vss.n1108 0.0661418
R46085 vss.n1108 vss.n1107 0.0661418
R46086 vss.n1113 vss.n1109 0.0661418
R46087 vss.n1109 vss.n813 0.0661418
R46088 vss.n1127 vss.n1124 0.0661418
R46089 vss.n1127 vss.n730 0.0661418
R46090 vss.n1187 vss.n1186 0.0661418
R46091 vss.n1186 vss.n1165 0.0661418
R46092 vss.n1166 vss.n1159 0.0661418
R46093 vss.n1166 vss.n1164 0.0661418
R46094 vss.n1174 vss.n1172 0.0661418
R46095 vss.n1172 vss.n1171 0.0661418
R46096 vss.n1177 vss.n1173 0.0661418
R46097 vss.n1173 vss.n814 0.0661418
R46098 vss.n1191 vss.n1188 0.0661418
R46099 vss.n1191 vss.n733 0.0661418
R46100 vss.n1386 vss.n1385 0.0661418
R46101 vss.n1385 vss.n1364 0.0661418
R46102 vss.n1365 vss.n1358 0.0661418
R46103 vss.n1365 vss.n1363 0.0661418
R46104 vss.n1373 vss.n1371 0.0661418
R46105 vss.n1371 vss.n1370 0.0661418
R46106 vss.n1376 vss.n1372 0.0661418
R46107 vss.n1372 vss.n815 0.0661418
R46108 vss.n1390 vss.n1387 0.0661418
R46109 vss.n1390 vss.n736 0.0661418
R46110 vss.n1681 vss.n1680 0.0661418
R46111 vss.n1680 vss.n1659 0.0661418
R46112 vss.n1660 vss.n1653 0.0661418
R46113 vss.n1660 vss.n1658 0.0661418
R46114 vss.n1668 vss.n1666 0.0661418
R46115 vss.n1666 vss.n1665 0.0661418
R46116 vss.n1671 vss.n1667 0.0661418
R46117 vss.n1667 vss.n816 0.0661418
R46118 vss.n1685 vss.n1682 0.0661418
R46119 vss.n1685 vss.n739 0.0661418
R46120 vss.n13222 vss.n13221 0.0661418
R46121 vss.n13221 vss.n800 0.0661418
R46122 vss.n801 vss.n794 0.0661418
R46123 vss.n801 vss.n799 0.0661418
R46124 vss.n809 vss.n807 0.0661418
R46125 vss.n807 vss.n806 0.0661418
R46126 vss.n13212 vss.n808 0.0661418
R46127 vss.n13211 vss.n808 0.0661418
R46128 vss.n13226 vss.n13223 0.0661418
R46129 vss.n13226 vss.n742 0.0661418
R46130 vss.n607 vss.n606 0.0661418
R46131 vss.n606 vss.n601 0.0661418
R46132 vss.n602 vss.n595 0.0661418
R46133 vss.n602 vss.n600 0.0661418
R46134 vss.n824 vss.n821 0.0661418
R46135 vss.n824 vss.n823 0.0661418
R46136 vss.n832 vss.n831 0.0661418
R46137 vss.n833 vss.n832 0.0661418
R46138 vss.n13944 vss.n608 0.0661418
R46139 vss.n13944 vss.n13943 0.0661418
R46140 vss.n847 vss.n844 0.0661418
R46141 vss.n847 vss.n846 0.0661418
R46142 vss.n841 vss.n840 0.0661418
R46143 vss.n842 vss.n841 0.0661418
R46144 vss.n850 vss.n837 0.0661418
R46145 vss.n850 vss.n849 0.0661418
R46146 vss.n873 vss.n872 0.0661418
R46147 vss.n874 vss.n873 0.0661418
R46148 vss.n861 vss.n845 0.0661418
R46149 vss.n861 vss.n613 0.0661418
R46150 vss.n887 vss.n884 0.0661418
R46151 vss.n887 vss.n886 0.0661418
R46152 vss.n889 vss.n881 0.0661418
R46153 vss.n882 vss.n881 0.0661418
R46154 vss.n894 vss.n878 0.0661418
R46155 vss.n894 vss.n893 0.0661418
R46156 vss.n917 vss.n916 0.0661418
R46157 vss.n918 vss.n917 0.0661418
R46158 vss.n905 vss.n885 0.0661418
R46159 vss.n905 vss.n612 0.0661418
R46160 vss.n1551 vss.n1550 0.0661418
R46161 vss.n1550 vss.n1529 0.0661418
R46162 vss.n1530 vss.n1523 0.0661418
R46163 vss.n1530 vss.n1528 0.0661418
R46164 vss.n1538 vss.n1536 0.0661418
R46165 vss.n1536 vss.n1535 0.0661418
R46166 vss.n1541 vss.n1537 0.0661418
R46167 vss.n1537 vss.n919 0.0661418
R46168 vss.n1556 vss.n1552 0.0661418
R46169 vss.n1556 vss.n1555 0.0661418
R46170 vss.n1634 vss.n1633 0.0661418
R46171 vss.n1633 vss.n1612 0.0661418
R46172 vss.n1613 vss.n1606 0.0661418
R46173 vss.n1613 vss.n1611 0.0661418
R46174 vss.n1621 vss.n1619 0.0661418
R46175 vss.n1619 vss.n1618 0.0661418
R46176 vss.n1624 vss.n1620 0.0661418
R46177 vss.n1620 vss.n920 0.0661418
R46178 vss.n1638 vss.n1635 0.0661418
R46179 vss.n1638 vss.n741 0.0661418
R46180 vss.n1471 vss.n1470 0.0661418
R46181 vss.n1470 vss.n1449 0.0661418
R46182 vss.n1450 vss.n1443 0.0661418
R46183 vss.n1450 vss.n1448 0.0661418
R46184 vss.n1458 vss.n1456 0.0661418
R46185 vss.n1456 vss.n1455 0.0661418
R46186 vss.n1461 vss.n1457 0.0661418
R46187 vss.n1457 vss.n921 0.0661418
R46188 vss.n1475 vss.n1472 0.0661418
R46189 vss.n1475 vss.n738 0.0661418
R46190 vss.n1339 vss.n1338 0.0661418
R46191 vss.n1338 vss.n1317 0.0661418
R46192 vss.n1318 vss.n1311 0.0661418
R46193 vss.n1318 vss.n1316 0.0661418
R46194 vss.n1326 vss.n1324 0.0661418
R46195 vss.n1324 vss.n1323 0.0661418
R46196 vss.n1329 vss.n1325 0.0661418
R46197 vss.n1325 vss.n922 0.0661418
R46198 vss.n1343 vss.n1340 0.0661418
R46199 vss.n1343 vss.n735 0.0661418
R46200 vss.n1078 vss.n1077 0.0661418
R46201 vss.n1077 vss.n1056 0.0661418
R46202 vss.n1057 vss.n1050 0.0661418
R46203 vss.n1057 vss.n1055 0.0661418
R46204 vss.n1065 vss.n1063 0.0661418
R46205 vss.n1063 vss.n1062 0.0661418
R46206 vss.n1068 vss.n1064 0.0661418
R46207 vss.n1064 vss.n923 0.0661418
R46208 vss.n1082 vss.n1079 0.0661418
R46209 vss.n1082 vss.n732 0.0661418
R46210 vss.n2013 vss.n2012 0.0661418
R46211 vss.n2012 vss.n1991 0.0661418
R46212 vss.n1992 vss.n1985 0.0661418
R46213 vss.n1992 vss.n1990 0.0661418
R46214 vss.n2000 vss.n1998 0.0661418
R46215 vss.n1998 vss.n1997 0.0661418
R46216 vss.n2003 vss.n1999 0.0661418
R46217 vss.n1999 vss.n924 0.0661418
R46218 vss.n2017 vss.n2014 0.0661418
R46219 vss.n2017 vss.n729 0.0661418
R46220 vss.n9601 vss.n9599 0.0661418
R46221 vss.n9599 vss.n9598 0.0661418
R46222 vss.n9593 vss.n9586 0.0661418
R46223 vss.n9593 vss.n9591 0.0661418
R46224 vss.n9615 vss.n9614 0.0661418
R46225 vss.n9614 vss.n9592 0.0661418
R46226 vss.n9617 vss.n9616 0.0661418
R46227 vss.n9617 vss.n495 0.0661418
R46228 vss.n9605 vss.n9600 0.0661418
R46229 vss.n9604 vss.n9600 0.0661418
R46230 vss.n8023 vss.n8022 0.0661418
R46231 vss.n8023 vss.n8019 0.0661418
R46232 vss.n8028 vss.n8025 0.0661418
R46233 vss.n8028 vss.n8027 0.0661418
R46234 vss.n8020 vss.n8016 0.0661418
R46235 vss.n8020 vss.n8012 0.0661418
R46236 vss.n8015 vss.n8011 0.0661418
R46237 vss.n8051 vss.n8011 0.0661418
R46238 vss.n8035 vss.n8026 0.0661418
R46239 vss.n8035 vss.n7323 0.0661418
R46240 vss.n5983 vss.n5977 0.0661418
R46241 vss.n5983 vss.n5981 0.0661418
R46242 vss.n5988 vss.n5987 0.0661418
R46243 vss.n5987 vss.n5982 0.0661418
R46244 vss.n9655 vss.n9654 0.0661418
R46245 vss.n9656 vss.n9655 0.0661418
R46246 vss.n9650 vss.n5994 0.0661418
R46247 vss.n9650 vss.n9649 0.0661418
R46248 vss.n9667 vss.n9666 0.0661418
R46249 vss.n9668 vss.n9667 0.0661418
R46250 vss.n8126 vss.n6002 0.0661418
R46251 vss.n8129 vss.n8126 0.0661418
R46252 vss.n8134 vss.n8131 0.0661418
R46253 vss.n8131 vss.n8130 0.0661418
R46254 vss.n9646 vss.n5998 0.0661418
R46255 vss.n9647 vss.n9646 0.0661418
R46256 vss.n8151 vss.n8150 0.0661418
R46257 vss.n8152 vss.n8151 0.0661418
R46258 vss.n8138 vss.n8132 0.0661418
R46259 vss.n8132 vss.n8052 0.0661418
R46260 vss.n8121 vss.n8120 0.0661418
R46261 vss.n8123 vss.n8121 0.0661418
R46262 vss.n7277 vss.n7271 0.0661418
R46263 vss.n7277 vss.n7275 0.0661418
R46264 vss.n7282 vss.n7281 0.0661418
R46265 vss.n7281 vss.n7276 0.0661418
R46266 vss.n9024 vss.n9023 0.0661418
R46267 vss.n9025 vss.n9024 0.0661418
R46268 vss.n9019 vss.n7288 0.0661418
R46269 vss.n9019 vss.n9018 0.0661418
R46270 vss.n9010 vss.n7295 0.0661418
R46271 vss.n9010 vss.n9009 0.0661418
R46272 vss.n8265 vss.n7903 0.0661418
R46273 vss.n8265 vss.n8263 0.0661418
R46274 vss.n8270 vss.n8269 0.0661418
R46275 vss.n8269 vss.n8264 0.0661418
R46276 vss.n9015 vss.n9014 0.0661418
R46277 vss.n9016 vss.n9015 0.0661418
R46278 vss.n8281 vss.n8280 0.0661418
R46279 vss.n8282 vss.n8281 0.0661418
R46280 vss.n7899 vss.n7898 0.0661418
R46281 vss.n7899 vss.n6574 0.0661418
R46282 vss.n7897 vss.n7896 0.0661418
R46283 vss.n7896 vss.n7894 0.0661418
R46284 vss.n7891 vss.n7890 0.0661418
R46285 vss.n7890 vss.n7885 0.0661418
R46286 vss.n7888 vss.n7881 0.0661418
R46287 vss.n7888 vss.n7886 0.0661418
R46288 vss.n8302 vss.n8301 0.0661418
R46289 vss.n8303 vss.n8302 0.0661418
R46290 vss.n8708 vss.n8707 0.0661418
R46291 vss.n8709 vss.n8708 0.0661418
R46292 vss.n8316 vss.n8315 0.0661418
R46293 vss.n8315 vss.n8313 0.0661418
R46294 vss.n8310 vss.n8309 0.0661418
R46295 vss.n8309 vss.n7877 0.0661418
R46296 vss.n8307 vss.n7870 0.0661418
R46297 vss.n8307 vss.n8305 0.0661418
R46298 vss.n8318 vss.n8317 0.0661418
R46299 vss.n8689 vss.n8318 0.0661418
R46300 vss.n8325 vss.n8322 0.0661418
R46301 vss.n8325 vss.n6572 0.0661418
R46302 vss.n8686 vss.n8685 0.0661418
R46303 vss.n8687 vss.n8686 0.0661418
R46304 vss.n8338 vss.n8331 0.0661418
R46305 vss.n8334 vss.n8331 0.0661418
R46306 vss.n8343 vss.n8342 0.0661418
R46307 vss.n8342 vss.n8335 0.0661418
R46308 vss.n8345 vss.n8344 0.0661418
R46309 vss.n8674 vss.n8345 0.0661418
R46310 vss.n8666 vss.n8663 0.0661418
R46311 vss.n8666 vss.n7681 0.0661418
R46312 vss.n8361 vss.n8360 0.0661418
R46313 vss.n8360 vss.n8356 0.0661418
R46314 vss.n8653 vss.n8353 0.0661418
R46315 vss.n8357 vss.n8353 0.0661418
R46316 vss.n8671 vss.n8670 0.0661418
R46317 vss.n8672 vss.n8671 0.0661418
R46318 vss.n8363 vss.n8362 0.0661418
R46319 vss.n8646 vss.n8363 0.0661418
R46320 vss.n8370 vss.n8367 0.0661418
R46321 vss.n8370 vss.n6570 0.0661418
R46322 vss.n8643 vss.n8642 0.0661418
R46323 vss.n8644 vss.n8643 0.0661418
R46324 vss.n8388 vss.n8381 0.0661418
R46325 vss.n8384 vss.n8381 0.0661418
R46326 vss.n8393 vss.n8392 0.0661418
R46327 vss.n8392 vss.n8385 0.0661418
R46328 vss.n8395 vss.n8394 0.0661418
R46329 vss.n8631 vss.n8395 0.0661418
R46330 vss.n8623 vss.n8619 0.0661418
R46331 vss.n8623 vss.n8622 0.0661418
R46332 vss.n8414 vss.n8413 0.0661418
R46333 vss.n8413 vss.n8409 0.0661418
R46334 vss.n8609 vss.n8406 0.0661418
R46335 vss.n8410 vss.n8406 0.0661418
R46336 vss.n8628 vss.n8627 0.0661418
R46337 vss.n8629 vss.n8628 0.0661418
R46338 vss.n8416 vss.n8415 0.0661418
R46339 vss.n8602 vss.n8416 0.0661418
R46340 vss.n8423 vss.n8420 0.0661418
R46341 vss.n8423 vss.n6568 0.0661418
R46342 vss.n8599 vss.n8598 0.0661418
R46343 vss.n8600 vss.n8599 0.0661418
R46344 vss.n8436 vss.n8429 0.0661418
R46345 vss.n8432 vss.n8429 0.0661418
R46346 vss.n8441 vss.n8440 0.0661418
R46347 vss.n8440 vss.n8433 0.0661418
R46348 vss.n8443 vss.n8442 0.0661418
R46349 vss.n8587 vss.n8443 0.0661418
R46350 vss.n8579 vss.n8576 0.0661418
R46351 vss.n8579 vss.n7538 0.0661418
R46352 vss.n8459 vss.n8458 0.0661418
R46353 vss.n8458 vss.n8454 0.0661418
R46354 vss.n8566 vss.n8451 0.0661418
R46355 vss.n8455 vss.n8451 0.0661418
R46356 vss.n8584 vss.n8583 0.0661418
R46357 vss.n8585 vss.n8584 0.0661418
R46358 vss.n8461 vss.n8460 0.0661418
R46359 vss.n8559 vss.n8461 0.0661418
R46360 vss.n8468 vss.n8465 0.0661418
R46361 vss.n8468 vss.n6556 0.0661418
R46362 vss.n8556 vss.n8555 0.0661418
R46363 vss.n8557 vss.n8556 0.0661418
R46364 vss.n8486 vss.n8479 0.0661418
R46365 vss.n8482 vss.n8479 0.0661418
R46366 vss.n8491 vss.n8490 0.0661418
R46367 vss.n8490 vss.n8483 0.0661418
R46368 vss.n8493 vss.n8492 0.0661418
R46369 vss.n8544 vss.n8493 0.0661418
R46370 vss.n8514 vss.n8504 0.0661418
R46371 vss.n8506 vss.n8504 0.0661418
R46372 vss.n8541 vss.n8540 0.0661418
R46373 vss.n8542 vss.n8541 0.0661418
R46374 vss.n8512 vss.n8507 0.0661418
R46375 vss.n8512 vss.n8511 0.0661418
R46376 vss.n8509 vss.n8508 0.0661418
R46377 vss.n8510 vss.n8509 0.0661418
R46378 vss.n8536 vss.n8532 0.0661418
R46379 vss.n8536 vss.n8535 0.0661418
R46380 vss.n6068 vss.n6056 0.0661418
R46381 vss.n6068 vss.n6061 0.0661418
R46382 vss.n6073 vss.n6071 0.0661418
R46383 vss.n6071 vss.n6070 0.0661418
R46384 vss.n9569 vss.n6063 0.0661418
R46385 vss.n9570 vss.n9569 0.0661418
R46386 vss.n9565 vss.n6065 0.0661418
R46387 vss.n6065 vss.n6064 0.0661418
R46388 vss.n9552 vss.n6072 0.0661418
R46389 vss.n6076 vss.n6072 0.0661418
R46390 vss.n6091 vss.n6090 0.0661418
R46391 vss.n6090 vss.n6085 0.0661418
R46392 vss.n6086 vss.n6080 0.0661418
R46393 vss.n6086 vss.n6084 0.0661418
R46394 vss.n7257 vss.n7252 0.0661418
R46395 vss.n7257 vss.n7256 0.0661418
R46396 vss.n9549 vss.n9548 0.0661418
R46397 vss.n9550 vss.n9549 0.0661418
R46398 vss.n7265 vss.n7264 0.0661418
R46399 vss.n7266 vss.n7265 0.0661418
R46400 vss.n6107 vss.n6096 0.0661418
R46401 vss.n6107 vss.n6101 0.0661418
R46402 vss.n6112 vss.n6110 0.0661418
R46403 vss.n6110 vss.n6109 0.0661418
R46404 vss.n9534 vss.n6103 0.0661418
R46405 vss.n9535 vss.n9534 0.0661418
R46406 vss.n9530 vss.n6104 0.0661418
R46407 vss.n7254 vss.n6104 0.0661418
R46408 vss.n9517 vss.n6111 0.0661418
R46409 vss.n6115 vss.n6111 0.0661418
R46410 vss.n6130 vss.n6129 0.0661418
R46411 vss.n6129 vss.n6124 0.0661418
R46412 vss.n6125 vss.n6119 0.0661418
R46413 vss.n6125 vss.n6123 0.0661418
R46414 vss.n7238 vss.n6579 0.0661418
R46415 vss.n7238 vss.n7237 0.0661418
R46416 vss.n9514 vss.n9513 0.0661418
R46417 vss.n9515 vss.n9514 0.0661418
R46418 vss.n7246 vss.n7245 0.0661418
R46419 vss.n7247 vss.n7246 0.0661418
R46420 vss.n6594 vss.n6593 0.0661418
R46421 vss.n6593 vss.n6588 0.0661418
R46422 vss.n6754 vss.n6751 0.0661418
R46423 vss.n6751 vss.n6747 0.0661418
R46424 vss.n6591 vss.n6584 0.0661418
R46425 vss.n6591 vss.n6589 0.0661418
R46426 vss.n7234 vss.n7233 0.0661418
R46427 vss.n7235 vss.n7234 0.0661418
R46428 vss.n6755 vss.n6749 0.0661418
R46429 vss.n6749 vss.n6169 0.0661418
R46430 vss.n6738 vss.n6737 0.0661418
R46431 vss.n6737 vss.n6735 0.0661418
R46432 vss.n6744 vss.n6743 0.0661418
R46433 vss.n6743 vss.n6741 0.0661418
R46434 vss.n6733 vss.n6730 0.0661418
R46435 vss.n6733 vss.n6726 0.0661418
R46436 vss.n6746 vss.n6745 0.0661418
R46437 vss.n6764 vss.n6746 0.0661418
R46438 vss.n6783 vss.n6782 0.0661418
R46439 vss.n6783 vss.n6573 0.0661418
R46440 vss.n6790 vss.n6718 0.0661418
R46441 vss.n6790 vss.n6723 0.0661418
R46442 vss.n6795 vss.n6793 0.0661418
R46443 vss.n6793 vss.n6792 0.0661418
R46444 vss.n7079 vss.n6725 0.0661418
R46445 vss.n7080 vss.n7079 0.0661418
R46446 vss.n7075 vss.n6787 0.0661418
R46447 vss.n6787 vss.n6786 0.0661418
R46448 vss.n7062 vss.n6794 0.0661418
R46449 vss.n6794 vss.n6172 0.0661418
R46450 vss.n6812 vss.n6811 0.0661418
R46451 vss.n6811 vss.n6806 0.0661418
R46452 vss.n6807 vss.n6801 0.0661418
R46453 vss.n6807 vss.n6805 0.0661418
R46454 vss.n6820 vss.n6816 0.0661418
R46455 vss.n7046 vss.n6816 0.0661418
R46456 vss.n7059 vss.n7058 0.0661418
R46457 vss.n7060 vss.n7059 0.0661418
R46458 vss.n6825 vss.n6824 0.0661418
R46459 vss.n6825 vss.n6571 0.0661418
R46460 vss.n6840 vss.n6839 0.0661418
R46461 vss.n6839 vss.n6834 0.0661418
R46462 vss.n6846 vss.n6845 0.0661418
R46463 vss.n6845 vss.n6843 0.0661418
R46464 vss.n6837 vss.n6830 0.0661418
R46465 vss.n6837 vss.n6835 0.0661418
R46466 vss.n7043 vss.n7042 0.0661418
R46467 vss.n7044 vss.n7043 0.0661418
R46468 vss.n6848 vss.n6847 0.0661418
R46469 vss.n6848 vss.n6175 0.0661418
R46470 vss.n6863 vss.n6862 0.0661418
R46471 vss.n6862 vss.n6857 0.0661418
R46472 vss.n6858 vss.n6852 0.0661418
R46473 vss.n6858 vss.n6856 0.0661418
R46474 vss.n6871 vss.n6867 0.0661418
R46475 vss.n6880 vss.n6867 0.0661418
R46476 vss.n6891 vss.n6890 0.0661418
R46477 vss.n6892 vss.n6891 0.0661418
R46478 vss.n6876 vss.n6875 0.0661418
R46479 vss.n6876 vss.n6569 0.0661418
R46480 vss.n6501 vss.n6490 0.0661418
R46481 vss.n6501 vss.n6495 0.0661418
R46482 vss.n6506 vss.n6504 0.0661418
R46483 vss.n6504 vss.n6503 0.0661418
R46484 vss.n9242 vss.n6497 0.0661418
R46485 vss.n9243 vss.n9242 0.0661418
R46486 vss.n9238 vss.n6498 0.0661418
R46487 vss.n6878 vss.n6498 0.0661418
R46488 vss.n9225 vss.n6505 0.0661418
R46489 vss.n6505 vss.n6178 0.0661418
R46490 vss.n6523 vss.n6522 0.0661418
R46491 vss.n6522 vss.n6517 0.0661418
R46492 vss.n6518 vss.n6512 0.0661418
R46493 vss.n6518 vss.n6516 0.0661418
R46494 vss.n6561 vss.n6527 0.0661418
R46495 vss.n9209 vss.n6527 0.0661418
R46496 vss.n9222 vss.n9221 0.0661418
R46497 vss.n9223 vss.n9222 0.0661418
R46498 vss.n6566 vss.n6565 0.0661418
R46499 vss.n6567 vss.n6566 0.0661418
R46500 vss.n6541 vss.n6540 0.0661418
R46501 vss.n6540 vss.n6535 0.0661418
R46502 vss.n9072 vss.n9069 0.0661418
R46503 vss.n9069 vss.n9065 0.0661418
R46504 vss.n6538 vss.n6531 0.0661418
R46505 vss.n6538 vss.n6536 0.0661418
R46506 vss.n9206 vss.n9205 0.0661418
R46507 vss.n9207 vss.n9206 0.0661418
R46508 vss.n9073 vss.n9067 0.0661418
R46509 vss.n9067 vss.n6181 0.0661418
R46510 vss.n9057 vss.n6547 0.0661418
R46511 vss.n9057 vss.n6552 0.0661418
R46512 vss.n9062 vss.n9060 0.0661418
R46513 vss.n9060 vss.n9059 0.0661418
R46514 vss.n9054 vss.n6554 0.0661418
R46515 vss.n9141 vss.n6554 0.0661418
R46516 vss.n9083 vss.n9061 0.0661418
R46517 vss.n9082 vss.n9061 0.0661418
R46518 vss.n9096 vss.n9095 0.0661418
R46519 vss.n9096 vss.n9050 0.0661418
R46520 vss.n9111 vss.n9110 0.0661418
R46521 vss.n9110 vss.n9105 0.0661418
R46522 vss.n9117 vss.n9116 0.0661418
R46523 vss.n9116 vss.n9114 0.0661418
R46524 vss.n9108 vss.n9101 0.0661418
R46525 vss.n9108 vss.n9106 0.0661418
R46526 vss.n9138 vss.n9137 0.0661418
R46527 vss.n9139 vss.n9138 0.0661418
R46528 vss.n9119 vss.n9118 0.0661418
R46529 vss.n9119 vss.n6184 0.0661418
R46530 vss.n9374 vss.n6188 0.0661418
R46531 vss.n9374 vss.n9373 0.0661418
R46532 vss.n6196 vss.n6192 0.0661418
R46533 vss.n6197 vss.n6196 0.0661418
R46534 vss.n6200 vss.n6199 0.0661418
R46535 vss.n6199 vss.n6195 0.0661418
R46536 vss.n6202 vss.n6201 0.0661418
R46537 vss.n6203 vss.n6202 0.0661418
R46538 vss.n9381 vss.n9380 0.0661418
R46539 vss.n9382 vss.n9381 0.0661418
R46540 vss.n9179 vss.n9178 0.0661418
R46541 vss.n9178 vss.n9156 0.0661418
R46542 vss.n9157 vss.n9150 0.0661418
R46543 vss.n9157 vss.n9155 0.0661418
R46544 vss.n9165 vss.n9163 0.0661418
R46545 vss.n9163 vss.n9162 0.0661418
R46546 vss.n9169 vss.n9164 0.0661418
R46547 vss.n9168 vss.n9164 0.0661418
R46548 vss.n9183 vss.n9180 0.0661418
R46549 vss.n9183 vss.n6182 0.0661418
R46550 vss.n6476 vss.n6475 0.0661418
R46551 vss.n6475 vss.n6453 0.0661418
R46552 vss.n6454 vss.n6447 0.0661418
R46553 vss.n6454 vss.n6452 0.0661418
R46554 vss.n6462 vss.n6460 0.0661418
R46555 vss.n6460 vss.n6459 0.0661418
R46556 vss.n6466 vss.n6461 0.0661418
R46557 vss.n6465 vss.n6461 0.0661418
R46558 vss.n6480 vss.n6477 0.0661418
R46559 vss.n6480 vss.n6179 0.0661418
R46560 vss.n7016 vss.n7015 0.0661418
R46561 vss.n7015 vss.n6993 0.0661418
R46562 vss.n6994 vss.n6987 0.0661418
R46563 vss.n6994 vss.n6992 0.0661418
R46564 vss.n7002 vss.n7000 0.0661418
R46565 vss.n7000 vss.n6999 0.0661418
R46566 vss.n7006 vss.n7001 0.0661418
R46567 vss.n7005 vss.n7001 0.0661418
R46568 vss.n7020 vss.n7017 0.0661418
R46569 vss.n7020 vss.n6176 0.0661418
R46570 vss.n6702 vss.n6701 0.0661418
R46571 vss.n6701 vss.n6679 0.0661418
R46572 vss.n6680 vss.n6673 0.0661418
R46573 vss.n6680 vss.n6678 0.0661418
R46574 vss.n6688 vss.n6686 0.0661418
R46575 vss.n6686 vss.n6685 0.0661418
R46576 vss.n6692 vss.n6687 0.0661418
R46577 vss.n6691 vss.n6687 0.0661418
R46578 vss.n6706 vss.n6703 0.0661418
R46579 vss.n6706 vss.n6173 0.0661418
R46580 vss.n7207 vss.n7206 0.0661418
R46581 vss.n7206 vss.n7184 0.0661418
R46582 vss.n7185 vss.n7178 0.0661418
R46583 vss.n7185 vss.n7183 0.0661418
R46584 vss.n7193 vss.n7191 0.0661418
R46585 vss.n7191 vss.n7190 0.0661418
R46586 vss.n7197 vss.n7192 0.0661418
R46587 vss.n7196 vss.n7192 0.0661418
R46588 vss.n7211 vss.n7208 0.0661418
R46589 vss.n7211 vss.n6170 0.0661418
R46590 vss.n6164 vss.n6163 0.0661418
R46591 vss.n6163 vss.n6141 0.0661418
R46592 vss.n6142 vss.n6135 0.0661418
R46593 vss.n6142 vss.n6140 0.0661418
R46594 vss.n6150 vss.n6148 0.0661418
R46595 vss.n6148 vss.n6147 0.0661418
R46596 vss.n6154 vss.n6149 0.0661418
R46597 vss.n6153 vss.n6149 0.0661418
R46598 vss.n9493 vss.n6165 0.0661418
R46599 vss.n9493 vss.n9492 0.0661418
R46600 vss.n9478 vss.n9448 0.0661418
R46601 vss.n9478 vss.n9477 0.0661418
R46602 vss.n9452 vss.n9451 0.0661418
R46603 vss.n9456 vss.n9452 0.0661418
R46604 vss.n9459 vss.n9458 0.0661418
R46605 vss.n9458 vss.n9455 0.0661418
R46606 vss.n9461 vss.n9460 0.0661418
R46607 vss.n9462 vss.n9461 0.0661418
R46608 vss.n9485 vss.n9484 0.0661418
R46609 vss.n9486 vss.n9485 0.0661418
R46610 vss.n6037 vss.n6036 0.0661418
R46611 vss.n6036 vss.n6014 0.0661418
R46612 vss.n6015 vss.n6008 0.0661418
R46613 vss.n6015 vss.n6013 0.0661418
R46614 vss.n6023 vss.n6021 0.0661418
R46615 vss.n6021 vss.n6020 0.0661418
R46616 vss.n6027 vss.n6022 0.0661418
R46617 vss.n6026 vss.n6022 0.0661418
R46618 vss.n6042 vss.n6038 0.0661418
R46619 vss.n6042 vss.n6041 0.0661418
R46620 vss.n9436 vss.n9403 0.0661418
R46621 vss.n9436 vss.n9435 0.0661418
R46622 vss.n9411 vss.n9407 0.0661418
R46623 vss.n9412 vss.n9411 0.0661418
R46624 vss.n9415 vss.n9414 0.0661418
R46625 vss.n9414 vss.n9410 0.0661418
R46626 vss.n9417 vss.n9416 0.0661418
R46627 vss.n9418 vss.n9417 0.0661418
R46628 vss.n9443 vss.n9442 0.0661418
R46629 vss.n9444 vss.n9443 0.0661418
R46630 vss.n7156 vss.n7155 0.0661418
R46631 vss.n7155 vss.n7133 0.0661418
R46632 vss.n7134 vss.n7127 0.0661418
R46633 vss.n7134 vss.n7132 0.0661418
R46634 vss.n7142 vss.n7140 0.0661418
R46635 vss.n7140 vss.n7139 0.0661418
R46636 vss.n7146 vss.n7141 0.0661418
R46637 vss.n7145 vss.n7141 0.0661418
R46638 vss.n7160 vss.n7157 0.0661418
R46639 vss.n7160 vss.n6168 0.0661418
R46640 vss.n6658 vss.n6657 0.0661418
R46641 vss.n6657 vss.n6635 0.0661418
R46642 vss.n6636 vss.n6629 0.0661418
R46643 vss.n6636 vss.n6634 0.0661418
R46644 vss.n6644 vss.n6642 0.0661418
R46645 vss.n6642 vss.n6641 0.0661418
R46646 vss.n6648 vss.n6643 0.0661418
R46647 vss.n6647 vss.n6643 0.0661418
R46648 vss.n6662 vss.n6659 0.0661418
R46649 vss.n6662 vss.n6171 0.0661418
R46650 vss.n6967 vss.n6966 0.0661418
R46651 vss.n6966 vss.n6944 0.0661418
R46652 vss.n6945 vss.n6938 0.0661418
R46653 vss.n6945 vss.n6943 0.0661418
R46654 vss.n6953 vss.n6951 0.0661418
R46655 vss.n6951 vss.n6950 0.0661418
R46656 vss.n6957 vss.n6952 0.0661418
R46657 vss.n6956 vss.n6952 0.0661418
R46658 vss.n6971 vss.n6968 0.0661418
R46659 vss.n6971 vss.n6174 0.0661418
R46660 vss.n6431 vss.n6430 0.0661418
R46661 vss.n6430 vss.n6408 0.0661418
R46662 vss.n6409 vss.n6402 0.0661418
R46663 vss.n6409 vss.n6407 0.0661418
R46664 vss.n6417 vss.n6415 0.0661418
R46665 vss.n6415 vss.n6414 0.0661418
R46666 vss.n6421 vss.n6416 0.0661418
R46667 vss.n6420 vss.n6416 0.0661418
R46668 vss.n6435 vss.n6432 0.0661418
R46669 vss.n6435 vss.n6177 0.0661418
R46670 vss.n6353 vss.n6352 0.0661418
R46671 vss.n6352 vss.n6330 0.0661418
R46672 vss.n6331 vss.n6324 0.0661418
R46673 vss.n6331 vss.n6329 0.0661418
R46674 vss.n6339 vss.n6337 0.0661418
R46675 vss.n6337 vss.n6336 0.0661418
R46676 vss.n6343 vss.n6338 0.0661418
R46677 vss.n6342 vss.n6338 0.0661418
R46678 vss.n6357 vss.n6354 0.0661418
R46679 vss.n6357 vss.n6180 0.0661418
R46680 vss.n9349 vss.n9348 0.0661418
R46681 vss.n9348 vss.n9326 0.0661418
R46682 vss.n9327 vss.n9320 0.0661418
R46683 vss.n9327 vss.n9325 0.0661418
R46684 vss.n9335 vss.n9333 0.0661418
R46685 vss.n9333 vss.n9332 0.0661418
R46686 vss.n9339 vss.n9334 0.0661418
R46687 vss.n9338 vss.n9334 0.0661418
R46688 vss.n9353 vss.n9350 0.0661418
R46689 vss.n9353 vss.n6183 0.0661418
R46690 vss.n5952 vss.n5950 0.0661418
R46691 vss.n5950 vss.n5949 0.0661418
R46692 vss.n5944 vss.n5937 0.0661418
R46693 vss.n5944 vss.n5942 0.0661418
R46694 vss.n5965 vss.n5964 0.0661418
R46695 vss.n5964 vss.n5943 0.0661418
R46696 vss.n5967 vss.n5966 0.0661418
R46697 vss.n9673 vss.n5967 0.0661418
R46698 vss.n5955 vss.n5951 0.0661418
R46699 vss.n5951 vss.n2784 0.0661418
R46700 vss.n2573 vss.n2571 0.0661418
R46701 vss.n2571 vss.n2570 0.0661418
R46702 vss.n2565 vss.n2558 0.0661418
R46703 vss.n2565 vss.n2563 0.0661418
R46704 vss.n2586 vss.n2585 0.0661418
R46705 vss.n2585 vss.n2564 0.0661418
R46706 vss.n2588 vss.n2587 0.0661418
R46707 vss.n10001 vss.n2588 0.0661418
R46708 vss.n2576 vss.n2572 0.0661418
R46709 vss.n2572 vss.n2160 0.0661418
R46710 vss.n9757 vss.n9744 0.0661418
R46711 vss.n9758 vss.n9757 0.0661418
R46712 vss.n9751 vss.n9748 0.0661418
R46713 vss.n9749 vss.n9748 0.0661418
R46714 vss.n9764 vss.n9759 0.0661418
R46715 vss.n9759 vss.n9756 0.0661418
R46716 vss.n9763 vss.n9760 0.0661418
R46717 vss.n9760 vss.n2740 0.0661418
R46718 vss.n9778 vss.n9750 0.0661418
R46719 vss.n9750 vss.n2768 0.0661418
R46720 vss.n3197 vss.n3184 0.0661418
R46721 vss.n3198 vss.n3197 0.0661418
R46722 vss.n3191 vss.n3188 0.0661418
R46723 vss.n3189 vss.n3188 0.0661418
R46724 vss.n3204 vss.n3199 0.0661418
R46725 vss.n3199 vss.n3196 0.0661418
R46726 vss.n3203 vss.n3200 0.0661418
R46727 vss.n3200 vss.n2741 0.0661418
R46728 vss.n3218 vss.n3190 0.0661418
R46729 vss.n3190 vss.n2769 0.0661418
R46730 vss.n3008 vss.n3007 0.0661418
R46731 vss.n3007 vss.n3001 0.0661418
R46732 vss.n3013 vss.n3010 0.0661418
R46733 vss.n3011 vss.n3010 0.0661418
R46734 vss.n3002 vss.n2998 0.0661418
R46735 vss.n3002 vss.n2994 0.0661418
R46736 vss.n2997 vss.n2993 0.0661418
R46737 vss.n9802 vss.n2993 0.0661418
R46738 vss.n3020 vss.n3012 0.0661418
R46739 vss.n3012 vss.n2770 0.0661418
R46740 vss.n5227 vss.n5214 0.0661418
R46741 vss.n5228 vss.n5227 0.0661418
R46742 vss.n5221 vss.n5218 0.0661418
R46743 vss.n5219 vss.n5218 0.0661418
R46744 vss.n5234 vss.n5229 0.0661418
R46745 vss.n5229 vss.n5226 0.0661418
R46746 vss.n5233 vss.n5230 0.0661418
R46747 vss.n5230 vss.n2990 0.0661418
R46748 vss.n5248 vss.n5220 0.0661418
R46749 vss.n5220 vss.n2771 0.0661418
R46750 vss.n3040 vss.n3027 0.0661418
R46751 vss.n3041 vss.n3040 0.0661418
R46752 vss.n3034 vss.n3031 0.0661418
R46753 vss.n3032 vss.n3031 0.0661418
R46754 vss.n3047 vss.n3042 0.0661418
R46755 vss.n3042 vss.n3039 0.0661418
R46756 vss.n3046 vss.n3043 0.0661418
R46757 vss.n3043 vss.n2991 0.0661418
R46758 vss.n3061 vss.n3033 0.0661418
R46759 vss.n3033 vss.n2772 0.0661418
R46760 vss.n5097 vss.n5084 0.0661418
R46761 vss.n5098 vss.n5097 0.0661418
R46762 vss.n5091 vss.n5088 0.0661418
R46763 vss.n5089 vss.n5088 0.0661418
R46764 vss.n5104 vss.n5099 0.0661418
R46765 vss.n5099 vss.n5096 0.0661418
R46766 vss.n5103 vss.n5100 0.0661418
R46767 vss.n5100 vss.n2987 0.0661418
R46768 vss.n5118 vss.n5090 0.0661418
R46769 vss.n5090 vss.n2773 0.0661418
R46770 vss.n5286 vss.n5273 0.0661418
R46771 vss.n5287 vss.n5286 0.0661418
R46772 vss.n5280 vss.n5277 0.0661418
R46773 vss.n5278 vss.n5277 0.0661418
R46774 vss.n5293 vss.n5288 0.0661418
R46775 vss.n5288 vss.n5285 0.0661418
R46776 vss.n5292 vss.n5289 0.0661418
R46777 vss.n5289 vss.n2984 0.0661418
R46778 vss.n5307 vss.n5279 0.0661418
R46779 vss.n5279 vss.n2774 0.0661418
R46780 vss.n5014 vss.n5001 0.0661418
R46781 vss.n5015 vss.n5014 0.0661418
R46782 vss.n5008 vss.n5005 0.0661418
R46783 vss.n5006 vss.n5005 0.0661418
R46784 vss.n5021 vss.n5016 0.0661418
R46785 vss.n5016 vss.n5013 0.0661418
R46786 vss.n5020 vss.n5017 0.0661418
R46787 vss.n5017 vss.n2985 0.0661418
R46788 vss.n5035 vss.n5007 0.0661418
R46789 vss.n5007 vss.n2775 0.0661418
R46790 vss.n4895 vss.n4882 0.0661418
R46791 vss.n4896 vss.n4895 0.0661418
R46792 vss.n4889 vss.n4886 0.0661418
R46793 vss.n4887 vss.n4886 0.0661418
R46794 vss.n4902 vss.n4897 0.0661418
R46795 vss.n4897 vss.n4894 0.0661418
R46796 vss.n4901 vss.n4898 0.0661418
R46797 vss.n4898 vss.n2981 0.0661418
R46798 vss.n4916 vss.n4888 0.0661418
R46799 vss.n4888 vss.n2776 0.0661418
R46800 vss.n2718 vss.n2712 0.0661418
R46801 vss.n2718 vss.n2716 0.0661418
R46802 vss.n2723 vss.n2722 0.0661418
R46803 vss.n2722 vss.n2717 0.0661418
R46804 vss.n9916 vss.n9915 0.0661418
R46805 vss.n9917 vss.n9916 0.0661418
R46806 vss.n9911 vss.n2729 0.0661418
R46807 vss.n9911 vss.n9910 0.0661418
R46808 vss.n9902 vss.n2736 0.0661418
R46809 vss.n9902 vss.n9901 0.0661418
R46810 vss.n4649 vss.n4640 0.0661418
R46811 vss.n4649 vss.n4647 0.0661418
R46812 vss.n4654 vss.n4653 0.0661418
R46813 vss.n4653 vss.n4648 0.0661418
R46814 vss.n9907 vss.n9906 0.0661418
R46815 vss.n9908 vss.n9907 0.0661418
R46816 vss.n4665 vss.n4664 0.0661418
R46817 vss.n4666 vss.n4665 0.0661418
R46818 vss.n5630 vss.n5629 0.0661418
R46819 vss.n5631 vss.n5630 0.0661418
R46820 vss.n4670 vss.n4631 0.0661418
R46821 vss.n4670 vss.n4668 0.0661418
R46822 vss.n4675 vss.n4674 0.0661418
R46823 vss.n4674 vss.n4669 0.0661418
R46824 vss.n5618 vss.n5617 0.0661418
R46825 vss.n5619 vss.n5618 0.0661418
R46826 vss.n5613 vss.n4681 0.0661418
R46827 vss.n5613 vss.n5612 0.0661418
R46828 vss.n5604 vss.n5601 0.0661418
R46829 vss.n5604 vss.n2992 0.0661418
R46830 vss.n4696 vss.n4695 0.0661418
R46831 vss.n4695 vss.n4691 0.0661418
R46832 vss.n5591 vss.n4688 0.0661418
R46833 vss.n4692 vss.n4688 0.0661418
R46834 vss.n5609 vss.n5608 0.0661418
R46835 vss.n5610 vss.n5609 0.0661418
R46836 vss.n4698 vss.n4697 0.0661418
R46837 vss.n5584 vss.n4698 0.0661418
R46838 vss.n4705 vss.n4702 0.0661418
R46839 vss.n4705 vss.n3630 0.0661418
R46840 vss.n5581 vss.n5580 0.0661418
R46841 vss.n5582 vss.n5581 0.0661418
R46842 vss.n4716 vss.n4709 0.0661418
R46843 vss.n4712 vss.n4709 0.0661418
R46844 vss.n4721 vss.n4720 0.0661418
R46845 vss.n4720 vss.n4713 0.0661418
R46846 vss.n4723 vss.n4722 0.0661418
R46847 vss.n5569 vss.n4723 0.0661418
R46848 vss.n5561 vss.n5558 0.0661418
R46849 vss.n5561 vss.n2989 0.0661418
R46850 vss.n4739 vss.n4738 0.0661418
R46851 vss.n4738 vss.n4734 0.0661418
R46852 vss.n5548 vss.n4731 0.0661418
R46853 vss.n4735 vss.n4731 0.0661418
R46854 vss.n5566 vss.n5565 0.0661418
R46855 vss.n5567 vss.n5566 0.0661418
R46856 vss.n4741 vss.n4740 0.0661418
R46857 vss.n5541 vss.n4741 0.0661418
R46858 vss.n4748 vss.n4745 0.0661418
R46859 vss.n4748 vss.n3628 0.0661418
R46860 vss.n5538 vss.n5537 0.0661418
R46861 vss.n5539 vss.n5538 0.0661418
R46862 vss.n4759 vss.n4752 0.0661418
R46863 vss.n4755 vss.n4752 0.0661418
R46864 vss.n4764 vss.n4763 0.0661418
R46865 vss.n4763 vss.n4756 0.0661418
R46866 vss.n4766 vss.n4765 0.0661418
R46867 vss.n5526 vss.n4766 0.0661418
R46868 vss.n5518 vss.n5515 0.0661418
R46869 vss.n5518 vss.n2986 0.0661418
R46870 vss.n4782 vss.n4781 0.0661418
R46871 vss.n4781 vss.n4777 0.0661418
R46872 vss.n5505 vss.n4774 0.0661418
R46873 vss.n4778 vss.n4774 0.0661418
R46874 vss.n5523 vss.n5522 0.0661418
R46875 vss.n5524 vss.n5523 0.0661418
R46876 vss.n4784 vss.n4783 0.0661418
R46877 vss.n5498 vss.n4784 0.0661418
R46878 vss.n4791 vss.n4788 0.0661418
R46879 vss.n4791 vss.n3626 0.0661418
R46880 vss.n5495 vss.n5494 0.0661418
R46881 vss.n5496 vss.n5495 0.0661418
R46882 vss.n4802 vss.n4795 0.0661418
R46883 vss.n4798 vss.n4795 0.0661418
R46884 vss.n4807 vss.n4806 0.0661418
R46885 vss.n4806 vss.n4799 0.0661418
R46886 vss.n4809 vss.n4808 0.0661418
R46887 vss.n5483 vss.n4809 0.0661418
R46888 vss.n5475 vss.n5472 0.0661418
R46889 vss.n5475 vss.n2983 0.0661418
R46890 vss.n4825 vss.n4824 0.0661418
R46891 vss.n4824 vss.n4820 0.0661418
R46892 vss.n5462 vss.n4817 0.0661418
R46893 vss.n4821 vss.n4817 0.0661418
R46894 vss.n5480 vss.n5479 0.0661418
R46895 vss.n5481 vss.n5480 0.0661418
R46896 vss.n4827 vss.n4826 0.0661418
R46897 vss.n5455 vss.n4827 0.0661418
R46898 vss.n4834 vss.n4831 0.0661418
R46899 vss.n4834 vss.n3624 0.0661418
R46900 vss.n5452 vss.n5451 0.0661418
R46901 vss.n5453 vss.n5452 0.0661418
R46902 vss.n4845 vss.n4838 0.0661418
R46903 vss.n4841 vss.n4838 0.0661418
R46904 vss.n4850 vss.n4849 0.0661418
R46905 vss.n4849 vss.n4842 0.0661418
R46906 vss.n4852 vss.n4851 0.0661418
R46907 vss.n5440 vss.n4852 0.0661418
R46908 vss.n5432 vss.n5429 0.0661418
R46909 vss.n5432 vss.n2980 0.0661418
R46910 vss.n4868 vss.n4867 0.0661418
R46911 vss.n4867 vss.n4863 0.0661418
R46912 vss.n5419 vss.n4860 0.0661418
R46913 vss.n4864 vss.n4860 0.0661418
R46914 vss.n5437 vss.n5436 0.0661418
R46915 vss.n5438 vss.n5437 0.0661418
R46916 vss.n4870 vss.n4869 0.0661418
R46917 vss.n5412 vss.n4870 0.0661418
R46918 vss.n4877 vss.n4874 0.0661418
R46919 vss.n4877 vss.n3612 0.0661418
R46920 vss.n5409 vss.n5408 0.0661418
R46921 vss.n5410 vss.n5409 0.0661418
R46922 vss.n5339 vss.n5332 0.0661418
R46923 vss.n5335 vss.n5332 0.0661418
R46924 vss.n5344 vss.n5343 0.0661418
R46925 vss.n5343 vss.n5336 0.0661418
R46926 vss.n5346 vss.n5345 0.0661418
R46927 vss.n5397 vss.n5346 0.0661418
R46928 vss.n5367 vss.n5357 0.0661418
R46929 vss.n5359 vss.n5357 0.0661418
R46930 vss.n5394 vss.n5393 0.0661418
R46931 vss.n5395 vss.n5394 0.0661418
R46932 vss.n5365 vss.n5360 0.0661418
R46933 vss.n5365 vss.n5364 0.0661418
R46934 vss.n5362 vss.n5361 0.0661418
R46935 vss.n5363 vss.n5362 0.0661418
R46936 vss.n5389 vss.n5385 0.0661418
R46937 vss.n5389 vss.n5388 0.0661418
R46938 vss.n2885 vss.n2872 0.0661418
R46939 vss.n2886 vss.n2885 0.0661418
R46940 vss.n2879 vss.n2876 0.0661418
R46941 vss.n2877 vss.n2876 0.0661418
R46942 vss.n9823 vss.n2887 0.0661418
R46943 vss.n2887 vss.n2884 0.0661418
R46944 vss.n9822 vss.n2888 0.0661418
R46945 vss.n9819 vss.n2888 0.0661418
R46946 vss.n9837 vss.n2878 0.0661418
R46947 vss.n2878 vss.n2777 0.0661418
R46948 vss.n2951 vss.n2950 0.0661418
R46949 vss.n2950 vss.n2944 0.0661418
R46950 vss.n2956 vss.n2953 0.0661418
R46951 vss.n2954 vss.n2953 0.0661418
R46952 vss.n2945 vss.n2941 0.0661418
R46953 vss.n2945 vss.n2937 0.0661418
R46954 vss.n2940 vss.n2936 0.0661418
R46955 vss.n2979 vss.n2936 0.0661418
R46956 vss.n2963 vss.n2955 0.0661418
R46957 vss.n2955 vss.n2778 0.0661418
R46958 vss.n2904 vss.n2903 0.0661418
R46959 vss.n2903 vss.n2897 0.0661418
R46960 vss.n2909 vss.n2906 0.0661418
R46961 vss.n2907 vss.n2906 0.0661418
R46962 vss.n2898 vss.n2894 0.0661418
R46963 vss.n2898 vss.n2890 0.0661418
R46964 vss.n2893 vss.n2889 0.0661418
R46965 vss.n2933 vss.n2889 0.0661418
R46966 vss.n2916 vss.n2908 0.0661418
R46967 vss.n2908 vss.n2779 0.0661418
R46968 vss.n4936 vss.n4923 0.0661418
R46969 vss.n4937 vss.n4936 0.0661418
R46970 vss.n4930 vss.n4927 0.0661418
R46971 vss.n4928 vss.n4927 0.0661418
R46972 vss.n4943 vss.n4938 0.0661418
R46973 vss.n4938 vss.n4935 0.0661418
R46974 vss.n4942 vss.n4939 0.0661418
R46975 vss.n4939 vss.n2982 0.0661418
R46976 vss.n4957 vss.n4929 0.0661418
R46977 vss.n4929 vss.n2780 0.0661418
R46978 vss.n5138 vss.n5125 0.0661418
R46979 vss.n5139 vss.n5138 0.0661418
R46980 vss.n5132 vss.n5129 0.0661418
R46981 vss.n5130 vss.n5129 0.0661418
R46982 vss.n5145 vss.n5140 0.0661418
R46983 vss.n5140 vss.n5137 0.0661418
R46984 vss.n5144 vss.n5141 0.0661418
R46985 vss.n5141 vss.n2988 0.0661418
R46986 vss.n5159 vss.n5131 0.0661418
R46987 vss.n5131 vss.n2781 0.0661418
R46988 vss.n3118 vss.n3105 0.0661418
R46989 vss.n3119 vss.n3118 0.0661418
R46990 vss.n3112 vss.n3109 0.0661418
R46991 vss.n3110 vss.n3109 0.0661418
R46992 vss.n3126 vss.n3120 0.0661418
R46993 vss.n3120 vss.n3117 0.0661418
R46994 vss.n3125 vss.n3121 0.0661418
R46995 vss.n3122 vss.n3121 0.0661418
R46996 vss.n3140 vss.n3111 0.0661418
R46997 vss.n3111 vss.n2782 0.0661418
R46998 vss.n4472 vss.n4461 0.0661418
R46999 vss.n4472 vss.n4466 0.0661418
R47000 vss.n4477 vss.n4475 0.0661418
R47001 vss.n4475 vss.n4474 0.0661418
R47002 vss.n4498 vss.n4468 0.0661418
R47003 vss.n4499 vss.n4498 0.0661418
R47004 vss.n4494 vss.n4469 0.0661418
R47005 vss.n4469 vss.n2703 0.0661418
R47006 vss.n4481 vss.n4476 0.0661418
R47007 vss.n4480 vss.n4476 0.0661418
R47008 vss.n4380 vss.n4369 0.0661418
R47009 vss.n4380 vss.n4374 0.0661418
R47010 vss.n4385 vss.n4383 0.0661418
R47011 vss.n4383 vss.n4382 0.0661418
R47012 vss.n4406 vss.n4376 0.0661418
R47013 vss.n4407 vss.n4406 0.0661418
R47014 vss.n4402 vss.n4377 0.0661418
R47015 vss.n4377 vss.n2700 0.0661418
R47016 vss.n4389 vss.n4384 0.0661418
R47017 vss.n4388 vss.n4384 0.0661418
R47018 vss.n4332 vss.n4321 0.0661418
R47019 vss.n4332 vss.n4326 0.0661418
R47020 vss.n4337 vss.n4335 0.0661418
R47021 vss.n4335 vss.n4334 0.0661418
R47022 vss.n4358 vss.n4328 0.0661418
R47023 vss.n4359 vss.n4358 0.0661418
R47024 vss.n4354 vss.n4329 0.0661418
R47025 vss.n4329 vss.n2702 0.0661418
R47026 vss.n4341 vss.n4336 0.0661418
R47027 vss.n4340 vss.n4336 0.0661418
R47028 vss.n3732 vss.n3721 0.0661418
R47029 vss.n3732 vss.n3726 0.0661418
R47030 vss.n3737 vss.n3735 0.0661418
R47031 vss.n3735 vss.n3734 0.0661418
R47032 vss.n3758 vss.n3728 0.0661418
R47033 vss.n3759 vss.n3758 0.0661418
R47034 vss.n3754 vss.n3729 0.0661418
R47035 vss.n3729 vss.n2697 0.0661418
R47036 vss.n3741 vss.n3736 0.0661418
R47037 vss.n3740 vss.n3736 0.0661418
R47038 vss.n4034 vss.n4023 0.0661418
R47039 vss.n4034 vss.n4028 0.0661418
R47040 vss.n4039 vss.n4037 0.0661418
R47041 vss.n4037 vss.n4036 0.0661418
R47042 vss.n4060 vss.n4030 0.0661418
R47043 vss.n4061 vss.n4060 0.0661418
R47044 vss.n4056 vss.n4031 0.0661418
R47045 vss.n4031 vss.n2694 0.0661418
R47046 vss.n4043 vss.n4038 0.0661418
R47047 vss.n4042 vss.n4038 0.0661418
R47048 vss.n3687 vss.n3676 0.0661418
R47049 vss.n3687 vss.n3681 0.0661418
R47050 vss.n3692 vss.n3690 0.0661418
R47051 vss.n3690 vss.n3689 0.0661418
R47052 vss.n3713 vss.n3683 0.0661418
R47053 vss.n3714 vss.n3713 0.0661418
R47054 vss.n3709 vss.n3684 0.0661418
R47055 vss.n3684 vss.n2696 0.0661418
R47056 vss.n3696 vss.n3691 0.0661418
R47057 vss.n3695 vss.n3691 0.0661418
R47058 vss.n4088 vss.n4077 0.0661418
R47059 vss.n4088 vss.n4082 0.0661418
R47060 vss.n4093 vss.n4091 0.0661418
R47061 vss.n4091 vss.n4090 0.0661418
R47062 vss.n4114 vss.n4084 0.0661418
R47063 vss.n4115 vss.n4114 0.0661418
R47064 vss.n4110 vss.n4085 0.0661418
R47065 vss.n4085 vss.n2691 0.0661418
R47066 vss.n4097 vss.n4092 0.0661418
R47067 vss.n4096 vss.n4092 0.0661418
R47068 vss.n3512 vss.n3501 0.0661418
R47069 vss.n3512 vss.n3506 0.0661418
R47070 vss.n3517 vss.n3515 0.0661418
R47071 vss.n3515 vss.n3514 0.0661418
R47072 vss.n3538 vss.n3508 0.0661418
R47073 vss.n3539 vss.n3538 0.0661418
R47074 vss.n3534 vss.n3509 0.0661418
R47075 vss.n3509 vss.n2688 0.0661418
R47076 vss.n3521 vss.n3516 0.0661418
R47077 vss.n3520 vss.n3516 0.0661418
R47078 vss.n3467 vss.n3456 0.0661418
R47079 vss.n3467 vss.n3461 0.0661418
R47080 vss.n3472 vss.n3470 0.0661418
R47081 vss.n3470 vss.n3469 0.0661418
R47082 vss.n3493 vss.n3463 0.0661418
R47083 vss.n3494 vss.n3493 0.0661418
R47084 vss.n3489 vss.n3464 0.0661418
R47085 vss.n3464 vss.n2690 0.0661418
R47086 vss.n3476 vss.n3471 0.0661418
R47087 vss.n3475 vss.n3471 0.0661418
R47088 vss.n5755 vss.n5744 0.0661418
R47089 vss.n5755 vss.n5749 0.0661418
R47090 vss.n5760 vss.n5758 0.0661418
R47091 vss.n5758 vss.n5757 0.0661418
R47092 vss.n5781 vss.n5751 0.0661418
R47093 vss.n5782 vss.n5781 0.0661418
R47094 vss.n5777 vss.n5752 0.0661418
R47095 vss.n5752 vss.n2685 0.0661418
R47096 vss.n5764 vss.n5759 0.0661418
R47097 vss.n5763 vss.n5759 0.0661418
R47098 vss.n4514 vss.n4452 0.0661418
R47099 vss.n4531 vss.n4452 0.0661418
R47100 vss.n4516 vss.n4447 0.0661418
R47101 vss.n4447 vss.n4443 0.0661418
R47102 vss.n4512 vss.n4509 0.0661418
R47103 vss.n4512 vss.n4455 0.0661418
R47104 vss.n4511 vss.n4510 0.0661418
R47105 vss.n4511 vss.n2707 0.0661418
R47106 vss.n4517 vss.n4445 0.0661418
R47107 vss.n4445 vss.n2704 0.0661418
R47108 vss.n4434 vss.n4433 0.0661418
R47109 vss.n4433 vss.n4431 0.0661418
R47110 vss.n4440 vss.n4439 0.0661418
R47111 vss.n4439 vss.n4437 0.0661418
R47112 vss.n4429 vss.n4426 0.0661418
R47113 vss.n4429 vss.n4421 0.0661418
R47114 vss.n4442 vss.n4441 0.0661418
R47115 vss.n4536 vss.n4442 0.0661418
R47116 vss.n4555 vss.n4554 0.0661418
R47117 vss.n4555 vss.n4422 0.0661418
R47118 vss.n4562 vss.n4413 0.0661418
R47119 vss.n4562 vss.n4418 0.0661418
R47120 vss.n4567 vss.n4565 0.0661418
R47121 vss.n4565 vss.n4564 0.0661418
R47122 vss.n4605 vss.n4420 0.0661418
R47123 vss.n4606 vss.n4605 0.0661418
R47124 vss.n4601 vss.n4559 0.0661418
R47125 vss.n4559 vss.n4558 0.0661418
R47126 vss.n4588 vss.n4566 0.0661418
R47127 vss.n4566 vss.n2701 0.0661418
R47128 vss.n3644 vss.n3643 0.0661418
R47129 vss.n3643 vss.n3638 0.0661418
R47130 vss.n4577 vss.n4574 0.0661418
R47131 vss.n4577 vss.n4576 0.0661418
R47132 vss.n3641 vss.n3634 0.0661418
R47133 vss.n3641 vss.n3639 0.0661418
R47134 vss.n4585 vss.n4584 0.0661418
R47135 vss.n4586 vss.n4585 0.0661418
R47136 vss.n4626 vss.n4625 0.0661418
R47137 vss.n4627 vss.n4626 0.0661418
R47138 vss.n3776 vss.n3763 0.0661418
R47139 vss.n3776 vss.n3768 0.0661418
R47140 vss.n3781 vss.n3779 0.0661418
R47141 vss.n3779 vss.n3778 0.0661418
R47142 vss.n4202 vss.n3770 0.0661418
R47143 vss.n4203 vss.n4202 0.0661418
R47144 vss.n4198 vss.n3773 0.0661418
R47145 vss.n3773 vss.n3772 0.0661418
R47146 vss.n4185 vss.n3780 0.0661418
R47147 vss.n3780 vss.n2698 0.0661418
R47148 vss.n3798 vss.n3797 0.0661418
R47149 vss.n3797 vss.n3792 0.0661418
R47150 vss.n3793 vss.n3787 0.0661418
R47151 vss.n3793 vss.n3791 0.0661418
R47152 vss.n3817 vss.n3816 0.0661418
R47153 vss.n3817 vss.n3811 0.0661418
R47154 vss.n4182 vss.n4181 0.0661418
R47155 vss.n4183 vss.n4182 0.0661418
R47156 vss.n3825 vss.n3824 0.0661418
R47157 vss.n3825 vss.n3629 0.0661418
R47158 vss.n3832 vss.n3803 0.0661418
R47159 vss.n3832 vss.n3808 0.0661418
R47160 vss.n3837 vss.n3835 0.0661418
R47161 vss.n3835 vss.n3834 0.0661418
R47162 vss.n4167 vss.n3810 0.0661418
R47163 vss.n4168 vss.n4167 0.0661418
R47164 vss.n4163 vss.n3829 0.0661418
R47165 vss.n3829 vss.n3828 0.0661418
R47166 vss.n4150 vss.n3836 0.0661418
R47167 vss.n3836 vss.n2695 0.0661418
R47168 vss.n3854 vss.n3853 0.0661418
R47169 vss.n3853 vss.n3848 0.0661418
R47170 vss.n3849 vss.n3843 0.0661418
R47171 vss.n3849 vss.n3847 0.0661418
R47172 vss.n3863 vss.n3859 0.0661418
R47173 vss.n4136 vss.n3859 0.0661418
R47174 vss.n4147 vss.n4146 0.0661418
R47175 vss.n4148 vss.n4147 0.0661418
R47176 vss.n3868 vss.n3867 0.0661418
R47177 vss.n3868 vss.n3627 0.0661418
R47178 vss.n3883 vss.n3882 0.0661418
R47179 vss.n3882 vss.n3877 0.0661418
R47180 vss.n3889 vss.n3888 0.0661418
R47181 vss.n3888 vss.n3886 0.0661418
R47182 vss.n3880 vss.n3873 0.0661418
R47183 vss.n3880 vss.n3878 0.0661418
R47184 vss.n4133 vss.n4132 0.0661418
R47185 vss.n4134 vss.n4133 0.0661418
R47186 vss.n3891 vss.n3890 0.0661418
R47187 vss.n3891 vss.n2692 0.0661418
R47188 vss.n3906 vss.n3905 0.0661418
R47189 vss.n3905 vss.n3900 0.0661418
R47190 vss.n3901 vss.n3895 0.0661418
R47191 vss.n3901 vss.n3899 0.0661418
R47192 vss.n3914 vss.n3910 0.0661418
R47193 vss.n3923 vss.n3910 0.0661418
R47194 vss.n3934 vss.n3933 0.0661418
R47195 vss.n3935 vss.n3934 0.0661418
R47196 vss.n3919 vss.n3918 0.0661418
R47197 vss.n3919 vss.n3625 0.0661418
R47198 vss.n3555 vss.n3544 0.0661418
R47199 vss.n3555 vss.n3549 0.0661418
R47200 vss.n3560 vss.n3558 0.0661418
R47201 vss.n3558 vss.n3557 0.0661418
R47202 vss.n5834 vss.n3551 0.0661418
R47203 vss.n5835 vss.n5834 0.0661418
R47204 vss.n5830 vss.n3552 0.0661418
R47205 vss.n3921 vss.n3552 0.0661418
R47206 vss.n5817 vss.n3559 0.0661418
R47207 vss.n3559 vss.n2689 0.0661418
R47208 vss.n3577 vss.n3576 0.0661418
R47209 vss.n3576 vss.n3571 0.0661418
R47210 vss.n3572 vss.n3566 0.0661418
R47211 vss.n3572 vss.n3570 0.0661418
R47212 vss.n3617 vss.n3583 0.0661418
R47213 vss.n5803 vss.n3583 0.0661418
R47214 vss.n5814 vss.n5813 0.0661418
R47215 vss.n5815 vss.n5814 0.0661418
R47216 vss.n3622 vss.n3621 0.0661418
R47217 vss.n3623 vss.n3622 0.0661418
R47218 vss.n3597 vss.n3596 0.0661418
R47219 vss.n3596 vss.n3591 0.0661418
R47220 vss.n5666 vss.n5663 0.0661418
R47221 vss.n5663 vss.n5659 0.0661418
R47222 vss.n3594 vss.n3587 0.0661418
R47223 vss.n3594 vss.n3592 0.0661418
R47224 vss.n5800 vss.n5799 0.0661418
R47225 vss.n5801 vss.n5800 0.0661418
R47226 vss.n5667 vss.n5661 0.0661418
R47227 vss.n5661 vss.n2686 0.0661418
R47228 vss.n5651 vss.n3603 0.0661418
R47229 vss.n5651 vss.n3608 0.0661418
R47230 vss.n5656 vss.n5654 0.0661418
R47231 vss.n5654 vss.n5653 0.0661418
R47232 vss.n5648 vss.n3610 0.0661418
R47233 vss.n5735 vss.n3610 0.0661418
R47234 vss.n5677 vss.n5655 0.0661418
R47235 vss.n5676 vss.n5655 0.0661418
R47236 vss.n5690 vss.n5689 0.0661418
R47237 vss.n5690 vss.n5644 0.0661418
R47238 vss.n5705 vss.n5704 0.0661418
R47239 vss.n5704 vss.n5699 0.0661418
R47240 vss.n5711 vss.n5710 0.0661418
R47241 vss.n5710 vss.n5708 0.0661418
R47242 vss.n5702 vss.n5695 0.0661418
R47243 vss.n5702 vss.n5700 0.0661418
R47244 vss.n5732 vss.n5731 0.0661418
R47245 vss.n5733 vss.n5732 0.0661418
R47246 vss.n5713 vss.n5712 0.0661418
R47247 vss.n5713 vss.n2639 0.0661418
R47248 vss.n9959 vss.n2631 0.0661418
R47249 vss.n9959 vss.n2636 0.0661418
R47250 vss.n9964 vss.n9962 0.0661418
R47251 vss.n9962 vss.n9961 0.0661418
R47252 vss.n9985 vss.n2638 0.0661418
R47253 vss.n9986 vss.n9985 0.0661418
R47254 vss.n9981 vss.n9956 0.0661418
R47255 vss.n9956 vss.n9955 0.0661418
R47256 vss.n9968 vss.n9963 0.0661418
R47257 vss.n9967 vss.n9963 0.0661418
R47258 vss.n2653 vss.n2652 0.0661418
R47259 vss.n2652 vss.n2647 0.0661418
R47260 vss.n2659 vss.n2658 0.0661418
R47261 vss.n2658 vss.n2656 0.0661418
R47262 vss.n2650 vss.n2643 0.0661418
R47263 vss.n2650 vss.n2648 0.0661418
R47264 vss.n2683 vss.n2682 0.0661418
R47265 vss.n2684 vss.n2683 0.0661418
R47266 vss.n2661 vss.n2660 0.0661418
R47267 vss.n2662 vss.n2661 0.0661418
R47268 vss.n3392 vss.n3381 0.0661418
R47269 vss.n3392 vss.n3386 0.0661418
R47270 vss.n3397 vss.n3395 0.0661418
R47271 vss.n3395 vss.n3394 0.0661418
R47272 vss.n3418 vss.n3388 0.0661418
R47273 vss.n3419 vss.n3418 0.0661418
R47274 vss.n3414 vss.n3389 0.0661418
R47275 vss.n3389 vss.n2687 0.0661418
R47276 vss.n3401 vss.n3396 0.0661418
R47277 vss.n3400 vss.n3396 0.0661418
R47278 vss.n3989 vss.n3978 0.0661418
R47279 vss.n3989 vss.n3983 0.0661418
R47280 vss.n3994 vss.n3992 0.0661418
R47281 vss.n3992 vss.n3991 0.0661418
R47282 vss.n4015 vss.n3985 0.0661418
R47283 vss.n4016 vss.n4015 0.0661418
R47284 vss.n4011 vss.n3986 0.0661418
R47285 vss.n3986 vss.n2693 0.0661418
R47286 vss.n3998 vss.n3993 0.0661418
R47287 vss.n3997 vss.n3993 0.0661418
R47288 vss.n4256 vss.n4245 0.0661418
R47289 vss.n4256 vss.n4250 0.0661418
R47290 vss.n4261 vss.n4259 0.0661418
R47291 vss.n4259 vss.n4258 0.0661418
R47292 vss.n4282 vss.n4252 0.0661418
R47293 vss.n4283 vss.n4282 0.0661418
R47294 vss.n4278 vss.n4253 0.0661418
R47295 vss.n4253 vss.n2699 0.0661418
R47296 vss.n4265 vss.n4260 0.0661418
R47297 vss.n4264 vss.n4260 0.0661418
R47298 vss.n5918 vss.n5917 0.0661418
R47299 vss.n5917 vss.n5895 0.0661418
R47300 vss.n5896 vss.n5889 0.0661418
R47301 vss.n5896 vss.n5894 0.0661418
R47302 vss.n5904 vss.n5902 0.0661418
R47303 vss.n5902 vss.n5901 0.0661418
R47304 vss.n5908 vss.n5903 0.0661418
R47305 vss.n5907 vss.n5903 0.0661418
R47306 vss.n5922 vss.n5919 0.0661418
R47307 vss.n5922 vss.n2705 0.0661418
R47308 vss.n9928 vss.n9927 0.0661418
R47309 vss.n9929 vss.n9928 0.0661418
R47310 vss.n3278 vss.n3276 0.0661418
R47311 vss.n3276 vss.n3275 0.0661418
R47312 vss.n3270 vss.n3263 0.0661418
R47313 vss.n3270 vss.n3268 0.0661418
R47314 vss.n3295 vss.n3292 0.0661418
R47315 vss.n3296 vss.n3295 0.0661418
R47316 vss.n3294 vss.n3293 0.0661418
R47317 vss.n3294 vss.n2742 0.0661418
R47318 vss.n3283 vss.n3277 0.0661418
R47319 vss.n3282 vss.n3277 0.0661418
R47320 vss.n9700 vss.n9698 0.0661418
R47321 vss.n9698 vss.n9697 0.0661418
R47322 vss.n9692 vss.n9685 0.0661418
R47323 vss.n9692 vss.n9690 0.0661418
R47324 vss.n9715 vss.n9714 0.0661418
R47325 vss.n9714 vss.n9691 0.0661418
R47326 vss.n9717 vss.n9716 0.0661418
R47327 vss.n9720 vss.n9717 0.0661418
R47328 vss.n9705 vss.n9699 0.0661418
R47329 vss.n9704 vss.n9699 0.0661418
R47330 vss.n2753 vss.n2747 0.0661418
R47331 vss.n2753 vss.n2751 0.0661418
R47332 vss.n2758 vss.n2757 0.0661418
R47333 vss.n2757 vss.n2752 0.0661418
R47334 vss.n9882 vss.n9881 0.0661418
R47335 vss.n9883 vss.n9882 0.0661418
R47336 vss.n9877 vss.n2764 0.0661418
R47337 vss.n9877 vss.n9876 0.0661418
R47338 vss.n9894 vss.n9893 0.0661418
R47339 vss.n9895 vss.n9894 0.0661418
R47340 vss.n9036 vss.n9035 0.0661418
R47341 vss.n9037 vss.n9036 0.0661418
R47342 vss.n8075 vss.n8074 0.0661418
R47343 vss.n8074 vss.n8072 0.0661418
R47344 vss.n8069 vss.n8068 0.0661418
R47345 vss.n8068 vss.n8063 0.0661418
R47346 vss.n8066 vss.n8056 0.0661418
R47347 vss.n8066 vss.n8064 0.0661418
R47348 vss.n8077 vss.n8076 0.0661418
R47349 vss.n8079 vss.n8077 0.0661418
R47350 vss.n8098 vss.n8097 0.0661418
R47351 vss.n8099 vss.n8098 0.0661418
R47352 vss.n8119 vss.n8118 0.0661418
R47353 vss.n8118 vss.n8116 0.0661418
R47354 vss.n8113 vss.n8112 0.0661418
R47355 vss.n8112 vss.n8107 0.0661418
R47356 vss.n8110 vss.n8103 0.0661418
R47357 vss.n8110 vss.n8108 0.0661418
R47358 vss.n8172 vss.n8171 0.0661418
R47359 vss.n8173 vss.n8172 0.0661418
R47360 vss.n7488 vss.n7486 0.0661418
R47361 vss.n7486 vss.n7485 0.0661418
R47362 vss.n7480 vss.n7473 0.0661418
R47363 vss.n7480 vss.n7478 0.0661418
R47364 vss.n8961 vss.n8960 0.0661418
R47365 vss.n8960 vss.n7479 0.0661418
R47366 vss.n8963 vss.n8962 0.0661418
R47367 vss.n8963 vss.n7325 0.0661418
R47368 vss.n8951 vss.n7487 0.0661418
R47369 vss.n8950 vss.n7487 0.0661418
R47370 vss.n8869 vss.n7543 0.0661418
R47371 vss.n8869 vss.n8867 0.0661418
R47372 vss.n8874 vss.n8873 0.0661418
R47373 vss.n8873 vss.n8868 0.0661418
R47374 vss.n8888 vss.n8887 0.0661418
R47375 vss.n8889 vss.n8888 0.0661418
R47376 vss.n8883 vss.n8880 0.0661418
R47377 vss.n8883 vss.n7326 0.0661418
R47378 vss.n8900 vss.n8899 0.0661418
R47379 vss.n8901 vss.n8900 0.0661418
R47380 vss.n7677 vss.n7675 0.0661418
R47381 vss.n7675 vss.n7674 0.0661418
R47382 vss.n7669 vss.n7662 0.0661418
R47383 vss.n7669 vss.n7667 0.0661418
R47384 vss.n8842 vss.n8841 0.0661418
R47385 vss.n8841 vss.n7668 0.0661418
R47386 vss.n8844 vss.n8843 0.0661418
R47387 vss.n8844 vss.n7327 0.0661418
R47388 vss.n8832 vss.n7676 0.0661418
R47389 vss.n8831 vss.n7676 0.0661418
R47390 vss.n8750 vss.n7686 0.0661418
R47391 vss.n8750 vss.n8748 0.0661418
R47392 vss.n8755 vss.n8754 0.0661418
R47393 vss.n8754 vss.n8749 0.0661418
R47394 vss.n8769 vss.n8768 0.0661418
R47395 vss.n8770 vss.n8769 0.0661418
R47396 vss.n8764 vss.n8761 0.0661418
R47397 vss.n8764 vss.n7328 0.0661418
R47398 vss.n8781 vss.n8780 0.0661418
R47399 vss.n8782 vss.n8781 0.0661418
R47400 vss.n7864 vss.n7862 0.0661418
R47401 vss.n7862 vss.n7861 0.0661418
R47402 vss.n7856 vss.n7849 0.0661418
R47403 vss.n7856 vss.n7854 0.0661418
R47404 vss.n8723 vss.n8722 0.0661418
R47405 vss.n8722 vss.n7855 0.0661418
R47406 vss.n8725 vss.n8724 0.0661418
R47407 vss.n8725 vss.n7329 0.0661418
R47408 vss.n8713 vss.n7863 0.0661418
R47409 vss.n8712 vss.n7863 0.0661418
R47410 vss.n7309 vss.n7303 0.0661418
R47411 vss.n7309 vss.n7307 0.0661418
R47412 vss.n7314 vss.n7313 0.0661418
R47413 vss.n7313 vss.n7308 0.0661418
R47414 vss.n8993 vss.n8992 0.0661418
R47415 vss.n8994 vss.n8993 0.0661418
R47416 vss.n8988 vss.n7320 0.0661418
R47417 vss.n8988 vss.n8987 0.0661418
R47418 vss.n9005 vss.n9004 0.0661418
R47419 vss.n9006 vss.n9005 0.0661418
R47420 vss.n8007 vss.n8005 0.0661418
R47421 vss.n8005 vss.n8004 0.0661418
R47422 vss.n7999 vss.n7992 0.0661418
R47423 vss.n7999 vss.n7997 0.0661418
R47424 vss.n8232 vss.n8231 0.0661418
R47425 vss.n8231 vss.n7998 0.0661418
R47426 vss.n8234 vss.n8233 0.0661418
R47427 vss.n8234 vss.n7330 0.0661418
R47428 vss.n8222 vss.n8006 0.0661418
R47429 vss.n8221 vss.n8006 0.0661418
R47430 vss.n8186 vss.n8178 0.0661418
R47431 vss.n8186 vss.n8184 0.0661418
R47432 vss.n8191 vss.n8190 0.0661418
R47433 vss.n8190 vss.n8185 0.0661418
R47434 vss.n8205 vss.n8204 0.0661418
R47435 vss.n8206 vss.n8205 0.0661418
R47436 vss.n8200 vss.n8197 0.0661418
R47437 vss.n8200 vss.n7331 0.0661418
R47438 vss.n8217 vss.n8216 0.0661418
R47439 vss.n8218 vss.n8217 0.0661418
R47440 vss.n7924 vss.n7922 0.0661418
R47441 vss.n7922 vss.n7921 0.0661418
R47442 vss.n7916 vss.n7909 0.0661418
R47443 vss.n7916 vss.n7914 0.0661418
R47444 vss.n7938 vss.n7937 0.0661418
R47445 vss.n7937 vss.n7915 0.0661418
R47446 vss.n7940 vss.n7939 0.0661418
R47447 vss.n7940 vss.n7333 0.0661418
R47448 vss.n7928 vss.n7923 0.0661418
R47449 vss.n7927 vss.n7923 0.0661418
R47450 vss.n7783 vss.n7781 0.0661418
R47451 vss.n7781 vss.n7780 0.0661418
R47452 vss.n7775 vss.n7768 0.0661418
R47453 vss.n7775 vss.n7773 0.0661418
R47454 vss.n7797 vss.n7796 0.0661418
R47455 vss.n7796 vss.n7774 0.0661418
R47456 vss.n7799 vss.n7798 0.0661418
R47457 vss.n7799 vss.n7334 0.0661418
R47458 vss.n7787 vss.n7782 0.0661418
R47459 vss.n7786 vss.n7782 0.0661418
R47460 vss.n7703 vss.n7701 0.0661418
R47461 vss.n7701 vss.n7700 0.0661418
R47462 vss.n7695 vss.n7688 0.0661418
R47463 vss.n7695 vss.n7693 0.0661418
R47464 vss.n7717 vss.n7716 0.0661418
R47465 vss.n7716 vss.n7694 0.0661418
R47466 vss.n7719 vss.n7718 0.0661418
R47467 vss.n7719 vss.n7335 0.0661418
R47468 vss.n7707 vss.n7702 0.0661418
R47469 vss.n7706 vss.n7702 0.0661418
R47470 vss.n8796 vss.n8788 0.0661418
R47471 vss.n8796 vss.n8794 0.0661418
R47472 vss.n8801 vss.n8800 0.0661418
R47473 vss.n8800 vss.n8795 0.0661418
R47474 vss.n8815 vss.n8814 0.0661418
R47475 vss.n8816 vss.n8815 0.0661418
R47476 vss.n8810 vss.n8807 0.0661418
R47477 vss.n8810 vss.n7336 0.0661418
R47478 vss.n8827 vss.n8826 0.0661418
R47479 vss.n8828 vss.n8827 0.0661418
R47480 vss.n7560 vss.n7558 0.0661418
R47481 vss.n7558 vss.n7557 0.0661418
R47482 vss.n7552 vss.n7545 0.0661418
R47483 vss.n7552 vss.n7550 0.0661418
R47484 vss.n7574 vss.n7573 0.0661418
R47485 vss.n7573 vss.n7551 0.0661418
R47486 vss.n7576 vss.n7575 0.0661418
R47487 vss.n7576 vss.n7337 0.0661418
R47488 vss.n7564 vss.n7559 0.0661418
R47489 vss.n7563 vss.n7559 0.0661418
R47490 vss.n8915 vss.n8907 0.0661418
R47491 vss.n8915 vss.n8913 0.0661418
R47492 vss.n8920 vss.n8919 0.0661418
R47493 vss.n8919 vss.n8914 0.0661418
R47494 vss.n8934 vss.n8933 0.0661418
R47495 vss.n8935 vss.n8934 0.0661418
R47496 vss.n8929 vss.n8926 0.0661418
R47497 vss.n8929 vss.n7338 0.0661418
R47498 vss.n8946 vss.n8945 0.0661418
R47499 vss.n8947 vss.n8946 0.0661418
R47500 vss.n7503 vss.n7494 0.0661418
R47501 vss.n7503 vss.n7501 0.0661418
R47502 vss.n7508 vss.n7507 0.0661418
R47503 vss.n7507 vss.n7502 0.0661418
R47504 vss.n7522 vss.n7521 0.0661418
R47505 vss.n7523 vss.n7522 0.0661418
R47506 vss.n7517 vss.n7514 0.0661418
R47507 vss.n7517 vss.n7339 0.0661418
R47508 vss.n7534 vss.n7533 0.0661418
R47509 vss.n7535 vss.n7534 0.0661418
R47510 vss.n650 vss.n617 0.0661418
R47511 vss.n650 vss.n649 0.0661418
R47512 vss.n625 vss.n621 0.0661418
R47513 vss.n626 vss.n625 0.0661418
R47514 vss.n629 vss.n628 0.0661418
R47515 vss.n628 vss.n624 0.0661418
R47516 vss.n631 vss.n630 0.0661418
R47517 vss.n631 vss.n512 0.0661418
R47518 vss.n657 vss.n656 0.0661418
R47519 vss.n658 vss.n657 0.0661418
R47520 vss.n462 vss.n460 0.0661418
R47521 vss.n460 vss.n458 0.0661418
R47522 vss.n454 vss.n453 0.0661418
R47523 vss.n453 vss.n451 0.0661418
R47524 vss.n448 vss.n447 0.0661418
R47525 vss.n447 vss.n441 0.0661418
R47526 vss.n445 vss.n437 0.0661418
R47527 vss.n445 vss.n444 0.0661418
R47528 vss.n14174 vss.n14173 0.0661418
R47529 vss.n14175 vss.n14174 0.0661418
R47530 vss.n456 vss.n455 0.0661418
R47531 vss.n14155 vss.n456 0.0661418
R47532 vss.n490 vss.n475 0.0661418
R47533 vss.n491 vss.n490 0.0661418
R47534 vss.n484 vss.n479 0.0661418
R47535 vss.n480 vss.n479 0.0661418
R47536 vss.n14067 vss.n492 0.0661418
R47537 vss.n492 vss.n489 0.0661418
R47538 vss.n14066 vss.n493 0.0661418
R47539 vss.n14063 vss.n493 0.0661418
R47540 vss.n14081 vss.n483 0.0661418
R47541 vss.n483 vss.n482 0.0661418
R47542 vss.n10115 vss.n10102 0.0661418
R47543 vss.n10116 vss.n10115 0.0661418
R47544 vss.n10109 vss.n10106 0.0661418
R47545 vss.n10107 vss.n10106 0.0661418
R47546 vss.n10122 vss.n10117 0.0661418
R47547 vss.n10117 vss.n10114 0.0661418
R47548 vss.n10121 vss.n10118 0.0661418
R47549 vss.n10118 vss.n2363 0.0661418
R47550 vss.n10136 vss.n10108 0.0661418
R47551 vss.n10108 vss.n2146 0.0661418
R47552 vss.n12873 vss.n12860 0.0661418
R47553 vss.n12874 vss.n12873 0.0661418
R47554 vss.n12867 vss.n12864 0.0661418
R47555 vss.n12865 vss.n12864 0.0661418
R47556 vss.n12880 vss.n12875 0.0661418
R47557 vss.n12875 vss.n12872 0.0661418
R47558 vss.n12879 vss.n12876 0.0661418
R47559 vss.n12876 vss.n2360 0.0661418
R47560 vss.n12894 vss.n12866 0.0661418
R47561 vss.n12866 vss.n2147 0.0661418
R47562 vss.n10156 vss.n10143 0.0661418
R47563 vss.n10157 vss.n10156 0.0661418
R47564 vss.n10150 vss.n10147 0.0661418
R47565 vss.n10148 vss.n10147 0.0661418
R47566 vss.n10163 vss.n10158 0.0661418
R47567 vss.n10158 vss.n10155 0.0661418
R47568 vss.n10162 vss.n10159 0.0661418
R47569 vss.n10159 vss.n2361 0.0661418
R47570 vss.n10177 vss.n10149 0.0661418
R47571 vss.n10149 vss.n2148 0.0661418
R47572 vss.n12422 vss.n12409 0.0661418
R47573 vss.n12423 vss.n12422 0.0661418
R47574 vss.n12416 vss.n12413 0.0661418
R47575 vss.n12414 vss.n12413 0.0661418
R47576 vss.n12429 vss.n12424 0.0661418
R47577 vss.n12424 vss.n12421 0.0661418
R47578 vss.n12428 vss.n12425 0.0661418
R47579 vss.n12425 vss.n2357 0.0661418
R47580 vss.n12443 vss.n12415 0.0661418
R47581 vss.n12415 vss.n2149 0.0661418
R47582 vss.n11751 vss.n11738 0.0661418
R47583 vss.n11752 vss.n11751 0.0661418
R47584 vss.n11745 vss.n11742 0.0661418
R47585 vss.n11743 vss.n11742 0.0661418
R47586 vss.n11758 vss.n11753 0.0661418
R47587 vss.n11753 vss.n11750 0.0661418
R47588 vss.n11757 vss.n11754 0.0661418
R47589 vss.n11754 vss.n2354 0.0661418
R47590 vss.n11772 vss.n11744 0.0661418
R47591 vss.n11744 vss.n2150 0.0661418
R47592 vss.n12467 vss.n12454 0.0661418
R47593 vss.n12468 vss.n12467 0.0661418
R47594 vss.n12461 vss.n12458 0.0661418
R47595 vss.n12459 vss.n12458 0.0661418
R47596 vss.n12474 vss.n12469 0.0661418
R47597 vss.n12469 vss.n12466 0.0661418
R47598 vss.n12473 vss.n12470 0.0661418
R47599 vss.n12470 vss.n2355 0.0661418
R47600 vss.n12488 vss.n12460 0.0661418
R47601 vss.n12460 vss.n2151 0.0661418
R47602 vss.n2321 vss.n2320 0.0661418
R47603 vss.n2320 vss.n2314 0.0661418
R47604 vss.n2326 vss.n2323 0.0661418
R47605 vss.n2324 vss.n2323 0.0661418
R47606 vss.n2315 vss.n2311 0.0661418
R47607 vss.n2315 vss.n2307 0.0661418
R47608 vss.n2310 vss.n2306 0.0661418
R47609 vss.n2349 vss.n2306 0.0661418
R47610 vss.n2333 vss.n2325 0.0661418
R47611 vss.n2325 vss.n2152 0.0661418
R47612 vss.n12292 vss.n12279 0.0661418
R47613 vss.n12293 vss.n12292 0.0661418
R47614 vss.n12286 vss.n12283 0.0661418
R47615 vss.n12284 vss.n12283 0.0661418
R47616 vss.n12299 vss.n12294 0.0661418
R47617 vss.n12294 vss.n12291 0.0661418
R47618 vss.n12298 vss.n12295 0.0661418
R47619 vss.n12295 vss.n2351 0.0661418
R47620 vss.n12313 vss.n12285 0.0661418
R47621 vss.n12285 vss.n2153 0.0661418
R47622 vss.n12337 vss.n12324 0.0661418
R47623 vss.n12338 vss.n12337 0.0661418
R47624 vss.n12331 vss.n12328 0.0661418
R47625 vss.n12329 vss.n12328 0.0661418
R47626 vss.n12344 vss.n12339 0.0661418
R47627 vss.n12339 vss.n12336 0.0661418
R47628 vss.n12343 vss.n12340 0.0661418
R47629 vss.n12340 vss.n2352 0.0661418
R47630 vss.n12358 vss.n12330 0.0661418
R47631 vss.n12330 vss.n2154 0.0661418
R47632 vss.n10233 vss.n10220 0.0661418
R47633 vss.n10234 vss.n10233 0.0661418
R47634 vss.n10227 vss.n10224 0.0661418
R47635 vss.n10225 vss.n10224 0.0661418
R47636 vss.n10240 vss.n10235 0.0661418
R47637 vss.n10235 vss.n10232 0.0661418
R47638 vss.n10239 vss.n10236 0.0661418
R47639 vss.n10236 vss.n2358 0.0661418
R47640 vss.n10254 vss.n10226 0.0661418
R47641 vss.n10226 vss.n2155 0.0661418
R47642 vss.n2413 vss.n2400 0.0661418
R47643 vss.n2414 vss.n2413 0.0661418
R47644 vss.n2407 vss.n2404 0.0661418
R47645 vss.n2405 vss.n2404 0.0661418
R47646 vss.n2420 vss.n2415 0.0661418
R47647 vss.n2415 vss.n2412 0.0661418
R47648 vss.n2419 vss.n2416 0.0661418
R47649 vss.n2416 vss.n2364 0.0661418
R47650 vss.n2434 vss.n2406 0.0661418
R47651 vss.n2406 vss.n2156 0.0661418
R47652 vss.n2381 vss.n2380 0.0661418
R47653 vss.n2380 vss.n2374 0.0661418
R47654 vss.n2386 vss.n2383 0.0661418
R47655 vss.n2384 vss.n2383 0.0661418
R47656 vss.n2375 vss.n2371 0.0661418
R47657 vss.n2375 vss.n2367 0.0661418
R47658 vss.n2370 vss.n2366 0.0661418
R47659 vss.n12974 vss.n2366 0.0661418
R47660 vss.n2393 vss.n2385 0.0661418
R47661 vss.n2385 vss.n2157 0.0661418
R47662 vss.n10043 vss.n10031 0.0661418
R47663 vss.n10035 vss.n10031 0.0661418
R47664 vss.n10040 vss.n10039 0.0661418
R47665 vss.n10041 vss.n10040 0.0661418
R47666 vss.n2492 vss.n2479 0.0661418
R47667 vss.n2493 vss.n2492 0.0661418
R47668 vss.n2486 vss.n2483 0.0661418
R47669 vss.n2484 vss.n2483 0.0661418
R47670 vss.n2500 vss.n2494 0.0661418
R47671 vss.n2494 vss.n2491 0.0661418
R47672 vss.n2499 vss.n2495 0.0661418
R47673 vss.n2496 vss.n2495 0.0661418
R47674 vss.n2514 vss.n2485 0.0661418
R47675 vss.n2485 vss.n2158 0.0661418
R47676 vss.n2129 vss.n2123 0.0661418
R47677 vss.n2129 vss.n2127 0.0661418
R47678 vss.n2134 vss.n2133 0.0661418
R47679 vss.n2133 vss.n2128 0.0661418
R47680 vss.n13063 vss.n13062 0.0661418
R47681 vss.n13064 vss.n13063 0.0661418
R47682 vss.n13058 vss.n2140 0.0661418
R47683 vss.n13058 vss.n13057 0.0661418
R47684 vss.n13075 vss.n13074 0.0661418
R47685 vss.n13076 vss.n13075 0.0661418
R47686 vss.n11841 vss.n11840 0.0661418
R47687 vss.n11840 vss.n11838 0.0661418
R47688 vss.n12113 vss.n11832 0.0661418
R47689 vss.n12113 vss.n11826 0.0661418
R47690 vss.n11847 vss.n11846 0.0661418
R47691 vss.n11846 vss.n11844 0.0661418
R47692 vss.n11849 vss.n11848 0.0661418
R47693 vss.n12100 vss.n11849 0.0661418
R47694 vss.n12119 vss.n11830 0.0661418
R47695 vss.n11830 vss.n11828 0.0661418
R47696 vss.n12125 vss.n11824 0.0661418
R47697 vss.n11825 vss.n11824 0.0661418
R47698 vss.n11822 vss.n11821 0.0661418
R47699 vss.n11821 vss.n11815 0.0661418
R47700 vss.n11816 vss.n11812 0.0661418
R47701 vss.n11816 vss.n11806 0.0661418
R47702 vss.n12132 vss.n12124 0.0661418
R47703 vss.n12124 vss.n12123 0.0661418
R47704 vss.n11811 vss.n11809 0.0661418
R47705 vss.n11809 vss.n11807 0.0661418
R47706 vss.n11797 vss.n11796 0.0661418
R47707 vss.n11796 vss.n11794 0.0661418
R47708 vss.n12166 vss.n11791 0.0661418
R47709 vss.n12166 vss.n11786 0.0661418
R47710 vss.n11803 vss.n11802 0.0661418
R47711 vss.n11802 vss.n11800 0.0661418
R47712 vss.n11805 vss.n11804 0.0661418
R47713 vss.n12153 vss.n11805 0.0661418
R47714 vss.n12172 vss.n11789 0.0661418
R47715 vss.n11789 vss.n2350 0.0661418
R47716 vss.n12178 vss.n11784 0.0661418
R47717 vss.n11785 vss.n11784 0.0661418
R47718 vss.n12184 vss.n11780 0.0661418
R47719 vss.n12185 vss.n12184 0.0661418
R47720 vss.n12258 vss.n12257 0.0661418
R47721 vss.n12258 vss.n12183 0.0661418
R47722 vss.n12269 vss.n12177 0.0661418
R47723 vss.n12177 vss.n12176 0.0661418
R47724 vss.n12254 vss.n12253 0.0661418
R47725 vss.n12253 vss.n12252 0.0661418
R47726 vss.n12204 vss.n12203 0.0661418
R47727 vss.n12203 vss.n12197 0.0661418
R47728 vss.n12229 vss.n12206 0.0661418
R47729 vss.n12209 vss.n12206 0.0661418
R47730 vss.n12198 vss.n12194 0.0661418
R47731 vss.n12198 vss.n12190 0.0661418
R47732 vss.n12193 vss.n12189 0.0661418
R47733 vss.n12250 vss.n12189 0.0661418
R47734 vss.n12233 vss.n12208 0.0661418
R47735 vss.n12208 vss.n2353 0.0661418
R47736 vss.n12221 vss.n12220 0.0661418
R47737 vss.n12220 vss.n12219 0.0661418
R47738 vss.n11734 vss.n11733 0.0661418
R47739 vss.n11733 vss.n11727 0.0661418
R47740 vss.n11728 vss.n11724 0.0661418
R47741 vss.n11728 vss.n11719 0.0661418
R47742 vss.n12225 vss.n12224 0.0661418
R47743 vss.n12226 vss.n12225 0.0661418
R47744 vss.n11723 vss.n11721 0.0661418
R47745 vss.n11721 vss.n10615 0.0661418
R47746 vss.n11710 vss.n11709 0.0661418
R47747 vss.n11709 vss.n11707 0.0661418
R47748 vss.n12562 vss.n11704 0.0661418
R47749 vss.n12562 vss.n11699 0.0661418
R47750 vss.n11716 vss.n11715 0.0661418
R47751 vss.n11715 vss.n11713 0.0661418
R47752 vss.n11718 vss.n11717 0.0661418
R47753 vss.n12549 vss.n11718 0.0661418
R47754 vss.n12568 vss.n11702 0.0661418
R47755 vss.n11702 vss.n2356 0.0661418
R47756 vss.n11636 vss.n11633 0.0661418
R47757 vss.n11636 vss.n11635 0.0661418
R47758 vss.n11638 vss.n11630 0.0661418
R47759 vss.n11631 vss.n11630 0.0661418
R47760 vss.n11688 vss.n11627 0.0661418
R47761 vss.n11688 vss.n11687 0.0661418
R47762 vss.n12573 vss.n11634 0.0661418
R47763 vss.n12573 vss.n12572 0.0661418
R47764 vss.n12585 vss.n12584 0.0661418
R47765 vss.n12586 vss.n12585 0.0661418
R47766 vss.n11655 vss.n11654 0.0661418
R47767 vss.n11654 vss.n11648 0.0661418
R47768 vss.n11664 vss.n11657 0.0661418
R47769 vss.n11660 vss.n11657 0.0661418
R47770 vss.n11649 vss.n11645 0.0661418
R47771 vss.n11649 vss.n11641 0.0661418
R47772 vss.n11644 vss.n11640 0.0661418
R47773 vss.n11685 vss.n11640 0.0661418
R47774 vss.n11668 vss.n11659 0.0661418
R47775 vss.n11659 vss.n2359 0.0661418
R47776 vss.n10310 vss.n10307 0.0661418
R47777 vss.n10308 vss.n10307 0.0661418
R47778 vss.n10316 vss.n10303 0.0661418
R47779 vss.n10317 vss.n10316 0.0661418
R47780 vss.n12838 vss.n12837 0.0661418
R47781 vss.n12838 vss.n10315 0.0661418
R47782 vss.n12849 vss.n10309 0.0661418
R47783 vss.n11661 vss.n10309 0.0661418
R47784 vss.n12834 vss.n12833 0.0661418
R47785 vss.n12833 vss.n12832 0.0661418
R47786 vss.n12786 vss.n12785 0.0661418
R47787 vss.n12785 vss.n12779 0.0661418
R47788 vss.n12811 vss.n12788 0.0661418
R47789 vss.n12791 vss.n12788 0.0661418
R47790 vss.n12780 vss.n12776 0.0661418
R47791 vss.n12780 vss.n12772 0.0661418
R47792 vss.n12775 vss.n12771 0.0661418
R47793 vss.n12830 vss.n12771 0.0661418
R47794 vss.n12815 vss.n12790 0.0661418
R47795 vss.n12790 vss.n2362 0.0661418
R47796 vss.n12803 vss.n12802 0.0661418
R47797 vss.n12802 vss.n12801 0.0661418
R47798 vss.n10099 vss.n10098 0.0661418
R47799 vss.n10098 vss.n10092 0.0661418
R47800 vss.n10093 vss.n10089 0.0661418
R47801 vss.n10093 vss.n10083 0.0661418
R47802 vss.n12807 vss.n12806 0.0661418
R47803 vss.n12808 vss.n12807 0.0661418
R47804 vss.n10088 vss.n10086 0.0661418
R47805 vss.n10086 vss.n10084 0.0661418
R47806 vss.n10080 vss.n10079 0.0661418
R47807 vss.n10079 vss.n10077 0.0661418
R47808 vss.n10074 vss.n10073 0.0661418
R47809 vss.n10073 vss.n10071 0.0661418
R47810 vss.n10069 vss.n10063 0.0661418
R47811 vss.n10069 vss.n10058 0.0661418
R47812 vss.n10082 vss.n10081 0.0661418
R47813 vss.n12922 vss.n10082 0.0661418
R47814 vss.n10032 vss.n10030 0.0661418
R47815 vss.n10030 vss.n10029 0.0661418
R47816 vss.n10024 vss.n10017 0.0661418
R47817 vss.n10024 vss.n10022 0.0661418
R47818 vss.n10053 vss.n10052 0.0661418
R47819 vss.n10052 vss.n10023 0.0661418
R47820 vss.n10055 vss.n10054 0.0661418
R47821 vss.n12943 vss.n10055 0.0661418
R47822 vss.n12939 vss.n10061 0.0661418
R47823 vss.n10061 vss.n2365 0.0661418
R47824 vss.n13090 vss.n13089 0.0661418
R47825 vss.n13091 vss.n13090 0.0661418
R47826 vss.n2108 vss.n2101 0.0661418
R47827 vss.n2104 vss.n2101 0.0661418
R47828 vss.n2113 vss.n2112 0.0661418
R47829 vss.n2112 vss.n2105 0.0661418
R47830 vss.n2115 vss.n2114 0.0661418
R47831 vss.n13078 vss.n2115 0.0661418
R47832 vss.n2082 vss.n2076 0.0661418
R47833 vss.n2082 vss.n2080 0.0661418
R47834 vss.n2087 vss.n2086 0.0661418
R47835 vss.n2086 vss.n2081 0.0661418
R47836 vss.n13099 vss.n13098 0.0661418
R47837 vss.n13100 vss.n13099 0.0661418
R47838 vss.n13094 vss.n2093 0.0661418
R47839 vss.n13094 vss.n13093 0.0661418
R47840 vss.n13111 vss.n13110 0.0661418
R47841 vss.n13112 vss.n13111 0.0661418
R47842 vss.n12096 vss.n12095 0.0661418
R47843 vss.n12097 vss.n12096 0.0661418
R47844 vss.n11871 vss.n11870 0.0661418
R47845 vss.n11870 vss.n11865 0.0661418
R47846 vss.n11877 vss.n11876 0.0661418
R47847 vss.n11876 vss.n11874 0.0661418
R47848 vss.n11868 vss.n11861 0.0661418
R47849 vss.n11868 vss.n11866 0.0661418
R47850 vss.n12085 vss.n12084 0.0661418
R47851 vss.n12086 vss.n12085 0.0661418
R47852 vss.n11879 vss.n11878 0.0661418
R47853 vss.n11879 vss.n2048 0.0661418
R47854 vss.n10472 vss.n10461 0.0661418
R47855 vss.n10472 vss.n10466 0.0661418
R47856 vss.n10477 vss.n10475 0.0661418
R47857 vss.n10475 vss.n10474 0.0661418
R47858 vss.n10497 vss.n10468 0.0661418
R47859 vss.n10498 vss.n10497 0.0661418
R47860 vss.n10493 vss.n10469 0.0661418
R47861 vss.n10469 vss.n2052 0.0661418
R47862 vss.n10480 vss.n10476 0.0661418
R47863 vss.n10476 vss.n10420 0.0661418
R47864 vss.n10693 vss.n10682 0.0661418
R47865 vss.n10693 vss.n10687 0.0661418
R47866 vss.n10698 vss.n10696 0.0661418
R47867 vss.n10696 vss.n10695 0.0661418
R47868 vss.n10718 vss.n10689 0.0661418
R47869 vss.n10719 vss.n10718 0.0661418
R47870 vss.n10714 vss.n10690 0.0661418
R47871 vss.n10690 vss.n2058 0.0661418
R47872 vss.n10701 vss.n10697 0.0661418
R47873 vss.n10697 vss.n10421 0.0661418
R47874 vss.n11007 vss.n10996 0.0661418
R47875 vss.n11007 vss.n11001 0.0661418
R47876 vss.n11012 vss.n11010 0.0661418
R47877 vss.n11010 vss.n11009 0.0661418
R47878 vss.n11032 vss.n11003 0.0661418
R47879 vss.n11033 vss.n11032 0.0661418
R47880 vss.n11028 vss.n11004 0.0661418
R47881 vss.n11004 vss.n2064 0.0661418
R47882 vss.n11015 vss.n11011 0.0661418
R47883 vss.n11011 vss.n10422 0.0661418
R47884 vss.n11133 vss.n11132 0.0661418
R47885 vss.n11132 vss.n11111 0.0661418
R47886 vss.n11112 vss.n11105 0.0661418
R47887 vss.n11112 vss.n11110 0.0661418
R47888 vss.n11120 vss.n11118 0.0661418
R47889 vss.n11118 vss.n11117 0.0661418
R47890 vss.n11123 vss.n11119 0.0661418
R47891 vss.n11119 vss.n10423 0.0661418
R47892 vss.n11137 vss.n11134 0.0661418
R47893 vss.n11137 vss.n2070 0.0661418
R47894 vss.n13549 vss 0.0465526
R47895 vss.n13650 vss 0.0465526
R47896 vss.n13702 vss 0.0465526
R47897 vss.n13755 vss 0.0465526
R47898 vss.n13807 vss 0.0465526
R47899 vss.n13860 vss 0.0465526
R47900 vss.n13318 vss 0.0465526
R47901 vss.n14139 vss 0.0465526
R47902 vss.n8057 vss 0.0465526
R47903 vss.n7871 vss 0.0465526
R47904 vss.n8402 vss 0.0465526
R47905 vss.n8500 vss 0.0465526
R47906 vss.n8471 vss 0.0465526
R47907 vss.n8373 vss 0.0465526
R47908 vss.n8255 vss 0.0465526
R47909 vss.n9638 vss 0.0465526
R47910 vss.n3262 vss 0.0465526
R47911 vss.n5205 vss 0.0465526
R47912 vss.n5081 vss 0.0465526
R47913 vss.n5353 vss 0.0465526
R47914 vss.n5324 vss 0.0465526
R47915 vss.n5265 vss 0.0465526
R47916 vss.n5206 vss 0.0465526
R47917 vss.n9736 vss 0.0465526
R47918 vss.n10299 vss 0.0465526
R47919 vss.n11737 vss 0.0465526
R47920 vss.n11779 vss 0.0465526
R47921 vss.n12405 vss 0.0465526
R47922 vss.n10101 vss 0.0465526
R47923 vss.n12956 vss 0.0465526
R47924 vss.n10064 vss 0.0465526
R47925 vss.n11833 vss 0.0465526
R47926 vss vss.n11400 0.0416184
R47927 vss vss.n10768 0.0416184
R47928 vss vss.n10547 0.0416184
R47929 vss.n12013 vss 0.0416184
R47930 vss.n10843 vss 0.0416184
R47931 vss.n11450 vss 0.0416184
R47932 vss.n641 vss 0.0416184
R47933 vss.n1807 vss 0.0416184
R47934 vss vss.n1648 0.0416184
R47935 vss.n1911 vss 0.0416184
R47936 vss vss.n1353 0.0416184
R47937 vss vss.n1093 0.0416184
R47938 vss vss.n1355 0.0416184
R47939 vss vss.n1400 0.0416184
R47940 vss vss.n1407 0.0416184
R47941 vss vss.n1486 0.0416184
R47942 vss.n1651 vss 0.0416184
R47943 vss.n1695 vss 0.0416184
R47944 vss vss.n1488 0.0416184
R47945 vss vss.n1567 0.0416184
R47946 vss.n553 vss 0.0416184
R47947 vss.n13955 vss 0.0416184
R47948 vss vss.n1568 0.0416184
R47949 vss.n890 vss 0.0416184
R47950 vss vss.n14031 0.0416184
R47951 vss vss.n1136 0.0416184
R47952 vss vss.n1983 0.0416184
R47953 vss vss.n2027 0.0416184
R47954 vss vss.n13202 0.0416184
R47955 vss vss.n6053 0.0416184
R47956 vss.n7049 vss 0.0416184
R47957 vss vss.n6672 0.0416184
R47958 vss.n9212 vss 0.0416184
R47959 vss vss.n6445 0.0416184
R47960 vss vss.n6368 0.0416184
R47961 vss vss.n9254 0.0416184
R47962 vss vss.n6904 0.0416184
R47963 vss.n6985 vss 0.0416184
R47964 vss vss.n6982 0.0416184
R47965 vss vss.n7091 0.0416184
R47966 vss.n6715 vss 0.0416184
R47967 vss.n7176 vss 0.0416184
R47968 vss vss.n7171 0.0416184
R47969 vss.n6093 vss 0.0416184
R47970 vss.n9504 vss 0.0416184
R47971 vss vss.n7172 0.0416184
R47972 vss.n9428 vss 0.0416184
R47973 vss vss.n9580 0.0416184
R47974 vss vss.n9147 0.0416184
R47975 vss.n9148 vss 0.0416184
R47976 vss vss.n9363 0.0416184
R47977 vss.n9365 vss 0.0416184
R47978 vss vss.n4364 0.0416184
R47979 vss vss.n3719 0.0416184
R47980 vss vss.n3499 0.0416184
R47981 vss.n3578 vss 0.0416184
R47982 vss vss.n4065 0.0416184
R47983 vss.n4615 vss 0.0416184
R47984 vss.n2672 vss 0.0416184
R47985 vss vss.n9992 0.0416184
R47986 vss vss.n5741 0.0416184
R47987 vss.n5742 vss 0.0416184
R47988 vss vss.n3425 0.0416184
R47989 vss vss.n5846 0.0416184
R47990 vss vss.n3947 0.0416184
R47991 vss.n4075 vss 0.0416184
R47992 vss vss.n4022 0.0416184
R47993 vss vss.n4071 0.0416184
R47994 vss.n3800 vss 0.0416184
R47995 vss vss.n4213 0.0416184
R47996 vss vss.n4289 0.0416184
R47997 vss.n4367 vss 0.0416184
R47998 vss vss.n4458 0.0416184
R47999 vss.n4459 vss 0.0416184
R48000 vss vss.n5933 0.0416184
R48001 vss vss.n11923 0.0416184
R48002 vss.n11924 vss 0.0416184
R48003 vss vss.n10504 0.0416184
R48004 vss vss.n12617 0.0416184
R48005 vss vss.n10680 0.0416184
R48006 vss.n11550 vss 0.0416184
R48007 vss vss.n10725 0.0416184
R48008 vss vss.n11546 0.0416184
R48009 vss vss.n10975 0.0416184
R48010 vss vss.n10994 0.0416184
R48011 vss vss.n11039 0.0416184
R48012 vss.n11403 vss 0.0416184
R48013 vss vss.n10372 0.0416184
R48014 vss vss.n11041 0.0416184
R48015 vss vss.n11148 0.0416184
R48016 vss vss.n12663 0.0416184
R48017 vss vss.n12664 0.0416184
R48018 vss.n11970 vss.n11969 0.0284605
R48019 vss.n11596 vss.n11595 0.0284605
R48020 vss.n10990 vss.n10989 0.0284605
R48021 vss.n12699 vss.n12698 0.0284605
R48022 vss.n1979 vss.n1978 0.0284605
R48023 vss.n13550 vss.n13549 0.0284605
R48024 vss.n13651 vss.n13650 0.0284605
R48025 vss.n13703 vss.n13702 0.0284605
R48026 vss.n13756 vss.n13755 0.0284605
R48027 vss.n13808 vss.n13807 0.0284605
R48028 vss.n13861 vss.n13860 0.0284605
R48029 vss.n13319 vss.n13318 0.0284605
R48030 vss.n14140 vss.n14139 0.0284605
R48031 vss.n13238 vss.n13237 0.0284605
R48032 vss.n1403 vss.n1402 0.0284605
R48033 vss.n1909 vss.n1908 0.0284605
R48034 vss.n1805 vss.n1804 0.0284605
R48035 vss.n593 vss.n592 0.0284605
R48036 vss.n14027 vss.n14026 0.0284605
R48037 vss.n13157 vss.n13156 0.0284605
R48038 vss.n9195 vss.n9194 0.0284605
R48039 vss.n8058 vss.n8057 0.0284605
R48040 vss.n7872 vss.n7871 0.0284605
R48041 vss.n8403 vss.n8402 0.0284605
R48042 vss.n8501 vss.n8500 0.0284605
R48043 vss.n8472 vss.n8471 0.0284605
R48044 vss.n8374 vss.n8373 0.0284605
R48045 vss.n8256 vss.n8255 0.0284605
R48046 vss.n9639 vss.n9638 0.0284605
R48047 vss.n7223 vss.n7222 0.0284605
R48048 vss.n7032 vss.n7031 0.0284605
R48049 vss.n9250 vss.n9249 0.0284605
R48050 vss.n7087 vss.n7086 0.0284605
R48051 vss.n6133 vss.n6132 0.0284605
R48052 vss.n9576 vss.n9575 0.0284605
R48053 vss.n6544 vss.n6543 0.0284605
R48054 vss.n4641 vss.n3262 0.0284605
R48055 vss.n5205 vss.n5204 0.0284605
R48056 vss.n5081 vss.n5080 0.0284605
R48057 vss.n5354 vss.n5353 0.0284605
R48058 vss.n5325 vss.n5324 0.0284605
R48059 vss.n5266 vss.n5265 0.0284605
R48060 vss.n5207 vss.n5206 0.0284605
R48061 vss.n9737 vss.n9736 0.0284605
R48062 vss.n5789 vss.n5788 0.0284605
R48063 vss.n4122 vss.n4121 0.0284605
R48064 vss.n4209 vss.n4208 0.0284605
R48065 vss.n4506 vss.n4505 0.0284605
R48066 vss.n3600 vss.n3599 0.0284605
R48067 vss.n5842 vss.n5841 0.0284605
R48068 vss.n4067 vss.n4066 0.0284605
R48069 vss.n4613 vss.n4612 0.0284605
R48070 vss.n11675 vss.n10299 0.0284605
R48071 vss.n12240 vss.n11737 0.0284605
R48072 vss.n12138 vss.n11779 0.0284605
R48073 vss.n12405 vss.n12404 0.0284605
R48074 vss.n10300 vss.n10101 0.0284605
R48075 vss.n12956 vss.n12955 0.0284605
R48076 vss.n10065 vss.n10064 0.0284605
R48077 vss.n11834 vss.n11833 0.0284605
R48078 vss.n11889 vss.n2030 0.0284605
R48079 vss.n12613 vss.n12612 0.0284605
R48080 vss.n11542 vss.n11541 0.0284605
R48081 vss.n11448 vss.n11447 0.0284605
R48082 vss.n11401 vss.n11357 0.021882
R48083 vss.n11231 vss.n10769 0.021882
R48084 vss.n11292 vss.n10548 0.021882
R48085 vss.n412 vss.n411 0.021882
R48086 vss.n289 vss.n288 0.021882
R48087 vss.n14446 vss.n14445 0.021882
R48088 vss.n230 vss.n229 0.021882
R48089 vss.n14641 vss.n14640 0.021882
R48090 vss.n153 vss.n152 0.021882
R48091 vss.n14251 vss.n380 0.021882
R48092 vss.n7373 vss.n6006 0.021882
R48093 vss.n7847 vss.n7846 0.021882
R48094 vss.n7660 vss.n7659 0.021882
R48095 vss.n7471 vss.n7470 0.021882
R48096 vss.n8979 vss.n8978 0.021882
R48097 vss.n8859 vss.n7624 0.021882
R48098 vss.n8740 vss.n7767 0.021882
R48099 vss.n8249 vss.n7988 0.021882
R48100 vss.n3261 vss.n3260 0.021882
R48101 vss.n3104 vss.n3103 0.021882
R48102 vss.n5078 vss.n5077 0.021882
R48103 vss.n2870 vss.n2869 0.021882
R48104 vss.n9849 vss.n9848 0.021882
R48105 vss.n5318 vss.n5000 0.021882
R48106 vss.n5259 vss.n5202 0.021882
R48107 vss.n9789 vss.n3183 0.021882
R48108 vss.n12905 vss.n10219 0.021882
R48109 vss.n12531 vss.n12530 0.021882
R48110 vss.n2239 vss.n2238 0.021882
R48111 vss.n12402 vss.n12401 0.021882
R48112 vss.n10298 vss.n10297 0.021882
R48113 vss.n2478 vss.n2477 0.021882
R48114 vss.n12961 vss.n2556 0.021882
R48115 vss.n13023 vss.n13022 0.021882
R48116 vss.n12619 vss.n10460 0.021882
R48117 vss.n11548 vss.n10681 0.021882
R48118 vss.n11200 vss.n11040 0.021882
R48119 vss.n11150 vss.n11149 0.021882
R48120 vss.n12666 vss.n12665 0.021882
R48121 vss.n14762 vss.n14761 0.021882
R48122 vss.n11969 vss 0.0136579
R48123 vss.n11595 vss 0.0136579
R48124 vss.n10990 vss 0.0136579
R48125 vss.n12698 vss 0.0136579
R48126 vss.n1979 vss 0.0136579
R48127 vss.n13237 vss 0.0136579
R48128 vss.n1403 vss 0.0136579
R48129 vss.n1909 vss 0.0136579
R48130 vss.n1805 vss 0.0136579
R48131 vss.n593 vss 0.0136579
R48132 vss.n14027 vss 0.0136579
R48133 vss.n13157 vss 0.0136579
R48134 vss.n9194 vss 0.0136579
R48135 vss.n7222 vss 0.0136579
R48136 vss.n7031 vss 0.0136579
R48137 vss.n9250 vss 0.0136579
R48138 vss.n7087 vss 0.0136579
R48139 vss.n6133 vss 0.0136579
R48140 vss.n9576 vss 0.0136579
R48141 vss.n6543 vss 0.0136579
R48142 vss.n5788 vss 0.0136579
R48143 vss.n4121 vss 0.0136579
R48144 vss.n4209 vss 0.0136579
R48145 vss.n4505 vss 0.0136579
R48146 vss.n3599 vss 0.0136579
R48147 vss.n5842 vss 0.0136579
R48148 vss.n4067 vss 0.0136579
R48149 vss.n4613 vss 0.0136579
R48150 vss.n2030 vss 0.0136579
R48151 vss.n12613 vss 0.0136579
R48152 vss.n11542 vss 0.0136579
R48153 vss.n11448 vss 0.0136579
R48154 vss.n14768 vss.n14767 0.0126193
R48155 vss.n14767 vss.t26 0.0126193
R48156 vss.n108 vss.n107 0.0126193
R48157 vss.n107 vss.t26 0.0126193
R48158 vss.n119 vss.n118 0.0126193
R48159 vss.n118 vss.t26 0.0126193
R48160 vss.n113 vss.n112 0.0126193
R48161 vss.n112 vss.t26 0.0126193
R48162 vss.n102 vss.n100 0.0126193
R48163 vss.n100 vss.t26 0.0126193
R48164 vss.n131 vss.n130 0.0126193
R48165 vss.n130 vss.t26 0.0126193
R48166 vss.n148 vss.t26 0.0126193
R48167 vss.n127 vss.n126 0.0126193
R48168 vss.n126 vss.t26 0.0126193
R48169 vss.n149 vss.n148 0.0126193
R48170 vss.n143 vss.n142 0.0126193
R48171 vss.n142 vss.t26 0.0126193
R48172 vss.n136 vss.n135 0.0126193
R48173 vss.n135 vss.t26 0.0126193
R48174 vss.n14619 vss.n14618 0.0126193
R48175 vss.n14618 vss.t26 0.0126193
R48176 vss.n14636 vss.t26 0.0126193
R48177 vss.n14615 vss.n14614 0.0126193
R48178 vss.n14614 vss.t26 0.0126193
R48179 vss.n14637 vss.n14636 0.0126193
R48180 vss.n14631 vss.n14630 0.0126193
R48181 vss.n14630 vss.t26 0.0126193
R48182 vss.n14624 vss.n14623 0.0126193
R48183 vss.n14623 vss.t26 0.0126193
R48184 vss.n208 vss.n207 0.0126193
R48185 vss.n207 vss.t26 0.0126193
R48186 vss.n225 vss.t26 0.0126193
R48187 vss.n204 vss.n203 0.0126193
R48188 vss.n203 vss.t26 0.0126193
R48189 vss.n226 vss.n225 0.0126193
R48190 vss.n220 vss.n219 0.0126193
R48191 vss.n219 vss.t26 0.0126193
R48192 vss.n213 vss.n212 0.0126193
R48193 vss.n212 vss.t26 0.0126193
R48194 vss.n14424 vss.n14423 0.0126193
R48195 vss.n14423 vss.t26 0.0126193
R48196 vss.n14441 vss.t26 0.0126193
R48197 vss.n14420 vss.n14419 0.0126193
R48198 vss.n14419 vss.t26 0.0126193
R48199 vss.n14442 vss.n14441 0.0126193
R48200 vss.n14436 vss.n14435 0.0126193
R48201 vss.n14435 vss.t26 0.0126193
R48202 vss.n14429 vss.n14428 0.0126193
R48203 vss.n14428 vss.t26 0.0126193
R48204 vss.n267 vss.n266 0.0126193
R48205 vss.n266 vss.t26 0.0126193
R48206 vss.n284 vss.t26 0.0126193
R48207 vss.n263 vss.n262 0.0126193
R48208 vss.n262 vss.t26 0.0126193
R48209 vss.n285 vss.n284 0.0126193
R48210 vss.n279 vss.n278 0.0126193
R48211 vss.n278 vss.t26 0.0126193
R48212 vss.n272 vss.n271 0.0126193
R48213 vss.n271 vss.t26 0.0126193
R48214 vss.n390 vss.n389 0.0126193
R48215 vss.n389 vss.t26 0.0126193
R48216 vss.n407 vss.t26 0.0126193
R48217 vss.n386 vss.n385 0.0126193
R48218 vss.n385 vss.t26 0.0126193
R48219 vss.n408 vss.n407 0.0126193
R48220 vss.n402 vss.n401 0.0126193
R48221 vss.n401 vss.t26 0.0126193
R48222 vss.n395 vss.n394 0.0126193
R48223 vss.n394 vss.t26 0.0126193
R48224 vss.n14780 vss.n14779 0.0126193
R48225 vss.n14780 vss.t26 0.0126193
R48226 vss.n364 vss.n363 0.0126193
R48227 vss.n363 vss.t26 0.0126193
R48228 vss.n368 vss.n367 0.0126193
R48229 vss.n367 vss.t26 0.0126193
R48230 vss.n374 vss.n369 0.0126193
R48231 vss.n369 vss.t26 0.0126193
R48232 vss.n14775 vss.t26 0.0126193
R48233 vss.n14776 vss.n14775 0.0126193
R48234 vss.n9316 vss.n9315 0.0126193
R48235 vss.t27 vss.n9316 0.0126193
R48236 vss.t27 vss.n9302 0.0126193
R48237 vss.n9312 vss.n9302 0.0126193
R48238 vss.n9318 vss.n9317 0.0126193
R48239 vss.n9317 vss.t27 0.0126193
R48240 vss.t27 vss.n9301 0.0126193
R48241 vss.n9301 vss.n9300 0.0126193
R48242 vss.n9297 vss.n9287 0.0126193
R48243 vss.t27 vss.n9287 0.0126193
R48244 vss.n9286 vss.n9285 0.0126193
R48245 vss.t27 vss.n9286 0.0126193
R48246 vss.t27 vss.n6319 0.0126193
R48247 vss.n6323 vss.n6319 0.0126193
R48248 vss.n9266 vss.n6318 0.0126193
R48249 vss.t27 vss.n6318 0.0126193
R48250 vss.t27 vss.n6317 0.0126193
R48251 vss.n9276 vss.n6317 0.0126193
R48252 vss.n9263 vss.n6316 0.0126193
R48253 vss.t27 vss.n6316 0.0126193
R48254 vss.n6379 vss.n6315 0.0126193
R48255 vss.t27 vss.n6315 0.0126193
R48256 vss.t27 vss.n6314 0.0126193
R48257 vss.n6380 vss.n6314 0.0126193
R48258 vss.n6400 vss.n6313 0.0126193
R48259 vss.t27 vss.n6313 0.0126193
R48260 vss.t27 vss.n6312 0.0126193
R48261 vss.n6375 vss.n6312 0.0126193
R48262 vss.n6391 vss.n6311 0.0126193
R48263 vss.t27 vss.n6311 0.0126193
R48264 vss.n6915 vss.n6310 0.0126193
R48265 vss.t27 vss.n6310 0.0126193
R48266 vss.t27 vss.n6309 0.0126193
R48267 vss.n6916 vss.n6309 0.0126193
R48268 vss.n6936 vss.n6308 0.0126193
R48269 vss.t27 vss.n6308 0.0126193
R48270 vss.t27 vss.n6307 0.0126193
R48271 vss.n6911 vss.n6307 0.0126193
R48272 vss.n6927 vss.n6306 0.0126193
R48273 vss.t27 vss.n6306 0.0126193
R48274 vss.n6606 vss.n6305 0.0126193
R48275 vss.t27 vss.n6305 0.0126193
R48276 vss.t27 vss.n6304 0.0126193
R48277 vss.n6607 vss.n6304 0.0126193
R48278 vss.n6627 vss.n6303 0.0126193
R48279 vss.t27 vss.n6303 0.0126193
R48280 vss.t27 vss.n6302 0.0126193
R48281 vss.n6602 vss.n6302 0.0126193
R48282 vss.n6618 vss.n6301 0.0126193
R48283 vss.t27 vss.n6301 0.0126193
R48284 vss.n7104 vss.n6300 0.0126193
R48285 vss.t27 vss.n6300 0.0126193
R48286 vss.t27 vss.n6299 0.0126193
R48287 vss.n7105 vss.n6299 0.0126193
R48288 vss.n7125 vss.n6298 0.0126193
R48289 vss.t27 vss.n6298 0.0126193
R48290 vss.t27 vss.n6297 0.0126193
R48291 vss.n7100 vss.n6297 0.0126193
R48292 vss.n7116 vss.n6296 0.0126193
R48293 vss.t27 vss.n6296 0.0126193
R48294 vss.n6295 vss.n6294 0.0126193
R48295 vss.t27 vss.n6295 0.0126193
R48296 vss.t27 vss.n6261 0.0126193
R48297 vss.n6265 vss.n6261 0.0126193
R48298 vss.n6275 vss.n6260 0.0126193
R48299 vss.t27 vss.n6260 0.0126193
R48300 vss.t27 vss.n6259 0.0126193
R48301 vss.n6285 vss.n6259 0.0126193
R48302 vss.n6272 vss.n6258 0.0126193
R48303 vss.t27 vss.n6258 0.0126193
R48304 vss.n6257 vss.n6256 0.0126193
R48305 vss.t27 vss.n6257 0.0126193
R48306 vss.t27 vss.n6224 0.0126193
R48307 vss.n6228 vss.n6224 0.0126193
R48308 vss.n6237 vss.n6223 0.0126193
R48309 vss.t27 vss.n6223 0.0126193
R48310 vss.t27 vss.n6222 0.0126193
R48311 vss.n6247 vss.n6222 0.0126193
R48312 vss.n6234 vss.n6221 0.0126193
R48313 vss.t27 vss.n6221 0.0126193
R48314 vss.n3235 vss.n2796 0.0126193
R48315 vss.t77 vss.n2796 0.0126193
R48316 vss.n3233 vss.n2795 0.0126193
R48317 vss.t77 vss.n2795 0.0126193
R48318 vss.n3230 vss.n2792 0.0126193
R48319 vss.t77 vss.n2792 0.0126193
R48320 vss.n3254 vss.n2794 0.0126193
R48321 vss.t77 vss.n2794 0.0126193
R48322 vss.n3242 vss.n2797 0.0126193
R48323 vss.t77 vss.n2797 0.0126193
R48324 vss.n3158 vss.n2800 0.0126193
R48325 vss.t77 vss.n2800 0.0126193
R48326 vss.n3156 vss.n2799 0.0126193
R48327 vss.t77 vss.n2799 0.0126193
R48328 vss.n3153 vss.n2791 0.0126193
R48329 vss.t77 vss.n2791 0.0126193
R48330 vss.n3177 vss.n2798 0.0126193
R48331 vss.t77 vss.n2798 0.0126193
R48332 vss.n3165 vss.n2801 0.0126193
R48333 vss.t77 vss.n2801 0.0126193
R48334 vss.n3078 vss.n2804 0.0126193
R48335 vss.t77 vss.n2804 0.0126193
R48336 vss.n3076 vss.n2803 0.0126193
R48337 vss.t77 vss.n2803 0.0126193
R48338 vss.n3073 vss.n2790 0.0126193
R48339 vss.t77 vss.n2790 0.0126193
R48340 vss.n3097 vss.n2802 0.0126193
R48341 vss.t77 vss.n2802 0.0126193
R48342 vss.n3085 vss.n2805 0.0126193
R48343 vss.t77 vss.n2805 0.0126193
R48344 vss.n5177 vss.n2808 0.0126193
R48345 vss.t77 vss.n2808 0.0126193
R48346 vss.n5175 vss.n2807 0.0126193
R48347 vss.t77 vss.n2807 0.0126193
R48348 vss.n5172 vss.n2789 0.0126193
R48349 vss.t77 vss.n2789 0.0126193
R48350 vss.n5196 vss.n2806 0.0126193
R48351 vss.t77 vss.n2806 0.0126193
R48352 vss.n5184 vss.n2809 0.0126193
R48353 vss.t77 vss.n2809 0.0126193
R48354 vss.n5052 vss.n2812 0.0126193
R48355 vss.t77 vss.n2812 0.0126193
R48356 vss.n5050 vss.n2811 0.0126193
R48357 vss.t77 vss.n2811 0.0126193
R48358 vss.n5047 vss.n2788 0.0126193
R48359 vss.t77 vss.n2788 0.0126193
R48360 vss.n5071 vss.n2810 0.0126193
R48361 vss.t77 vss.n2810 0.0126193
R48362 vss.n5059 vss.n2813 0.0126193
R48363 vss.t77 vss.n2813 0.0126193
R48364 vss.n4975 vss.n2816 0.0126193
R48365 vss.t77 vss.n2816 0.0126193
R48366 vss.n4973 vss.n2815 0.0126193
R48367 vss.t77 vss.n2815 0.0126193
R48368 vss.n4970 vss.n2787 0.0126193
R48369 vss.t77 vss.n2787 0.0126193
R48370 vss.n4994 vss.n2814 0.0126193
R48371 vss.t77 vss.n2814 0.0126193
R48372 vss.n4982 vss.n2817 0.0126193
R48373 vss.t77 vss.n2817 0.0126193
R48374 vss.n2844 vss.n2820 0.0126193
R48375 vss.t77 vss.n2820 0.0126193
R48376 vss.n2842 vss.n2819 0.0126193
R48377 vss.t77 vss.n2819 0.0126193
R48378 vss.n2839 vss.n2786 0.0126193
R48379 vss.t77 vss.n2786 0.0126193
R48380 vss.n2863 vss.n2818 0.0126193
R48381 vss.t77 vss.n2818 0.0126193
R48382 vss.n2851 vss.n2821 0.0126193
R48383 vss.t77 vss.n2821 0.0126193
R48384 vss.n2828 vss.n2824 0.0126193
R48385 vss.t77 vss.n2824 0.0126193
R48386 vss.n9852 vss.n2823 0.0126193
R48387 vss.t77 vss.n2823 0.0126193
R48388 vss.n9862 vss.n2785 0.0126193
R48389 vss.t77 vss.n2785 0.0126193
R48390 vss.n2834 vss.n2822 0.0126193
R48391 vss.t77 vss.n2822 0.0126193
R48392 vss.n9872 vss.n9871 0.0126193
R48393 vss.t77 vss.n9872 0.0126193
R48394 vss.n988 vss.n986 0.0126193
R48395 vss.n986 vss.t83 0.0126193
R48396 vss.n992 vss.t83 0.0126193
R48397 vss.n992 vss.n989 0.0126193
R48398 vss.n1015 vss.n1014 0.0126193
R48399 vss.n1014 vss.t83 0.0126193
R48400 vss.n1007 vss.t83 0.0126193
R48401 vss.n1008 vss.n1007 0.0126193
R48402 vss.n1003 vss.n1002 0.0126193
R48403 vss.n1002 vss.t83 0.0126193
R48404 vss.n1023 vss.n1022 0.0126193
R48405 vss.n1022 vss.t83 0.0126193
R48406 vss.n1027 vss.t83 0.0126193
R48407 vss.n1028 vss.n1027 0.0126193
R48408 vss.n1048 vss.n1047 0.0126193
R48409 vss.n1047 vss.t83 0.0126193
R48410 vss.n1040 vss.t83 0.0126193
R48411 vss.n1041 vss.n1040 0.0126193
R48412 vss.n1036 vss.n1035 0.0126193
R48413 vss.n1035 vss.t83 0.0126193
R48414 vss.n1284 vss.n1283 0.0126193
R48415 vss.n1283 vss.t83 0.0126193
R48416 vss.n1288 vss.t83 0.0126193
R48417 vss.n1289 vss.n1288 0.0126193
R48418 vss.n1309 vss.n1308 0.0126193
R48419 vss.n1308 vss.t83 0.0126193
R48420 vss.n1301 vss.t83 0.0126193
R48421 vss.n1302 vss.n1301 0.0126193
R48422 vss.n1297 vss.n1296 0.0126193
R48423 vss.n1296 vss.t83 0.0126193
R48424 vss.n1416 vss.n1415 0.0126193
R48425 vss.n1415 vss.t83 0.0126193
R48426 vss.n1420 vss.t83 0.0126193
R48427 vss.n1421 vss.n1420 0.0126193
R48428 vss.n1441 vss.n1440 0.0126193
R48429 vss.n1440 vss.t83 0.0126193
R48430 vss.n1433 vss.t83 0.0126193
R48431 vss.n1434 vss.n1433 0.0126193
R48432 vss.n1429 vss.n1428 0.0126193
R48433 vss.n1428 vss.t83 0.0126193
R48434 vss.n1579 vss.n1578 0.0126193
R48435 vss.n1578 vss.t83 0.0126193
R48436 vss.n1583 vss.t83 0.0126193
R48437 vss.n1584 vss.n1583 0.0126193
R48438 vss.n1604 vss.n1603 0.0126193
R48439 vss.n1603 vss.t83 0.0126193
R48440 vss.n1596 vss.t83 0.0126193
R48441 vss.n1597 vss.n1596 0.0126193
R48442 vss.n1592 vss.n1591 0.0126193
R48443 vss.n1591 vss.t83 0.0126193
R48444 vss.n1496 vss.n1495 0.0126193
R48445 vss.n1495 vss.t83 0.0126193
R48446 vss.n1500 vss.t83 0.0126193
R48447 vss.n1501 vss.n1500 0.0126193
R48448 vss.n1521 vss.n1520 0.0126193
R48449 vss.n1520 vss.t83 0.0126193
R48450 vss.n1513 vss.t83 0.0126193
R48451 vss.n1514 vss.n1513 0.0126193
R48452 vss.n1509 vss.n1508 0.0126193
R48453 vss.n1508 vss.t83 0.0126193
R48454 vss.n936 vss.n934 0.0126193
R48455 vss.n934 vss.t83 0.0126193
R48456 vss.n940 vss.t83 0.0126193
R48457 vss.n940 vss.n937 0.0126193
R48458 vss.n963 vss.n962 0.0126193
R48459 vss.n962 vss.t83 0.0126193
R48460 vss.n955 vss.t83 0.0126193
R48461 vss.n956 vss.n955 0.0126193
R48462 vss.n951 vss.n950 0.0126193
R48463 vss.n950 vss.t83 0.0126193
R48464 vss.n505 vss.n503 0.0126193
R48465 vss.t83 vss.n503 0.0126193
R48466 vss.n7352 vss.n7344 0.0126193
R48467 vss.n7352 vss.t25 0.0126193
R48468 vss.n7343 vss.n7341 0.0126193
R48469 vss.n7341 vss.t25 0.0126193
R48470 vss.n7972 vss.n7971 0.0126193
R48471 vss.n7972 vss.t25 0.0126193
R48472 vss.n7961 vss.n7960 0.0126193
R48473 vss.n7960 vss.t25 0.0126193
R48474 vss.n7985 vss.n7984 0.0126193
R48475 vss.n7984 vss.t25 0.0126193
R48476 vss.n7980 vss.n7979 0.0126193
R48477 vss.n7979 vss.t25 0.0126193
R48478 vss.n7967 vss.n7966 0.0126193
R48479 vss.n7966 vss.t25 0.0126193
R48480 vss.n7830 vss.n7829 0.0126193
R48481 vss.n7830 vss.t25 0.0126193
R48482 vss.n7819 vss.n7818 0.0126193
R48483 vss.n7818 vss.t25 0.0126193
R48484 vss.n7843 vss.n7842 0.0126193
R48485 vss.n7842 vss.t25 0.0126193
R48486 vss.n7838 vss.n7837 0.0126193
R48487 vss.n7837 vss.t25 0.0126193
R48488 vss.n7825 vss.n7824 0.0126193
R48489 vss.n7824 vss.t25 0.0126193
R48490 vss.n7751 vss.n7750 0.0126193
R48491 vss.n7751 vss.t25 0.0126193
R48492 vss.n7740 vss.n7739 0.0126193
R48493 vss.n7739 vss.t25 0.0126193
R48494 vss.n7764 vss.n7763 0.0126193
R48495 vss.n7763 vss.t25 0.0126193
R48496 vss.n7759 vss.n7758 0.0126193
R48497 vss.n7758 vss.t25 0.0126193
R48498 vss.n7746 vss.n7745 0.0126193
R48499 vss.n7745 vss.t25 0.0126193
R48500 vss.n7643 vss.n7642 0.0126193
R48501 vss.n7643 vss.t25 0.0126193
R48502 vss.n7632 vss.n7631 0.0126193
R48503 vss.n7631 vss.t25 0.0126193
R48504 vss.n7656 vss.n7655 0.0126193
R48505 vss.n7655 vss.t25 0.0126193
R48506 vss.n7651 vss.n7650 0.0126193
R48507 vss.n7650 vss.t25 0.0126193
R48508 vss.n7638 vss.n7637 0.0126193
R48509 vss.n7637 vss.t25 0.0126193
R48510 vss.n7608 vss.n7607 0.0126193
R48511 vss.n7608 vss.t25 0.0126193
R48512 vss.n7597 vss.n7596 0.0126193
R48513 vss.n7596 vss.t25 0.0126193
R48514 vss.n7621 vss.n7620 0.0126193
R48515 vss.n7620 vss.t25 0.0126193
R48516 vss.n7616 vss.n7615 0.0126193
R48517 vss.n7615 vss.t25 0.0126193
R48518 vss.n7603 vss.n7602 0.0126193
R48519 vss.n7602 vss.t25 0.0126193
R48520 vss.n7454 vss.n7453 0.0126193
R48521 vss.n7454 vss.t25 0.0126193
R48522 vss.n7443 vss.n7442 0.0126193
R48523 vss.n7442 vss.t25 0.0126193
R48524 vss.n7467 vss.n7466 0.0126193
R48525 vss.n7466 vss.t25 0.0126193
R48526 vss.n7462 vss.n7461 0.0126193
R48527 vss.n7461 vss.t25 0.0126193
R48528 vss.n7449 vss.n7448 0.0126193
R48529 vss.n7448 vss.t25 0.0126193
R48530 vss.n7420 vss.n7409 0.0126193
R48531 vss.n7420 vss.t25 0.0126193
R48532 vss.n7415 vss.n7410 0.0126193
R48533 vss.n7415 vss.t25 0.0126193
R48534 vss.n7433 vss.n7432 0.0126193
R48535 vss.n7432 vss.t25 0.0126193
R48536 vss.n7428 vss.n7427 0.0126193
R48537 vss.n7427 vss.t25 0.0126193
R48538 vss.n7408 vss.n7406 0.0126193
R48539 vss.n7406 vss.t25 0.0126193
R48540 vss.n14055 vss.n14054 0.0126193
R48541 vss.n14054 vss.t242 0.0126193
R48542 vss.n14038 vss.n14037 0.0126193
R48543 vss.n14037 vss.t242 0.0126193
R48544 vss.n14046 vss.t242 0.0126193
R48545 vss.n14047 vss.n14046 0.0126193
R48546 vss.n14042 vss.n14041 0.0126193
R48547 vss.n14041 vss.t242 0.0126193
R48548 vss.n7369 vss.t257 0.0126193
R48549 vss.n7351 vss.n7345 0.0126193
R48550 vss.n7351 vss.t257 0.0126193
R48551 vss.n7369 vss.n7368 0.0126193
R48552 vss.n7364 vss.n7363 0.0126193
R48553 vss.n7364 vss.t257 0.0126193
R48554 vss.n2531 vss.n2174 0.0126193
R48555 vss.t76 vss.n2174 0.0126193
R48556 vss.n2529 vss.n2173 0.0126193
R48557 vss.t76 vss.n2173 0.0126193
R48558 vss.n2526 vss.n2170 0.0126193
R48559 vss.t76 vss.n2170 0.0126193
R48560 vss.n2550 vss.n2172 0.0126193
R48561 vss.t76 vss.n2172 0.0126193
R48562 vss.n2538 vss.n2175 0.0126193
R48563 vss.t76 vss.n2175 0.0126193
R48564 vss.n2452 vss.n2178 0.0126193
R48565 vss.t76 vss.n2178 0.0126193
R48566 vss.n2450 vss.n2177 0.0126193
R48567 vss.t76 vss.n2177 0.0126193
R48568 vss.n2447 vss.n2169 0.0126193
R48569 vss.t76 vss.n2169 0.0126193
R48570 vss.n2471 vss.n2176 0.0126193
R48571 vss.t76 vss.n2176 0.0126193
R48572 vss.n2459 vss.n2179 0.0126193
R48573 vss.t76 vss.n2179 0.0126193
R48574 vss.n10194 vss.n2182 0.0126193
R48575 vss.t76 vss.n2182 0.0126193
R48576 vss.n10192 vss.n2181 0.0126193
R48577 vss.t76 vss.n2181 0.0126193
R48578 vss.n10189 vss.n2168 0.0126193
R48579 vss.t76 vss.n2168 0.0126193
R48580 vss.n10213 vss.n2180 0.0126193
R48581 vss.t76 vss.n2180 0.0126193
R48582 vss.n10201 vss.n2183 0.0126193
R48583 vss.t76 vss.n2183 0.0126193
R48584 vss.n10272 vss.n2186 0.0126193
R48585 vss.t76 vss.n2186 0.0126193
R48586 vss.n10270 vss.n2185 0.0126193
R48587 vss.t76 vss.n2185 0.0126193
R48588 vss.n10267 vss.n2167 0.0126193
R48589 vss.t76 vss.n2167 0.0126193
R48590 vss.n10291 vss.n2184 0.0126193
R48591 vss.t76 vss.n2184 0.0126193
R48592 vss.n10279 vss.n2187 0.0126193
R48593 vss.t76 vss.n2187 0.0126193
R48594 vss.n12505 vss.n2190 0.0126193
R48595 vss.t76 vss.n2190 0.0126193
R48596 vss.n12503 vss.n2189 0.0126193
R48597 vss.t76 vss.n2189 0.0126193
R48598 vss.n12500 vss.n2166 0.0126193
R48599 vss.t76 vss.n2166 0.0126193
R48600 vss.n12524 vss.n2188 0.0126193
R48601 vss.t76 vss.n2188 0.0126193
R48602 vss.n12512 vss.n2191 0.0126193
R48603 vss.t76 vss.n2191 0.0126193
R48604 vss.n12376 vss.n2194 0.0126193
R48605 vss.t76 vss.n2194 0.0126193
R48606 vss.n12374 vss.n2193 0.0126193
R48607 vss.t76 vss.n2193 0.0126193
R48608 vss.n12371 vss.n2165 0.0126193
R48609 vss.t76 vss.n2165 0.0126193
R48610 vss.n12395 vss.n2192 0.0126193
R48611 vss.t76 vss.n2192 0.0126193
R48612 vss.n12383 vss.n2195 0.0126193
R48613 vss.t76 vss.n2195 0.0126193
R48614 vss.n2213 vss.n2198 0.0126193
R48615 vss.t76 vss.n2198 0.0126193
R48616 vss.n2211 vss.n2197 0.0126193
R48617 vss.t76 vss.n2197 0.0126193
R48618 vss.n2208 vss.n2164 0.0126193
R48619 vss.t76 vss.n2164 0.0126193
R48620 vss.n2232 vss.n2196 0.0126193
R48621 vss.t76 vss.n2196 0.0126193
R48622 vss.n2220 vss.n2199 0.0126193
R48623 vss.t76 vss.n2199 0.0126193
R48624 vss.n2626 vss.n2624 0.0126193
R48625 vss.n2624 vss.t90 0.0126193
R48626 vss.n5864 vss.t90 0.0126193
R48627 vss.n5864 vss.n2627 0.0126193
R48628 vss.n5861 vss.n2629 0.0126193
R48629 vss.n5861 vss.t90 0.0126193
R48630 vss.n5873 vss.t90 0.0126193
R48631 vss.n5874 vss.n5873 0.0126193
R48632 vss.n5868 vss.n5867 0.0126193
R48633 vss.n5867 vss.t90 0.0126193
R48634 vss.n3361 vss.n3359 0.0126193
R48635 vss.n3359 vss.t90 0.0126193
R48636 vss.n5853 vss.t90 0.0126193
R48637 vss.n5854 vss.n5853 0.0126193
R48638 vss.n3380 vss.n3379 0.0126193
R48639 vss.n3379 vss.t90 0.0126193
R48640 vss.n3372 vss.t90 0.0126193
R48641 vss.n3373 vss.n3372 0.0126193
R48642 vss.n3367 vss.n3366 0.0126193
R48643 vss.n3366 vss.t90 0.0126193
R48644 vss.n3441 vss.n3440 0.0126193
R48645 vss.n3440 vss.t90 0.0126193
R48646 vss.n3446 vss.t90 0.0126193
R48647 vss.n3447 vss.n3446 0.0126193
R48648 vss.n3454 vss.n3453 0.0126193
R48649 vss.n3453 vss.t90 0.0126193
R48650 vss.n3435 vss.t90 0.0126193
R48651 vss.n3436 vss.n3435 0.0126193
R48652 vss.n3430 vss.n3429 0.0126193
R48653 vss.n3429 vss.t90 0.0126193
R48654 vss.n3963 vss.n3962 0.0126193
R48655 vss.n3962 vss.t90 0.0126193
R48656 vss.n3968 vss.t90 0.0126193
R48657 vss.n3969 vss.n3968 0.0126193
R48658 vss.n3976 vss.n3975 0.0126193
R48659 vss.n3975 vss.t90 0.0126193
R48660 vss.n3957 vss.t90 0.0126193
R48661 vss.n3958 vss.n3957 0.0126193
R48662 vss.n3952 vss.n3951 0.0126193
R48663 vss.n3951 vss.t90 0.0126193
R48664 vss.n3661 vss.n3660 0.0126193
R48665 vss.n3660 vss.t90 0.0126193
R48666 vss.n3666 vss.t90 0.0126193
R48667 vss.n3667 vss.n3666 0.0126193
R48668 vss.n3674 vss.n3673 0.0126193
R48669 vss.n3673 vss.t90 0.0126193
R48670 vss.n3655 vss.t90 0.0126193
R48671 vss.n3656 vss.n3655 0.0126193
R48672 vss.n3650 vss.n3649 0.0126193
R48673 vss.n3649 vss.t90 0.0126193
R48674 vss.n4230 vss.n4229 0.0126193
R48675 vss.n4229 vss.t90 0.0126193
R48676 vss.n4235 vss.t90 0.0126193
R48677 vss.n4236 vss.n4235 0.0126193
R48678 vss.n4243 vss.n4242 0.0126193
R48679 vss.n4242 vss.t90 0.0126193
R48680 vss.n4224 vss.t90 0.0126193
R48681 vss.n4225 vss.n4224 0.0126193
R48682 vss.n4219 vss.n4218 0.0126193
R48683 vss.n4218 vss.t90 0.0126193
R48684 vss.n4306 vss.n4305 0.0126193
R48685 vss.n4305 vss.t90 0.0126193
R48686 vss.n4311 vss.t90 0.0126193
R48687 vss.n4312 vss.n4311 0.0126193
R48688 vss.n4319 vss.n4318 0.0126193
R48689 vss.n4318 vss.t90 0.0126193
R48690 vss.n4300 vss.t90 0.0126193
R48691 vss.n4301 vss.n4300 0.0126193
R48692 vss.n4295 vss.n4294 0.0126193
R48693 vss.n4294 vss.t90 0.0126193
R48694 vss.n3326 vss.n3324 0.0126193
R48695 vss.n3324 vss.t90 0.0126193
R48696 vss.n3331 vss.t90 0.0126193
R48697 vss.n3332 vss.n3331 0.0126193
R48698 vss.n5887 vss.n5886 0.0126193
R48699 vss.n5886 vss.t90 0.0126193
R48700 vss.n3317 vss.t90 0.0126193
R48701 vss.n3318 vss.n3317 0.0126193
R48702 vss.n3321 vss.n3314 0.0126193
R48703 vss.n3314 vss.t90 0.0126193
R48704 vss.n13053 vss.n2202 0.0126193
R48705 vss.t76 vss.n13053 0.0126193
R48706 vss.n13039 vss.n2163 0.0126193
R48707 vss.t76 vss.n2163 0.0126193
R48708 vss.n13026 vss.n2162 0.0126193
R48709 vss.t76 vss.n2162 0.0126193
R48710 vss.n13030 vss.n2161 0.0126193
R48711 vss.t76 vss.n2161 0.0126193
R48712 vss.n13049 vss.n2200 0.0126193
R48713 vss.t76 vss.n2200 0.0126193
R48714 vss.n11327 vss.n11326 0.0126193
R48715 vss.t79 vss.n11327 0.0126193
R48716 vss.n11322 vss.n11053 0.0126193
R48717 vss.t79 vss.n11053 0.0126193
R48718 vss.n11307 vss.n11300 0.0126193
R48719 vss.t79 vss.n11300 0.0126193
R48720 vss.n11306 vss.n11055 0.0126193
R48721 vss.t79 vss.n11055 0.0126193
R48722 vss.n11312 vss.n11298 0.0126193
R48723 vss.t79 vss.n11298 0.0126193
R48724 vss.n11297 vss.n11296 0.0126193
R48725 vss.t79 vss.n11297 0.0126193
R48726 vss.n11272 vss.n11057 0.0126193
R48727 vss.t79 vss.n11057 0.0126193
R48728 vss.n11273 vss.n11269 0.0126193
R48729 vss.t79 vss.n11269 0.0126193
R48730 vss.n11274 vss.n11059 0.0126193
R48731 vss.t79 vss.n11059 0.0126193
R48732 vss.n11287 vss.n11267 0.0126193
R48733 vss.t79 vss.n11267 0.0126193
R48734 vss.n11266 vss.n11265 0.0126193
R48735 vss.t79 vss.n11266 0.0126193
R48736 vss.n11261 vss.n11061 0.0126193
R48737 vss.t79 vss.n11061 0.0126193
R48738 vss.n11246 vss.n11239 0.0126193
R48739 vss.t79 vss.n11239 0.0126193
R48740 vss.n11245 vss.n11063 0.0126193
R48741 vss.t79 vss.n11063 0.0126193
R48742 vss.n11251 vss.n11237 0.0126193
R48743 vss.t79 vss.n11237 0.0126193
R48744 vss.n11236 vss.n11235 0.0126193
R48745 vss.t79 vss.n11236 0.0126193
R48746 vss.n11211 vss.n11065 0.0126193
R48747 vss.t79 vss.n11065 0.0126193
R48748 vss.n11212 vss.n11208 0.0126193
R48749 vss.t79 vss.n11208 0.0126193
R48750 vss.n11213 vss.n11067 0.0126193
R48751 vss.t79 vss.n11067 0.0126193
R48752 vss.n11226 vss.n11206 0.0126193
R48753 vss.t79 vss.n11206 0.0126193
R48754 vss.n11205 vss.n11204 0.0126193
R48755 vss.t79 vss.n11205 0.0126193
R48756 vss.n11180 vss.n11069 0.0126193
R48757 vss.t79 vss.n11069 0.0126193
R48758 vss.n11181 vss.n11177 0.0126193
R48759 vss.t79 vss.n11177 0.0126193
R48760 vss.n11182 vss.n11071 0.0126193
R48761 vss.t79 vss.n11071 0.0126193
R48762 vss.n11195 vss.n11175 0.0126193
R48763 vss.t79 vss.n11175 0.0126193
R48764 vss.n11174 vss.n11173 0.0126193
R48765 vss.t79 vss.n11174 0.0126193
R48766 vss.n11170 vss.n11073 0.0126193
R48767 vss.t79 vss.n11073 0.0126193
R48768 vss.n11157 vss.n11044 0.0126193
R48769 vss.t79 vss.n11157 0.0126193
R48770 vss.n11075 vss.n11045 0.0126193
R48771 vss.t79 vss.n11075 0.0126193
R48772 vss.n11352 vss.n11351 0.0126193
R48773 vss.n11351 vss.t79 0.0126193
R48774 vss.n11155 vss.n11154 0.0126193
R48775 vss.t79 vss.n11155 0.0126193
R48776 vss.n11085 vss.n11077 0.0126193
R48777 vss.t79 vss.n11077 0.0126193
R48778 vss.n11086 vss.n11082 0.0126193
R48779 vss.t79 vss.n11082 0.0126193
R48780 vss.n11087 vss.n11079 0.0126193
R48781 vss.t79 vss.n11079 0.0126193
R48782 vss.n11100 vss.n11080 0.0126193
R48783 vss.t79 vss.n11080 0.0126193
R48784 vss.n11350 vss.n11348 0.0126193
R48785 vss.t79 vss.n11350 0.0126193
R48786 vss.n11330 vss.n11051 0.0126193
R48787 vss.t79 vss.n11051 0.0126193
R48788 vss.n11049 vss.n10458 0.0126193
R48789 vss.t79 vss.n11049 0.0126193
R48790 vss.n10457 vss.n10455 0.0126193
R48791 vss.t79 vss.n10455 0.0126193
R48792 vss.n11345 vss.n11328 0.0126193
R48793 vss.t79 vss.n11328 0.0126193
R48794 vss.n14256 vss.n14255 0.000501408
R48795 vss.n14366 vss.n14365 0.000501408
R48796 vss.n14412 vss.n14411 0.000501408
R48797 vss.n14451 vss.n14450 0.000501408
R48798 vss.n14561 vss.n14560 0.000501408
R48799 vss.n14607 vss.n14606 0.000501408
R48800 vss.n14646 vss.n14645 0.000501408
R48801 vss.n14756 vss.n14755 0.000501408
R48802 vss.n13859 vss.n13330 0.000501408
R48803 vss.n13864 vss.n13863 0.000501408
R48804 vss.n13754 vss.n13410 0.000501408
R48805 vss.n13759 vss.n13758 0.000501408
R48806 vss.n13649 vss.n13490 0.000501408
R48807 vss.n13654 vss.n13653 0.000501408
R48808 vss.n359 vss.n358 0.000501408
R48809 vss.n14247 vss.n14246 0.000501408
R48810 vss.n14146 vss.n14145 0.000501408
R48811 vss.n14142 vss.n438 0.000501408
R48812 vss.n14138 vss.n14137 0.000501408
R48813 vss.n644 vss.n643 0.000501408
R48814 vss.n1091 vss.n1090 0.000501408
R48815 vss.n1200 vss.n1199 0.000501408
R48816 vss.n1405 vss.n1398 0.000501408
R48817 vss.n1484 vss.n1483 0.000501408
R48818 vss.n1694 vss.n1693 0.000501408
R48819 vss.n13235 vss.n13234 0.000501408
R48820 vss.n1565 vss.n1564 0.000501408
R48821 vss.n13953 vss.n13952 0.000501408
R48822 vss.n14029 vss.n516 0.000501408
R48823 vss.n13992 vss.n13991 0.000501408
R48824 vss.n13990 vss.n13989 0.000501408
R48825 vss.n1738 vss.n1697 0.000501408
R48826 vss.n1802 vss.n1801 0.000501408
R48827 vss.n1842 vss.n1201 0.000501408
R48828 vss.n1906 vss.n1905 0.000501408
R48829 vss.n13289 vss.n13288 0.000501408
R48830 vss.n13291 vss.n13290 0.000501408
R48831 vss.n1981 vss.n1135 0.000501408
R48832 vss.n13200 vss.n13199 0.000501408
R48833 vss.n7498 vss.n7497 0.000501408
R48834 vss.n8974 vss.n8973 0.000501408
R48835 vss.n8478 vss.n8477 0.000501408
R48836 vss.n8474 vss.n8450 0.000501408
R48837 vss.n8864 vss.n8863 0.000501408
R48838 vss.n7587 vss.n7586 0.000501408
R48839 vss.n8855 vss.n8854 0.000501408
R48840 vss.n8380 vss.n8379 0.000501408
R48841 vss.n8376 vss.n8352 0.000501408
R48842 vss.n8745 vss.n8744 0.000501408
R48843 vss.n7730 vss.n7729 0.000501408
R48844 vss.n8736 vss.n8735 0.000501408
R48845 vss.n7906 vss.n7882 0.000501408
R48846 vss.n8259 vss.n8258 0.000501408
R48847 vss.n8253 vss.n7304 0.000501408
R48848 vss.n7951 vss.n7950 0.000501408
R48849 vss.n8245 vss.n8244 0.000501408
R48850 vss.n8104 vss.n6004 0.000501408
R48851 vss.n9642 vss.n9641 0.000501408
R48852 vss.n9637 vss.n6005 0.000501408
R48853 vss.n6051 vss.n6050 0.000501408
R48854 vss.n6366 vss.n6365 0.000501408
R48855 vss.n9252 vss.n6488 0.000501408
R48856 vss.n7029 vss.n7028 0.000501408
R48857 vss.n6980 vss.n6979 0.000501408
R48858 vss.n7089 vss.n6714 0.000501408
R48859 vss.n7220 vss.n7219 0.000501408
R48860 vss.n7169 vss.n7168 0.000501408
R48861 vss.n9502 vss.n9501 0.000501408
R48862 vss.n9578 vss.n6055 0.000501408
R48863 vss.n9541 vss.n9540 0.000501408
R48864 vss.n9539 vss.n9538 0.000501408
R48865 vss.n6774 vss.n6717 0.000501408
R48866 vss.n7084 vss.n7083 0.000501408
R48867 vss.n6883 vss.n6489 0.000501408
R48868 vss.n9247 vss.n9246 0.000501408
R48869 vss.n9129 vss.n6546 0.000501408
R48870 vss.n9145 vss.n9144 0.000501408
R48871 vss.n9192 vss.n9191 0.000501408
R48872 vss.n9368 vss.n9367 0.000501408
R48873 vss.n2925 vss.n2924 0.000501408
R48874 vss.n9844 vss.n9843 0.000501408
R48875 vss.n5331 vss.n5330 0.000501408
R48876 vss.n5327 vss.n4859 0.000501408
R48877 vss.n5322 vss.n4922 0.000501408
R48878 vss.n4964 vss.n4963 0.000501408
R48879 vss.n5314 vss.n5313 0.000501408
R48880 vss.n5269 vss.n4794 0.000501408
R48881 vss.n5268 vss.n4773 0.000501408
R48882 vss.n5263 vss.n5124 0.000501408
R48883 vss.n5166 vss.n5165 0.000501408
R48884 vss.n5255 vss.n5254 0.000501408
R48885 vss.n5210 vss.n4708 0.000501408
R48886 vss.n5209 vss.n4687 0.000501408
R48887 vss.n9794 vss.n9793 0.000501408
R48888 vss.n3147 vss.n3146 0.000501408
R48889 vss.n9785 vss.n9784 0.000501408
R48890 vss.n9740 vss.n2713 0.000501408
R48891 vss.n9739 vss.n3306 0.000501408
R48892 vss.n9735 vss.n2748 0.000501408
R48893 vss.n9990 vss.n9989 0.000501408
R48894 vss.n5723 vss.n3602 0.000501408
R48895 vss.n5739 vss.n5738 0.000501408
R48896 vss.n5786 vss.n5785 0.000501408
R48897 vss.n3423 vss.n3422 0.000501408
R48898 vss.n5844 vss.n3542 0.000501408
R48899 vss.n5839 vss.n5838 0.000501408
R48900 vss.n3926 vss.n3543 0.000501408
R48901 vss.n4119 vss.n4118 0.000501408
R48902 vss.n4020 vss.n4019 0.000501408
R48903 vss.n4069 vss.n4064 0.000501408
R48904 vss.n4172 vss.n4171 0.000501408
R48905 vss.n4174 vss.n4173 0.000501408
R48906 vss.n4211 vss.n3762 0.000501408
R48907 vss.n4287 vss.n4286 0.000501408
R48908 vss.n4411 vss.n4410 0.000501408
R48909 vss.n4610 vss.n4609 0.000501408
R48910 vss.n4546 vss.n4412 0.000501408
R48911 vss.n4503 vss.n4502 0.000501408
R48912 vss.n5931 vss.n5930 0.000501408
R48913 vss.n14090 vss.n14087 0.000501408
R48914 vss.n10013 vss.n2077 0.000501408
R48915 vss.n10010 vss.n10009 0.000501408
R48916 vss.n9729 vss.n9728 0.000501408
R48917 vss.n9682 vss.n9681 0.000501408
R48918 vss.n9631 vss.n5978 0.000501408
R48919 vss.n9628 vss.n9627 0.000501408
R48920 vss.n12320 vss.n12319 0.000501408
R48921 vss.n12365 vss.n12364 0.000501408
R48922 vss.n12535 vss.n11778 0.000501408
R48923 vss.n12450 vss.n12449 0.000501408
R48924 vss.n10261 vss.n10260 0.000501408
R48925 vss.n12901 vss.n12900 0.000501408
R48926 vss.n12909 vss.n10142 0.000501408
R48927 vss.n2441 vss.n2440 0.000501408
R48928 vss.n12953 vss.n2100 0.000501408
R48929 vss.n12952 vss.n12951 0.000501408
R48930 vss.n12966 vss.n12965 0.000501408
R48931 vss.n12957 vss.n2124 0.000501408
R48932 vss.n2266 vss.n2265 0.000501408
R48933 vss.n13018 vss.n13017 0.000501408
R48934 vss.n12144 vss.n12143 0.000501408
R48935 vss.n12140 vss.n11792 0.000501408
R48936 vss.n12540 vss.n12539 0.000501408
R48937 vss.n11736 vss.n11705 0.000501408
R48938 vss.n12856 vss.n12855 0.000501408
R48939 vss.n12822 vss.n10302 0.000501408
R48940 vss.n12076 vss.n12075 0.000501408
R48941 vss.n12074 vss.n12073 0.000501408
R48942 vss.n11967 vss.n11966 0.000501408
R48943 vss.n10502 vss.n10501 0.000501408
R48944 vss.n12615 vss.n10589 0.000501408
R48945 vss.n12610 vss.n12609 0.000501408
R48946 vss.n10658 vss.n10590 0.000501408
R48947 vss.n11593 vss.n11592 0.000501408
R48948 vss.n10723 vss.n10722 0.000501408
R48949 vss.n11544 vss.n10810 0.000501408
R48950 vss.n11539 vss.n11538 0.000501408
R48951 vss.n11500 vss.n10811 0.000501408
R48952 vss.n10992 vss.n10973 0.000501408
R48953 vss.n11037 vss.n11036 0.000501408
R48954 vss.n11446 vss.n11445 0.000501408
R48955 vss.n12741 vss.n12740 0.000501408
R48956 vss.n12739 vss.n12738 0.000501408
R48957 vss.n12696 vss.n12695 0.000501408
R48958 vss.n11146 vss.n11145 0.000501408
R48959 vss.n13148 vss.n13147 0.000501408
R48960 vss.n14793 vss.n14792 0.000501408
R48961 X2.X2.X3.vin1.n0 X2.X2.X3.vin1.t2 43.0572
R48962 X2.X2.X3.vin1.t1 X2.X2.X3.vin1.t0 28.6406
R48963 X2.X2.X3.vin1 X2.X2.X3.vin1.t3 28.5751
R48964 X2.X2.X3.vin1 X2.X2.X3.vin1.n0 26.802
R48965 X2.X2.X3.vin1.n0 X2.X2.X3.vin1 1.29627
R48966 X2.X2.X3.vin1 X2.X2.X3.vin1.t1 0.959305
R48967 d0.n0 d0.t245 40.0866
R48968 d0.n314 d0.t160 40.0866
R48969 d0.n1 d0.t135 40.0866
R48970 d0.n310 d0.t66 40.0866
R48971 d0.n3 d0.t174 40.0866
R48972 d0.n306 d0.t106 40.0866
R48973 d0.n5 d0.t216 40.0866
R48974 d0.n302 d0.t76 40.0866
R48975 d0.n7 d0.t125 40.0866
R48976 d0.n298 d0.t228 40.0866
R48977 d0.n9 d0.t165 40.0866
R48978 d0.n294 d0.t14 40.0866
R48979 d0.n11 d0.t128 40.0866
R48980 d0.n290 d0.t167 40.0866
R48981 d0.n13 d0.t15 40.0866
R48982 d0.n286 d0.t204 40.0866
R48983 d0.n283 d0.t96 40.0866
R48984 d0.n281 d0.t235 40.0866
R48985 d0.n279 d0.t54 40.0866
R48986 d0.n277 d0.t190 40.0866
R48987 d0.n275 d0.t223 40.0866
R48988 d0.n273 d0.t47 40.0866
R48989 d0.n271 d0.t197 40.0866
R48990 d0.n269 d0.t4 40.0866
R48991 d0.n267 d0.t157 40.0866
R48992 d0.n265 d0.t183 40.0866
R48993 d0.n263 d0.t251 40.0866
R48994 d0.n261 d0.t144 40.0866
R48995 d0.n259 d0.t207 40.0866
R48996 d0.n257 d0.t89 40.0866
R48997 d0.n254 d0.t188 40.0866
R48998 d0.n255 d0.t115 40.0866
R48999 d0.n247 d0.t184 40.0866
R49000 d0.n241 d0.t52 40.0866
R49001 d0.n235 d0.t88 40.0866
R49002 d0.n229 d0.t51 40.0866
R49003 d0.n223 d0.t150 40.0866
R49004 d0.n217 d0.t98 40.0866
R49005 d0.n211 d0.t59 40.0866
R49006 d0.n206 d0.t169 40.0866
R49007 d0.n208 d0.t83 40.0866
R49008 d0.n214 d0.t240 40.0866
R49009 d0.n220 d0.t22 40.0866
R49010 d0.n226 d0.t253 40.0866
R49011 d0.n232 d0.t159 40.0866
R49012 d0.n238 d0.t199 40.0866
R49013 d0.n244 d0.t72 40.0866
R49014 d0.n250 d0.t111 40.0866
R49015 d0.n203 d0.t170 40.0866
R49016 d0.n201 d0.t62 40.0866
R49017 d0.n199 d0.t130 40.0866
R49018 d0.n197 d0.t5 40.0866
R49019 d0.n195 d0.t103 40.0866
R49020 d0.n193 d0.t171 40.0866
R49021 d0.n191 d0.t64 40.0866
R49022 d0.n189 d0.t132 40.0866
R49023 d0.n187 d0.t19 40.0866
R49024 d0.n185 d0.t48 40.0866
R49025 d0.n183 d0.t116 40.0866
R49026 d0.n181 d0.t7 40.0866
R49027 d0.n179 d0.t78 40.0866
R49028 d0.n177 d0.t210 40.0866
R49029 d0.n174 d0.t55 40.0866
R49030 d0.n175 d0.t237 40.0866
R49031 d0.n167 d0.t220 40.0866
R49032 d0.n161 d0.t31 40.0866
R49033 d0.n155 d0.t68 40.0866
R49034 d0.n149 d0.t25 40.0866
R49035 d0.n143 d0.t122 40.0866
R49036 d0.n137 d0.t73 40.0866
R49037 d0.n131 d0.t35 40.0866
R49038 d0.n126 d0.t149 40.0866
R49039 d0.n128 d0.t65 40.0866
R49040 d0.n134 d0.t213 40.0866
R49041 d0.n140 d0.t255 40.0866
R49042 d0.n146 d0.t226 40.0866
R49043 d0.n152 d0.t138 40.0866
R49044 d0.n158 d0.t178 40.0866
R49045 d0.n164 d0.t120 40.0866
R49046 d0.n170 d0.t158 40.0866
R49047 d0.n123 d0.t155 40.0866
R49048 d0.n121 d0.t41 40.0866
R49049 d0.n119 d0.t113 40.0866
R49050 d0.n117 d0.t246 40.0866
R49051 d0.n115 d0.t163 40.0866
R49052 d0.n113 d0.t225 40.0866
R49053 d0.n111 d0.t121 40.0866
R49054 d0.n109 d0.t198 40.0866
R49055 d0.n107 d0.t85 40.0866
R49056 d0.n105 d0.t112 40.0866
R49057 d0.n103 d0.t185 40.0866
R49058 d0.n101 d0.t74 40.0866
R49059 d0.n99 d0.t147 40.0866
R49060 d0.n97 d0.t20 40.0866
R49061 d0.n94 d0.t117 40.0866
R49062 d0.n95 d0.t49 40.0866
R49063 d0.n87 d0.t239 40.0866
R49064 d0.n81 d0.t236 40.0866
R49065 d0.n75 d0.t18 40.0866
R49066 d0.n69 d0.t234 40.0866
R49067 d0.n63 d0.t79 40.0866
R49068 d0.n57 d0.t26 40.0866
R49069 d0.n51 d0.t243 40.0866
R49070 d0.n46 d0.t105 40.0866
R49071 d0.n48 d0.t10 40.0866
R49072 d0.n54 d0.t177 40.0866
R49073 d0.n60 d0.t211 40.0866
R49074 d0.n66 d0.t191 40.0866
R49075 d0.n72 d0.t93 40.0866
R49076 d0.n78 d0.t131 40.0866
R49077 d0.n84 d0.t134 40.0866
R49078 d0.n90 d0.t173 40.0866
R49079 d0.n44 d0.t146 40.0866
R49080 d0.n42 d0.t33 40.0866
R49081 d0.n40 d0.t107 40.0866
R49082 d0.n38 d0.t229 40.0866
R49083 d0.n36 d0.t63 40.0866
R49084 d0.n34 d0.t129 40.0866
R49085 d0.n32 d0.t17 40.0866
R49086 d0.n30 d0.t92 40.0866
R49087 d0.n28 d0.t233 40.0866
R49088 d0.n26 d0.t6 40.0866
R49089 d0.n24 d0.t77 40.0866
R49090 d0.n22 d0.t218 40.0866
R49091 d0.n20 d0.t38 40.0866
R49092 d0.n18 d0.t176 40.0866
R49093 d0.n15 d0.t9 40.0866
R49094 d0.n16 d0.t200 40.0866
R49095 d0.n93 d0.n45 26.0319
R49096 d0.n288 d0.n285 25.885
R49097 d0.n314 d0.t58 23.8528
R49098 d0.n1 d0.t28 23.8528
R49099 d0.n310 d0.t219 23.8528
R49100 d0.n3 d0.t81 23.8528
R49101 d0.n306 d0.t193 23.8528
R49102 d0.n5 d0.t119 23.8528
R49103 d0.n302 d0.t95 23.8528
R49104 d0.n7 d0.t21 23.8528
R49105 d0.n298 d0.t133 23.8528
R49106 d0.n9 d0.t238 23.8528
R49107 d0.n294 d0.t172 23.8528
R49108 d0.n11 d0.t136 23.8528
R49109 d0.n290 d0.t75 23.8528
R49110 d0.n13 d0.t186 23.8528
R49111 d0.n286 d0.t104 23.8528
R49112 d0.n283 d0.t217 23.8528
R49113 d0.n281 d0.t108 23.8528
R49114 d0.n279 d0.t175 23.8528
R49115 d0.n277 d0.t212 23.8528
R49116 d0.n275 d0.t109 23.8528
R49117 d0.n273 d0.t179 23.8528
R49118 d0.n271 d0.t69 23.8528
R49119 d0.n269 d0.t141 23.8528
R49120 d0.n267 d0.t166 23.8528
R49121 d0.n265 d0.t60 23.8528
R49122 d0.n263 d0.t126 23.8528
R49123 d0.n261 d0.t208 23.8528
R49124 d0.n259 d0.t8 23.8528
R49125 d0.n257 d0.t161 23.8528
R49126 d0.n254 d0.t254 23.8528
R49127 d0.n255 d0.t189 23.8528
R49128 d0.n247 d0.t90 23.8528
R49129 d0.n241 d0.t36 23.8528
R49130 d0.n235 d0.t164 23.8528
R49131 d0.n229 d0.t202 23.8528
R49132 d0.n223 d0.t42 23.8528
R49133 d0.n217 d0.t0 23.8528
R49134 d0.n211 d0.t205 23.8528
R49135 d0.n206 d0.t50 23.8528
R49136 d0.n208 d0.t227 23.8528
R49137 d0.n214 d0.t153 23.8528
R49138 d0.n220 d0.t114 23.8528
R49139 d0.n226 d0.t12 23.8528
R49140 d0.n232 d0.t57 23.8528
R49141 d0.n238 d0.t97 23.8528
R49142 d0.n244 d0.t230 23.8528
R49143 d0.n250 d0.t1 23.8528
R49144 d0.n203 d0.t45 23.8528
R49145 d0.n201 d0.t181 23.8528
R49146 d0.n199 d0.t248 23.8528
R49147 d0.n197 d0.t84 23.8528
R49148 d0.n195 d0.t222 23.8528
R49149 d0.n193 d0.t46 23.8528
R49150 d0.n191 d0.t196 23.8528
R49151 d0.n189 d0.t3 23.8528
R49152 d0.n187 d0.t34 23.8528
R49153 d0.n185 d0.t182 23.8528
R49154 d0.n183 d0.t250 23.8528
R49155 d0.n181 d0.t80 23.8528
R49156 d0.n179 d0.t139 23.8528
R49157 d0.n177 d0.t27 23.8528
R49158 d0.n174 d0.t123 23.8528
R49159 d0.n175 d0.t56 23.8528
R49160 d0.n167 d0.t140 23.8528
R49161 d0.n161 d0.t86 23.8528
R49162 d0.n155 d0.t145 23.8528
R49163 d0.n149 d0.t180 23.8528
R49164 d0.n143 d0.t16 23.8528
R49165 d0.n137 d0.t231 23.8528
R49166 d0.n131 d0.t187 23.8528
R49167 d0.n126 d0.t24 23.8528
R49168 d0.n128 d0.t209 23.8528
R49169 d0.n134 d0.t127 23.8528
R49170 d0.n140 d0.t91 23.8528
R49171 d0.n146 d0.t247 23.8528
R49172 d0.n152 d0.t32 23.8528
R49173 d0.n158 d0.t71 23.8528
R49174 d0.n164 d0.t29 23.8528
R49175 d0.n170 d0.t53 23.8528
R49176 d0.n123 d0.t30 23.8528
R49177 d0.n121 d0.t162 23.8528
R49178 d0.n119 d0.t224 23.8528
R49179 d0.n117 d0.t151 23.8528
R49180 d0.n115 d0.t37 23.8528
R49181 d0.n113 d0.t110 23.8528
R49182 d0.n111 d0.t252 23.8528
R49183 d0.n109 d0.t70 23.8528
R49184 d0.n107 d0.t102 23.8528
R49185 d0.n105 d0.t244 23.8528
R49186 d0.n103 d0.t61 23.8528
R49187 d0.n101 d0.t148 23.8528
R49188 d0.n99 d0.t201 23.8528
R49189 d0.n97 d0.t94 23.8528
R49190 d0.n94 d0.t192 23.8528
R49191 d0.n95 d0.t118 23.8528
R49192 d0.n87 d0.t152 23.8528
R49193 d0.n81 d0.t101 23.8528
R49194 d0.n75 d0.t99 23.8528
R49195 d0.n69 d0.t137 23.8528
R49196 d0.n63 d0.t221 23.8528
R49197 d0.n57 d0.t194 23.8528
R49198 d0.n51 d0.t142 23.8528
R49199 d0.n46 d0.t232 23.8528
R49200 d0.n48 d0.t168 23.8528
R49201 d0.n54 d0.t82 23.8528
R49202 d0.n60 d0.t44 23.8528
R49203 d0.n66 d0.t203 23.8528
R49204 d0.n72 d0.t241 23.8528
R49205 d0.n78 d0.t23 23.8528
R49206 d0.n84 d0.t40 23.8528
R49207 d0.n90 d0.t67 23.8528
R49208 d0.n44 d0.t13 23.8528
R49209 d0.n42 d0.t154 23.8528
R49210 d0.n40 d0.t214 23.8528
R49211 d0.n38 d0.t43 23.8528
R49212 d0.n36 d0.t195 23.8528
R49213 d0.n34 d0.t2 23.8528
R49214 d0.n32 d0.t156 23.8528
R49215 d0.n30 d0.t215 23.8528
R49216 d0.n28 d0.t249 23.8528
R49217 d0.n26 d0.t143 23.8528
R49218 d0.n24 d0.t206 23.8528
R49219 d0.n22 d0.t39 23.8528
R49220 d0.n20 d0.t100 23.8528
R49221 d0.n18 d0.t242 23.8528
R49222 d0.n15 d0.t87 23.8528
R49223 d0.n16 d0.t11 23.8528
R49224 d0.n0 d0.t124 23.8528
R49225 d0.n173 d0.n125 20.6255
R49226 d0.n253 d0.n205 20.6255
R49227 d0.n258 d0.n256 7.54113
R49228 d0.n262 d0.n260 7.54113
R49229 d0.n266 d0.n264 7.54113
R49230 d0.n270 d0.n268 7.54113
R49231 d0.n274 d0.n272 7.54113
R49232 d0.n278 d0.n276 7.54113
R49233 d0.n282 d0.n280 7.54113
R49234 d0.n213 d0.n210 7.54113
R49235 d0.n219 d0.n216 7.54113
R49236 d0.n225 d0.n222 7.54113
R49237 d0.n231 d0.n228 7.54113
R49238 d0.n237 d0.n234 7.54113
R49239 d0.n243 d0.n240 7.54113
R49240 d0.n249 d0.n246 7.54113
R49241 d0.n178 d0.n176 7.54113
R49242 d0.n182 d0.n180 7.54113
R49243 d0.n186 d0.n184 7.54113
R49244 d0.n190 d0.n188 7.54113
R49245 d0.n194 d0.n192 7.54113
R49246 d0.n198 d0.n196 7.54113
R49247 d0.n202 d0.n200 7.54113
R49248 d0.n133 d0.n130 7.54113
R49249 d0.n139 d0.n136 7.54113
R49250 d0.n145 d0.n142 7.54113
R49251 d0.n151 d0.n148 7.54113
R49252 d0.n157 d0.n154 7.54113
R49253 d0.n163 d0.n160 7.54113
R49254 d0.n169 d0.n166 7.54113
R49255 d0.n98 d0.n96 7.54113
R49256 d0.n102 d0.n100 7.54113
R49257 d0.n106 d0.n104 7.54113
R49258 d0.n110 d0.n108 7.54113
R49259 d0.n114 d0.n112 7.54113
R49260 d0.n118 d0.n116 7.54113
R49261 d0.n122 d0.n120 7.54113
R49262 d0.n53 d0.n50 7.54113
R49263 d0.n59 d0.n56 7.54113
R49264 d0.n65 d0.n62 7.54113
R49265 d0.n71 d0.n68 7.54113
R49266 d0.n77 d0.n74 7.54113
R49267 d0.n83 d0.n80 7.54113
R49268 d0.n89 d0.n86 7.54113
R49269 d0.n19 d0.n17 7.54113
R49270 d0.n23 d0.n21 7.54113
R49271 d0.n27 d0.n25 7.54113
R49272 d0.n31 d0.n29 7.54113
R49273 d0.n35 d0.n33 7.54113
R49274 d0.n39 d0.n37 7.54113
R49275 d0.n43 d0.n41 7.54113
R49276 d0.n292 d0.n289 7.54113
R49277 d0.n296 d0.n293 7.54113
R49278 d0.n300 d0.n297 7.54113
R49279 d0.n304 d0.n301 7.54113
R49280 d0.n308 d0.n305 7.54113
R49281 d0.n312 d0.n309 7.54113
R49282 d0.n316 d0.n313 7.54113
R49283 d0.n285 d0.n284 5.40687
R49284 d0.n205 d0.n204 5.40687
R49285 d0.n125 d0.n124 5.40687
R49286 d0.n253 d0.n252 5.25999
R49287 d0.n173 d0.n172 5.25999
R49288 d0.n93 d0.n92 5.25999
R49289 d0.n256 d0 2.97874
R49290 d0.n176 d0 2.97874
R49291 d0.n96 d0 2.97874
R49292 d0.n17 d0 2.97874
R49293 d0.n210 d0.n207 2.91624
R49294 d0.n130 d0.n127 2.91624
R49295 d0.n50 d0.n47 2.91624
R49296 d0.n317 d0.n316 2.91624
R49297 d0.n260 d0.n258 2.91613
R49298 d0.n264 d0.n262 2.91613
R49299 d0.n268 d0.n266 2.91613
R49300 d0.n272 d0.n270 2.91613
R49301 d0.n276 d0.n274 2.91613
R49302 d0.n280 d0.n278 2.91613
R49303 d0.n284 d0.n282 2.91613
R49304 d0.n216 d0.n213 2.91613
R49305 d0.n222 d0.n219 2.91613
R49306 d0.n228 d0.n225 2.91613
R49307 d0.n234 d0.n231 2.91613
R49308 d0.n240 d0.n237 2.91613
R49309 d0.n246 d0.n243 2.91613
R49310 d0.n252 d0.n249 2.91613
R49311 d0.n180 d0.n178 2.91613
R49312 d0.n184 d0.n182 2.91613
R49313 d0.n188 d0.n186 2.91613
R49314 d0.n192 d0.n190 2.91613
R49315 d0.n196 d0.n194 2.91613
R49316 d0.n200 d0.n198 2.91613
R49317 d0.n204 d0.n202 2.91613
R49318 d0.n136 d0.n133 2.91613
R49319 d0.n142 d0.n139 2.91613
R49320 d0.n148 d0.n145 2.91613
R49321 d0.n154 d0.n151 2.91613
R49322 d0.n160 d0.n157 2.91613
R49323 d0.n166 d0.n163 2.91613
R49324 d0.n172 d0.n169 2.91613
R49325 d0.n100 d0.n98 2.91613
R49326 d0.n104 d0.n102 2.91613
R49327 d0.n108 d0.n106 2.91613
R49328 d0.n112 d0.n110 2.91613
R49329 d0.n116 d0.n114 2.91613
R49330 d0.n120 d0.n118 2.91613
R49331 d0.n124 d0.n122 2.91613
R49332 d0.n56 d0.n53 2.91613
R49333 d0.n62 d0.n59 2.91613
R49334 d0.n68 d0.n65 2.91613
R49335 d0.n74 d0.n71 2.91613
R49336 d0.n80 d0.n77 2.91613
R49337 d0.n86 d0.n83 2.91613
R49338 d0.n92 d0.n89 2.91613
R49339 d0.n21 d0.n19 2.91613
R49340 d0.n25 d0.n23 2.91613
R49341 d0.n29 d0.n27 2.91613
R49342 d0.n33 d0.n31 2.91613
R49343 d0.n37 d0.n35 2.91613
R49344 d0.n41 d0.n39 2.91613
R49345 d0.n45 d0.n43 2.91613
R49346 d0.n289 d0.n288 2.91613
R49347 d0.n293 d0.n292 2.91613
R49348 d0.n297 d0.n296 2.91613
R49349 d0.n301 d0.n300 2.91613
R49350 d0.n305 d0.n304 2.91613
R49351 d0.n309 d0.n308 2.91613
R49352 d0.n313 d0.n312 2.91613
R49353 d0.n125 d0.n93 2.2505
R49354 d0.n205 d0.n173 2.2505
R49355 d0.n285 d0.n253 2.2505
R49356 d0.n315 d0.n314 0.2505
R49357 d0.n2 d0.n1 0.2505
R49358 d0.n311 d0.n310 0.2505
R49359 d0.n4 d0.n3 0.2505
R49360 d0.n307 d0.n306 0.2505
R49361 d0.n6 d0.n5 0.2505
R49362 d0.n303 d0.n302 0.2505
R49363 d0.n8 d0.n7 0.2505
R49364 d0.n299 d0.n298 0.2505
R49365 d0.n10 d0.n9 0.2505
R49366 d0.n295 d0.n294 0.2505
R49367 d0.n12 d0.n11 0.2505
R49368 d0.n291 d0.n290 0.2505
R49369 d0.n14 d0.n13 0.2505
R49370 d0.n287 d0.n286 0.2505
R49371 d0 d0.n279 0.2505
R49372 d0 d0.n277 0.2505
R49373 d0 d0.n275 0.2505
R49374 d0 d0.n271 0.2505
R49375 d0 d0.n269 0.2505
R49376 d0 d0.n267 0.2505
R49377 d0 d0.n263 0.2505
R49378 d0 d0.n261 0.2505
R49379 d0 d0.n259 0.2505
R49380 d0 d0.n254 0.2505
R49381 d0 d0.n255 0.2505
R49382 d0.n248 d0.n247 0.2505
R49383 d0.n242 d0.n241 0.2505
R49384 d0.n236 d0.n235 0.2505
R49385 d0.n230 d0.n229 0.2505
R49386 d0.n224 d0.n223 0.2505
R49387 d0.n218 d0.n217 0.2505
R49388 d0.n212 d0.n211 0.2505
R49389 d0.n207 d0.n206 0.2505
R49390 d0.n209 d0.n208 0.2505
R49391 d0.n215 d0.n214 0.2505
R49392 d0.n221 d0.n220 0.2505
R49393 d0.n227 d0.n226 0.2505
R49394 d0.n233 d0.n232 0.2505
R49395 d0.n239 d0.n238 0.2505
R49396 d0.n245 d0.n244 0.2505
R49397 d0.n251 d0.n250 0.2505
R49398 d0 d0.n199 0.2505
R49399 d0 d0.n197 0.2505
R49400 d0 d0.n195 0.2505
R49401 d0 d0.n191 0.2505
R49402 d0 d0.n189 0.2505
R49403 d0 d0.n187 0.2505
R49404 d0 d0.n183 0.2505
R49405 d0 d0.n181 0.2505
R49406 d0 d0.n179 0.2505
R49407 d0 d0.n174 0.2505
R49408 d0 d0.n175 0.2505
R49409 d0.n168 d0.n167 0.2505
R49410 d0.n162 d0.n161 0.2505
R49411 d0.n156 d0.n155 0.2505
R49412 d0.n150 d0.n149 0.2505
R49413 d0.n144 d0.n143 0.2505
R49414 d0.n138 d0.n137 0.2505
R49415 d0.n132 d0.n131 0.2505
R49416 d0.n127 d0.n126 0.2505
R49417 d0.n129 d0.n128 0.2505
R49418 d0.n135 d0.n134 0.2505
R49419 d0.n141 d0.n140 0.2505
R49420 d0.n147 d0.n146 0.2505
R49421 d0.n153 d0.n152 0.2505
R49422 d0.n159 d0.n158 0.2505
R49423 d0.n165 d0.n164 0.2505
R49424 d0.n171 d0.n170 0.2505
R49425 d0 d0.n119 0.2505
R49426 d0 d0.n117 0.2505
R49427 d0 d0.n115 0.2505
R49428 d0 d0.n111 0.2505
R49429 d0 d0.n109 0.2505
R49430 d0 d0.n107 0.2505
R49431 d0 d0.n103 0.2505
R49432 d0 d0.n101 0.2505
R49433 d0 d0.n99 0.2505
R49434 d0 d0.n94 0.2505
R49435 d0 d0.n95 0.2505
R49436 d0.n88 d0.n87 0.2505
R49437 d0.n82 d0.n81 0.2505
R49438 d0.n76 d0.n75 0.2505
R49439 d0.n70 d0.n69 0.2505
R49440 d0.n64 d0.n63 0.2505
R49441 d0.n58 d0.n57 0.2505
R49442 d0.n52 d0.n51 0.2505
R49443 d0.n47 d0.n46 0.2505
R49444 d0.n49 d0.n48 0.2505
R49445 d0.n55 d0.n54 0.2505
R49446 d0.n61 d0.n60 0.2505
R49447 d0.n67 d0.n66 0.2505
R49448 d0.n73 d0.n72 0.2505
R49449 d0.n79 d0.n78 0.2505
R49450 d0.n85 d0.n84 0.2505
R49451 d0.n91 d0.n90 0.2505
R49452 d0 d0.n40 0.2505
R49453 d0 d0.n38 0.2505
R49454 d0 d0.n36 0.2505
R49455 d0 d0.n32 0.2505
R49456 d0 d0.n30 0.2505
R49457 d0 d0.n28 0.2505
R49458 d0 d0.n24 0.2505
R49459 d0 d0.n22 0.2505
R49460 d0 d0.n20 0.2505
R49461 d0 d0.n15 0.2505
R49462 d0 d0.n16 0.2505
R49463 d0.n317 d0.n0 0.2505
R49464 d0 d0.n283 0.188
R49465 d0 d0.n281 0.188
R49466 d0 d0.n273 0.188
R49467 d0 d0.n265 0.188
R49468 d0 d0.n257 0.188
R49469 d0 d0.n203 0.188
R49470 d0 d0.n201 0.188
R49471 d0 d0.n193 0.188
R49472 d0 d0.n185 0.188
R49473 d0 d0.n177 0.188
R49474 d0 d0.n123 0.188
R49475 d0 d0.n121 0.188
R49476 d0 d0.n113 0.188
R49477 d0 d0.n105 0.188
R49478 d0 d0.n97 0.188
R49479 d0 d0.n44 0.188
R49480 d0 d0.n42 0.188
R49481 d0 d0.n34 0.188
R49482 d0 d0.n26 0.188
R49483 d0 d0.n18 0.188
R49484 d0.n315 d0 0.063
R49485 d0.n2 d0 0.063
R49486 d0.n311 d0 0.063
R49487 d0.n4 d0 0.063
R49488 d0.n307 d0 0.063
R49489 d0.n6 d0 0.063
R49490 d0.n303 d0 0.063
R49491 d0.n8 d0 0.063
R49492 d0.n299 d0 0.063
R49493 d0.n10 d0 0.063
R49494 d0.n295 d0 0.063
R49495 d0.n12 d0 0.063
R49496 d0.n291 d0 0.063
R49497 d0.n14 d0 0.063
R49498 d0.n287 d0 0.063
R49499 d0.n248 d0 0.063
R49500 d0.n242 d0 0.063
R49501 d0.n236 d0 0.063
R49502 d0.n230 d0 0.063
R49503 d0.n224 d0 0.063
R49504 d0.n218 d0 0.063
R49505 d0.n212 d0 0.063
R49506 d0.n207 d0 0.063
R49507 d0.n209 d0 0.063
R49508 d0.n215 d0 0.063
R49509 d0.n221 d0 0.063
R49510 d0.n227 d0 0.063
R49511 d0.n233 d0 0.063
R49512 d0.n239 d0 0.063
R49513 d0.n245 d0 0.063
R49514 d0.n251 d0 0.063
R49515 d0.n168 d0 0.063
R49516 d0.n162 d0 0.063
R49517 d0.n156 d0 0.063
R49518 d0.n150 d0 0.063
R49519 d0.n144 d0 0.063
R49520 d0.n138 d0 0.063
R49521 d0.n132 d0 0.063
R49522 d0.n129 d0 0.063
R49523 d0.n135 d0 0.063
R49524 d0.n141 d0 0.063
R49525 d0.n147 d0 0.063
R49526 d0.n153 d0 0.063
R49527 d0.n159 d0 0.063
R49528 d0.n165 d0 0.063
R49529 d0.n171 d0 0.063
R49530 d0.n88 d0 0.063
R49531 d0.n82 d0 0.063
R49532 d0.n76 d0 0.063
R49533 d0.n70 d0 0.063
R49534 d0.n64 d0 0.063
R49535 d0.n58 d0 0.063
R49536 d0.n52 d0 0.063
R49537 d0.n47 d0 0.063
R49538 d0.n49 d0 0.063
R49539 d0.n55 d0 0.063
R49540 d0.n61 d0 0.063
R49541 d0.n67 d0 0.063
R49542 d0.n73 d0 0.063
R49543 d0.n79 d0 0.063
R49544 d0.n85 d0 0.063
R49545 d0.n91 d0 0.063
R49546 d0.n127 d0 0.03175
R49547 d0 d0.n317 0.03175
R49548 d0.n256 d0 0.000617139
R49549 d0.n258 d0 0.000617139
R49550 d0.n260 d0 0.000617139
R49551 d0.n262 d0 0.000617139
R49552 d0.n264 d0 0.000617139
R49553 d0.n266 d0 0.000617139
R49554 d0.n268 d0 0.000617139
R49555 d0.n270 d0 0.000617139
R49556 d0.n272 d0 0.000617139
R49557 d0.n274 d0 0.000617139
R49558 d0.n276 d0 0.000617139
R49559 d0.n278 d0 0.000617139
R49560 d0.n280 d0 0.000617139
R49561 d0.n282 d0 0.000617139
R49562 d0.n284 d0 0.000617139
R49563 d0.n210 d0.n209 0.000617139
R49564 d0.n213 d0.n212 0.000617139
R49565 d0.n216 d0.n215 0.000617139
R49566 d0.n219 d0.n218 0.000617139
R49567 d0.n222 d0.n221 0.000617139
R49568 d0.n225 d0.n224 0.000617139
R49569 d0.n228 d0.n227 0.000617139
R49570 d0.n231 d0.n230 0.000617139
R49571 d0.n234 d0.n233 0.000617139
R49572 d0.n237 d0.n236 0.000617139
R49573 d0.n240 d0.n239 0.000617139
R49574 d0.n243 d0.n242 0.000617139
R49575 d0.n246 d0.n245 0.000617139
R49576 d0.n249 d0.n248 0.000617139
R49577 d0.n252 d0.n251 0.000617139
R49578 d0.n176 d0 0.000617139
R49579 d0.n178 d0 0.000617139
R49580 d0.n180 d0 0.000617139
R49581 d0.n182 d0 0.000617139
R49582 d0.n184 d0 0.000617139
R49583 d0.n186 d0 0.000617139
R49584 d0.n188 d0 0.000617139
R49585 d0.n190 d0 0.000617139
R49586 d0.n192 d0 0.000617139
R49587 d0.n194 d0 0.000617139
R49588 d0.n196 d0 0.000617139
R49589 d0.n198 d0 0.000617139
R49590 d0.n200 d0 0.000617139
R49591 d0.n202 d0 0.000617139
R49592 d0.n204 d0 0.000617139
R49593 d0.n130 d0.n129 0.000617139
R49594 d0.n133 d0.n132 0.000617139
R49595 d0.n136 d0.n135 0.000617139
R49596 d0.n139 d0.n138 0.000617139
R49597 d0.n142 d0.n141 0.000617139
R49598 d0.n145 d0.n144 0.000617139
R49599 d0.n148 d0.n147 0.000617139
R49600 d0.n151 d0.n150 0.000617139
R49601 d0.n154 d0.n153 0.000617139
R49602 d0.n157 d0.n156 0.000617139
R49603 d0.n160 d0.n159 0.000617139
R49604 d0.n163 d0.n162 0.000617139
R49605 d0.n166 d0.n165 0.000617139
R49606 d0.n169 d0.n168 0.000617139
R49607 d0.n172 d0.n171 0.000617139
R49608 d0.n96 d0 0.000617139
R49609 d0.n98 d0 0.000617139
R49610 d0.n100 d0 0.000617139
R49611 d0.n102 d0 0.000617139
R49612 d0.n104 d0 0.000617139
R49613 d0.n106 d0 0.000617139
R49614 d0.n108 d0 0.000617139
R49615 d0.n110 d0 0.000617139
R49616 d0.n112 d0 0.000617139
R49617 d0.n114 d0 0.000617139
R49618 d0.n116 d0 0.000617139
R49619 d0.n118 d0 0.000617139
R49620 d0.n120 d0 0.000617139
R49621 d0.n122 d0 0.000617139
R49622 d0.n124 d0 0.000617139
R49623 d0.n50 d0.n49 0.000617139
R49624 d0.n53 d0.n52 0.000617139
R49625 d0.n56 d0.n55 0.000617139
R49626 d0.n59 d0.n58 0.000617139
R49627 d0.n62 d0.n61 0.000617139
R49628 d0.n65 d0.n64 0.000617139
R49629 d0.n68 d0.n67 0.000617139
R49630 d0.n71 d0.n70 0.000617139
R49631 d0.n74 d0.n73 0.000617139
R49632 d0.n77 d0.n76 0.000617139
R49633 d0.n80 d0.n79 0.000617139
R49634 d0.n83 d0.n82 0.000617139
R49635 d0.n86 d0.n85 0.000617139
R49636 d0.n89 d0.n88 0.000617139
R49637 d0.n92 d0.n91 0.000617139
R49638 d0.n17 d0 0.000617139
R49639 d0.n19 d0 0.000617139
R49640 d0.n21 d0 0.000617139
R49641 d0.n23 d0 0.000617139
R49642 d0.n25 d0 0.000617139
R49643 d0.n27 d0 0.000617139
R49644 d0.n29 d0 0.000617139
R49645 d0.n31 d0 0.000617139
R49646 d0.n33 d0 0.000617139
R49647 d0.n35 d0 0.000617139
R49648 d0.n37 d0 0.000617139
R49649 d0.n39 d0 0.000617139
R49650 d0.n41 d0 0.000617139
R49651 d0.n43 d0 0.000617139
R49652 d0.n45 d0 0.000617139
R49653 d0.n288 d0.n287 0.000617139
R49654 d0.n289 d0.n14 0.000617139
R49655 d0.n292 d0.n291 0.000617139
R49656 d0.n293 d0.n12 0.000617139
R49657 d0.n296 d0.n295 0.000617139
R49658 d0.n297 d0.n10 0.000617139
R49659 d0.n300 d0.n299 0.000617139
R49660 d0.n301 d0.n8 0.000617139
R49661 d0.n304 d0.n303 0.000617139
R49662 d0.n305 d0.n6 0.000617139
R49663 d0.n308 d0.n307 0.000617139
R49664 d0.n309 d0.n4 0.000617139
R49665 d0.n312 d0.n311 0.000617139
R49666 d0.n313 d0.n2 0.000617139
R49667 d0.n316 d0.n315 0.000617139
R49668 d1.n1 d1.t44 40.0866
R49669 d1.n13 d1.t11 40.0866
R49670 d1.n11 d1.t120 40.0866
R49671 d1.n109 d1.t62 40.0866
R49672 d1.n110 d1.t10 40.0866
R49673 d1.n112 d1.t37 40.0866
R49674 d1.n114 d1.t59 40.0866
R49675 d1.n116 d1.t100 40.0866
R49676 d1.n118 d1.t117 40.0866
R49677 d1.n120 d1.t93 40.0866
R49678 d1.n122 d1.t118 40.0866
R49679 d1.n124 d1.t4 40.0866
R49680 d1.n126 d1.t86 40.0866
R49681 d1.n129 d1.t109 40.0866
R49682 d1.n132 d1.t94 40.0866
R49683 d1.n135 d1.t43 40.0866
R49684 d1.n138 d1.t66 40.0866
R49685 d1.n141 d1.t71 40.0866
R49686 d1.n144 d1.t92 40.0866
R49687 d1.n69 d1.t52 40.0866
R49688 d1.n70 d1.t1 40.0866
R49689 d1.n72 d1.t23 40.0866
R49690 d1.n74 d1.t47 40.0866
R49691 d1.n76 d1.t91 40.0866
R49692 d1.n78 d1.t111 40.0866
R49693 d1.n80 d1.t58 40.0866
R49694 d1.n82 d1.t82 40.0866
R49695 d1.n84 d1.t126 40.0866
R49696 d1.n86 d1.t73 40.0866
R49697 d1.n89 d1.t95 40.0866
R49698 d1.n92 d1.t83 40.0866
R49699 d1.n95 d1.t30 40.0866
R49700 d1.n98 d1.t56 40.0866
R49701 d1.n101 d1.t98 40.0866
R49702 d1.n104 d1.t116 40.0866
R49703 d1.n30 d1.t40 40.0866
R49704 d1.n31 d1.t119 40.0866
R49705 d1.n33 d1.t18 40.0866
R49706 d1.n35 d1.t36 40.0866
R49707 d1.n37 d1.t76 40.0866
R49708 d1.n39 d1.t99 40.0866
R49709 d1.n41 d1.t80 40.0866
R49710 d1.n43 d1.t108 40.0866
R49711 d1.n45 d1.t103 40.0866
R49712 d1.n47 d1.t54 40.0866
R49713 d1.n50 d1.t69 40.0866
R49714 d1.n53 d1.t61 40.0866
R49715 d1.n56 d1.t9 40.0866
R49716 d1.n59 d1.t27 40.0866
R49717 d1.n62 d1.t105 40.0866
R49718 d1.n65 d1.t124 40.0866
R49719 d1.n15 d1.t102 40.0866
R49720 d1.n16 d1.t53 40.0866
R49721 d1.n18 d1.t77 40.0866
R49722 d1.n20 d1.t101 40.0866
R49723 d1.n22 d1.t8 40.0866
R49724 d1.n24 d1.t26 40.0866
R49725 d1.n26 d1.t79 40.0866
R49726 d1.n28 d1.t107 40.0866
R49727 d1.n9 d1.t104 40.0866
R49728 d1.n7 d1.t85 40.0866
R49729 d1.n5 d1.t2 40.0866
R49730 d1.n3 d1.t15 40.0866
R49731 d1.n0 d1.t127 40.0866
R49732 d1.n108 d1.n68 25.9475
R49733 d1.n149 d1.n148 25.9475
R49734 d1.n13 d1.t87 23.8528
R49735 d1.n11 d1.t72 23.8528
R49736 d1.n109 d1.t96 23.8528
R49737 d1.n110 d1.t45 23.8528
R49738 d1.n112 d1.t70 23.8528
R49739 d1.n114 d1.t125 23.8528
R49740 d1.n116 d1.t32 23.8528
R49741 d1.n118 d1.t57 23.8528
R49742 d1.n120 d1.t28 23.8528
R49743 d1.n122 d1.t50 23.8528
R49744 d1.n124 d1.t84 23.8528
R49745 d1.n126 d1.t41 23.8528
R49746 d1.n129 d1.t19 23.8528
R49747 d1.n132 d1.t42 23.8528
R49748 d1.n135 d1.t121 23.8528
R49749 d1.n138 d1.t12 23.8528
R49750 d1.n141 d1.t21 23.8528
R49751 d1.n144 d1.t39 23.8528
R49752 d1.n69 d1.t89 23.8528
R49753 d1.n70 d1.t38 23.8528
R49754 d1.n72 d1.t65 23.8528
R49755 d1.n74 d1.t114 23.8528
R49756 d1.n76 d1.t22 23.8528
R49757 d1.n78 d1.t46 23.8528
R49758 d1.n80 d1.t123 23.8528
R49759 d1.n82 d1.t13 23.8528
R49760 d1.n84 d1.t68 23.8528
R49761 d1.n86 d1.t24 23.8528
R49762 d1.n89 d1.t7 23.8528
R49763 d1.n92 d1.t25 23.8528
R49764 d1.n95 d1.t112 23.8528
R49765 d1.n98 d1.t0 23.8528
R49766 d1.n101 d1.t51 23.8528
R49767 d1.n104 d1.t64 23.8528
R49768 d1.n30 d1.t74 23.8528
R49769 d1.n31 d1.t20 23.8528
R49770 d1.n33 d1.t55 23.8528
R49771 d1.n35 d1.t106 23.8528
R49772 d1.n37 d1.t14 23.8528
R49773 d1.n39 d1.t31 23.8528
R49774 d1.n41 d1.t17 23.8528
R49775 d1.n43 d1.t35 23.8528
R49776 d1.n45 d1.t48 23.8528
R49777 d1.n47 d1.t3 23.8528
R49778 d1.n50 d1.t115 23.8528
R49779 d1.n53 d1.t5 23.8528
R49780 d1.n56 d1.t88 23.8528
R49781 d1.n59 d1.t110 23.8528
R49782 d1.n62 d1.t60 23.8528
R49783 d1.n65 d1.t67 23.8528
R49784 d1.n15 d1.t6 23.8528
R49785 d1.n16 d1.t90 23.8528
R49786 d1.n18 d1.t113 23.8528
R49787 d1.n20 d1.t33 23.8528
R49788 d1.n22 d1.t75 23.8528
R49789 d1.n24 d1.t97 23.8528
R49790 d1.n26 d1.t16 23.8528
R49791 d1.n28 d1.t34 23.8528
R49792 d1.n9 d1.t49 23.8528
R49793 d1.n7 d1.t29 23.8528
R49794 d1.n5 d1.t81 23.8528
R49795 d1.n3 d1.t63 23.8528
R49796 d1.n0 d1.t78 23.8528
R49797 d1.n1 d1.t122 23.8528
R49798 d1.n148 d1.n108 22.8755
R49799 d1.n147 d1.n146 10.6976
R49800 d1.n107 d1.n106 10.6976
R49801 d1.n68 d1.n67 10.6976
R49802 d1.n150 d1.n149 10.6976
R49803 d1.n111 d1 5.95687
R49804 d1.n128 d1.n125 5.95687
R49805 d1.n71 d1 5.95687
R49806 d1.n88 d1.n85 5.95687
R49807 d1.n32 d1 5.95687
R49808 d1.n49 d1.n46 5.95687
R49809 d1.n17 d1 5.95687
R49810 d1.n156 d1.n2 5.95687
R49811 d1.n115 d1.n113 5.95675
R49812 d1.n117 d1.n115 5.95675
R49813 d1.n119 d1.n117 5.95675
R49814 d1.n134 d1.n131 5.95675
R49815 d1.n137 d1.n134 5.95675
R49816 d1.n140 d1.n137 5.95675
R49817 d1.n146 d1.n143 5.95675
R49818 d1.n123 d1.n121 5.95675
R49819 d1.n75 d1.n73 5.95675
R49820 d1.n77 d1.n75 5.95675
R49821 d1.n79 d1.n77 5.95675
R49822 d1.n94 d1.n91 5.95675
R49823 d1.n97 d1.n94 5.95675
R49824 d1.n100 d1.n97 5.95675
R49825 d1.n106 d1.n103 5.95675
R49826 d1.n83 d1.n81 5.95675
R49827 d1.n36 d1.n34 5.95675
R49828 d1.n38 d1.n36 5.95675
R49829 d1.n40 d1.n38 5.95675
R49830 d1.n55 d1.n52 5.95675
R49831 d1.n58 d1.n55 5.95675
R49832 d1.n61 d1.n58 5.95675
R49833 d1.n67 d1.n64 5.95675
R49834 d1.n44 d1.n42 5.95675
R49835 d1.n21 d1.n19 5.95675
R49836 d1.n23 d1.n21 5.95675
R49837 d1.n25 d1.n23 5.95675
R49838 d1.n29 d1.n27 5.95675
R49839 d1.n151 d1.n150 5.95675
R49840 d1.n155 d1.n154 5.95675
R49841 d1.n154 d1.n153 5.95675
R49842 d1.n153 d1.n152 5.95675
R49843 d1.n113 d1.n111 5.36034
R49844 d1.n121 d1.n119 5.36034
R49845 d1.n73 d1.n71 5.36034
R49846 d1.n81 d1.n79 5.36034
R49847 d1.n34 d1.n32 5.36034
R49848 d1.n42 d1.n40 5.36034
R49849 d1.n19 d1.n17 5.36034
R49850 d1.n27 d1.n25 5.36034
R49851 d1.n152 d1.n151 5.36034
R49852 d1.n156 d1.n155 5.36034
R49853 d1.n131 d1.n128 5.36034
R49854 d1.n143 d1.n140 5.36034
R49855 d1.n91 d1.n88 5.36034
R49856 d1.n103 d1.n100 5.36034
R49857 d1.n52 d1.n49 5.36034
R49858 d1.n64 d1.n61 5.36034
R49859 d1.n148 d1.n147 3.07249
R49860 d1.n108 d1.n107 3.07249
R49861 d1.n147 d1.n123 1.82237
R49862 d1.n107 d1.n83 1.82237
R49863 d1.n68 d1.n44 1.82237
R49864 d1.n149 d1.n29 1.82237
R49865 d1.n14 d1.n13 0.2505
R49866 d1.n12 d1.n11 0.2505
R49867 d1 d1.n109 0.2505
R49868 d1 d1.n112 0.2505
R49869 d1 d1.n116 0.2505
R49870 d1 d1.n120 0.2505
R49871 d1.n125 d1.n124 0.2505
R49872 d1.n127 d1.n126 0.2505
R49873 d1.n130 d1.n129 0.2505
R49874 d1.n133 d1.n132 0.2505
R49875 d1.n136 d1.n135 0.2505
R49876 d1.n139 d1.n138 0.2505
R49877 d1.n142 d1.n141 0.2505
R49878 d1.n145 d1.n144 0.2505
R49879 d1 d1.n69 0.2505
R49880 d1 d1.n72 0.2505
R49881 d1 d1.n76 0.2505
R49882 d1 d1.n80 0.2505
R49883 d1.n85 d1.n84 0.2505
R49884 d1.n87 d1.n86 0.2505
R49885 d1.n90 d1.n89 0.2505
R49886 d1.n93 d1.n92 0.2505
R49887 d1.n96 d1.n95 0.2505
R49888 d1.n99 d1.n98 0.2505
R49889 d1.n102 d1.n101 0.2505
R49890 d1.n105 d1.n104 0.2505
R49891 d1 d1.n30 0.2505
R49892 d1 d1.n33 0.2505
R49893 d1 d1.n37 0.2505
R49894 d1 d1.n41 0.2505
R49895 d1.n46 d1.n45 0.2505
R49896 d1.n48 d1.n47 0.2505
R49897 d1.n51 d1.n50 0.2505
R49898 d1.n54 d1.n53 0.2505
R49899 d1.n57 d1.n56 0.2505
R49900 d1.n60 d1.n59 0.2505
R49901 d1.n63 d1.n62 0.2505
R49902 d1.n66 d1.n65 0.2505
R49903 d1 d1.n15 0.2505
R49904 d1 d1.n18 0.2505
R49905 d1 d1.n22 0.2505
R49906 d1 d1.n26 0.2505
R49907 d1.n10 d1.n9 0.2505
R49908 d1.n8 d1.n7 0.2505
R49909 d1.n6 d1.n5 0.2505
R49910 d1.n4 d1.n3 0.2505
R49911 d1.n157 d1.n0 0.2505
R49912 d1.n2 d1.n1 0.2505
R49913 d1 d1.n110 0.188
R49914 d1 d1.n114 0.188
R49915 d1 d1.n118 0.188
R49916 d1 d1.n122 0.188
R49917 d1 d1.n70 0.188
R49918 d1 d1.n74 0.188
R49919 d1 d1.n78 0.188
R49920 d1 d1.n82 0.188
R49921 d1 d1.n31 0.188
R49922 d1 d1.n35 0.188
R49923 d1 d1.n39 0.188
R49924 d1 d1.n43 0.188
R49925 d1 d1.n16 0.188
R49926 d1 d1.n20 0.188
R49927 d1 d1.n24 0.188
R49928 d1 d1.n28 0.188
R49929 d1.n14 d1 0.063
R49930 d1.n12 d1 0.063
R49931 d1.n125 d1 0.063
R49932 d1.n127 d1 0.063
R49933 d1.n130 d1 0.063
R49934 d1.n133 d1 0.063
R49935 d1.n136 d1 0.063
R49936 d1.n139 d1 0.063
R49937 d1.n142 d1 0.063
R49938 d1.n145 d1 0.063
R49939 d1.n85 d1 0.063
R49940 d1.n87 d1 0.063
R49941 d1.n90 d1 0.063
R49942 d1.n93 d1 0.063
R49943 d1.n96 d1 0.063
R49944 d1.n99 d1 0.063
R49945 d1.n102 d1 0.063
R49946 d1.n105 d1 0.063
R49947 d1.n46 d1 0.063
R49948 d1.n48 d1 0.063
R49949 d1.n51 d1 0.063
R49950 d1.n54 d1 0.063
R49951 d1.n57 d1 0.063
R49952 d1.n60 d1 0.063
R49953 d1.n63 d1 0.063
R49954 d1.n66 d1 0.063
R49955 d1.n10 d1 0.063
R49956 d1.n8 d1 0.063
R49957 d1.n6 d1 0.063
R49958 d1.n4 d1 0.063
R49959 d1 d1.n157 0.063
R49960 d1.n2 d1 0.063
R49961 d1.n111 d1 0.000617139
R49962 d1.n119 d1 0.000617139
R49963 d1.n117 d1 0.000617139
R49964 d1.n115 d1 0.000617139
R49965 d1.n113 d1 0.000617139
R49966 d1.n128 d1.n127 0.000617139
R49967 d1.n140 d1.n139 0.000617139
R49968 d1.n137 d1.n136 0.000617139
R49969 d1.n134 d1.n133 0.000617139
R49970 d1.n131 d1.n130 0.000617139
R49971 d1.n146 d1.n145 0.000617139
R49972 d1.n143 d1.n142 0.000617139
R49973 d1.n123 d1 0.000617139
R49974 d1.n121 d1 0.000617139
R49975 d1.n71 d1 0.000617139
R49976 d1.n79 d1 0.000617139
R49977 d1.n77 d1 0.000617139
R49978 d1.n75 d1 0.000617139
R49979 d1.n73 d1 0.000617139
R49980 d1.n88 d1.n87 0.000617139
R49981 d1.n100 d1.n99 0.000617139
R49982 d1.n97 d1.n96 0.000617139
R49983 d1.n94 d1.n93 0.000617139
R49984 d1.n91 d1.n90 0.000617139
R49985 d1.n106 d1.n105 0.000617139
R49986 d1.n103 d1.n102 0.000617139
R49987 d1.n83 d1 0.000617139
R49988 d1.n81 d1 0.000617139
R49989 d1.n32 d1 0.000617139
R49990 d1.n40 d1 0.000617139
R49991 d1.n38 d1 0.000617139
R49992 d1.n36 d1 0.000617139
R49993 d1.n34 d1 0.000617139
R49994 d1.n49 d1.n48 0.000617139
R49995 d1.n61 d1.n60 0.000617139
R49996 d1.n58 d1.n57 0.000617139
R49997 d1.n55 d1.n54 0.000617139
R49998 d1.n52 d1.n51 0.000617139
R49999 d1.n67 d1.n66 0.000617139
R50000 d1.n64 d1.n63 0.000617139
R50001 d1.n44 d1 0.000617139
R50002 d1.n42 d1 0.000617139
R50003 d1.n17 d1 0.000617139
R50004 d1.n25 d1 0.000617139
R50005 d1.n23 d1 0.000617139
R50006 d1.n21 d1 0.000617139
R50007 d1.n19 d1 0.000617139
R50008 d1.n29 d1 0.000617139
R50009 d1.n27 d1 0.000617139
R50010 d1.n151 d1.n12 0.000617139
R50011 d1.n150 d1.n14 0.000617139
R50012 d1.n155 d1.n4 0.000617139
R50013 d1.n154 d1.n6 0.000617139
R50014 d1.n153 d1.n8 0.000617139
R50015 d1.n152 d1.n10 0.000617139
R50016 d1.n157 d1.n156 0.000617139
R50017 vrefl.n0 vrefl.t2 41.5062
R50018 vrefl.n1 vrefl.t1 31.2889
R50019 vrefl vrefl.t0 30.1295
R50020 vrefl.n2 vrefl.n1 3.51937
R50021 vrefl.n1 vrefl.n0 0.211106
R50022 vrefl vrefl.n2 0.0363796
R50023 vrefl.n2 vrefl 0.016125
R50024 vrefl.n0 vrefl 0.0133913
R50025 d3.n64 d3.t1 40.0866
R50026 d3.n51 d3.t0 40.0866
R50027 d3.n41 d3.t20 40.0866
R50028 d3.n15 d3.t19 40.0866
R50029 d3.n1 d3.t13 40.0866
R50030 d3.n10 d3.t23 40.0866
R50031 d3.n0 d3.t17 40.0866
R50032 d3.n20 d3.t25 40.0866
R50033 d3.n35 d3.t21 40.0866
R50034 d3.n30 d3.t18 40.0866
R50035 d3.n21 d3.t26 40.0866
R50036 d3.n56 d3.t28 40.0795
R50037 d3.n42 d3.t15 40.0795
R50038 d3.n62 d3.t3 40.0795
R50039 d3.n81 d3.t7 40.0322
R50040 d3.n74 d3.t29 40.0251
R50041 d3.n40 d3.n19 31.476
R50042 d3.n63 d3.n61 31.4135
R50043 d3.n56 d3.t5 23.8528
R50044 d3.n42 d3.t2 23.8528
R50045 d3.n51 d3.t14 23.8528
R50046 d3.n15 d3.t27 23.8528
R50047 d3.n1 d3.t30 23.8528
R50048 d3.n10 d3.t8 23.8528
R50049 d3.n0 d3.t6 23.8528
R50050 d3.n20 d3.t31 23.8528
R50051 d3.n30 d3.t4 23.8528
R50052 d3.n21 d3.t10 23.8528
R50053 d3.n62 d3.t11 23.8528
R50054 d3.n41 d3.t9 23.8457
R50055 d3.n35 d3.t12 23.8457
R50056 d3.n64 d3.t24 23.8457
R50057 d3.n81 d3.t22 23.7914
R50058 d3.n74 d3.t16 23.7914
R50059 d3.n61 d3.n40 21.8199
R50060 d3.n61 d3.n60 12.6287
R50061 d3.n40 d3.n39 12.5662
R50062 d3.n58 d3.n50 6.088
R50063 d3.n59 d3.n46 6.088
R50064 d3.n57 d3.n55 6.088
R50065 d3.n17 d3.n9 6.088
R50066 d3.n18 d3.n5 6.088
R50067 d3.n16 d3.n14 6.088
R50068 d3.n37 d3.n29 6.088
R50069 d3.n36 d3.n34 6.088
R50070 d3.n38 d3.n25 6.088
R50071 d3.n68 d3.n67 6.088
R50072 d3.n54 d3.n53 5.88488
R50073 d3.n45 d3.n44 5.88488
R50074 d3.n49 d3.n48 5.88488
R50075 d3.n13 d3.n12 5.88488
R50076 d3.n4 d3.n3 5.88488
R50077 d3.n8 d3.n7 5.88488
R50078 d3.n24 d3.n23 5.88488
R50079 d3.n33 d3.n32 5.88488
R50080 d3.n28 d3.n27 5.88488
R50081 d3.n70 d3.n69 5.88488
R50082 d3.n77 d3.n76 5.88488
R50083 d3.n73 d3.n72 5.88488
R50084 d3.n53 d3.n52 5.65675
R50085 d3.n48 d3.n47 5.65675
R50086 d3.n44 d3.n43 5.65675
R50087 d3.n12 d3.n11 5.65675
R50088 d3.n7 d3.n6 5.65675
R50089 d3.n3 d3.n2 5.65675
R50090 d3.n23 d3.n22 5.65675
R50091 d3.n27 d3.n26 5.65675
R50092 d3.n32 d3.n31 5.65675
R50093 d3.n80 d3.n70 5.65675
R50094 d3.n79 d3.n73 5.65675
R50095 d3.n78 d3.n77 5.65675
R50096 d3.n55 d3.n54 5.51612
R50097 d3.n50 d3.n49 5.51612
R50098 d3.n46 d3.n45 5.51612
R50099 d3.n14 d3.n13 5.51612
R50100 d3.n9 d3.n8 5.51612
R50101 d3.n5 d3.n4 5.51612
R50102 d3.n25 d3.n24 5.51612
R50103 d3.n29 d3.n28 5.51612
R50104 d3.n34 d3.n33 5.51612
R50105 d3.n69 d3.n68 5.51612
R50106 d3.n72 d3.n71 5.51612
R50107 d3.n76 d3.n75 5.51612
R50108 d3.n52 d3.n51 1.59714
R50109 d3.n11 d3.n10 1.59714
R50110 d3.n36 d3.n35 1.59714
R50111 d3.n22 d3.n21 1.59714
R50112 d3.n81 d3.n80 1.59714
R50113 d3.n65 d3.n64 1.59714
R50114 d3.n60 d3.n41 1.59703
R50115 d3.n19 d3.n0 1.59703
R50116 d3.n57 d3.n56 1.45966
R50117 d3.n43 d3.n42 1.45966
R50118 d3.n16 d3.n15 1.45966
R50119 d3.n2 d3.n1 1.45966
R50120 d3.n31 d3.n30 1.45966
R50121 d3.n78 d3.n74 1.45966
R50122 d3.n39 d3.n20 1.27758
R50123 d3.n63 d3.n62 1.27758
R50124 d3.n74 d3 0.384875
R50125 d3.n58 d3.n57 0.332778
R50126 d3.n59 d3.n58 0.332778
R50127 d3.n17 d3.n16 0.332778
R50128 d3.n18 d3.n17 0.332778
R50129 d3.n38 d3.n37 0.332778
R50130 d3.n37 d3.n36 0.332778
R50131 d3.n80 d3.n79 0.332778
R50132 d3.n79 d3.n78 0.332778
R50133 d3.n67 d3.n66 0.332778
R50134 d3.n66 d3.n65 0.332778
R50135 d3.n42 d3 0.313
R50136 d3.n41 d3 0.313
R50137 d3.n1 d3 0.313
R50138 d3.n0 d3 0.313
R50139 d3.n35 d3 0.313
R50140 d3.n30 d3 0.313
R50141 d3.n64 d3 0.313
R50142 d3 d3.n81 0.259875
R50143 d3.n56 d3 0.2505
R50144 d3.n15 d3 0.2505
R50145 d3.n20 d3 0.2505
R50146 d3.n62 d3 0.2505
R50147 d3.n51 d3 0.188
R50148 d3.n10 d3 0.188
R50149 d3.n21 d3 0.188
R50150 d3.n39 d3.n38 0.182579
R50151 d3.n67 d3.n63 0.182579
R50152 d3.n60 d3.n59 0.000617139
R50153 d3.n19 d3.n18 0.000617139
R50154 d5.n4 d5.t4 40.0866
R50155 d5.n2 d5.t3 40.0866
R50156 d5.n1 d5.t6 40.0866
R50157 d5.n0 d5.t5 40.0866
R50158 d5.n3 d5 24.7257
R50159 d5.n5 d5 24.4414
R50160 d5.n2 d5.t2 23.8528
R50161 d5.n1 d5.t1 23.8528
R50162 d5.n0 d5.t7 23.8528
R50163 d5.n4 d5.t0 23.8528
R50164 d5.n5 d5.n3 23.1567
R50165 d5 d5.n5 2.13198
R50166 d5.n3 d5 1.84761
R50167 d5 d5.n2 0.313
R50168 d5 d5.n1 0.313
R50169 d5 d5.n0 0.313
R50170 d5 d5.n4 0.313
R50171 X2.X2.X2.vrefh.n0 X2.X2.X2.vrefh.t1 41.5063
R50172 X2.X2.X2.vrefh.n1 X2.X2.X2.vrefh.t2 31.2889
R50173 X2.X2.X2.vrefh.n2 X2.X2.X2.vrefh.t0 30.264
R50174 X2.X2.X2.vrefh X2.X2.X2.vrefh.t3 30.0196
R50175 X2.X2.X2.vrefh.n2 X2.X2.X2.vrefh.n1 3.51937
R50176 X2.X2.X2.vrefh.n1 X2.X2.X2.vrefh.n0 0.211107
R50177 X2.X2.X2.vrefh.n0 X2.X2.X2.vrefh 0.0729068
R50178 X2.X2.X2.vrefh X2.X2.X2.vrefh.n2 0.0195972
R50179 X1.X2.X3.vin1.n0 X1.X2.X3.vin1.t2 43.0572
R50180 X1.X2.X3.vin1.t0 X1.X2.X3.vin1.t3 28.6406
R50181 X1.X2.X3.vin1 X1.X2.X3.vin1.t1 28.5751
R50182 X1.X2.X3.vin1 X1.X2.X3.vin1.n0 26.802
R50183 X1.X2.X3.vin1.n0 X1.X2.X3.vin1 1.29627
R50184 X1.X2.X3.vin1 X1.X2.X3.vin1.t0 0.959305
R50185 d4.n8 d4.n3 45.8392
R50186 d4.n15 d4.n13 45.8392
R50187 d4.n14 d4.t13 40.0866
R50188 d4.n11 d4.t7 40.0866
R50189 d4.n6 d4.t10 40.0866
R50190 d4.n2 d4.t4 40.0866
R50191 d4.n10 d4.t11 40.0322
R50192 d4.n5 d4.t9 40.0322
R50193 d4.n1 d4.t6 40.0322
R50194 d4.n16 d4.t12 40.0322
R50195 d4.n13 d4.n12 24.8948
R50196 d4.n8 d4.n7 24.8948
R50197 d4.n9 d4.t3 23.8528
R50198 d4.n11 d4.t1 23.8528
R50199 d4.n4 d4.t0 23.8528
R50200 d4.n6 d4.t2 23.8528
R50201 d4.n0 d4.t14 23.8528
R50202 d4.n2 d4.t15 23.8528
R50203 d4.n17 d4.t5 23.8528
R50204 d4.n14 d4.t8 23.8528
R50205 d4.n13 d4.n8 19.7227
R50206 d4.n12 d4.n11 1.76105
R50207 d4.n3 d4.n2 1.76105
R50208 d4.n7 d4.n5 1.74408
R50209 d4.n16 d4.n15 1.74408
R50210 d4.n15 d4.n14 1.51486
R50211 d4.n7 d4.n6 1.51486
R50212 d4.n12 d4.n10 1.49789
R50213 d4.n3 d4.n1 1.49789
R50214 d4.n11 d4 0.313
R50215 d4.n6 d4 0.313
R50216 d4.n2 d4 0.313
R50217 d4.n14 d4 0.313
R50218 d4.n9 d4 0.188
R50219 d4.n4 d4 0.188
R50220 d4.n0 d4 0.188
R50221 d4 d4.n17 0.188
R50222 d4.n10 d4.n9 0.0548478
R50223 d4.n5 d4.n4 0.0548478
R50224 d4.n1 d4.n0 0.0548478
R50225 d4.n17 d4.n16 0.0548478
R50226 d2.n66 d2.t42 40.0866
R50227 d2.n55 d2.t13 40.0866
R50228 d2.n56 d2.t2 40.0866
R50229 d2.n53 d2.t32 40.0866
R50230 d2.n47 d2.t38 40.0866
R50231 d2.n48 d2.t39 40.0866
R50232 d2.n49 d2.t18 40.0866
R50233 d2.n58 d2.t57 40.0866
R50234 d2.n60 d2.t5 40.0866
R50235 d2.n37 d2.t15 40.0866
R50236 d2.n38 d2.t58 40.0866
R50237 d2.n35 d2.t22 40.0866
R50238 d2.n29 d2.t27 40.0866
R50239 d2.n30 d2.t28 40.0866
R50240 d2.n31 d2.t24 40.0866
R50241 d2.n40 d2.t60 40.0866
R50242 d2.n42 d2.t8 40.0866
R50243 d2.n20 d2.t9 40.0866
R50244 d2.n21 d2.t61 40.0866
R50245 d2.n18 d2.t12 40.0866
R50246 d2.n12 d2.t19 40.0866
R50247 d2.n13 d2.t20 40.0866
R50248 d2.n14 d2.t35 40.0866
R50249 d2.n23 d2.t47 40.0866
R50250 d2.n25 d2.t63 40.0866
R50251 d2.n2 d2.t3 40.0866
R50252 d2.n10 d2.t48 40.0866
R50253 d2.n6 d2.t52 40.0866
R50254 d2.n7 d2.t53 40.0866
R50255 d2.n0 d2.t34 40.0866
R50256 d2.n4 d2.t14 40.0866
R50257 d2.n69 d2.t30 40.0866
R50258 d2.n65 d2.n64 25.7145
R50259 d2.n46 d2.n28 25.7131
R50260 d2.n55 d2.t21 23.8528
R50261 d2.n56 d2.t41 23.8528
R50262 d2.n53 d2.t37 23.8528
R50263 d2.n47 d2.t7 23.8528
R50264 d2.n48 d2.t59 23.8528
R50265 d2.n49 d2.t50 23.8528
R50266 d2.n58 d2.t26 23.8528
R50267 d2.n60 d2.t43 23.8528
R50268 d2.n37 d2.t23 23.8528
R50269 d2.n38 d2.t31 23.8528
R50270 d2.n35 d2.t25 23.8528
R50271 d2.n29 d2.t62 23.8528
R50272 d2.n30 d2.t44 23.8528
R50273 d2.n31 d2.t55 23.8528
R50274 d2.n40 d2.t29 23.8528
R50275 d2.n42 d2.t46 23.8528
R50276 d2.n20 d2.t10 23.8528
R50277 d2.n21 d2.t36 23.8528
R50278 d2.n18 d2.t17 23.8528
R50279 d2.n12 d2.t56 23.8528
R50280 d2.n13 d2.t40 23.8528
R50281 d2.n14 d2.t1 23.8528
R50282 d2.n23 d2.t11 23.8528
R50283 d2.n25 d2.t33 23.8528
R50284 d2.n2 d2.t45 23.8528
R50285 d2.n10 d2.t51 23.8528
R50286 d2.n6 d2.t16 23.8528
R50287 d2.n7 d2.t4 23.8528
R50288 d2.n0 d2.t0 23.8528
R50289 d2.n4 d2.t54 23.8528
R50290 d2.n69 d2.t6 23.8528
R50291 d2.n66 d2.t49 23.8528
R50292 d2.n64 d2.n46 20.7519
R50293 d2.n59 d2.n57 9.35243
R50294 d2.n41 d2.n39 9.35243
R50295 d2.n24 d2.n22 9.35243
R50296 d2.n5 d2.n3 9.35243
R50297 d2.n62 d2.n61 9.35243
R50298 d2.n44 d2.n43 9.35243
R50299 d2.n27 d2.n26 9.35243
R50300 d2.n68 d2.n67 9.35243
R50301 d2.n54 d2.n52 9.33579
R50302 d2.n36 d2.n34 9.33579
R50303 d2.n19 d2.n17 9.33579
R50304 d2.n11 d2.n9 9.33579
R50305 d2.n51 d2.n50 9.32359
R50306 d2.n33 d2.n32 9.32359
R50307 d2.n16 d2.n15 9.32359
R50308 d2.n52 d2.n51 9.24786
R50309 d2.n61 d2.n59 9.24786
R50310 d2.n34 d2.n33 9.24786
R50311 d2.n43 d2.n41 9.24786
R50312 d2.n17 d2.n16 9.24786
R50313 d2.n26 d2.n24 9.24786
R50314 d2.n9 d2.n8 9.24786
R50315 d2.n68 d2.n5 9.24786
R50316 d2.n46 d2.n45 5.79918
R50317 d2.n64 d2.n63 5.7978
R50318 d2.n3 d2.n1 2.79465
R50319 d2.n45 d2.n44 1.51198
R50320 d2.n67 d2.n65 1.51198
R50321 d2.n63 d2.n54 1.39016
R50322 d2.n28 d2.n19 1.39016
R50323 d2.n63 d2.n62 1.35282
R50324 d2.n28 d2.n27 1.35282
R50325 d2.n45 d2.n36 1.231
R50326 d2.n65 d2.n11 1.231
R50327 d2.n52 d2.n47 0.624393
R50328 d2.n51 d2.n48 0.624393
R50329 d2.n59 d2.n58 0.624393
R50330 d2.n61 d2.n60 0.624393
R50331 d2.n34 d2.n29 0.624393
R50332 d2.n33 d2.n30 0.624393
R50333 d2.n41 d2.n40 0.624393
R50334 d2.n43 d2.n42 0.624393
R50335 d2.n17 d2.n12 0.624393
R50336 d2.n16 d2.n13 0.624393
R50337 d2.n24 d2.n23 0.624393
R50338 d2.n26 d2.n25 0.624393
R50339 d2.n9 d2.n6 0.624393
R50340 d2.n8 d2.n7 0.624393
R50341 d2.n5 d2.n4 0.624393
R50342 d2.n69 d2.n68 0.624393
R50343 d2.n55 d2 0.313
R50344 d2.n56 d2 0.313
R50345 d2.n58 d2 0.313
R50346 d2.n60 d2 0.313
R50347 d2.n37 d2 0.313
R50348 d2.n38 d2 0.313
R50349 d2.n40 d2 0.313
R50350 d2.n42 d2 0.313
R50351 d2.n20 d2 0.313
R50352 d2.n21 d2 0.313
R50353 d2.n23 d2 0.313
R50354 d2.n25 d2 0.313
R50355 d2.n2 d2 0.313
R50356 d2.n4 d2 0.313
R50357 d2 d2.n69 0.313
R50358 d2.n66 d2 0.313
R50359 d2.n62 d2.n55 0.301802
R50360 d2.n57 d2.n56 0.301802
R50361 d2.n54 d2.n53 0.301802
R50362 d2.n50 d2.n49 0.301802
R50363 d2.n44 d2.n37 0.301802
R50364 d2.n39 d2.n38 0.301802
R50365 d2.n36 d2.n35 0.301802
R50366 d2.n32 d2.n31 0.301802
R50367 d2.n27 d2.n20 0.301802
R50368 d2.n22 d2.n21 0.301802
R50369 d2.n19 d2.n18 0.301802
R50370 d2.n15 d2.n14 0.301802
R50371 d2.n3 d2.n2 0.301802
R50372 d2.n11 d2.n10 0.301802
R50373 d2.n1 d2.n0 0.301802
R50374 d2.n67 d2.n66 0.301802
R50375 d2.n53 d2 0.188
R50376 d2.n47 d2 0.188
R50377 d2.n48 d2 0.188
R50378 d2.n49 d2 0.188
R50379 d2.n35 d2 0.188
R50380 d2.n29 d2 0.188
R50381 d2.n30 d2 0.188
R50382 d2.n31 d2 0.188
R50383 d2.n18 d2 0.188
R50384 d2.n12 d2 0.188
R50385 d2.n13 d2 0.188
R50386 d2.n14 d2 0.188
R50387 d2.n10 d2 0.188
R50388 d2.n6 d2 0.188
R50389 d2.n7 d2 0.188
R50390 d2.n0 d2 0.188
R50391 X1.X1.X3.vin2.t0 X1.X1.X3.vin2.t3 41.6232
R50392 X1.X1.X3.vin2 X1.X1.X3.vin2.t2 41.5063
R50393 X1.X1.X3.vin2.n0 X1.X1.X3.vin2.t1 30.1014
R50394 X1.X1.X3.vin2 X1.X1.X3.vin2.n0 28.8475
R50395 X1.X1.X3.vin2.n0 X1.X1.X3.vin2 1.39861
R50396 X1.X1.X3.vin2 X1.X1.X3.vin2.t0 0.958436
R50397 d6.n1 d6.t0 40.0866
R50398 d6.n0 d6.t3 40.0866
R50399 d6.n0 d6.t1 23.8528
R50400 d6.n1 d6.t2 23.8528
R50401 d6 d6.n0 0.313
R50402 d6 d6.n1 0.313
R50403 vout.n1 vout.t3 41.6232
R50404 vout.n1 vout.t0 41.6232
R50405 vout.n0 vout.t2 28.6406
R50406 vout.n0 vout.t1 28.6406
R50407 vout vout.n0 0.515744
R50408 vout vout.n1 0.439524
R50409 X3.vin1 X3.vin1.t3 44.0416
R50410 X3.vin1.t0 X3.vin1.t2 28.6406
R50411 X3.vin1 X3.vin1.t1 28.5751
R50412 X3.vin1 X3.vin1.t0 0.698671
R50413 X2.X2.X3.vin2.t0 X2.X2.X3.vin2.t1 41.6232
R50414 X2.X2.X3.vin2 X2.X2.X3.vin2.t3 41.5063
R50415 X2.X2.X3.vin2.n0 X2.X2.X3.vin2.t2 30.1014
R50416 X2.X2.X3.vin2 X2.X2.X3.vin2.n0 28.8475
R50417 X2.X2.X3.vin2.n0 X2.X2.X3.vin2 1.39861
R50418 X2.X2.X3.vin2 X2.X2.X3.vin2.t0 0.958436
R50419 X1.X2.X3.vin2.t0 X1.X2.X3.vin2.t1 41.6232
R50420 X1.X2.X3.vin2 X1.X2.X3.vin2.t2 41.5063
R50421 X1.X2.X3.vin2.n0 X1.X2.X3.vin2.t3 30.1014
R50422 X1.X2.X3.vin2 X1.X2.X3.vin2.n0 28.8475
R50423 X1.X2.X3.vin2.n0 X1.X2.X3.vin2 1.39861
R50424 X1.X2.X3.vin2 X1.X2.X3.vin2.t0 0.958436
R50425 X2.X1.X3.vin2.t2 X2.X1.X3.vin2.t1 41.6232
R50426 X2.X1.X3.vin2 X2.X1.X3.vin2.t4 41.5063
R50427 X2.X1.X3.vin2.n0 X2.X1.X3.vin2.t3 30.1014
R50428 X2.X1.X3.vin2 X2.X1.X3.vin2.n0 28.8475
R50429 X2.X1.X3.vin2 X2.X1.X3.vin2.t0 28.6406
R50430 X2.X1.X3.vin2.n0 X2.X1.X3.vin2 1.39861
R50431 X2.X1.X3.vin2 X2.X1.X3.vin2.t2 0.958436
R50432 X3.vin2 X3.vin2.t0 41.5063
R50433 X3.vin2.n0 X3.vin2.t3 30.1014
R50434 X3.vin2.t1 X3.vin2.t2 28.6406
R50435 X3.vin2 X3.vin2.n0 24.251
R50436 X3.vin2.n0 X3.vin2 1.39861
R50437 X3.vin2 X3.vin2.t1 0.698671
R50438 X1.X1.X3.vin1.n0 X1.X1.X3.vin1.t1 43.0572
R50439 X1.X1.X3.vin1.t0 X1.X1.X3.vin1.t3 28.6406
R50440 X1.X1.X3.vin1 X1.X1.X3.vin1.t2 28.5751
R50441 X1.X1.X3.vin1 X1.X1.X3.vin1.n0 26.802
R50442 X1.X1.X3.vin1.n0 X1.X1.X3.vin1 1.29627
R50443 X1.X1.X3.vin1 X1.X1.X3.vin1.t0 0.959305
R50444 X2.X1.X3.vin1.n0 X2.X1.X3.vin1.t2 43.0572
R50445 X2.X1.X3.vin1.t1 X2.X1.X3.vin1.t0 28.6406
R50446 X2.X1.X3.vin1 X2.X1.X3.vin1.t3 28.5751
R50447 X2.X1.X3.vin1 X2.X1.X3.vin1.n0 26.802
R50448 X2.X1.X3.vin1.n0 X2.X1.X3.vin1 1.29627
R50449 X2.X1.X3.vin1 X2.X1.X3.vin1.t1 0.959305
R50450 X2.X1.X2.vrefh.n0 X2.X1.X2.vrefh.t0 41.5063
R50451 X2.X1.X2.vrefh.n1 X2.X1.X2.vrefh.t3 31.2889
R50452 X2.X1.X2.vrefh.n2 X2.X1.X2.vrefh.t2 30.264
R50453 X2.X1.X2.vrefh X2.X1.X2.vrefh.t1 30.0201
R50454 X2.X1.X2.vrefh.n2 X2.X1.X2.vrefh.n1 3.51937
R50455 X2.X1.X2.vrefh.n1 X2.X1.X2.vrefh.n0 0.211107
R50456 X2.X1.X2.vrefh.n0 X2.X1.X2.vrefh 0.0729068
R50457 X2.X1.X2.vrefh X2.X1.X2.vrefh.n2 0.0195972
R50458 X1.X2.X2.vrefh.n0 X1.X2.X2.vrefh.t3 41.5063
R50459 X1.X2.X2.vrefh.n1 X1.X2.X2.vrefh.t1 31.2889
R50460 X1.X2.X2.vrefh.n2 X1.X2.X2.vrefh.t2 30.264
R50461 X1.X2.X2.vrefh X1.X2.X2.vrefh.t0 30.0201
R50462 X1.X2.X2.vrefh.n2 X1.X2.X2.vrefh.n1 3.51937
R50463 X1.X2.X2.vrefh.n1 X1.X2.X2.vrefh.n0 0.211107
R50464 X1.X2.X2.vrefh.n0 X1.X2.X2.vrefh 0.0729068
R50465 X1.X2.X2.vrefh X1.X2.X2.vrefh.n2 0.0195972
R50466 d7.n0 d7.t1 40.0866
R50467 d7.n0 d7.t0 23.8528
R50468 d7 d7.n0 0.313
R50469 X1.X1.X2.vrefh.n0 X1.X1.X2.vrefh.t3 41.5063
R50470 X1.X1.X2.vrefh.n1 X1.X1.X2.vrefh.t1 31.2889
R50471 X1.X1.X2.vrefh.n2 X1.X1.X2.vrefh.t0 30.264
R50472 X1.X1.X2.vrefh X1.X1.X2.vrefh.t2 30.0196
R50473 X1.X1.X2.vrefh.n2 X1.X1.X2.vrefh.n1 3.51937
R50474 X1.X1.X2.vrefh.n1 X1.X1.X2.vrefh.n0 0.211107
R50475 X1.X1.X2.vrefh.n0 X1.X1.X2.vrefh 0.0729068
R50476 X1.X1.X2.vrefh X1.X1.X2.vrefh.n2 0.0195972
R50477 vrefh vrefh.t0 30.0562
C0 X1.X1.X1.X2.X2.X2.vrefh X1.X1.X1.X2.X2.X2.X1.vin1 0.267f
C1 a_17222_19446# a_19336_18540# 4.72e-20
C2 a_17222_13728# X1.X2.X1.X2.X1.X2.X1.vin2 0.273f
C3 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.vout 0.326f
C4 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X3.vin1 0.00836f
C5 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 0.234f
C6 X1.X2.X1.X2.X2.X2.X3.vin1 a_17222_4198# 0.00207f
C7 X1.X2.X1.X1.X2.X2.vout X1.X2.X1.X1.X2.X2.X3.vin1 0.335f
C8 X2.X1.X1.X1.X2.X1.X2.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 0.234f
C9 a_46116_13728# a_46116_11822# 0.00396f
C10 a_54606_7922# a_54992_7922# 0.419f
C11 X1.X2.X2.X2.X2.X1.vout X1.X2.X2.X2.X3.vin2 0.399f
C12 a_54606_13640# a_52406_12640# 4.77e-21
C13 a_8186_22210# X1.X1.X2.X2.X1.X1.X3.vin2 0.00815f
C14 a_49002_29936# a_48702_28070# 5.55e-20
C15 X1.X2.X2.X1.X2.X1.vout X1.X2.X2.X1.X2.X1.X3.vin2 0.326f
C16 X2.X1.X1.X2.X1.X2.vrefh X1.X2.X2.X1.X2.X2.vrefh 0.117f
C17 X2.X1.X2.X2.X2.X2.X3.vin1 a_37466_29834# 0.00874f
C18 a_31476_21352# a_31476_19446# 0.00396f
C19 a_37852_25982# X2.X1.X2.X2.X1.X2.X3.vin2 0.00535f
C20 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X1.X2.X2.X1.X1.X1.vin1 0.668f
C21 X2.X2.X2.X2.X2.X1.X3.vin1 a_52792_27888# 0.199f
C22 a_23126_24076# a_25326_23170# 4.2e-20
C23 X2.X2.X2.X1.X1.X2.X2.vin1 a_54992_7922# 1.78e-19
C24 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 0.216f
C25 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X1.vin1 2.23e-19
C26 X2.X1.X1.X2.X1.X2.X3.vin2 a_31862_9916# 8.07e-19
C27 a_2196_30882# X1.X1.X1.X1.X1.X2.X1.vin1 1.64e-19
C28 a_2582_30882# a_2582_28976# 0.00198f
C29 X2.X1.X2.X3.vin1 a_37466_10734# 0.509f
C30 X2.X1.X3.vin2 X2.X1.X1.X2.X3.vin2 0.00254f
C31 a_31476_6104# a_31862_6104# 0.419f
C32 X1.X2.X2.X1.X1.X1.X2.vin1 X2.X1.X1.X2.X2.X2.X1.vin2 0.00232f
C33 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X1.vin2 0.076f
C34 X1.X2.X2.X1.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X1.vin2 8.93e-19
C35 X1.X2.X2.X1.X2.X1.X2.vin1 a_25326_11734# 8.88e-20
C36 X2.X1.X2.X2.X2.X1.X3.vin2 a_40352_28888# 0.354f
C37 X1.X1.X2.X1.X2.X1.X3.vin1 a_8872_12640# 0.199f
C38 a_46116_23258# a_46502_23258# 0.419f
C39 X1.X2.X1.X1.X2.vrefh a_16836_25164# 1.64e-19
C40 X2.X1.X1.X2.X2.X2.vrefh X1.X2.X2.X1.X1.X2.vrefh 0.117f
C41 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X2.X3.vin1 0.206f
C42 a_2582_28976# a_4396_28070# 1.06e-19
C43 X2.X1.X1.X2.X2.X1.X1.vin2 a_31862_8010# 8.88e-20
C44 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X2.vin1 0.0689f
C45 X1.X2.X2.X2.X2.X1.vout a_23126_27888# 0.422f
C46 X2.X1.X3.vin1 a_34362_14688# 3.28e-19
C47 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X3.vin2 0.161f
C48 X1.X1.X3.vin2 X1.X1.X2.X1.X3.vin1 0.0361f
C49 X1.X1.X2.X3.vin1 a_8572_10734# 0.356f
C50 a_10686_21264# X1.X1.X2.X2.X1.X1.X1.vin2 8.88e-20
C51 a_28482_892# X3.vin2 0.263f
C52 a_33676_28070# X2.X1.X1.X1.X1.X2.X3.vin2 0.101f
C53 a_17222_19446# X1.X2.X1.X2.X1.X1.X1.vin1 8.22e-20
C54 d7 a_28096_892# 0.502f
C55 a_52492_18358# a_52792_16452# 6.48e-19
C56 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.vrefh 2.33e-19
C57 a_39966_17452# X2.X1.X2.X1.X2.X2.X3.vin1 0.00207f
C58 X1.X1.X1.X1.X1.X2.vout a_4782_28070# 0.418f
C59 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.vout 0.0857f
C60 X2.X1.X2.X1.X1.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X1.vin1 2.23e-19
C61 X2.X1.X2.X1.X1.X1.X2.vin1 a_40352_4110# 1.78e-19
C62 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 2.23e-19
C63 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X2.X3.vin1 0.00789f
C64 a_10686_30794# X1.X1.X2.X2.X2.X2.X1.vin1 0.417f
C65 X1.X1.X2.X2.X2.X2.X1.vin2 a_11072_30794# 0.12f
C66 X2.X2.X1.X1.X1.X2.vrefh a_46116_30882# 0.118f
C67 a_52406_31700# a_52106_29834# 5.55e-20
C68 a_17222_9916# X1.X2.X1.X2.X2.X1.X2.vin1 8.88e-20
C69 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X2.vrefh 0.076f
C70 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X2.vin1 0.564f
C71 X1.X2.X2.X1.X2.X2.X3.vin2 a_23512_16452# 0.101f
C72 a_54606_32700# vrefl 0.3f
C73 X2.X2.X2.X2.X2.X2.X2.vin1 a_54992_32700# 0.197f
C74 a_23126_20264# X1.X2.X3.vin2 7.93e-20
C75 X1.X1.X2.X2.X2.X2.vout a_8872_31700# 0.36f
C76 X1.X1.X3.vin1 X1.X1.X2.X1.X1.X1.vout 5.53e-20
C77 X2.X1.X2.vrefh a_35312_892# 7.3e-19
C78 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.vrefh 2.33e-19
C79 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.X1.vin1 5.19e-19
C80 X2.X2.X1.X2.X2.X1.vout X2.X2.X1.X2.X2.X2.vout 0.514f
C81 a_4396_28070# a_5082_26164# 3.08e-19
C82 a_4782_28070# a_4696_26164# 3.3e-19
C83 a_46502_32788# X2.X2.X1.X1.X1.X1.X3.vin1 0.52f
C84 a_39966_28888# a_37766_27888# 4.77e-21
C85 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin1 0.195f
C86 X1.X2.X3.vin1 a_19422_12822# 2.12e-19
C87 X2.X1.X2.X2.X2.vrefh a_39966_25076# 0.3f
C88 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.vout 0.399f
C89 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X2.X3.vin1 0.0131f
C90 X1.X2.X2.X2.X1.X2.X1.vin2 X2.X1.X1.X1.X2.X1.X2.vin1 0.00232f
C91 X2.X1.X2.X1.X2.X1.vout a_37852_10734# 1.64e-19
C92 X1.X1.X1.X2.X1.X1.X3.vin1 a_2582_15634# 0.00207f
C93 X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X3.vin1 0.546f
C94 a_33976_7064# a_33676_5198# 6.71e-19
C95 X2.X1.X2.X1.X1.X1.X1.vin1 X2.X2.X2.vrefh 0.00437f
C96 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X2.vin1 0.0689f
C97 a_17222_6104# a_19036_5198# 1.06e-19
C98 a_19336_10916# a_19722_10916# 0.414f
C99 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X3.vin1 0.0131f
C100 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.vout 0.2f
C101 X2.X2.X1.X1.X3.vin2 a_49002_22312# 0.423f
C102 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X1.X3.vin2 5.19e-19
C103 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X3.vin1 0.00118f
C104 a_54992_9828# X2.X2.X2.X1.X1.X2.X1.vin2 1.78e-19
C105 X2.X1.X2.X2.X2.X1.vout X2.X1.X2.X2.X2.X1.X3.vin1 0.118f
C106 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.vout 0.118f
C107 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.vout 0.398f
C108 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.X1.X3.vin1 1.22e-19
C109 a_10686_7922# a_10686_6016# 0.00198f
C110 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X1.X1.vin2 8.93e-19
C111 X1.X1.X2.X2.X2.X1.X2.vin1 a_10686_26982# 8.88e-20
C112 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.vrefh 2.33e-19
C113 X1.X1.X2.X1.X2.X1.X3.vin1 a_10686_11734# 0.52f
C114 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X2.vrefh 0.267f
C115 X1.X1.X2.X3.vin1 a_8486_16452# 5.31e-19
C116 X1.X2.X1.X2.X2.X1.X3.vin2 a_19336_7064# 0.00546f
C117 a_54606_9828# a_54992_9828# 0.419f
C118 X2.X2.X2.X1.X2.X1.X3.vin1 a_54606_11734# 0.52f
C119 X2.X2.X1.X1.X2.X2.X2.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 0.234f
C120 X1.X2.X2.X1.X1.X1.X1.vin1 X2.X1.X2.vrefh 0.00437f
C121 a_48316_20446# a_48702_20446# 0.419f
C122 a_8186_25982# X1.X1.X2.X2.X1.X2.X3.vin2 0.00846f
C123 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X1.vin2 0.668f
C124 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin1 0.267f
C125 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 2.23e-19
C126 a_46502_9916# X2.X2.X1.X2.X2.X1.X1.vin1 0.417f
C127 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin2 0.12f
C128 a_8186_14586# a_8572_14586# 0.419f
C129 a_46116_9916# X2.X2.X1.X2.X2.X1.X3.vin1 0.354f
C130 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X1.vin1 0.206f
C131 X2.X2.X3.vin2 X2.X3.vin2 0.147f
C132 X2.X2.X3.vin2 a_52406_12640# 2.33e-19
C133 a_37852_14586# a_37766_12640# 3.14e-19
C134 a_25326_28888# X1.X2.X2.X2.X2.X1.X3.vin2 0.567f
C135 X2.X2.X1.X1.X2.X1.X2.vin1 a_46502_23258# 0.402f
C136 X2.X2.X2.X2.X1.X2.vout a_52792_24076# 0.36f
C137 X2.X1.X1.X1.X2.X1.vout a_34362_22312# 0.383f
C138 a_19422_31882# a_17222_30882# 4.77e-21
C139 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X3.vin1 2.33e-19
C140 a_23512_12640# a_22826_10734# 2.97e-19
C141 X1.X1.X1.X1.X1.X1.vout a_5082_29936# 0.386f
C142 a_4782_31882# X1.X1.X1.X1.X3.vin1 1.52e-19
C143 X2.X1.X3.vin1 a_34926_892# 0.17f
C144 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.vout 0.197f
C145 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X3.vin1 0.0131f
C146 X2.X1.X2.X1.X2.X1.X3.vin1 a_40352_11734# 0.354f
C147 a_40352_6016# X2.X1.X2.X1.X1.X1.X1.vin2 1.78e-19
C148 a_25326_19358# X1.X2.X2.X2.vrefh 8.22e-20
C149 a_33676_20446# a_33976_18540# 6.48e-19
C150 a_2196_15634# a_2582_15634# 0.419f
C151 X2.X1.X1.X1.X2.X2.X2.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 0.234f
C152 a_33676_20446# a_34062_20446# 0.419f
C153 X1.X2.X1.X2.X1.X2.vout X1.X2.X1.X2.X1.X2.X3.vin2 0.075f
C154 a_25326_9828# a_23126_8828# 4.77e-21
C155 X2.X2.X1.X1.X1.X2.X3.vin1 X2.X2.X1.X1.X1.X2.X3.vin2 0.587f
C156 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 0.242f
C157 a_25326_17452# a_25326_15546# 0.00198f
C158 a_48616_29936# X2.X2.X1.X1.X1.X2.vout 0.0929f
C159 X1.X1.X1.X1.X1.X2.vrefh a_2196_30882# 0.118f
C160 a_54992_26982# a_54992_25076# 0.00396f
C161 X2.X2.X1.X1.X1.X1.vout X2.X2.X1.X1.X3.vin1 0.13f
C162 X1.X1.X1.X2.X1.X1.X2.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 0.234f
C163 X2.X2.X1.X1.X1.X1.X2.vin1 X2.X2.X1.X1.X1.X2.vrefh 0.564f
C164 X1.X1.X1.X1.X2.X1.X3.vin1 a_4782_24258# 0.428f
C165 a_37766_24076# X2.X1.X2.X2.X1.X2.vout 0.418f
C166 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin1 0.267f
C167 X1.X1.X3.vin1 a_8486_5016# 8.66e-20
C168 a_4396_24258# a_4696_22312# 6.1e-19
C169 a_25712_7922# a_25712_6016# 0.00396f
C170 a_33976_14688# X2.X1.X1.X2.X1.X2.X3.vin1 0.00329f
C171 X2.X1.X2.X1.X1.X1.vout a_38152_5016# 0.359f
C172 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin1 0.267f
C173 a_39966_30794# a_40352_30794# 0.419f
C174 a_10686_19358# X1.X1.X2.X2.vrefh 8.22e-20
C175 X2.X1.X2.X2.X2.X2.vrefh X2.X1.X2.X2.X2.X1.X1.vin2 0.076f
C176 X1.X2.X1.X1.X2.X2.X2.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 0.234f
C177 a_19036_20446# a_19422_20446# 0.419f
C178 a_2196_8010# a_2582_8010# 0.419f
C179 X2.X2.X1.X1.X2.vrefh X2.X1.X2.X2.X2.vrefh 0.117f
C180 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X3.vin2 1.42e-20
C181 X1.X2.X3.vin2 a_23126_16452# 3.98e-19
C182 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin1 0.267f
C183 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 2.23e-19
C184 X2.X1.X1.X1.X2.X2.X3.vin1 a_34062_20446# 0.42f
C185 X2.X2.X1.X2.X1.X2.X3.vin2 a_48616_10916# 0.00535f
C186 a_48702_12822# a_49002_10916# 4.41e-20
C187 X2.X2.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X1.vout 0.13f
C188 X1.X1.X1.X1.X1.X1.X1.vin2 a_4396_31882# 0.00113f
C189 a_46116_9916# a_46116_8010# 0.00396f
C190 a_25326_11734# X1.X2.X2.X1.X1.X2.X3.vin2 8.07e-19
C191 X1.X2.X3.vin2 a_23126_8828# 2.33e-19
C192 X1.X2.X1.X1.X1.X2.vout a_19336_26164# 7.93e-20
C193 X2.X1.X3.vin1 a_34362_10916# 6.09e-19
C194 X1.X2.X1.X1.X1.X1.X3.vin2 a_19722_29936# 0.00815f
C195 X2.X1.X2.X3.vin2 a_37852_25982# 0.355f
C196 X2.X2.X1.X2.X2.vrefh a_46116_11822# 0.118f
C197 X1.X2.X2.X1.X3.vin1 a_23212_6962# 0.363f
C198 a_52106_25982# a_52792_24076# 3.08e-19
C199 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X3.vin2 0.161f
C200 X1.X1.X2.X1.X2.X2.X3.vin2 a_8186_14586# 3.85e-19
C201 a_10686_7922# a_8572_6962# 2.68e-20
C202 X1.X2.X2.X1.X1.X1.X1.vin2 X2.X1.X1.X2.X2.X2.X2.vin1 0.00232f
C203 X1.X1.X2.X2.X1.X2.X3.vin1 a_11072_23170# 0.354f
C204 a_40352_17452# a_40352_15546# 0.00396f
C205 a_2582_6104# X1.X1.X1.X2.X2.X2.X1.vin2 0.273f
C206 X1.X2.X2.X1.X1.X1.vout X1.X2.X2.X1.X1.X1.X3.vin2 0.342f
C207 X1.X2.X1.X2.X1.X1.vout X1.X2.X1.X2.X1.X1.X3.vin2 0.342f
C208 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin2 0.17f
C209 X1.X1.X3.vin1 a_8186_10734# 3.93e-19
C210 a_54606_13640# a_54992_13640# 0.419f
C211 X2.X2.X1.X2.X3.vin2 a_48702_9010# 0.00101f
C212 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.vrefh 0.161f
C213 X1.X2.X2.X2.X2.X1.X1.vin2 X2.X1.X1.X1.X2.vrefh 0.0128f
C214 a_4396_24258# a_2582_23258# 1.15e-20
C215 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X3.vin1 0.00118f
C216 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin2 7.84e-19
C217 a_16836_28976# a_17222_28976# 0.419f
C218 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X2.X1.X1.X1.X2.X1.vin2 0.00232f
C219 a_37466_18358# a_37852_18358# 0.416f
C220 X1.X1.X2.X2.vrefh a_11072_17452# 0.118f
C221 a_46116_13728# X2.X2.X1.X2.X1.X2.X3.vin1 0.354f
C222 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X1.X2.X2.X2.X2.vrefh 0.1f
C223 a_19336_7064# a_17222_6104# 2.68e-20
C224 a_46502_13728# X2.X2.X1.X2.X1.X2.X1.vin1 0.417f
C225 X2.X1.X2.X2.X2.X2.X2.vin1 a_38152_31700# 5.34e-19
C226 X1.X1.X1.X1.X2.X2.X3.vin1 a_4396_20446# 0.199f
C227 a_37852_25982# a_37766_24076# 3.3e-19
C228 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin2 7.84e-19
C229 a_19036_31882# X1.X2.X1.X1.X1.X1.vout 0.359f
C230 X2.X1.X2.X1.X2.X2.vout X2.X1.X2.X1.X3.vin2 0.0866f
C231 a_14082_892# X3.vin1 0.472f
C232 a_38152_12640# a_39966_11734# 1.06e-19
C233 X2.X1.X1.X2.X2.vrefh a_31862_11822# 0.3f
C234 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X2.vin1 0.0689f
C235 a_17222_25164# a_19036_24258# 1.06e-19
C236 a_37852_10734# a_39966_9828# 4.72e-20
C237 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.vrefh 2.33e-19
C238 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X3.vin2 8.93e-19
C239 a_31476_6104# a_31476_4198# 0.00396f
C240 a_39966_6016# a_37766_5016# 4.77e-21
C241 X1.X2.X2.X1.X2.X2.X3.vin1 a_23212_14586# 0.00329f
C242 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X2.vin1 0.242f
C243 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X1.vin2 0.216f
C244 X1.X1.X2.X1.X1.X1.vout a_8486_5016# 0.422f
C245 a_10686_9828# X1.X1.X2.X1.X1.X2.X1.vin2 8.88e-20
C246 X1.X2.X1.X2.X2.X1.vout X1.X2.X1.X2.X2.X1.X3.vin2 0.326f
C247 a_46502_27070# X2.X2.X1.X1.X2.X1.X1.vin1 8.22e-20
C248 a_52106_29834# a_52792_27888# 2.86e-19
C249 a_33976_29936# X2.X1.X1.X1.X3.vin1 0.363f
C250 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 1.22e-19
C251 X2.X2.X2.X2.X3.vin2 X2.X2.X2.X3.vin2 0.17f
C252 a_4696_14688# a_4396_12822# 6.71e-19
C253 X2.X2.X2.X2.X2.X1.vout a_52492_25982# 1.64e-19
C254 a_37852_6962# a_37766_5016# 3.14e-19
C255 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.X1.vin2 0.216f
C256 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X3.vin2 0.161f
C257 X2.X2.X2.X2.X2.X1.X1.vin2 a_54606_26982# 0.273f
C258 X3.vin2 a_34926_892# 4.87e-19
C259 a_17222_8010# X1.X2.X1.X2.X2.X2.X1.vin1 8.22e-20
C260 X1.X2.X1.X1.X1.X1.X3.vin2 X1.X2.X1.X1.X1.X2.X3.vin1 1.22e-19
C261 X1.X1.X1.X3.vin2 a_4782_9010# 7.93e-20
C262 X2.X1.X1.X1.X1.X1.X3.vin2 a_33976_29936# 0.00546f
C263 X1.X2.X2.X1.X2.vrefh a_25712_9828# 0.118f
C264 a_10686_11734# X1.X1.X2.X1.X2.vrefh 8.22e-20
C265 X2.X2.X2.X2.X1.X1.vout a_52406_20264# 0.422f
C266 a_10686_6016# a_10686_4110# 0.00198f
C267 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 0.242f
C268 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.vout 0.08f
C269 X1.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X3.vin2 0.0533f
C270 a_4396_20446# a_4696_18540# 6.48e-19
C271 X2.X1.X1.X2.X1.X2.X1.vin2 a_31862_11822# 8.88e-20
C272 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X2.vin1 0.242f
C273 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.vout 0.398f
C274 X1.X2.X3.vin1 a_20672_892# 0.386f
C275 a_31476_23258# a_31476_21352# 0.00396f
C276 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 2.23e-19
C277 X2.X1.X1.X2.X1.X2.X3.vin1 a_34062_12822# 0.42f
C278 a_4782_20446# a_2582_19446# 4.77e-21
C279 X2.X2.X2.X2.X2.X2.X3.vin2 a_54606_30794# 7.84e-19
C280 X2.X2.X2.X2.X2.X2.X2.vin1 X2.X2.X2.X2.X2.X2.X1.vin1 0.0689f
C281 X1.X1.X1.X1.X2.X2.X3.vin2 a_2196_19446# 0.354f
C282 a_25326_15546# X1.X2.X2.X1.X2.X2.X1.vin1 0.417f
C283 X1.X2.X2.X1.X2.X2.X1.vin2 a_25712_15546# 0.12f
C284 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X2.X1.X1.vin1 0.668f
C285 a_46116_9916# X2.X2.X1.X2.X2.X1.X2.vin1 1.78e-19
C286 X1.X1.X2.X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X3.vin1 0.00118f
C287 X1.X2.X2.X2.X1.X1.X3.vin2 a_23512_20264# 0.1f
C288 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X2.vrefh 0.076f
C289 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X2.vrefh 0.076f
C290 X1.X1.X2.X1.X1.X1.X3.vin1 a_11072_4110# 0.354f
C291 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X2.X1.X2.vrefh 0.0128f
C292 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X1.X3.vin1 0.0425f
C293 a_52792_16452# a_52106_14586# 3.31e-19
C294 a_17222_21352# a_19422_20446# 4.2e-20
C295 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X1.X2.X2.X2.vin1 0.00117f
C296 X1.X2.X1.X3.vin2 a_19336_10916# 0.355f
C297 X1.X1.X1.X1.X3.vin1 a_4696_26164# 0.169f
C298 a_42976_892# X2.X3.vin2 0.0927f
C299 a_19722_29936# a_19422_28070# 5.55e-20
C300 a_54606_6016# a_54606_4110# 0.00198f
C301 X1.X1.X2.X1.X3.vin1 a_8186_6962# 0.436f
C302 X1.X2.X2.X2.X3.vin1 a_23212_25982# 0.17f
C303 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 0.242f
C304 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.vrefh 0.00118f
C305 X2.X1.X1.X3.vin1 X2.X1.X3.vin2 7.53e-21
C306 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X2.vin1 0.564f
C307 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X1.vin1 5.19e-19
C308 X2.X2.X1.X1.X1.X2.vout X2.X2.X1.X1.X1.X2.X3.vin1 0.326f
C309 a_39966_32700# X2.X1.X2.X2.X2.X2.X1.vin2 8.88e-20
C310 X1.X1.X2.X2.X1.X2.X3.vin1 a_8872_24076# 0.199f
C311 X1.X2.X2.X2.X2.X1.X1.vin1 a_25712_26982# 0.195f
C312 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X1.vin2 0.668f
C313 a_8486_8828# a_10686_7922# 4.2e-20
C314 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 0.216f
C315 a_25326_25076# X1.X2.X2.X2.X1.X2.X3.vin1 0.00207f
C316 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.X1.X1.X1.vin2 3.94e-19
C317 X2.X1.X2.X2.X1.X1.X3.vin1 a_37466_18358# 0.00837f
C318 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.X1.vin2 0.216f
C319 a_37766_16452# a_37852_14586# 3.38e-19
C320 a_23512_24076# a_23212_22210# 6.71e-19
C321 X1.X2.X2.X1.X1.X2.X1.vin2 a_25712_7922# 0.12f
C322 a_25326_7922# X1.X2.X2.X1.X1.X2.X1.vin1 0.417f
C323 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X1.vin2 3.94e-19
C324 a_22826_18358# X1.X2.X3.vin2 0.451f
C325 X2.X1.X1.X2.X1.X2.X2.vin1 X2.X1.X1.X2.X2.vrefh 0.564f
C326 a_37766_12640# X2.X1.X2.X1.X2.X1.X3.vin1 0.428f
C327 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.X1.vin1 2.23e-19
C328 a_8486_16452# X1.X1.X2.X1.X2.X2.vout 0.418f
C329 X1.X2.X2.X2.X2.X2.X2.vin1 a_25712_30794# 1.78e-19
C330 X2.X1.X1.X1.X2.X1.X3.vin2 a_31862_23258# 0.567f
C331 a_52106_10734# X2.X2.X2.X1.X3.vin1 0.385f
C332 X1.X2.X2.X1.X1.X2.vrefh a_25712_6016# 0.118f
C333 X1.X1.X1.X2.X2.X1.X3.vin2 X1.X1.X1.X2.X2.X2.X1.vin1 5.19e-19
C334 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X2.vrefh 0.267f
C335 X2.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 8.36e-19
C336 X1.X1.X2.X2.X1.X2.X3.vin1 a_8186_22210# 0.00874f
C337 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X1.vout 0.0524f
C338 a_37466_14586# X2.X1.X2.X1.X2.X1.X3.vin2 0.00815f
C339 a_48702_31882# X2.X2.X1.X1.X1.X1.vout 0.422f
C340 X2.X2.X2.X1.X1.X1.X3.vin1 a_54606_4110# 0.52f
C341 X1.X2.X2.X2.X1.X2.X2.vin1 a_25712_25076# 0.197f
C342 X2.X2.X1.X2.X1.X2.vout a_48616_10916# 7.93e-20
C343 a_40352_32700# X2.X2.vrefh 0.118f
C344 a_22826_10734# a_23212_10734# 0.414f
C345 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin1 0.52f
C346 a_19036_12822# a_17222_11822# 1.15e-20
C347 a_54606_19358# a_54606_17452# 0.00198f
C348 X1.X1.X2.X2.X2.X2.X2.vin1 a_10686_30794# 8.88e-20
C349 X2.X1.X2.X1.X2.X2.X2.vin1 a_40352_17452# 0.197f
C350 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.X1.vin2 8.93e-19
C351 a_34062_16634# a_31862_15634# 4.77e-21
C352 X1.X2.X1.X1.X1.X2.X1.vin2 a_17222_27070# 8.88e-20
C353 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.vrefh 0.161f
C354 X2.X1.X2.X2.X1.X1.X3.vin2 a_37466_18358# 3.49e-19
C355 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.X1.vin2 0.23f
C356 X2.X2.X2.X2.X1.X1.X1.vin2 X2.X2.X2.X2.vrefh 0.1f
C357 X2.X1.X2.X2.X3.vin2 X2.X1.X2.X2.X3.vin1 0.552f
C358 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 0.049f
C359 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X1.vin2 0.668f
C360 a_2582_17540# X1.X1.X1.X2.X1.X1.X2.vin1 8.88e-20
C361 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X3.vin1 1.42e-20
C362 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin1 0.52f
C363 X1.X2.X2.X1.X1.X2.X3.vin2 a_22826_6962# 3.85e-19
C364 a_25326_30794# a_23212_29834# 2.68e-20
C365 X2.X1.X1.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X1.X2.vrefh 0.165f
C366 X1.X2.X1.X1.X1.X2.X3.vin1 a_19422_28070# 0.42f
C367 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X2.X3.vin2 2.23e-19
C368 a_34362_29936# X2.X1.X1.X1.X1.X2.X3.vin2 3.85e-19
C369 X2.X1.X1.X1.X3.vin1 a_34062_28070# 9.54e-19
C370 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X2.vrefh 0.267f
C371 X1.X2.X2.X2.X1.X1.X2.vin1 a_25712_19358# 1.78e-19
C372 X2.X1.X2.X1.X1.X1.X3.vin1 a_39966_4110# 0.52f
C373 X1.X2.X2.X2.X1.X1.X3.vin2 X1.X2.X2.X2.X1.X1.X1.vin1 2.23e-19
C374 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X2.vin1 0.242f
C375 X2.X2.X1.X1.X2.X2.X2.vin1 a_46502_19446# 0.402f
C376 a_54606_17452# a_54606_15546# 0.00198f
C377 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 0.242f
C378 a_23512_8828# a_22826_6962# 3.31e-19
C379 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X1.vin2 0.076f
C380 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.vrefh 2.33e-19
C381 a_8872_5016# a_10686_4110# 1.06e-19
C382 X1.X1.X2.vrefh a_2582_4198# 0.301f
C383 X1.X2.X1.X2.X2.vrefh a_16836_9916# 1.64e-19
C384 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X1.X3.vin2 0.0533f
C385 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X2.vout 0.0866f
C386 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X3.vin1 0.0131f
C387 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 2.23e-19
C388 X1.X1.X2.X2.X1.X2.X1.vin2 a_10686_23170# 0.273f
C389 X1.X2.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X2.X1.X3.vin1 0.00118f
C390 X2.X1.X2.X2.X1.X2.vout X2.X1.X2.X2.X1.X1.vout 0.507f
C391 a_39966_19358# a_40352_19358# 0.419f
C392 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X1.vin2 0.076f
C393 a_34062_9010# a_31862_8010# 4.77e-21
C394 a_39966_9828# a_38152_8828# 1.15e-20
C395 X1.X2.X3.vin2 X1.X2.X2.X1.X3.vin2 0.039f
C396 a_54992_7922# a_54992_6016# 0.00396f
C397 X1.X2.X2.X1.X1.X1.X3.vin1 X1.X2.X2.X1.X1.X1.X1.vin1 0.206f
C398 X2.X2.X2.X1.X2.X2.X1.vin2 X2.X2.X2.X1.X2.X2.vrefh 0.1f
C399 a_11072_23170# a_11072_21264# 0.00396f
C400 a_48616_7064# X2.X2.X1.X2.X2.X2.vout 0.0929f
C401 a_8572_29834# a_8486_27888# 3.14e-19
C402 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X3.vin2 0.449f
C403 X2.X1.X1.X1.X2.X2.X2.vin1 a_31476_19446# 0.197f
C404 X2.X1.X1.X2.X1.X1.X3.vin1 a_33676_16634# 0.199f
C405 a_49002_18540# X2.X2.X1.X2.X1.X1.X3.vin2 3.49e-19
C406 X2.X2.X1.X3.vin2 a_48702_16634# 5.21e-19
C407 a_52492_22210# a_54606_21264# 2.95e-20
C408 a_25326_21264# a_25712_21264# 0.419f
C409 a_37852_10734# a_38152_8828# 6.48e-19
C410 a_17222_9916# a_17222_8010# 0.00198f
C411 X1.X1.X2.X1.X1.X2.X2.vin1 a_11072_9828# 0.197f
C412 a_52792_31700# a_52492_29834# 6.71e-19
C413 a_17222_21352# X1.X2.X1.X1.X2.X2.X1.vin1 0.417f
C414 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 0.242f
C415 a_10686_25076# a_10686_23170# 0.00198f
C416 a_16836_21352# X1.X2.X1.X1.X2.X2.X3.vin1 0.354f
C417 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin1 0.52f
C418 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X2.vin1 0.564f
C419 a_25712_32700# X1.X2.X2.X2.X2.X2.X1.vin2 1.78e-19
C420 a_25326_19358# a_25712_19358# 0.419f
C421 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X1.vin2 0.216f
C422 X2.X2.X1.X1.X2.X2.X1.vin2 a_46116_19446# 1.78e-19
C423 X2.X2.X2.X1.X1.X2.X3.vin1 a_52492_6962# 0.00329f
C424 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X3.vin2 8.93e-19
C425 a_8186_18358# X1.X1.X2.X3.vin1 0.374f
C426 X1.X1.X1.X3.vin2 X1.X1.X3.vin2 3.82e-19
C427 X2.X2.X1.X3.vin2 a_48702_9010# 7.93e-20
C428 X1.X1.X2.X1.X2.X1.vout a_8486_12640# 0.422f
C429 X2.X1.X2.X1.X2.vrefh a_39966_9828# 0.3f
C430 X1.X2.X3.vin2 a_23126_12640# 2.33e-19
C431 a_34062_24258# X2.X1.X1.X1.X2.X1.X3.vin2 0.267f
C432 X2.X2.X2.vrefh a_46116_4198# 0.119f
C433 a_46502_13728# a_46502_11822# 0.00198f
C434 X2.X2.X2.X1.X1.X2.X1.vin2 X2.X2.X2.X1.X1.X2.vrefh 0.1f
C435 X1.X2.X1.X1.X2.X2.X2.vin1 a_16836_19446# 0.197f
C436 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X2.vrefh 0.00118f
C437 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X3.vin1 0.00117f
C438 a_10686_19358# a_8572_18358# 5.36e-21
C439 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X2.X3.vin2 0.0565f
C440 X2.X2.X2.X1.X2.X1.X3.vin2 a_52406_12640# 0.267f
C441 X1.X2.X1.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X1.vin2 0.1f
C442 a_52106_14586# a_52492_14586# 0.419f
C443 a_10686_17452# a_8486_16452# 4.77e-21
C444 a_31862_21352# a_31862_19446# 0.00198f
C445 a_33976_22312# X2.X1.X1.X1.X2.X2.vout 0.0929f
C446 X1.X1.X2.X2.X1.X1.X3.vin1 a_8186_18358# 0.00837f
C447 X1.X2.X2.X1.X2.X1.X3.vin1 a_23512_12640# 0.199f
C448 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X1.X3.vin2 1.22e-19
C449 a_10686_25076# X1.X1.X2.X2.X1.X2.X2.vin1 0.402f
C450 X1.X2.X2.X1.X2.X2.X1.vin2 X1.X2.X2.X1.X2.X2.vrefh 0.1f
C451 a_10686_19358# a_11072_19358# 0.419f
C452 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X1.vin1 0.206f
C453 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X3.vin1 1.22e-19
C454 a_33676_16634# X2.X1.X1.X2.X1.X1.vout 0.359f
C455 a_48316_28070# a_48702_28070# 0.419f
C456 X2.X1.X2.X2.X2.X2.X3.vin1 a_38152_31700# 0.199f
C457 X2.X2.X1.X1.X1.X2.X2.vin1 X2.X2.X1.X1.X1.X2.X3.vin2 0.234f
C458 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X2.X2.vin1 0.242f
C459 a_39966_6016# a_40352_6016# 0.419f
C460 X1.X2.X1.X1.X2.X1.X2.vin1 a_17222_23258# 0.402f
C461 a_25326_17452# X1.X2.X2.X1.X2.X2.X2.vin1 0.402f
C462 a_46502_25164# X2.X2.X1.X1.X2.X1.X2.vin1 8.88e-20
C463 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X3.vin1 0.00118f
C464 X2.X2.X1.X2.vrefh X2.X1.X2.X2.vrefh 0.117f
C465 a_25712_21264# X1.X2.X2.X2.X1.X1.X1.vin2 1.78e-19
C466 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.vrefh 2.33e-19
C467 X1.X2.X2.X2.X2.X2.X1.vin2 X2.X1.X1.X1.X1.X2.vrefh 0.0128f
C468 a_31476_6104# X2.X1.X1.X2.X2.X2.X3.vin1 0.354f
C469 a_31862_6104# X2.X1.X1.X2.X2.X2.X1.vin1 0.417f
C470 X1.X2.X2.X2.X2.X2.vout X1.X2.X2.X2.X2.X1.vout 0.514f
C471 X1.X1.X1.X1.X2.X2.X2.vin1 X1.X1.X1.X2.vrefh 0.564f
C472 a_8486_20264# X1.X1.X2.X2.X1.X1.X3.vin1 0.428f
C473 X1.X2.X2.X1.X2.X1.X2.vin1 a_25712_11734# 1.78e-19
C474 X1.X2.X2.X1.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X1.vin1 2.23e-19
C475 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin1 0.267f
C476 a_38152_27888# a_37852_25982# 6.2e-19
C477 X1.X1.X1.X1.X1.X2.X3.vin1 a_4396_28070# 0.199f
C478 X1.X2.X2.X2.X1.X1.vout a_23212_18358# 1.64e-19
C479 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin2 7.84e-19
C480 X1.X1.X1.X2.X1.X2.X2.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 0.234f
C481 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X1.vin1 5.19e-19
C482 a_4396_12822# a_4782_12822# 0.419f
C483 a_37766_24076# a_37852_22210# 3.38e-19
C484 a_25712_25076# a_25712_23170# 0.00396f
C485 X1.X1.X2.X2.X1.X1.X3.vin2 X1.X1.X2.X2.X1.X1.X1.vin2 8.93e-19
C486 X2.X2.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.vout 0.398f
C487 X1.X1.X2.X2.X1.X1.X2.vin1 a_10686_19358# 8.88e-20
C488 a_4696_14688# a_5082_14688# 0.419f
C489 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin2 7.84e-19
C490 X1.X1.X2.X2.X2.X2.X3.vin1 a_8186_29834# 0.00874f
C491 X1.X2.X2.X1.X1.X2.X1.vin2 X1.X2.X2.X1.X1.X2.vrefh 0.1f
C492 X2.X1.X1.X3.vin1 a_34362_18540# 0.389f
C493 X1.X2.X2.vrefh a_16836_4198# 0.119f
C494 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 0.139f
C495 a_46502_8010# X2.X2.X1.X2.X2.X2.X1.vin1 8.22e-20
C496 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X1.vin2 0.076f
C497 X1.X2.X1.X1.X1.X1.X2.vin1 X1.X2.X1.X1.X1.X2.vrefh 0.564f
C498 a_33676_9010# X2.X1.X1.X2.X2.X1.vout 0.359f
C499 a_23126_31700# X1.X2.X2.X2.X2.X2.X3.vin1 0.42f
C500 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.X3.vin1 0.587f
C501 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X2.X1.vin1 5.19e-19
C502 X1.X1.X1.X2.X1.X2.X1.vin2 a_2196_11822# 1.78e-19
C503 a_19036_12822# a_19722_10916# 3.08e-19
C504 a_19422_12822# a_19336_10916# 3.3e-19
C505 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X3.vin2 0.418f
C506 X1.X1.X3.vin2 X1.X1.X2.X1.X2.X1.vout 3.2e-19
C507 X2.X1.X3.vin2 a_37466_6962# 0.00111f
C508 a_2582_23258# X1.X1.X1.X1.X2.X2.X1.vin1 8.22e-20
C509 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X1.X2.X2.X1.X2.X1.vin1 0.668f
C510 X1.X1.X2.X2.X2.X2.X1.vin1 a_11072_30794# 0.195f
C511 X1.X2.X2.X2.X2.X1.X3.vin1 a_25326_26982# 0.52f
C512 a_11072_19358# a_11072_17452# 0.00396f
C513 X2.X2.X2.X2.X2.X1.X3.vin2 a_52106_25982# 3.49e-19
C514 a_34362_10916# X2.X1.X1.X2.X2.X1.X3.vin1 0.00837f
C515 a_52792_31700# a_54606_30794# 1.06e-19
C516 a_8872_12640# a_8186_10734# 2.97e-19
C517 X2.X2.X2.X1.X1.X1.vout a_52406_5016# 0.422f
C518 a_10686_15546# a_10686_13640# 0.00198f
C519 a_54992_11734# a_54992_9828# 0.00396f
C520 a_17222_9916# a_19422_9010# 4.2e-20
C521 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.X2.vin1 0.00117f
C522 a_2196_4198# a_2582_4198# 0.419f
C523 X2.X2.X2.X2.X2.X2.X3.vin2 vrefl 0.183f
C524 X1.X1.X1.X1.X1.X1.X3.vin2 a_2196_30882# 0.354f
C525 X1.X1.X1.X2.X1.X2.vrefh a_2582_13728# 8.22e-20
C526 a_16836_32788# a_16836_30882# 0.00396f
C527 X1.X1.X2.X1.X2.X1.X2.vin1 a_11072_13640# 0.197f
C528 a_4696_7064# a_5082_7064# 0.419f
C529 X1.X1.X1.X1.X1.X2.X3.vin2 a_5082_26164# 0.00846f
C530 a_4782_28070# X1.X1.X1.X3.vin1 1.64e-19
C531 X1.X2.X1.X2.X2.X2.X1.vin2 a_17222_4198# 8.88e-20
C532 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X1.X3.vin1 0.00117f
C533 X2.X1.X2.X2.X2.X1.X3.vin2 a_37766_27888# 0.267f
C534 a_25326_30794# a_25326_28888# 0.00198f
C535 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X3.vin2 0.161f
C536 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin1 0.52f
C537 X2.X1.X1.X2.X2.X2.vout a_33676_5198# 0.36f
C538 X1.X2.X1.X2.X2.X2.X3.vin1 a_19036_5198# 0.199f
C539 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin2 7.84e-19
C540 a_34362_7064# a_34062_5198# 5.55e-20
C541 X2.X1.X2.X2.X2.X2.vout a_37466_29834# 0.263f
C542 X2.X2.X1.X1.X2.X1.X3.vin2 a_46502_21352# 8.07e-19
C543 a_46116_13728# X2.X2.X1.X2.X1.X2.X2.vin1 1.78e-19
C544 a_19722_10916# X1.X2.X1.X2.X3.vin2 0.263f
C545 a_37766_8828# a_37466_6962# 5.55e-20
C546 X1.X2.X1.X1.X2.X2.vrefh X1.X1.X2.X2.X1.X2.vrefh 0.117f
C547 a_54606_25076# a_52406_24076# 4.77e-21
C548 X2.X2.X2.X3.vin1 a_52106_10734# 0.509f
C549 X2.X2.X3.vin2 X2.X2.X1.X2.X3.vin2 0.00254f
C550 a_37466_14586# X2.X1.X2.X1.X3.vin2 0.423f
C551 a_10686_7922# X1.X1.X2.X1.X1.X1.X3.vin2 8.07e-19
C552 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X1.X1.vin1 2.23e-19
C553 X1.X1.X2.X2.X2.X1.X2.vin1 a_11072_26982# 1.78e-19
C554 a_23126_31700# X1.X2.X2.X2.X3.vin2 9.7e-20
C555 X1.X1.X2.X1.X2.X1.X3.vin1 a_11072_11734# 0.354f
C556 a_16836_21352# a_16836_19446# 0.00396f
C557 X2.X2.X2.X1.X2.X1.X3.vin1 a_54992_11734# 0.354f
C558 X2.X2.X2.X1.X1.X2.X3.vin2 a_54992_9828# 0.354f
C559 a_25712_13640# X1.X2.X2.X1.X2.X1.X1.vin2 1.78e-19
C560 a_48702_20446# X2.X2.X1.X1.X2.X2.X3.vin2 0.277f
C561 X1.X2.X2.X3.vin1 a_23212_10734# 0.356f
C562 X1.X2.X3.vin2 X1.X2.X2.X1.X3.vin1 0.0361f
C563 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X3.vin1 0.206f
C564 a_22826_29834# a_23512_27888# 2.86e-19
C565 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X2.X1.vin2 0.668f
C566 a_33976_26164# X2.X1.X1.X1.X3.vin2 0.0927f
C567 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X2.vrefh 0.00118f
C568 a_23126_16452# a_23512_16452# 0.419f
C569 X1.X1.X2.X2.X1.X2.vrefh a_11072_21264# 0.118f
C570 a_52492_10734# a_52406_8828# 3.3e-19
C571 a_48702_24258# a_46502_23258# 4.77e-21
C572 a_25712_15546# a_25712_13640# 0.00396f
C573 X1.X2.X3.vin2 a_19722_14688# 2.04e-19
C574 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.vout 0.0857f
C575 X2.X1.X3.vin1 X2.X3.vin1 0.273f
C576 X1.X1.X1.X1.X2.vrefh a_2582_25164# 8.22e-20
C577 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X1.X1.vin2 0.242f
C578 a_54606_28888# a_54606_26982# 0.00198f
C579 a_40352_30794# a_40352_28888# 0.00396f
C580 a_33976_18540# a_34362_18540# 0.413f
C581 a_4696_18540# a_2582_17540# 5.36e-21
C582 a_25712_19358# X1.X2.X2.X2.vrefh 1.64e-19
C583 a_34062_20446# a_34362_18540# 4.41e-20
C584 X2.X1.X1.X1.X2.X2.X3.vin2 a_33976_18540# 0.00504f
C585 X2.X2.X2.X2.X2.X2.X1.vin2 a_54606_30794# 0.273f
C586 X2.X2.X2.vrefh X2.X3.vin2 4.75e-20
C587 a_34062_20446# X2.X1.X1.X1.X2.X2.X3.vin2 0.277f
C588 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X3.vin1 0.00117f
C589 X1.X2.X2.X1.X2.X2.X3.vin2 a_25326_15546# 7.84e-19
C590 X1.X2.X2.X1.X1.X2.X3.vin2 a_23126_8828# 0.277f
C591 a_54606_25076# X2.X2.X2.X2.X1.X2.X3.vin2 0.567f
C592 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X1.vin1 0.0689f
C593 X1.X2.X3.vin1 X1.X2.X2.X1.X1.X1.vout 5.53e-20
C594 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X2.vout 0.398f
C595 a_2582_19446# X1.X1.X1.X2.X1.X1.X1.vin1 8.22e-20
C596 a_19336_29936# a_17222_28976# 2.68e-20
C597 a_17222_15634# a_19336_14688# 2.95e-20
C598 a_4782_16634# X1.X1.X1.X2.X1.X1.X3.vin2 0.267f
C599 a_46502_11822# X2.X2.X1.X2.X2.X1.X1.vin1 8.22e-20
C600 a_23126_8828# a_23512_8828# 0.419f
C601 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 1.22e-19
C602 a_5082_18540# X1.X1.X1.X3.vin2 0.233f
C603 X2.X2.X2.X1.X3.vin2 X2.X2.X2.X1.X3.vin1 0.546f
C604 X2.X2.X2.X1.X2.X1.vout a_52492_10734# 1.64e-19
C605 a_46502_32788# X2.X2.X1.X1.X1.X1.X1.vin2 0.273f
C606 a_19722_26164# a_19036_24258# 2.97e-19
C607 X1.X1.X1.X1.X2.X1.vout a_4696_22312# 0.169f
C608 a_4782_24258# a_5082_22312# 4.19e-20
C609 a_19336_26164# a_19422_24258# 3.21e-19
C610 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X3.vin1 0.0174f
C611 a_4396_31882# a_4782_31882# 0.419f
C612 a_17222_32788# X1.X2.X1.X1.X1.X1.X2.vin1 8.88e-20
C613 a_2196_27070# a_2582_27070# 0.419f
C614 a_22826_29834# a_23212_29834# 0.419f
C615 a_31476_28976# X2.X1.X1.X1.X1.X2.X2.vin1 1.78e-19
C616 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 0.139f
C617 X1.X1.X1.X2.X1.X1.X1.vin2 a_2582_15634# 8.88e-20
C618 a_8572_22210# a_10686_21264# 2.95e-20
C619 a_11072_19358# X1.X1.X2.X2.vrefh 1.64e-19
C620 X1.X1.X3.vin2 a_8486_8828# 2.33e-19
C621 a_19422_20446# X1.X2.X1.X1.X2.X2.X3.vin2 0.277f
C622 X2.X2.X1.X1.X3.vin1 a_48616_26164# 0.169f
C623 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.vout 0.197f
C624 a_2582_32788# X1.X1.X1.X1.X1.X1.X2.vin1 8.88e-20
C625 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X1.vin2 0.076f
C626 X1.X2.X1.X2.X2.X2.vrefh a_16836_6104# 1.64e-19
C627 X2.X1.X2.X2.X1.X2.X1.vin1 a_40352_21264# 1.64e-19
C628 X2.vrefh X2.X1.X1.X1.X1.X1.X1.vin2 0.109f
C629 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 1.22e-19
C630 X1.X1.X1.X2.X2.X1.X3.vin2 X1.X1.X1.X2.X2.X2.vrefh 0.161f
C631 a_33976_26164# a_31862_25164# 5.36e-21
C632 X2.X1.X2.X2.X2.X1.vout a_38152_27888# 0.359f
C633 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.X1.X1.vin2 3.94e-19
C634 X1.X2.X2.X2.X1.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin2 0.0128f
C635 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X2.X1.X1.X2.vrefh 0.0128f
C636 a_46502_9916# a_46502_8010# 0.00198f
C637 a_11072_28888# X1.X1.X2.X2.X2.X1.X1.vin2 1.78e-19
C638 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X1.X3.vin2 0.546f
C639 a_39966_25076# X2.X1.X2.X2.X1.X2.X1.vin2 8.88e-20
C640 X1.X1.X1.X2.X2.vrefh a_2582_11822# 0.3f
C641 a_46116_11822# a_46502_11822# 0.419f
C642 a_22826_14586# X1.X2.X2.X1.X2.X1.vout 0.383f
C643 a_8872_12640# a_10686_11734# 1.06e-19
C644 a_37852_18358# a_39966_17452# 4.72e-20
C645 a_52792_12640# a_54606_11734# 1.06e-19
C646 a_37466_22210# a_37766_20264# 4.19e-20
C647 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin2 0.12f
C648 a_10686_32700# X1.X1.X2.X2.X2.X2.X2.vin1 0.402f
C649 a_16836_13728# a_16836_11822# 0.00396f
C650 X1.X1.X2.X2.X3.vin1 a_8186_22210# 0.436f
C651 a_25326_13640# X1.X2.X2.X1.X2.X1.X3.vin1 0.00207f
C652 a_10686_9828# a_8872_8828# 1.15e-20
C653 a_54606_21264# X2.X2.X2.X2.X1.X1.X2.vin1 0.402f
C654 a_52492_29834# a_54606_28888# 2.95e-20
C655 a_25326_28888# a_25712_28888# 0.419f
C656 a_39966_9828# X2.X1.X2.X1.X1.X2.X3.vin2 0.567f
C657 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.X1.vin2 0.22f
C658 X1.X2.X2.X2.X2.X1.X1.vin1 X2.X1.X1.X1.X2.vrefh 0.00437f
C659 X2.X2.X2.X1.X2.X1.X3.vin2 a_54992_13640# 0.354f
C660 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 0.581f
C661 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X1.vin2 0.1f
C662 X1.X2.X2.X1.X2.X1.X3.vin1 a_23212_10734# 0.00251f
C663 a_16836_28976# X1.X2.X1.X1.X1.X2.X3.vin1 0.354f
C664 X2.X2.X2.X1.X1.X1.vout a_52492_6962# 0.169f
C665 a_17222_28976# X1.X2.X1.X1.X1.X2.X1.vin1 0.417f
C666 a_19336_26164# X1.X2.X1.X3.vin1 0.356f
C667 a_17222_15634# X1.X2.X1.X2.X1.X2.X1.vin1 8.22e-20
C668 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X1.X2.X2.X1.X2.vrefh 0.1f
C669 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X1.X2.X2.X2.X2.vrefh 0.267f
C670 a_19336_7064# X1.X2.X1.X2.X2.X2.X3.vin1 0.00329f
C671 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X3.vin1 0.206f
C672 a_48316_24258# a_48702_24258# 0.419f
C673 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.vout 0.2f
C674 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 0.587f
C675 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.vout 0.197f
C676 X1.X2.X1.X1.X2.X1.X3.vin1 a_19036_24258# 0.199f
C677 X1.X1.X3.vin1 a_8186_14586# 2.24e-19
C678 a_37852_10734# X2.X1.X2.X1.X1.X2.X3.vin2 0.00535f
C679 a_33976_26164# a_33676_24258# 6.2e-19
C680 X2.X1.X3.vin1 a_37766_12640# 8.66e-20
C681 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X2.X3.vin2 8.93e-19
C682 a_31862_6104# a_31862_4198# 0.00198f
C683 X2.X2.X2.X1.X2.X2.X3.vin1 a_52792_16452# 0.199f
C684 a_49002_22312# X2.X2.X1.X1.X2.X2.X3.vin1 0.00874f
C685 a_31862_30882# X2.X1.X1.X1.X1.X2.X1.vin1 8.22e-20
C686 X2.X1.X2.X1.X1.X1.X3.vin2 a_37766_5016# 0.267f
C687 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X3.vin1 0.00117f
C688 X1.X2.X2.X1.X2.X1.X1.vin2 X1.X2.X2.X1.X2.vrefh 0.1f
C689 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X2.X1.X1.X2.X1.X1.vin2 0.00232f
C690 a_46116_25164# a_46502_25164# 0.419f
C691 a_23212_25982# X1.X2.X2.X2.X1.X2.vout 7.93e-20
C692 X1.X1.X2.X1.X1.X2.X2.vin1 a_10686_7922# 8.88e-20
C693 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.X1.vin2 8.93e-19
C694 X2.X2.X1.X2.X2.X1.X3.vin2 a_49002_7064# 0.00815f
C695 a_25326_32700# a_23126_31700# 4.77e-21
C696 a_5082_29936# X1.X1.X1.X1.X1.X2.X3.vin1 0.00874f
C697 a_19422_16634# a_19336_14688# 3.14e-19
C698 a_19036_16634# a_19722_14688# 2.86e-19
C699 X2.X2.X2.X2.X2.X1.X1.vin2 a_54992_26982# 0.12f
C700 a_5082_14688# a_4782_12822# 5.55e-20
C701 a_54606_26982# X2.X2.X2.X2.X2.X1.X1.vin1 0.417f
C702 X3.vin2 X2.X3.vin1 0.145f
C703 a_19722_10916# X1.X2.X1.X2.X2.X1.X3.vin2 3.49e-19
C704 a_54992_25076# a_54992_23170# 0.00396f
C705 X2.X1.X2.X2.X1.X1.vout a_37852_22210# 0.169f
C706 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X2.vin1 0.564f
C707 a_31862_8010# a_33976_7064# 2.95e-20
C708 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X2.X3.vin1 0.00836f
C709 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X1.vin2 0.076f
C710 a_8572_25982# a_8486_24076# 3.3e-19
C711 a_22826_18358# a_23512_16452# 3.08e-19
C712 X2.X1.X1.X1.X1.X1.vout X2.X1.X1.X1.X1.X2.vout 0.507f
C713 X1.X1.X2.X1.X2.X2.vout X1.X1.X2.X1.X3.vin2 0.0866f
C714 a_11072_11734# X1.X1.X2.X1.X2.vrefh 1.64e-19
C715 X1.X1.X1.X1.X1.X2.X2.vin1 X1.X1.X1.X1.X2.vrefh 0.564f
C716 X1.X1.X2.X1.X1.X2.vrefh a_10686_6016# 0.3f
C717 X1.X1.X2.X1.X1.X1.X3.vin2 a_10686_4110# 7.84e-19
C718 a_8486_27888# X1.X1.X2.X2.X2.X1.X3.vin1 0.428f
C719 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X1.vin1 0.0689f
C720 X2.X1.X1.X2.X1.X1.X2.vin1 X2.X1.X1.X2.X1.X2.vrefh 0.564f
C721 a_37766_16452# X2.X1.X2.X1.X2.X2.X3.vin1 0.42f
C722 a_4782_20446# a_5082_18540# 4.41e-20
C723 a_8186_29834# X1.X1.X2.X2.X3.vin2 0.422f
C724 X2.X2.X2.X1.X1.X2.X3.vin1 a_52792_8828# 0.199f
C725 X1.X1.X1.X1.X2.X2.X3.vin2 a_4696_18540# 0.00504f
C726 X1.X1.X2.X1.X1.X2.X3.vin1 a_8872_8828# 0.199f
C727 X2.X1.X2.X2.X3.vin2 a_37766_27888# 0.00101f
C728 a_31476_23258# X2.X1.X1.X1.X2.X2.X1.vin1 1.64e-19
C729 a_31862_23258# a_31862_21352# 0.00198f
C730 X2.X2.X3.vin1 a_49002_10916# 6.09e-19
C731 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X3.vin2 2.23e-19
C732 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X3.vin2 0.449f
C733 a_52492_14586# a_52792_12640# 6.1e-19
C734 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X1.X2.X1.X2.X1.X1.vin1 0.668f
C735 X1.X2.X2.X1.X2.X2.X1.vin1 a_25712_15546# 0.195f
C736 a_39966_26982# a_40352_26982# 0.419f
C737 a_19722_26164# X1.X2.X1.X1.X2.X1.X3.vin1 0.00837f
C738 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X2.vin1 0.0689f
C739 a_46502_9916# a_48316_9010# 1.06e-19
C740 a_2196_28976# a_2196_27070# 0.00396f
C741 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X2.X1.X2.vrefh 0.00437f
C742 X1.X2.X2.X1.X2.X2.vrefh a_25712_13640# 0.118f
C743 X2.X1.X1.X2.vrefh a_31862_17540# 8.22e-20
C744 X1.X2.X1.X1.X2.X2.X3.vin1 a_19422_20446# 0.42f
C745 X1.X1.X2.X2.X2.vrefh a_10686_25076# 0.3f
C746 X1.X2.X3.vin1 a_22826_10734# 3.93e-19
C747 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X3.vin2 0.17f
C748 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 2.23e-19
C749 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X3.vin1 0.199f
C750 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X2.X3.vin2 0.0565f
C751 X2.X1.X2.X3.vin2 a_37852_18358# 0.0927f
C752 X2.X2.X1.X2.X1.X2.X2.vin1 X2.X2.X1.X2.X2.vrefh 0.564f
C753 X2.X2.X2.X1.X1.X1.X3.vin2 a_54606_4110# 7.84e-19
C754 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X1.vin1 0.0689f
C755 a_54606_30794# a_54606_28888# 0.00198f
C756 a_52106_18358# X2.X2.X2.X3.vin1 0.374f
C757 X2.X2.X1.X3.vin2 X2.X2.X3.vin2 3.82e-19
C758 X2.X1.X1.X1.X2.X1.X3.vin2 a_33976_22312# 0.00546f
C759 a_37766_8828# X2.X1.X2.X1.X1.X2.X3.vin1 0.42f
C760 X2.X1.X1.X2.X2.X1.X2.vin1 X2.X1.X1.X2.X2.X2.vrefh 0.564f
C761 X2.X1.X2.X2.X2.X2.X2.vin1 a_39966_30794# 8.88e-20
C762 X2.X1.X2.X2.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X2.X1.vin2 8.93e-19
C763 X1.X2.X2.X1.X1.X2.X2.vin1 X2.X1.X1.X2.X2.X1.X1.vin2 0.00232f
C764 a_31476_9916# a_31862_9916# 0.419f
C765 X1.X1.X1.X1.X1.X1.X3.vin2 a_4696_29936# 0.00546f
C766 X1.X2.X2.X2.X2.X1.X1.vin2 X2.X1.X1.X1.X1.X2.X2.vin1 0.00232f
C767 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin2 0.12f
C768 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X3.vin1 0.587f
C769 X2.X2.X3.vin2 a_52406_16452# 3.98e-19
C770 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.X1.vin1 0.206f
C771 a_8572_10734# a_8872_8828# 6.48e-19
C772 X1.X2.X2.X1.X1.X2.X1.vin1 a_25712_7922# 0.195f
C773 a_37466_6962# X2.X1.X2.X1.X1.X1.vout 0.386f
C774 a_10686_13640# a_8486_12640# 4.77e-21
C775 a_39966_13640# X2.X1.X2.X1.X2.X1.X3.vin2 0.567f
C776 a_52406_16452# a_54606_15546# 4.2e-20
C777 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 0.216f
C778 X1.X1.X1.X2.X2.X1.X2.vin1 a_2582_8010# 0.402f
C779 X2.X1.X1.X3.vin2 a_34062_12822# 6.03e-19
C780 a_33676_16634# a_33976_14688# 6.1e-19
C781 X2.X1.X1.X2.X1.X2.X2.vin1 a_31862_11822# 0.402f
C782 X2.X1.X2.X1.X1.X2.X1.vin1 a_39966_6016# 8.22e-20
C783 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X1.X2.X1.X1.X1.X3.vin2 3.94e-19
C784 X2.X2.X3.vin2 a_52406_8828# 2.33e-19
C785 a_8186_6962# a_8572_6962# 0.419f
C786 a_31476_6104# X2.X1.X1.X2.X2.X2.X2.vin1 1.78e-19
C787 X1.X1.X1.X2.vrefh a_2196_17540# 1.64e-19
C788 X2.X2.X1.X1.X1.X1.X3.vin2 a_49002_29936# 0.00815f
C789 X1.X2.X2.X1.X2.X2.vout a_23212_14586# 0.0929f
C790 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin2 7.84e-19
C791 a_8186_6962# a_8872_5016# 2.86e-19
C792 X2.X2.X2.X1.X1.X1.X3.vin1 a_54992_4110# 0.354f
C793 X1.X2.X2.X1.X2.X1.X3.vin2 a_22826_10734# 3.49e-19
C794 X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X1.X3.vin1 0.0321f
C795 X2.X1.X2.X2.X1.X2.vrefh a_40352_21264# 0.118f
C796 a_54992_15546# a_54992_13640# 0.00396f
C797 a_54606_19358# X2.X2.X2.X1.X2.X2.X3.vin2 8.07e-19
C798 X1.X2.X1.X2.X1.X2.X3.vin2 a_17222_11822# 0.567f
C799 X1.X1.X2.X2.X2.X2.X2.vin1 a_11072_30794# 1.78e-19
C800 X1.X2.X1.X1.X1.X1.X3.vin2 X1.X2.X1.X1.X1.X2.X1.vin2 3.94e-19
C801 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.X1.vin1 2.23e-19
C802 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 0.216f
C803 a_52406_8828# a_54606_7922# 4.2e-20
C804 a_48616_14688# a_49002_14688# 0.419f
C805 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X2.vrefh 0.267f
C806 a_8486_16452# a_8572_14586# 3.38e-19
C807 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X2.vin1 0.00117f
C808 a_2582_17540# a_4782_16634# 4.2e-20
C809 a_52106_22210# a_52792_20264# 2.86e-19
C810 a_22826_22210# X1.X2.X2.X2.X1.X1.vout 0.387f
C811 a_34062_9010# a_33976_7064# 3.14e-19
C812 a_33676_9010# a_34362_7064# 2.86e-19
C813 X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X3.vin2 0.0011f
C814 a_52406_27888# a_52106_25982# 5.25e-20
C815 X2.X1.X2.X1.X1.X1.X3.vin1 a_40352_4110# 0.354f
C816 X2.X2.X3.vin2 X2.X2.X2.X1.X2.X1.vout 3.2e-19
C817 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin2 0.418f
C818 X2.X2.X2.X1.X2.X2.X3.vin2 a_54606_15546# 7.84e-19
C819 a_25712_26982# a_25712_25076# 0.00396f
C820 vrefl X2.X2.X2.X2.X2.X2.X1.vin2 0.0763f
C821 a_54606_9828# X2.X2.X2.X1.X1.X2.X3.vin1 0.00207f
C822 X2.X2.X1.X1.X2.X2.X3.vin2 a_46116_19446# 0.354f
C823 a_48702_20446# a_46502_19446# 4.77e-21
C824 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X1.vin1 0.0689f
C825 X2.X1.X1.X3.vin2 a_33976_10916# 0.355f
C826 a_19722_14688# X1.X2.X1.X2.X1.X2.vout 0.254f
C827 X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X1.vin2 0.096f
C828 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin1 0.267f
C829 X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 8.36e-19
C830 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X1.vout 0.0524f
C831 X2.X2.X2.X1.X2.X2.X3.vin1 a_52492_14586# 0.00329f
C832 X1.X1.X2.X2.X1.X2.X1.vin2 a_11072_23170# 0.12f
C833 a_10686_23170# X1.X1.X2.X2.X1.X2.X1.vin1 0.417f
C834 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X2.vin1 0.242f
C835 X2.X2.X1.X1.X2.X2.vrefh a_46116_23258# 0.118f
C836 X1.X2.X1.X1.X1.X2.vrefh a_17222_30882# 0.3f
C837 a_23512_31700# a_25326_30794# 1.06e-19
C838 X1.X1.X1.X3.vin1 a_5082_22312# 7.98e-19
C839 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X2.vrefh 0.076f
C840 X2.X1.X2.X1.X1.X2.X3.vin2 a_38152_8828# 0.101f
C841 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X3.vin2 0.102f
C842 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X1.X3.vin1 0.0425f
C843 X1.X1.X2.X2.X1.X2.vout a_8872_24076# 0.36f
C844 X2.X1.X1.X2.X1.X1.X1.vin2 a_31476_15634# 1.78e-19
C845 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X2.vrefh 0.267f
C846 a_25326_23170# a_23212_22210# 2.68e-20
C847 X1.X2.X2.X3.vin2 X1.X2.X3.vin2 0.171f
C848 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 1.22e-19
C849 a_33676_20446# a_31862_19446# 1.15e-20
C850 X2.X1.X3.vin1 X2.X1.X3.vin2 3.25f
C851 X2.X1.X1.X3.vin2 X2.X1.X2.X3.vin1 1.22e-19
C852 a_17222_27070# a_19336_26164# 4.72e-20
C853 a_38152_20264# a_37466_18358# 2.97e-19
C854 X2.X2.X1.X2.X2.X2.vrefh a_46116_6104# 1.64e-19
C855 X1.X2.X1.X1.X1.X1.X2.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 0.234f
C856 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.vout 0.118f
C857 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X3.vin2 0.0523f
C858 a_52492_22210# X2.X2.X2.X2.X1.X1.X3.vin2 0.00546f
C859 X1.X2.X2.X2.X1.X1.X3.vin2 a_25712_21264# 0.354f
C860 X1.X2.X1.X2.X2.X1.X3.vin1 a_17222_8010# 0.00207f
C861 a_31476_13728# a_31862_13728# 0.419f
C862 X1.X1.X2.X1.X2.X2.X3.vin1 a_10686_15546# 0.52f
C863 X1.X2.X2.X1.X2.X1.X2.vin1 X2.X1.X1.X2.X1.X2.X1.vin2 0.00232f
C864 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X1.vin1 0.0689f
C865 X1.X1.X2.X2.X1.X2.X3.vin2 a_10686_23170# 7.84e-19
C866 X1.X1.X1.X1.X1.X1.X2.vin1 a_2582_30882# 0.402f
C867 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X3.vin1 0.206f
C868 a_19036_24258# a_19336_22312# 6.1e-19
C869 a_37766_12640# a_38152_12640# 0.419f
C870 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X1.X3.vin2 1.22e-19
C871 X1.X1.X1.X2.X1.X1.X2.vin1 a_2196_15634# 0.197f
C872 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X2.vrefh 0.00118f
C873 a_40352_28888# a_40352_26982# 0.00396f
C874 a_4782_12822# a_4696_10916# 3.3e-19
C875 X2.X2.X1.X1.X1.X1.X3.vin2 a_46502_30882# 0.567f
C876 a_4396_12822# a_5082_10916# 3.08e-19
C877 a_8486_27888# X1.X1.X2.X3.vin2 7.93e-20
C878 X1.X1.X2.X2.X2.X1.vout X1.X1.X2.X2.X2.X1.X3.vin2 0.326f
C879 X2.X1.X3.vin1 a_37766_16452# 8.66e-20
C880 X1.X1.X2.X2.X1.X2.vout a_8186_22210# 0.254f
C881 X1.X1.X1.X2.X1.X1.X3.vin2 a_2582_13728# 8.07e-19
C882 a_52792_5016# a_54606_4110# 1.06e-19
C883 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X3.vin2 0.161f
C884 a_16836_17540# X1.X2.X1.X2.X1.X1.X2.vin1 1.78e-19
C885 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X1.X3.vin2 0.0943f
C886 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X2.vrefh 0.267f
C887 X2.X2.X1.X2.X1.X2.X3.vin1 a_46502_11822# 0.00207f
C888 a_19036_20446# a_17222_19446# 1.15e-20
C889 a_17222_25164# X1.X2.X1.X1.X2.X1.X1.vin2 0.273f
C890 a_8486_8828# a_8186_6962# 5.55e-20
C891 a_11072_32700# X1.X1.X2.X2.X2.X2.X1.vin2 1.78e-19
C892 a_5082_22312# X1.X1.X1.X1.X2.X2.X3.vin1 0.00874f
C893 X1.X2.X1.X2.X1.X2.vout X1.X2.X1.X2.X1.X2.X3.vin1 0.326f
C894 X2.X1.X1.X1.X2.X2.X3.vin1 a_31862_19446# 0.00207f
C895 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X3.vin1 0.00117f
C896 X1.X1.X2.X1.X2.X2.X3.vin2 a_8486_16452# 0.277f
C897 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X3.vin2 0.234f
C898 X2.X1.X3.vin1 a_37766_8828# 8.66e-20
C899 a_46502_15634# X2.X2.X1.X2.X1.X2.X1.vin1 8.22e-20
C900 X1.X1.X2.X2.X2.X2.X2.vin1 a_8872_31700# 5.34e-19
C901 a_31862_17540# X2.X1.X1.X2.X1.X1.X1.vin2 0.273f
C902 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X2.vrefh 0.267f
C903 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X1.X3.vin2 0.0943f
C904 a_19036_12822# a_19422_12822# 0.419f
C905 X1.X2.X1.X2.X1.X2.X2.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 0.234f
C906 a_46502_25164# a_48702_24258# 4.2e-20
C907 a_19422_24258# a_17222_23258# 4.77e-21
C908 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X2.vin1 0.00117f
C909 a_31476_4198# a_31862_4198# 0.419f
C910 X2.X1.X2.X1.X1.X1.X3.vin2 a_40352_6016# 0.354f
C911 a_48702_28070# X2.X2.X1.X1.X1.X2.X3.vin2 0.277f
C912 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 0.234f
C913 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 0.0565f
C914 a_38152_5016# a_39966_4110# 1.06e-19
C915 X2.X1.X2.vrefh a_31862_4198# 0.301f
C916 a_54606_28888# X2.X2.X2.X2.X2.X1.X2.vin1 0.402f
C917 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X3.vin1 0.206f
C918 X1.X2.X2.X2.X2.X2.X1.vin1 X2.X1.X1.X1.X1.X2.vrefh 0.00437f
C919 a_52106_6962# X2.X2.X2.X1.X1.X1.X3.vin2 0.00815f
C920 a_17222_27070# X1.X2.X1.X1.X2.X1.X1.vin1 8.22e-20
C921 X2.X1.X2.X1.X2.X1.X3.vin1 a_37466_10734# 0.00837f
C922 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X1.vout 0.038f
C923 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X1.X1.vin2 0.216f
C924 a_49566_892# a_49952_892# 0.406f
C925 a_37766_27888# a_39966_26982# 4.2e-20
C926 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 0.587f
C927 X1.X1.X1.X2.X2.X2.X2.vin1 a_2582_4198# 0.402f
C928 a_4782_12822# X1.X1.X1.X2.X1.X2.X3.vin2 0.277f
C929 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 0.242f
C930 a_39966_9828# a_39966_7922# 0.00198f
C931 X1.X1.X1.X1.X2.X2.vrefh a_2196_23258# 0.118f
C932 a_5082_14688# X1.X1.X1.X2.X3.vin1 0.436f
C933 X1.X1.X2.X2.X1.X1.X2.vin1 a_11072_19358# 1.78e-19
C934 X1.X1.X2.X2.X1.X1.X3.vin2 X1.X1.X2.X2.X1.X1.X1.vin1 2.23e-19
C935 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 0.581f
C936 a_49002_18540# X2.X2.X1.X3.vin2 0.233f
C937 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X2.vrefh 0.267f
C938 X2.X2.X1.X1.X2.X1.X2.vin1 X2.X2.X1.X1.X2.X2.vrefh 0.564f
C939 X1.X1.X1.X2.X2.vrefh a_2582_9916# 8.22e-20
C940 X2.X1.X1.X2.vrefh X1.X2.X2.X2.vrefh 0.117f
C941 X1.X2.X1.X2.X1.X2.X3.vin2 a_19722_10916# 0.00846f
C942 X1.X1.X1.X1.X1.X1.X1.vin2 vrefh 0.0964f
C943 X2.X1.X2.X1.X1.X2.vrefh a_39966_6016# 0.3f
C944 a_39966_23170# a_40352_23170# 0.419f
C945 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X2.X1.X1.X1.X1.X2.vin1 0.00232f
C946 X1.X2.X2.X2.X2.X1.X3.vin1 a_25712_26982# 0.354f
C947 X1.X1.X2.X3.vin2 X1.X1.X2.X3.vin1 0.559f
C948 X1.X2.X3.vin1 X1.X2.X2.X3.vin1 3.45e-19
C949 a_10686_15546# X1.X1.X2.X1.X2.X1.X3.vin2 8.07e-19
C950 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin2 0.12f
C951 a_2582_9916# X1.X1.X1.X2.X2.X1.X1.vin2 0.273f
C952 a_33976_10916# a_33676_9010# 6.2e-19
C953 X1.X2.X1.X2.X2.X1.X3.vin1 a_19422_9010# 0.428f
C954 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 0.0565f
C955 a_10686_25076# a_8872_24076# 1.15e-20
C956 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X3.vin1 2.33e-19
C957 a_10686_21264# X1.X1.X2.X2.X1.X1.X3.vin2 0.567f
C958 a_49002_14688# X2.X2.X1.X2.X1.X2.X3.vin1 0.00874f
C959 X2.X2.X2.X1.X1.X2.vout a_52492_6962# 0.0929f
C960 a_17222_32788# a_17222_30882# 0.00198f
C961 a_19336_10916# a_17222_9916# 5.36e-21
C962 a_5082_7064# X1.X1.X1.X2.X2.X2.vout 0.263f
C963 a_8186_14586# a_8872_12640# 2.86e-19
C964 a_48316_31882# X2.X2.X1.X1.X1.X1.X3.vin2 0.1f
C965 a_23212_10734# X1.X2.X2.X1.X1.X2.vout 7.93e-20
C966 a_25326_30794# X1.X2.X2.X2.X2.X1.X3.vin2 8.07e-19
C967 X1.X2.X1.X2.vrefh X1.X1.X2.X2.vrefh 0.117f
C968 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X1.X3.vin1 0.0425f
C969 X2.X1.X3.vin1 X2.X1.X2.vrefh 0.178f
C970 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X2.vrefh 0.076f
C971 X1.X1.X2.X2.X2.X2.vrefh X1.X2.X1.X1.X1.X2.X1.vin1 0.00437f
C972 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 0.587f
C973 X2.X1.X1.X2.X2.X2.vout X2.X1.X1.X2.X2.X2.X3.vin2 0.08f
C974 a_46502_13728# a_48316_12822# 1.06e-19
C975 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X3.vin1 1.22e-19
C976 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X2.vin1 0.0689f
C977 X2.X1.X3.vin2 X3.vin2 0.00486f
C978 X2.X1.X2.X2.X2.X1.X1.vin1 a_39966_25076# 8.22e-20
C979 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X1.X2.X3.vin2 3.94e-19
C980 X3.vin1 X3.vin2 0.514f
C981 a_19336_29936# a_19722_29936# 0.419f
C982 a_8872_20264# a_8186_18358# 2.97e-19
C983 X3.vin1 a_20672_892# 5.96e-19
C984 X2.X2.X2.X2.X1.X2.X3.vin2 a_52406_24076# 0.277f
C985 X2.X1.X2.X2.X2.X2.X3.vin1 a_39966_30794# 0.52f
C986 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X3.vin1 0.00117f
C987 a_2196_32788# a_2196_30882# 0.00396f
C988 a_54606_23170# a_52492_22210# 2.68e-20
C989 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X1.vin2 3.94e-19
C990 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin1 0.195f
C991 X2.X1.X1.X1.X1.X1.X2.vin1 a_31476_30882# 0.197f
C992 X2.X1.X2.X2.X2.X2.vout a_38152_31700# 0.36f
C993 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X1.X3.vin1 0.00789f
C994 X2.X1.X1.X1.X1.X2.vout a_33676_28070# 0.36f
C995 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 0.0903f
C996 X2.X2.X1.X2.X3.vin2 a_49002_7064# 0.422f
C997 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin2 0.12f
C998 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X1.X2.X2.X1.X2.vrefh 0.1f
C999 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin1 0.195f
C1000 X2.X2.X3.vin1 a_52106_14586# 2.24e-19
C1001 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X2.vout 0.197f
C1002 a_19036_24258# X1.X2.X1.X1.X2.X1.vout 0.359f
C1003 X2.X1.X2.X2.X1.X1.vout a_37852_18358# 1.64e-19
C1004 X1.X2.vrefh X1.X2.X1.X1.X1.X1.X1.vin1 0.108f
C1005 a_8486_20264# a_8872_20264# 0.419f
C1006 a_17222_21352# a_17222_19446# 0.00198f
C1007 a_25326_6016# X1.X2.X2.X1.X1.X1.X3.vin2 0.567f
C1008 X1.X2.X2.X2.X1.X2.X1.vin2 X1.X2.X2.X2.X1.X1.X3.vin2 3.94e-19
C1009 X1.X2.X2.X2.X1.X2.X1.vin1 a_25326_21264# 8.22e-20
C1010 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.vrefh 2.33e-19
C1011 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X3.vin2 0.418f
C1012 a_38152_24076# a_37466_22210# 3.31e-19
C1013 a_46502_32788# X2.X2.X1.X1.X1.X1.X2.vin1 8.88e-20
C1014 a_11072_21264# X1.X1.X2.X2.X1.X1.X1.vin2 1.78e-19
C1015 a_33676_28070# a_33976_26164# 6.48e-19
C1016 X2.X2.X3.vin2 a_52106_6962# 0.00111f
C1017 X1.X1.X2.X2.X2.X2.vout a_8186_29834# 0.263f
C1018 a_23126_31700# X1.X2.X2.X2.X2.X2.vout 0.418f
C1019 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.vout 0.08f
C1020 X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X2.X1.X3.vin1 2.33e-19
C1021 X1.X1.X2.X2.X2.X1.X3.vin1 X1.X1.X2.X2.X1.X2.X3.vin2 1.22e-19
C1022 a_8186_25982# a_8572_25982# 0.414f
C1023 X1.X2.X1.X2.X2.X2.X2.vin1 a_16836_4198# 0.197f
C1024 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X1.X1.vin1 0.0689f
C1025 X2.X2.X2.X2.X2.X1.X3.vin2 a_54606_26982# 7.84e-19
C1026 X1.X2.X1.X2.X1.X2.vrefh a_16836_13728# 1.64e-19
C1027 X1.X2.X1.X2.X2.X2.X2.vin1 X1.X2.X2.vrefh 0.564f
C1028 a_23126_5016# X1.X2.X2.X1.X1.X1.X3.vin1 0.428f
C1029 a_34362_18540# X2.X1.X3.vin1 0.47f
C1030 a_4696_18540# X1.X1.X1.X2.X1.X1.X3.vin1 0.00232f
C1031 a_23212_14586# a_23512_12640# 6.1e-19
C1032 X2.X2.X2.X2.X2.X2.X1.vin2 a_54992_30794# 0.12f
C1033 X1.X2.X2.X2.X1.X2.X3.vin1 a_22826_22210# 0.00874f
C1034 a_54606_30794# X2.X2.X2.X2.X2.X2.X1.vin1 0.417f
C1035 X1.X2.X1.X1.X2.vrefh a_17222_27070# 0.3f
C1036 a_23512_27888# a_25326_26982# 1.06e-19
C1037 X1.X1.X2.X1.X2.X1.X3.vin1 a_8572_10734# 0.00251f
C1038 a_52106_29834# X2.X2.X2.X2.X3.vin2 0.422f
C1039 a_52106_6962# a_52792_5016# 2.86e-19
C1040 X2.X1.X1.X1.X1.X2.vrefh a_31476_28976# 1.64e-19
C1041 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X2.vin1 0.242f
C1042 X2.X2.X2.X2.X2.X2.vout X2.X2.X2.X2.X2.X1.vout 0.514f
C1043 a_19336_29936# X1.X2.X1.X1.X1.X2.X3.vin1 0.00329f
C1044 a_54992_32700# vrefl 0.118f
C1045 X2.X2.X1.X1.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X1.X1.vin2 0.23f
C1046 a_2196_21352# a_2582_21352# 0.419f
C1047 X1.X2.X1.X3.vin1 a_19422_24258# 5.28e-19
C1048 X1.X1.X1.X1.X2.X1.vout X1.X1.X1.X1.X2.X2.vout 0.514f
C1049 X2.X1.X2.X2.X2.vrefh a_40352_25076# 0.118f
C1050 a_2582_13728# X1.X1.X1.X2.X1.X2.X1.vin2 0.273f
C1051 a_4782_31882# X1.X1.X1.X1.X1.X1.vout 0.422f
C1052 a_17222_32788# a_19422_31882# 4.2e-20
C1053 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.X2.vin1 0.00117f
C1054 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X2.X2.vin1 0.0689f
C1055 a_31862_28976# a_33676_28070# 1.06e-19
C1056 X2.X2.X1.X1.X1.X2.vout a_48702_28070# 0.418f
C1057 X2.X1.X1.X2.X1.X2.vrefh a_31862_15634# 0.3f
C1058 a_38152_16452# a_39966_15546# 1.06e-19
C1059 X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.vrefh 0.117f
C1060 a_8572_22210# X1.X1.X2.X2.X1.X1.X3.vin2 0.00546f
C1061 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X3.vin1 0.199f
C1062 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.X2.vin1 0.00117f
C1063 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin1 0.267f
C1064 X2.X1.X2.X2.vrefh a_39966_17452# 0.3f
C1065 a_33976_26164# X2.X1.X1.X1.X2.X1.X3.vin1 0.00251f
C1066 a_46116_19446# a_46502_19446# 0.419f
C1067 X2.X1.X1.X2.X1.X1.X2.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 0.234f
C1068 X1.X3.vin1 a_13696_892# 0.195f
C1069 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X2.X1.X1.X2.vrefh 0.00437f
C1070 X2.X2.X1.X2.X2.X1.X3.vin1 a_46502_8010# 0.00207f
C1071 a_48702_28070# a_48616_26164# 3.3e-19
C1072 X1.X2.X2.X2.X3.vin2 a_22826_25982# 0.263f
C1073 X2.X1.X2.X3.vin1 a_37852_10734# 0.356f
C1074 X2.X1.X3.vin2 X2.X1.X2.X1.X3.vin1 0.0361f
C1075 a_48316_28070# a_49002_26164# 3.08e-19
C1076 X2.X1.X2.X2.X1.X2.X2.vin1 a_39966_23170# 8.88e-20
C1077 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X1.vin2 8.93e-19
C1078 a_23512_31700# a_22826_29834# 3.31e-19
C1079 X1.X1.X1.X2.X3.vin1 a_4696_10916# 0.17f
C1080 a_37852_18358# X2.X1.X2.X1.X2.X2.X3.vin2 0.00517f
C1081 X1.X2.X2.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin2 0.0128f
C1082 X2.X1.X2.X2.X1.X1.vout X2.X1.X2.X2.X1.X1.X3.vin1 0.118f
C1083 X1.X1.X2.X1.X2.vrefh a_10686_9828# 0.3f
C1084 a_54606_32700# a_52406_31700# 4.77e-21
C1085 X2.X1.X2.vrefh X3.vin2 3.04e-19
C1086 a_23126_16452# a_25326_15546# 4.2e-20
C1087 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 0.216f
C1088 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X3.vin2 0.237f
C1089 a_17222_13728# a_17222_11822# 0.00198f
C1090 a_16836_6104# a_17222_6104# 0.419f
C1091 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X1.vin2 0.668f
C1092 X2.X1.X1.X2.X2.X2.vrefh a_31862_8010# 0.3f
C1093 a_38152_8828# a_39966_7922# 1.06e-19
C1094 X1.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X1.X3.vin1 0.0321f
C1095 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X2.X1.X2.X2.X2.X1.vin2 0.00232f
C1096 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X3.vin1 0.449f
C1097 X1.X2.X2.X1.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X3.vin1 0.581f
C1098 X2.X1.X3.vin1 X2.X1.X1.X2.X1.X2.vout 3.08e-19
C1099 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X2.vrefh 0.00118f
C1100 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X2.vrefh 0.076f
C1101 X1.X1.X2.X1.X1.X2.X3.vin2 a_8872_8828# 0.101f
C1102 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X3.vin2 0.234f
C1103 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X1.X2.X1.X2.vrefh 0.1f
C1104 a_52492_29834# X2.X2.X2.X2.X2.X1.X3.vin2 0.00546f
C1105 X1.X2.X2.X2.X2.X1.X3.vin2 a_25712_28888# 0.354f
C1106 a_52106_10734# a_52792_8828# 3.08e-19
C1107 X1.X1.X1.X2.X3.vin2 a_4696_7064# 0.363f
C1108 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X2.X3.vin1 0.206f
C1109 X1.X2.X1.X1.X2.X1.X1.vin2 a_16836_23258# 1.78e-19
C1110 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X2.vrefh 0.267f
C1111 X2.X1.X1.X1.X3.vin2 a_34062_20446# 9.7e-20
C1112 a_2196_21352# a_2196_19446# 0.00396f
C1113 X1.X2.X1.X2.X2.X2.vout X1.X2.X1.X2.X2.X2.X3.vin1 0.335f
C1114 X2.X1.X1.X2.X2.X1.X2.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 0.234f
C1115 a_48702_24258# X2.X2.X1.X1.X2.X1.vout 0.422f
C1116 X1.X1.X2.X1.X2.X2.vrefh a_10686_13640# 0.3f
C1117 a_46116_15634# a_46502_15634# 0.419f
C1118 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.vout 0.118f
C1119 X2.X1.X3.vin1 X2.X1.X2.X1.X1.X1.vout 5.53e-20
C1120 a_8186_6962# X1.X1.X2.X1.X1.X1.X3.vin2 0.00815f
C1121 a_23126_27888# a_22826_25982# 5.25e-20
C1122 X2.X1.X1.X2.X3.vin2 a_34062_5198# 9.7e-20
C1123 a_33976_26164# X2.X1.X1.X1.X2.X1.vout 1.64e-19
C1124 a_34362_26164# a_34062_24258# 5.25e-20
C1125 a_54606_25076# a_54992_25076# 0.419f
C1126 X2.X1.X1.X2.X2.X2.X3.vin1 a_31862_4198# 0.00207f
C1127 X2.X1.X2.X1.X3.vin1 a_37766_8828# 9.54e-19
C1128 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X2.vrefh 0.267f
C1129 X2.X2.X2.X1.X2.X1.vout X2.X2.X2.X1.X2.X1.X3.vin2 0.326f
C1130 a_46502_25164# X2.X2.X1.X1.X2.X1.X1.vin1 0.417f
C1131 a_46116_25164# X2.X2.X1.X1.X2.X1.X3.vin1 0.354f
C1132 a_23126_8828# a_25326_7922# 4.2e-20
C1133 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 0.216f
C1134 a_52406_31700# X2.X2.X2.X2.X3.vin2 9.7e-20
C1135 X1.X2.X2.X2.X2.X2.vrefh a_25326_28888# 0.3f
C1136 X2.X1.X2.X2.X1.X1.vout X2.X1.X2.X2.X1.X1.X3.vin2 0.342f
C1137 a_23126_27888# X1.X2.X2.X2.X2.X1.X3.vin1 0.428f
C1138 X1.X2.X1.X1.X1.X2.X2.vin1 X1.X2.X1.X1.X2.vrefh 0.564f
C1139 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.vout 0.335f
C1140 a_33976_22312# a_31862_21352# 2.68e-20
C1141 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.vrefh 0.161f
C1142 X1.X2.X2.X2.X1.X1.X3.vin1 a_23212_18358# 0.00255f
C1143 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.X1.vin1 2.23e-19
C1144 X1.X1.X2.X1.X1.X2.X2.vin1 a_11072_7922# 1.78e-19
C1145 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X3.vin1 0.00117f
C1146 a_37466_29834# X2.X1.X2.X2.X2.X1.vout 0.383f
C1147 a_48616_10916# X2.X2.X1.X2.X3.vin2 0.0927f
C1148 X1.X2.X2.X2.X2.X2.X3.vin2 a_23126_31700# 0.277f
C1149 X1.X2.X2.X1.X2.X1.X1.vin2 a_25326_11734# 0.273f
C1150 a_54606_21264# a_52406_20264# 4.77e-21
C1151 X1.X2.X1.X2.X1.X1.vout a_19722_14688# 0.387f
C1152 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X3.vin2 0.102f
C1153 a_5082_7064# a_4396_5198# 3.31e-19
C1154 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 0.0565f
C1155 a_19422_16634# X1.X2.X1.X2.X3.vin1 1.52e-19
C1156 a_4696_7064# a_4782_5198# 3.38e-19
C1157 X2.X2.X2.X2.X2.X1.X1.vin1 a_54992_26982# 0.195f
C1158 a_46116_8010# a_46502_8010# 0.419f
C1159 a_4782_9010# a_4696_7064# 3.14e-19
C1160 a_4396_9010# a_5082_7064# 2.86e-19
C1161 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X3.vin1 0.00118f
C1162 X1.X1.X2.X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X3.vin2 0.165f
C1163 a_39966_13640# a_39966_11734# 0.00198f
C1164 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 0.242f
C1165 a_4696_26164# a_4396_24258# 6.2e-19
C1166 a_49002_22312# a_48316_20446# 3.31e-19
C1167 a_48616_22312# a_48702_20446# 3.38e-19
C1168 a_10686_11734# a_11072_11734# 0.419f
C1169 a_25712_11734# a_25712_9828# 0.00396f
C1170 a_52406_24076# a_52106_22210# 5.55e-20
C1171 X1.X2.X2.X1.X2.X2.X1.vin2 X2.X1.X1.X2.X1.X1.X2.vin1 0.00232f
C1172 X2.X1.X2.X1.X2.X2.X1.vin1 a_39966_13640# 8.22e-20
C1173 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X1.X2.X1.X2.X1.X3.vin2 3.94e-19
C1174 X1.X2.X2.X2.X3.vin1 a_22826_22210# 0.436f
C1175 X2.X2.X1.X2.X2.X1.X3.vin1 a_48316_9010# 0.199f
C1176 a_2582_28976# a_2582_27070# 0.00198f
C1177 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X3.vin2 0.102f
C1178 X1.X1.X1.X2.X1.X2.X2.vin1 a_2582_11822# 0.402f
C1179 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 1.22e-19
C1180 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X3.vin1 2.33e-19
C1181 X1.X1.X2.X1.X3.vin2 a_8572_14586# 0.363f
C1182 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X3.vin2 0.161f
C1183 X2.X2.X1.X2.X1.X2.X2.vin1 a_46502_11822# 0.402f
C1184 a_52406_20264# a_52106_18358# 5.25e-20
C1185 a_25326_13640# a_23512_12640# 1.15e-20
C1186 X2.X1.X2.X2.X2.X1.X3.vin1 a_37466_25982# 0.00837f
C1187 a_48616_26164# a_48702_24258# 3.21e-19
C1188 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.X3.vin1 0.00789f
C1189 a_49002_26164# a_48316_24258# 2.97e-19
C1190 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin1 0.195f
C1191 a_54606_30794# X2.X2.X2.X2.X2.X1.X3.vin2 8.07e-19
C1192 a_39966_9828# a_40352_9828# 0.419f
C1193 X1.X2.X1.X1.X1.X1.X3.vin2 a_17222_30882# 0.567f
C1194 a_17222_13728# X1.X2.X1.X2.X1.X2.X2.vin1 8.88e-20
C1195 X2.X1.X2.X2.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X2.X1.vin1 2.23e-19
C1196 X2.X1.X2.X2.X2.X2.X2.vin1 a_40352_30794# 1.78e-19
C1197 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin1 0.195f
C1198 a_10686_26982# a_10686_25076# 0.00198f
C1199 X2.X1.X2.X2.X2.X2.vrefh X2.X2.X1.X1.X1.X2.X1.vin1 0.00437f
C1200 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X3.vin2 8.93e-19
C1201 a_23512_12640# a_23212_10734# 6.2e-19
C1202 a_31862_9916# X2.X1.X1.X2.X2.X1.X1.vin1 0.417f
C1203 a_31476_9916# X2.X1.X1.X2.X2.X1.X3.vin1 0.354f
C1204 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin2 0.12f
C1205 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X1.vin2 0.668f
C1206 X1.X1.X1.X1.X1.X1.vout X1.X1.X1.X1.X1.X2.vout 0.507f
C1207 X1.X2.X3.vin1 X1.X2.X1.X2.X3.vin1 7.18e-19
C1208 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X3.vin2 8.93e-19
C1209 a_8186_18358# X1.X1.X2.X1.X2.X2.X3.vin2 0.00846f
C1210 a_10686_28888# X1.X1.X2.X2.X2.X1.X3.vin2 0.567f
C1211 X1.X1.X2.X1.X2.X1.X3.vin2 a_8486_12640# 0.267f
C1212 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X3.vin1 0.00117f
C1213 X1.X2.X2.X1.X1.X2.X1.vin2 X2.X1.X1.X2.X2.X1.X2.vin1 0.00232f
C1214 a_4782_9010# a_2582_8010# 4.77e-21
C1215 X1.X2.X1.X3.vin1 a_19336_18540# 0.17f
C1216 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X1.vin1 0.206f
C1217 a_10686_6016# X1.X1.X2.X1.X1.X1.X3.vin1 0.00207f
C1218 a_34062_16634# a_34362_14688# 4.19e-20
C1219 X2.X1.X1.X2.X1.X1.vout a_33976_14688# 0.169f
C1220 a_34062_12822# a_31862_11822# 4.77e-21
C1221 X2.X1.X1.X2.X1.X2.X3.vin2 a_31476_11822# 0.354f
C1222 X2.X2.X2.X1.X2.X2.vout a_52792_16452# 0.36f
C1223 X2.X2.X1.X2.X1.X1.X2.vin1 a_46502_15634# 0.402f
C1224 X1.X1.X2.X2.X1.X1.vout a_8486_20264# 0.422f
C1225 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X1.X3.vin2 5.19e-19
C1226 a_22826_29834# X1.X2.X2.X2.X2.X1.X3.vin2 0.00815f
C1227 X2.X2.X2.X2.X1.X2.X3.vin2 a_52106_22210# 3.85e-19
C1228 a_31862_6104# a_33676_5198# 1.06e-19
C1229 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X2.vin1 0.0689f
C1230 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X1.vin1 0.267f
C1231 X2.X1.X3.vin2 X2.X1.X2.X1.X2.X2.vout 3.38e-19
C1232 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 0.581f
C1233 X2.X1.X2.X2.X1.X2.X3.vin1 a_38152_24076# 0.199f
C1234 a_11072_9828# X1.X1.X2.X1.X1.X2.X1.vin2 1.78e-19
C1235 X2.X2.X2.X2.X1.X2.X1.vin2 X2.X2.X2.X2.X1.X1.X3.vin2 3.94e-19
C1236 X2.X2.X2.X2.X1.X2.X1.vin1 a_54606_21264# 8.22e-20
C1237 X1.X2.X2.X2.X1.X2.X1.vin2 X2.X1.X1.X1.X2.X2.vrefh 0.0128f
C1238 X1.X1.X1.X2.X2.X2.X3.vin2 X1.X1.X2.vrefh 0.172f
C1239 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.X1.X1.vin1 5.19e-19
C1240 X1.X1.X1.X1.X3.vin2 a_4782_20446# 9.7e-20
C1241 a_23212_14586# a_25326_13640# 2.95e-20
C1242 X1.X2.X1.X1.X3.vin1 X1.X2.X2.X2.X3.vin2 0.0604f
C1243 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X2.vout 0.0898f
C1244 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X1.X1.vin2 0.242f
C1245 a_25326_28888# a_25326_26982# 0.00198f
C1246 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.X1.vin1 0.206f
C1247 a_49002_14688# X2.X2.X1.X2.X3.vin1 0.436f
C1248 a_37466_25982# X2.X1.X2.X2.X1.X2.X3.vin2 0.00846f
C1249 a_8486_27888# a_8872_27888# 0.419f
C1250 a_37766_16452# X2.X1.X2.X1.X2.X2.vout 0.418f
C1251 X1.X1.X1.X2.X1.X1.X3.vin1 a_4782_16634# 0.428f
C1252 X2.X1.X2.X2.X2.X2.vrefh X2.X1.X2.X2.X2.X1.X3.vin1 0.00118f
C1253 X2.X2.X2.X1.X1.X2.vout a_52792_8828# 0.36f
C1254 X2.X1.X1.X2.X2.X1.vout a_34362_7064# 0.383f
C1255 X2.X2.X1.X2.X2.X1.X2.vin1 a_46502_8010# 0.402f
C1256 X2.X2.X1.X2.X1.X2.vrefh a_46116_13728# 1.64e-19
C1257 a_4696_10916# a_5082_10916# 0.414f
C1258 X1.X2.X3.vin2 X1.X3.vin2 0.147f
C1259 X1.X1.X2.X1.X1.X2.vout a_8872_8828# 0.36f
C1260 a_4396_16634# a_4696_14688# 6.1e-19
C1261 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X3.vin1 0.00118f
C1262 a_22826_6962# a_23126_5016# 4.19e-20
C1263 X1.X2.X1.X1.X2.X1.X2.vin1 X1.X2.X1.X1.X2.X2.vrefh 0.564f
C1264 a_23126_24076# X1.X2.X2.X2.X1.X2.X3.vin1 0.42f
C1265 a_54992_32700# a_54992_30794# 0.00396f
C1266 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X3.vin1 0.587f
C1267 a_17222_11822# X1.X2.X1.X2.X2.X1.X1.vin1 8.22e-20
C1268 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X3.vin2 0.17f
C1269 a_31862_11822# a_33976_10916# 4.72e-20
C1270 a_48616_14688# a_48316_12822# 6.71e-19
C1271 X2.X1.X3.vin1 a_37466_10734# 3.93e-19
C1272 X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X1.vin1 0.142f
C1273 X2.X2.X2.X3.vin2 X2.X2.X2.X3.vin1 0.559f
C1274 a_52492_25982# X2.X2.X2.X2.X1.X2.vout 7.93e-20
C1275 X1.X1.X2.X2.X1.X2.X1.vin1 a_11072_23170# 0.195f
C1276 a_52792_24076# a_54606_23170# 1.06e-19
C1277 a_48316_16634# a_49002_14688# 2.86e-19
C1278 a_48702_16634# a_48616_14688# 3.14e-19
C1279 X1.X1.X2.X3.vin1 X1.X1.X1.X2.X3.vin2 7.46e-20
C1280 a_40352_32700# X2.X1.X2.X2.X2.X2.X1.vin2 1.78e-19
C1281 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X3.vin1 0.00118f
C1282 a_37766_8828# X2.X1.X2.X1.X1.X2.vout 0.418f
C1283 X1.X1.X1.X1.X2.X1.X3.vin2 a_2196_23258# 0.354f
C1284 X2.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X3.vin2 0.0533f
C1285 X2.X1.X3.vin2 a_37852_18358# 0.355f
C1286 a_20286_892# a_20672_892# 0.406f
C1287 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.vout 0.075f
C1288 X2.X1.X1.X1.X2.X2.X3.vin2 a_31862_19446# 0.567f
C1289 a_19422_31882# X1.X2.X1.X1.X1.X1.X3.vin2 0.267f
C1290 a_52106_18358# a_52792_16452# 3.08e-19
C1291 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin1 0.267f
C1292 X1.X2.X1.X2.vrefh a_17222_17540# 8.22e-20
C1293 a_39966_13640# a_40352_13640# 0.419f
C1294 a_2196_28976# a_2582_28976# 0.419f
C1295 a_4696_10916# a_4396_9010# 6.2e-19
C1296 a_31476_13728# X2.X1.X1.X2.X1.X2.X3.vin1 0.354f
C1297 X1.X1.X2.X1.X2.X2.X3.vin1 a_11072_15546# 0.354f
C1298 a_2196_13728# X1.X1.X1.X2.X1.X2.X2.vin1 1.78e-19
C1299 a_31862_13728# X2.X1.X1.X2.X1.X2.X1.vin1 0.417f
C1300 a_19422_24258# a_19722_22312# 4.19e-20
C1301 X1.X2.X1.X1.X2.X1.vout a_19336_22312# 0.169f
C1302 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.vrefh 0.161f
C1303 X1.X1.X1.X2.X1.X2.X3.vin2 a_5082_10916# 0.00846f
C1304 a_4396_16634# a_2582_15634# 1.15e-20
C1305 a_54606_21264# X2.X2.X2.X2.X1.X1.X1.vin2 8.88e-20
C1306 a_37852_18358# a_37766_16452# 3.3e-19
C1307 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X3.vin1 1.22e-19
C1308 X2.X2.X2.vrefh a_54606_4110# 4.89e-19
C1309 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X2.vin1 0.0689f
C1310 a_17222_17540# a_19036_16634# 1.06e-19
C1311 X1.X1.X2.X1.X1.X1.X3.vin1 a_8872_5016# 0.199f
C1312 a_34362_29936# X2.X1.X1.X1.X1.X2.vout 0.254f
C1313 a_2196_9916# a_2196_8010# 0.00396f
C1314 X1.X2.X1.X1.X2.X2.X3.vin2 a_17222_19446# 0.567f
C1315 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X1.vin2 0.216f
C1316 X2.X1.X2.X1.X2.X1.X1.vin1 a_39966_9828# 8.22e-20
C1317 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X1.X2.X1.X1.X2.X3.vin2 3.94e-19
C1318 X1.X1.X2.X2.X2.X1.X3.vin1 X1.X1.X2.X2.X2.X1.X1.vin2 0.216f
C1319 a_8486_27888# a_10686_26982# 4.2e-20
C1320 a_31476_30882# a_31862_30882# 0.419f
C1321 a_52406_27888# a_54606_26982# 4.2e-20
C1322 X2.X2.X1.X1.X2.X1.X1.vin2 a_46116_23258# 1.78e-19
C1323 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X1.X1.vin2 0.216f
C1324 a_19422_12822# X1.X2.X1.X2.X1.X2.X3.vin2 0.277f
C1325 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X1.vin2 0.216f
C1326 X1.X2.X2.X2.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin2 0.0128f
C1327 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X2.vin1 0.242f
C1328 X2.X1.X2.X1.X2.X2.X3.vin2 a_37466_14586# 3.85e-19
C1329 X2.X1.X2.X1.X2.X2.vrefh a_39966_13640# 0.3f
C1330 X2.X2.X1.X1.X2.X1.X3.vin1 a_48702_24258# 0.428f
C1331 X1.X2.X3.vin1 X1.X2.X2.vrefh 0.178f
C1332 X2.X2.X1.X3.vin2 a_48616_10916# 0.355f
C1333 a_52106_25982# a_52492_25982# 0.414f
C1334 X2.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X1.vin2 0.096f
C1335 a_25326_32700# X1.X2.X2.X2.X2.X2.X2.vin1 0.402f
C1336 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X1.X3.vin2 0.234f
C1337 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X1.X2.X1.X2.X2.X3.vin2 3.94e-19
C1338 X2.X1.X2.X2.X1.X1.X1.vin1 a_39966_17452# 8.22e-20
C1339 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X1.vout 0.13f
C1340 X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.vout 1.71e-19
C1341 X2.X2.X1.X3.vin1 a_48702_20446# 5.31e-19
C1342 X2.X2.X2.X2.X1.X2.X1.vin2 a_54606_23170# 0.273f
C1343 X1.X2.X1.X3.vin1 a_19722_22312# 7.98e-19
C1344 X1.X2.X2.X2.X2.X2.X1.vin2 X1.X2.X2.X2.X2.X2.X1.vin1 0.668f
C1345 X2.X2.X2.X1.X2.X2.vout a_52492_14586# 0.0929f
C1346 X1.X1.X3.vin1 a_8486_16452# 8.66e-20
C1347 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X1.X1.vin1 0.206f
C1348 X1.X1.X1.X2.X2.X2.X3.vin2 a_2196_4198# 0.354f
C1349 X2.X1.X2.X1.X1.X2.X3.vin2 a_39966_7922# 7.84e-19
C1350 a_4782_5198# a_2582_4198# 4.77e-21
C1351 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X1.vin1 0.0689f
C1352 X1.X2.X1.X1.X1.X2.vout a_19422_28070# 0.418f
C1353 a_37466_14586# a_37766_12640# 4.19e-20
C1354 X1.X1.X2.X1.X3.vin1 a_8572_6962# 0.363f
C1355 X1.X2.X2.vrefh a_25326_4110# 4.89e-19
C1356 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X3.vin1 2.33e-19
C1357 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 1.22e-19
C1358 a_54606_6016# a_52406_5016# 4.77e-21
C1359 a_10686_13640# X1.X1.X2.X1.X2.X1.X1.vin2 8.88e-20
C1360 a_31476_32788# a_31476_30882# 0.00396f
C1361 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X3.vin2 0.165f
C1362 a_4396_24258# a_4782_24258# 0.419f
C1363 X1.X2.X1.X2.X2.X1.X1.vin2 a_17222_8010# 8.88e-20
C1364 a_4696_26164# a_5082_26164# 0.414f
C1365 a_19036_28070# a_19722_26164# 3.08e-19
C1366 X1.X1.X2.X2.X2.X2.vrefh X1.X1.X2.X2.X2.X1.X1.vin2 0.076f
C1367 X1.X2.X2.X3.vin1 a_23212_18358# 0.17f
C1368 a_19422_28070# a_19336_26164# 3.3e-19
C1369 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X1.vin2 0.668f
C1370 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X1.vin2 0.216f
C1371 a_33976_10916# X2.X1.X1.X2.X2.X1.vout 1.64e-19
C1372 a_34362_10916# a_34062_9010# 5.25e-20
C1373 X1.X1.X2.X1.X2.X2.X3.vin1 a_8872_16452# 0.199f
C1374 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X2.vrefh 0.076f
C1375 X1.X1.X2.X2.X1.X2.X3.vin2 a_8872_24076# 0.101f
C1376 X2.X2.X2.X1.X3.vin1 a_52492_10734# 0.169f
C1377 a_48616_7064# a_48702_5198# 3.38e-19
C1378 X1.X2.X1.X1.X1.X1.X3.vin1 a_17222_30882# 0.00207f
C1379 a_31476_8010# a_31476_6104# 0.00396f
C1380 a_49002_7064# a_48316_5198# 3.31e-19
C1381 a_19336_10916# X1.X2.X1.X2.X2.X1.X3.vin1 0.00251f
C1382 a_25326_17452# X1.X2.X2.X1.X2.X2.X3.vin1 0.00207f
C1383 X1.X1.X2.X2.X1.X2.X3.vin1 a_8572_22210# 0.00329f
C1384 X1.X2.X2.X2.X3.vin1 a_23126_24076# 9.54e-19
C1385 X2.X1.X2.X1.X2.vrefh a_40352_9828# 0.118f
C1386 X2.X2.X1.X1.X1.X1.vout X2.X2.X1.X1.X1.X1.X3.vin2 0.342f
C1387 X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X3.vin2 0.0533f
C1388 a_25326_6016# a_25326_4110# 0.00198f
C1389 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 0.242f
C1390 X2.X2.X1.X2.X1.X2.X1.vin2 a_46502_11822# 8.88e-20
C1391 a_52492_29834# a_52406_27888# 3.14e-19
C1392 X2.X2.X1.X2.X2.X2.X2.vin1 a_46502_4198# 0.402f
C1393 a_52406_5016# X2.X2.X2.X1.X1.X1.X3.vin1 0.428f
C1394 X2.X2.X1.X2.X1.X2.X3.vin1 a_48316_12822# 0.199f
C1395 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin2 7.84e-19
C1396 X2.X1.X1.X1.X2.X2.X1.vin2 a_31862_19446# 8.88e-20
C1397 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 5.19e-19
C1398 X2.X1.X1.X2.X1.X1.X3.vin2 a_31862_15634# 0.567f
C1399 X1.X1.X2.X2.X1.X2.X2.vin1 a_11072_25076# 0.197f
C1400 a_19722_29936# X1.X2.X1.X1.X3.vin1 0.434f
C1401 X2.X1.X2.X2.X2.X2.X3.vin1 a_40352_30794# 0.354f
C1402 a_2582_32788# a_2582_30882# 0.00198f
C1403 X1.X1.X2.X3.vin1 a_8486_12640# 5.28e-19
C1404 X1.X2.X1.X2.X2.X1.X3.vin2 X1.X2.X1.X2.X2.X2.X1.vin1 5.19e-19
C1405 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin1 0.52f
C1406 X1.X1.X2.X2.X1.X2.X3.vin2 a_8186_22210# 3.85e-19
C1407 a_33676_31882# a_31862_30882# 1.15e-20
C1408 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X2.vin1 0.242f
C1409 X1.X2.X2.X1.X2.X2.X2.vin1 a_25712_17452# 0.197f
C1410 X2.X1.X1.X1.X1.X2.vout X2.X1.X1.X1.X1.X2.X3.vin2 0.075f
C1411 X2.X2.X2.X1.X2.X1.vout a_52406_12640# 0.422f
C1412 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X2.vrefh 0.267f
C1413 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X1.vin2 0.668f
C1414 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin1 0.52f
C1415 a_48316_24258# a_49002_22312# 2.86e-19
C1416 a_48702_24258# a_48616_22312# 3.14e-19
C1417 X2.X1.X1.X2.X2.X2.X2.vin1 a_31862_4198# 0.402f
C1418 X1.X2.X1.X1.X2.X2.X3.vin1 a_17222_19446# 0.00207f
C1419 a_23512_8828# a_23212_6962# 6.71e-19
C1420 X2.X2.X2.X2.X2.X2.X3.vin2 a_52106_29834# 3.85e-19
C1421 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin1 0.195f
C1422 a_38152_12640# a_37466_10734# 2.97e-19
C1423 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X1.X3.vin2 5.19e-19
C1424 a_37466_25982# X2.X1.X2.X3.vin2 0.452f
C1425 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X3.vin2 8.93e-19
C1426 X2.X1.X1.X1.X2.vrefh a_31476_27070# 0.118f
C1427 a_46502_32788# a_48702_31882# 4.2e-20
C1428 X2.X2.X1.X1.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X1.X2.vin1 0.00117f
C1429 X1.X2.X1.X1.X1.X2.X3.vin2 a_17222_25164# 8.07e-19
C1430 X1.X1.X1.X1.X3.vin2 a_4696_22312# 0.363f
C1431 X2.X3.vin1 a_42976_892# 0.195f
C1432 a_48316_20446# a_49002_18540# 3.08e-19
C1433 X2.X1.X1.X2.X2.X1.X3.vin2 a_31862_8010# 0.567f
C1434 a_48702_20446# a_48616_18540# 3.3e-19
C1435 a_34062_28070# a_34362_26164# 4.41e-20
C1436 X2.X1.X1.X1.X1.X2.X3.vin2 a_33976_26164# 0.00535f
C1437 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X3.vin2 8.93e-19
C1438 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X3.vin1 0.00118f
C1439 X1.X2.X2.X2.X1.X1.vout a_23126_20264# 0.422f
C1440 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.vrefh 2.33e-19
C1441 a_19036_5198# a_17222_4198# 1.15e-20
C1442 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin1 0.267f
C1443 a_37466_25982# a_37766_24076# 4.41e-20
C1444 X1.X1.X2.X1.X2.X2.X1.vin2 a_10686_15546# 0.273f
C1445 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 2.23e-19
C1446 X2.X2.X2.X2.X2.X2.X1.vin1 a_54992_30794# 0.195f
C1447 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X1.X3.vin2 0.0943f
C1448 X1.X1.X2.X1.X3.vin1 a_8486_8828# 9.54e-19
C1449 a_31862_32788# X2.X1.X1.X1.X1.X1.X2.vin1 8.88e-20
C1450 X2.X1.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X1.vin1 0.267f
C1451 a_10686_21264# a_11072_21264# 0.419f
C1452 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X2.X3.vin1 0.0174f
C1453 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X1.vin2 0.1f
C1454 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.vrefh 0.1f
C1455 X1.X1.X2.X3.vin1 X1.X1.X3.vin2 1.16f
C1456 X2.X1.X1.X1.X1.X2.X1.vin2 a_31476_27070# 1.78e-19
C1457 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X3.vin1 1.42e-20
C1458 a_2582_21352# X1.X1.X1.X1.X2.X2.X1.vin1 0.417f
C1459 a_2196_21352# X1.X1.X1.X1.X2.X2.X3.vin1 0.354f
C1460 X1.X2.X2.X1.X2.X2.X3.vin1 a_22826_14586# 0.00874f
C1461 X1.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X3.vin1 0.0321f
C1462 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X1.vin2 0.216f
C1463 a_37466_10734# X2.X1.X2.X1.X3.vin1 0.385f
C1464 X1.X2.X1.X1.X1.X1.X3.vin1 a_19422_31882# 0.428f
C1465 a_31862_28976# X2.X1.X1.X1.X1.X2.X3.vin2 7.84e-19
C1466 X2.X1.X1.X1.X1.X2.X3.vin1 a_33676_28070# 0.199f
C1467 X2.X2.X2.X1.X3.vin2 a_52492_14586# 0.363f
C1468 a_10686_17452# a_10686_15546# 0.00198f
C1469 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 0.242f
C1470 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X3.vin2 8.93e-19
C1471 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X1.vin2 3.94e-19
C1472 X1.X1.X2.X1.X1.X2.X1.vin2 a_10686_7922# 0.273f
C1473 X2.X1.X2.X1.X1.X2.vout X2.X1.X2.X1.X1.X1.vout 0.507f
C1474 a_8186_10734# a_8572_10734# 0.414f
C1475 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X3.vin2 0.161f
C1476 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X3.vin1 0.0131f
C1477 X1.X3.vin1 X3.vin1 0.143f
C1478 a_34062_16634# X2.X1.X1.X2.X1.X1.X3.vin2 0.267f
C1479 X2.X2.X2.X2.X1.X1.vout a_52492_18358# 1.64e-19
C1480 X2.X1.X1.X1.X2.X2.vrefh a_31862_21352# 8.22e-20
C1481 a_11072_7922# a_11072_6016# 0.00396f
C1482 X2.X2.X1.X1.X1.X2.X3.vin2 a_49002_26164# 0.00846f
C1483 a_48702_28070# X2.X2.X1.X3.vin1 1.64e-19
C1484 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X1.vin1 2.23e-19
C1485 X2.X1.X2.X2.X1.X2.X2.vin1 a_40352_23170# 1.78e-19
C1486 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X3.vin1 0.00118f
C1487 a_33676_31882# a_34062_31882# 0.419f
C1488 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X3.vin2 0.552f
C1489 a_52492_6962# a_54606_6016# 2.95e-20
C1490 a_25326_6016# a_25712_6016# 0.419f
C1491 a_10686_17452# X1.X1.X2.X1.X2.X2.X2.vin1 0.402f
C1492 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X3.vin2 0.161f
C1493 X2.X2.X2.X2.X2.X2.X2.vin1 X2.X2.X2.X2.X2.X2.X3.vin1 0.00117f
C1494 X2.X2.X2.X2.X2.X2.X3.vin2 a_52406_31700# 0.277f
C1495 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X1.vin1 0.206f
C1496 X2.X1.X3.vin2 a_37466_14586# 3.67e-19
C1497 X1.X2.X1.X2.X1.X2.X3.vin1 a_17222_11822# 0.00207f
C1498 a_33976_22312# a_33676_20446# 6.71e-19
C1499 a_17222_6104# X1.X2.X1.X2.X2.X2.X1.vin1 0.417f
C1500 a_16836_6104# X1.X2.X1.X2.X2.X2.X3.vin1 0.354f
C1501 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X2.vrefh 0.267f
C1502 a_46502_17540# X2.X2.X1.X2.X1.X1.X2.vin1 8.88e-20
C1503 X1.X2.X1.X2.X1.X1.X2.vin1 a_17222_15634# 0.402f
C1504 a_4696_14688# X1.X1.X1.X2.X1.X2.vout 0.0929f
C1505 a_10686_11734# a_10686_9828# 0.00198f
C1506 a_31476_19446# a_31862_19446# 0.419f
C1507 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X2.vout 0.0866f
C1508 X1.X2.X1.X1.X3.vin2 X1.X2.X2.X3.vin2 7.46e-20
C1509 a_22826_25982# X1.X2.X2.X2.X3.vin1 0.372f
C1510 X2.X1.X1.X3.vin1 X2.X1.X1.X3.vin2 0.552f
C1511 a_2582_21352# a_2582_19446# 0.00198f
C1512 a_34062_9010# X2.X1.X1.X2.X2.X1.X3.vin2 0.267f
C1513 X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X2.X1.X1.vin2 0.1f
C1514 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X3.vin2 0.161f
C1515 a_23126_5016# a_23512_5016# 0.419f
C1516 a_39966_32700# a_37766_31700# 4.77e-21
C1517 a_37766_16452# a_37466_14586# 5.55e-20
C1518 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X1.vout 0.038f
C1519 X1.X2.X2.X2.X1.X2.vout a_22826_22210# 0.254f
C1520 a_33976_7064# X2.X1.X1.X2.X2.X2.vout 0.0929f
C1521 X2.X2.X2.X2.X1.X2.X3.vin2 a_54992_25076# 0.354f
C1522 a_25712_17452# a_25712_15546# 0.00396f
C1523 a_8872_12640# a_8572_10734# 6.2e-19
C1524 a_19336_14688# a_19036_12822# 6.71e-19
C1525 a_19722_18540# X1.X2.X3.vin2 6.58e-20
C1526 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.X1.vin1 0.206f
C1527 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin2 7.84e-19
C1528 X1.X2.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X2.X1.X3.vin2 0.161f
C1529 X2.X2.X3.vin1 a_48702_5198# 2.12e-19
C1530 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X3.vin1 0.206f
C1531 X1.X2.X1.X1.X1.X2.X2.vin1 a_17222_27070# 0.402f
C1532 X1.X2.X1.X2.X2.X1.X2.vin1 a_17222_8010# 0.402f
C1533 a_33976_22312# X2.X1.X1.X1.X2.X2.X3.vin1 0.00329f
C1534 a_16836_19446# a_17222_19446# 0.419f
C1535 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X3.vin1 0.00117f
C1536 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X2.vrefh 0.00118f
C1537 X2.X2.X2.X2.X1.X1.X3.vin2 a_52406_20264# 0.267f
C1538 X1.X1.X3.vin1 X1.X1.X2.vrefh 0.178f
C1539 a_25326_11734# X1.X2.X2.X1.X2.X1.X1.vin1 0.417f
C1540 X1.X2.X2.X1.X2.X1.X1.vin2 a_25712_11734# 0.12f
C1541 X1.X1.X1.X2.X2.X2.vout a_4782_5198# 0.418f
C1542 a_5082_7064# X1.X1.X1.X2.X2.X2.X3.vin2 3.85e-19
C1543 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X1.vin1 5.19e-19
C1544 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X1.X2.X1.X2.X2.X1.vin1 0.668f
C1545 a_54606_26982# X2.X2.X2.X2.X2.vrefh 8.22e-20
C1546 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X2.vin1 0.242f
C1547 X2.X1.X2.X2.X2.X2.vout X2.X1.X2.X2.X3.vin2 0.0866f
C1548 X1.X1.X1.X2.X2.X1.vout a_5082_7064# 0.383f
C1549 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X2.vin1 0.242f
C1550 a_37766_8828# a_37852_6962# 3.38e-19
C1551 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X1.vin1 0.0689f
C1552 X2.X1.X2.X1.X2.X1.X3.vin2 a_39966_11734# 7.84e-19
C1553 X1.X2.X1.X1.X2.X2.vrefh a_17222_23258# 0.3f
C1554 a_23512_24076# a_25326_23170# 1.06e-19
C1555 X2.X1.X2.X1.X2.X1.vout a_37852_14586# 0.169f
C1556 X2.X2.X2.X3.vin1 a_52492_10734# 0.356f
C1557 X2.X2.X3.vin2 X2.X2.X2.X1.X3.vin1 0.0361f
C1558 X2.X1.X2.X2.X3.vin2 X2.X1.X1.X3.vin1 7.46e-20
C1559 a_31476_27070# a_31476_25164# 0.00396f
C1560 a_4696_26164# X1.X1.X1.X1.X2.X1.vout 1.64e-19
C1561 a_5082_26164# a_4782_24258# 5.25e-20
C1562 a_19336_22312# X1.X2.X1.X1.X2.X2.vout 0.0929f
C1563 X2.X2.X1.X1.X2.X2.vout a_48702_20446# 0.418f
C1564 a_49002_22312# X2.X2.X1.X1.X2.X2.X3.vin2 3.85e-19
C1565 X2.X1.X1.X1.X2.vrefh a_31862_25164# 8.22e-20
C1566 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.X1.X1.X1.vin1 5.19e-19
C1567 a_2196_19446# a_2582_19446# 0.419f
C1568 X2.X2.X1.X2.X2.X1.X1.vin2 a_46502_8010# 8.88e-20
C1569 X1.X2.X1.X2.X3.vin1 a_19336_10916# 0.17f
C1570 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X2.vin1 0.564f
C1571 X1.X2.X2.X2.X2.X2.X3.vin1 a_23212_29834# 0.00329f
C1572 a_40352_25076# X2.X1.X2.X2.X1.X2.X1.vin2 1.78e-19
C1573 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 5.19e-19
C1574 a_2582_8010# X1.X1.X1.X2.X2.X2.X1.vin1 8.22e-20
C1575 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.vout 0.118f
C1576 X1.X2.X1.X1.X2.X1.X2.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 0.234f
C1577 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X1.X2.X1.X1.X2.X1.vin1 0.668f
C1578 X1.X1.X1.X1.X1.X2.X3.vin1 a_2582_27070# 0.00207f
C1579 X2.X1.X2.X2.X1.X1.vout a_38152_20264# 0.359f
C1580 a_4782_12822# a_2582_11822# 4.77e-21
C1581 X1.X1.X1.X2.X1.X2.X3.vin2 a_2196_11822# 0.354f
C1582 a_48702_12822# a_46502_11822# 4.77e-21
C1583 X1.X2.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X2.X2.vrefh 0.117f
C1584 a_54606_17452# a_52406_16452# 4.77e-21
C1585 a_10686_32700# X1.X2.vrefh 0.3f
C1586 X1.X1.X2.X2.X2.X2.X2.vin1 a_11072_32700# 0.197f
C1587 X2.X2.X1.X2.X1.X2.X3.vin2 a_46116_11822# 0.354f
C1588 X1.X2.X2.X1.X2.X1.X3.vin2 a_23512_12640# 0.1f
C1589 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X2.vrefh 0.076f
C1590 X2.X2.X1.X3.vin1 a_48702_24258# 5.28e-19
C1591 X2.X2.X2.X2.X1.X1.X2.vin1 a_54992_21264# 0.197f
C1592 a_16836_23258# a_16836_21352# 0.00396f
C1593 X2.X1.X2.X1.X1.X2.X3.vin2 a_40352_9828# 0.354f
C1594 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin1 0.52f
C1595 X2.X2.X1.X1.X2.X1.X3.vin2 a_46502_23258# 0.567f
C1596 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X2.vin1 0.00117f
C1597 a_17222_13728# a_19422_12822# 4.2e-20
C1598 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin1 0.52f
C1599 X1.X2.X2.X3.vin1 a_22826_14586# 7.98e-19
C1600 a_10686_26982# X1.X1.X2.X2.X1.X2.X3.vin2 8.07e-19
C1601 a_33976_14688# a_34062_12822# 3.38e-19
C1602 a_34362_14688# a_33676_12822# 3.31e-19
C1603 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X2.X1.vin2 0.668f
C1604 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X3.vin1 0.206f
C1605 X1.X2.X1.X3.vin2 X1.X2.X2.X1.X3.vin2 7.46e-20
C1606 X2.X2.X3.vin1 X2.X2.X2.X1.X1.X1.vout 5.53e-20
C1607 X1.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin2 0.0128f
C1608 a_31476_9916# X2.X1.X1.X2.X2.X1.X2.vin1 1.78e-19
C1609 a_52106_10734# X2.X2.X2.X1.X1.X2.X3.vin2 0.00846f
C1610 a_8186_29834# a_8486_27888# 4.19e-20
C1611 X1.X1.X1.X3.vin1 X1.X1.X2.X3.vin2 1.22e-19
C1612 a_10686_11734# a_8572_10734# 5.36e-21
C1613 X1.X2.X1.X3.vin1 X1.X2.X3.vin1 0.188f
C1614 a_33976_18540# X2.X1.X1.X3.vin2 0.0927f
C1615 X2.X2.X1.X2.X2.X1.X3.vin2 a_46502_6104# 8.07e-19
C1616 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X2.vrefh 0.00118f
C1617 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X3.vin1 0.581f
C1618 X2.X1.X1.X2.X1.X1.vout X2.X1.X1.X2.X3.vin1 0.131f
C1619 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X2.vrefh 0.00118f
C1620 X2.X1.X1.X2.X2.X2.X1.vin2 a_31862_4198# 8.88e-20
C1621 a_54606_28888# X2.X2.X2.X2.X2.X1.X3.vin1 0.00207f
C1622 a_48702_16634# a_46502_15634# 4.77e-21
C1623 X1.X2.X1.X2.X2.X2.vrefh X1.X1.X2.X1.X1.X2.vrefh 0.117f
C1624 a_52792_31700# a_52106_29834# 3.31e-19
C1625 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin2 0.12f
C1626 a_23126_27888# a_23512_27888# 0.419f
C1627 X2.X1.X1.X2.X2.X2.X3.vin1 a_33676_5198# 0.199f
C1628 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin2 7.84e-19
C1629 a_23512_20264# a_23212_18358# 6.2e-19
C1630 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X2.vrefh 0.165f
C1631 a_39966_25076# X2.X1.X2.X2.X1.X2.X3.vin2 0.567f
C1632 X1.X1.X3.vin1 a_8186_18358# 5.87e-20
C1633 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X1.X3.vin2 5.19e-19
C1634 X1.X1.X1.X1.X2.X1.X3.vin2 a_5082_22312# 0.00815f
C1635 X1.X2.X2.X2.X1.X2.X1.vin1 X2.X1.X1.X1.X2.X2.vrefh 0.00437f
C1636 a_4396_31882# X1.X1.X1.X1.X1.X1.X3.vin2 0.1f
C1637 a_46116_21352# X2.X2.X1.X1.X2.X2.X2.vin1 1.78e-19
C1638 a_54606_17452# X2.X2.X2.X1.X2.X2.X3.vin2 0.567f
C1639 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X2.X1.X1.X1.X1.X1.vin2 0.00232f
C1640 X1.X2.X2.X2.X3.vin2 a_23212_29834# 0.363f
C1641 a_23212_14586# X1.X2.X2.X1.X2.X1.X3.vin2 0.00546f
C1642 a_37766_31700# a_37852_29834# 3.38e-19
C1643 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X2.vin1 0.564f
C1644 X1.X2.X2.X2.X2.X1.X3.vin2 a_25326_26982# 7.84e-19
C1645 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X1.X1.vin1 0.0689f
C1646 X1.X2.X2.X1.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin2 0.0128f
C1647 X1.X1.X2.X1.X1.X2.vrefh a_11072_6016# 0.118f
C1648 a_11072_6016# a_11072_4110# 0.00396f
C1649 a_48702_9010# a_46502_8010# 4.77e-21
C1650 a_39966_21264# a_37766_20264# 4.77e-21
C1651 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin1 0.267f
C1652 a_5082_10916# X1.X1.X1.X2.X3.vin2 0.263f
C1653 a_19722_18540# a_19036_16634# 2.97e-19
C1654 X1.X1.X1.X2.X1.X1.vout a_4696_14688# 0.169f
C1655 a_4782_16634# a_5082_14688# 4.19e-20
C1656 a_19336_18540# a_19422_16634# 3.21e-19
C1657 X1.X2.X2.X1.X1.X1.vout X1.X2.X2.X1.X1.X1.X3.vin1 0.118f
C1658 X2.X1.X2.X2.X3.vin1 a_37466_22210# 0.436f
C1659 a_8486_20264# a_10686_19358# 4.2e-20
C1660 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 0.216f
C1661 X2.X2.X2.X3.vin2 a_52406_20264# 5.21e-19
C1662 a_49002_14688# a_48702_12822# 5.55e-20
C1663 X1.X2.X2.X1.X2.X1.vout X1.X2.X2.X1.X3.vin2 0.399f
C1664 a_48616_26164# a_49002_26164# 0.414f
C1665 X1.X1.X3.vin2 X1.X1.X2.X1.X2.X2.vout 3.38e-19
C1666 X1.X1.X3.vin1 a_5646_892# 0.17f
C1667 a_31476_25164# a_31476_23258# 0.00396f
C1668 a_37852_22210# a_37766_20264# 3.14e-19
C1669 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin2 0.1f
C1670 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X2.X1.X1.X2.X1.X2.vin1 0.00232f
C1671 a_23212_29834# a_23126_27888# 3.14e-19
C1672 X1.X1.X2.X2.X2.vrefh a_11072_25076# 0.118f
C1673 a_33976_18540# a_31862_17540# 5.36e-21
C1674 X1.X1.X2.X2.X3.vin1 a_8572_22210# 0.363f
C1675 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X1.vout 0.0524f
C1676 X2.X2.X2.X1.X2.X1.X3.vin1 a_52792_12640# 0.199f
C1677 a_38152_27888# a_37466_25982# 2.97e-19
C1678 a_54992_6016# a_54992_4110# 0.00396f
C1679 a_48702_16634# X2.X2.X1.X2.X3.vin1 1.52e-19
C1680 X2.X2.X1.X2.X1.X1.vout a_49002_14688# 0.387f
C1681 a_39966_17452# X2.X1.X2.X1.X2.X2.X1.vin2 8.88e-20
C1682 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin2 0.12f
C1683 a_19722_26164# X1.X2.X1.X1.X3.vin2 0.241f
C1684 d7 X3.vin2 4.93e-19
C1685 a_28096_892# vout 0.349f
C1686 a_48616_29936# a_46502_28976# 2.68e-20
C1687 a_48316_24258# X2.X2.X1.X1.X2.X1.X3.vin2 0.1f
C1688 a_39966_21264# X2.X1.X2.X2.X1.X1.X2.vin1 0.402f
C1689 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 1.22e-19
C1690 a_10686_28888# a_11072_28888# 0.419f
C1691 a_25326_9828# X1.X2.X2.X1.X1.X2.X3.vin2 0.567f
C1692 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X3.vin1 2.33e-19
C1693 X2.X1.X2.X1.X2.X1.X3.vin2 a_40352_13640# 0.354f
C1694 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 2.23e-19
C1695 a_8572_6962# a_10686_6016# 2.95e-20
C1696 X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin1 4.41e-19
C1697 a_2196_28976# X1.X1.X1.X1.X1.X2.X3.vin1 0.354f
C1698 X1.X1.X3.vin1 X1.X1.X2.X1.X3.vin2 6.26e-19
C1699 a_2582_28976# X1.X1.X1.X1.X1.X2.X1.vin1 0.417f
C1700 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X1.X3.vin2 1.22e-19
C1701 a_5082_10916# a_4782_9010# 5.25e-20
C1702 a_10686_6016# a_8872_5016# 1.15e-20
C1703 a_4696_10916# X1.X1.X1.X2.X2.X1.vout 1.64e-19
C1704 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X3.vin1 0.206f
C1705 X1.X2.X2.X1.X2.X1.vout a_23126_12640# 0.422f
C1706 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X2.vin1 0.0689f
C1707 a_2582_13728# a_4396_12822# 1.06e-19
C1708 X1.X2.X1.X1.X2.X1.vout X1.X2.X1.X1.X2.X2.vout 0.514f
C1709 a_25326_9828# a_23512_8828# 1.15e-20
C1710 X2.X2.X2.vrefh X2.X3.vin1 0.00136f
C1711 X2.X1.X2.X1.X1.X2.X1.vin1 a_40352_6016# 1.64e-19
C1712 a_8186_22210# a_8872_20264# 2.86e-19
C1713 a_2582_6104# X1.X1.X1.X2.X2.X2.X2.vin1 8.88e-20
C1714 X2.X2.X2.X2.X1.X1.X3.vin2 X2.X2.X2.X2.X1.X1.X1.vin2 8.93e-19
C1715 X2.X2.X2.X2.X1.X1.X2.vin1 a_54606_19358# 8.88e-20
C1716 a_19336_18540# X1.X2.X3.vin1 0.354f
C1717 X2.X1.X2.X2.X1.X2.X3.vin1 a_39966_23170# 0.52f
C1718 X1.X2.X2.X1.X1.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin2 0.0128f
C1719 a_33676_12822# X2.X1.X1.X2.X1.X2.X3.vin2 0.101f
C1720 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X1.X2.X1.X2.X2.vrefh 0.1f
C1721 a_52406_31700# a_52792_31700# 0.419f
C1722 a_48316_16634# a_48702_16634# 0.419f
C1723 X2.X1.X1.X1.X2.X1.X2.vin1 a_31476_23258# 0.197f
C1724 X1.X1.X3.vin2 X1.X1.X1.X2.X2.X2.vout 1.5e-19
C1725 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X3.vin2 8.93e-19
C1726 X2.X1.X2.X2.X1.X2.vout a_38152_24076# 0.36f
C1727 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X2.vrefh 2.33e-19
C1728 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X1.vin2 0.076f
C1729 X2.X2.X2.vrefh a_54992_4110# 9.79e-19
C1730 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X2.X1.X1.X1.X2.vrefh 0.0128f
C1731 X1.X2.X1.X2.X1.X1.X3.vin1 a_19036_16634# 0.199f
C1732 X1.X1.X1.X1.X1.X2.vout X1.X1.X1.X1.X1.X2.X3.vin1 0.326f
C1733 a_31476_25164# a_31862_25164# 0.419f
C1734 X1.X2.X2.X2.X1.X2.X2.vin1 X2.X1.X1.X1.X2.X1.X1.vin2 0.00232f
C1735 a_2582_9916# a_2582_8010# 0.00198f
C1736 a_33976_18540# a_33676_16634# 6.2e-19
C1737 X1.X2.X1.X2.X1.X1.X3.vin2 a_19336_14688# 0.00546f
C1738 X1.X1.X1.X2.X1.X2.vout a_4782_12822# 0.418f
C1739 a_4396_5198# a_4782_5198# 0.419f
C1740 X1.X1.X1.X2.X2.X2.X2.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 0.234f
C1741 a_54992_19358# a_54992_17452# 0.00396f
C1742 X1.X1.X2.X2.X2.X1.X3.vin1 X1.X1.X2.X2.X2.X1.X1.vin1 0.206f
C1743 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 5.19e-19
C1744 X1.X1.X3.vin1 X1.X1.X2.X1.X1.X2.vout 1.71e-19
C1745 a_46116_17540# a_46502_17540# 0.419f
C1746 a_39966_32700# X2.X1.X2.X2.X2.X2.X3.vin2 0.567f
C1747 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X2.X1.X2.X1.X1.X1.vin2 0.00232f
C1748 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X1.X1.vin1 0.206f
C1749 a_23212_18358# X1.X2.X2.X1.X2.X2.vout 7.93e-20
C1750 a_54606_6016# X2.X2.X2.X1.X1.X1.X2.vin1 0.402f
C1751 X1.X1.X2.X2.X2.X1.vout a_8572_29834# 0.169f
C1752 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X3.vin2 0.161f
C1753 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X3.vin2 0.0523f
C1754 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X3.vin2 0.17f
C1755 X2.X1.X1.X1.X3.vin1 a_34362_26164# 0.385f
C1756 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X1.X2.X1.X1.X2.vrefh 0.1f
C1757 X2.X2.X3.vin1 a_52106_10734# 3.93e-19
C1758 X2.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X1.vin1 0.142f
C1759 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X3.vin2 0.237f
C1760 a_39966_13640# a_37766_12640# 4.77e-21
C1761 a_48316_9010# a_48702_9010# 0.419f
C1762 a_23126_24076# X1.X2.X2.X2.X1.X2.vout 0.418f
C1763 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.vout 0.075f
C1764 a_4396_9010# a_4782_9010# 0.419f
C1765 a_54992_17452# a_54992_15546# 0.00396f
C1766 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 5.19e-19
C1767 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X1.X3.vin1 0.0321f
C1768 a_8572_18358# a_8486_16452# 3.3e-19
C1769 X2.X2.X2.X2.X1.X2.X1.vin2 a_54992_23170# 0.12f
C1770 a_54606_23170# X2.X2.X2.X2.X1.X2.X1.vin1 0.417f
C1771 a_31476_15634# a_31476_13728# 0.00396f
C1772 a_25326_30794# a_25712_30794# 0.419f
C1773 a_49002_7064# X2.X2.X1.X2.X2.X2.X3.vin1 0.00874f
C1774 X1.X2.X2.X3.vin1 X1.X2.X1.X2.X3.vin2 7.46e-20
C1775 a_34062_12822# a_33976_10916# 3.3e-19
C1776 X1.X2.X1.X2.X1.X2.X3.vin2 a_17222_9916# 8.07e-19
C1777 a_33676_12822# a_34362_10916# 3.08e-19
C1778 a_31862_25164# X2.X1.X1.X1.X2.X1.X2.vin1 8.88e-20
C1779 X2.X2.X2.X3.vin1 X2.X2.X3.vin2 1.16f
C1780 X2.X1.X2.X1.X2.X1.vout X2.X1.X2.X1.X2.X1.X3.vin1 0.118f
C1781 X1.X2.X2.vrefh a_25712_4110# 9.79e-19
C1782 a_19722_18540# X1.X2.X1.X2.X1.X1.X3.vin1 0.00837f
C1783 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X2.vrefh 0.00118f
C1784 X2.X2.X2.X1.X1.X1.X3.vin2 a_52406_5016# 0.267f
C1785 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X3.vin1 0.00117f
C1786 X1.X1.X2.X1.X2.X1.X2.vin1 a_10686_11734# 8.88e-20
C1787 X1.X2.X1.X3.vin2 a_19722_14688# 0.00292f
C1788 X1.X1.X2.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X1.vin2 8.93e-19
C1789 a_31862_32788# a_31862_30882# 0.00198f
C1790 a_37852_25982# a_38152_24076# 6.48e-19
C1791 a_4782_24258# X1.X1.X1.X1.X2.X1.vout 0.422f
C1792 X2.X1.X2.X1.X1.X1.vout a_37852_6962# 0.169f
C1793 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X2.X1.X2.X2.X1.X1.vin2 0.00232f
C1794 a_16836_9916# a_17222_9916# 0.419f
C1795 a_34362_29936# X2.X1.X1.X1.X1.X2.X3.vin1 0.00874f
C1796 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X1.vin1 5.19e-19
C1797 a_5082_26164# X1.X1.X1.X3.vin1 0.509f
C1798 X1.X2.X1.X1.X1.X2.X3.vin2 a_19722_26164# 0.00846f
C1799 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin2 0.12f
C1800 a_19422_28070# X1.X2.X1.X3.vin1 1.64e-19
C1801 a_11072_25076# a_11072_23170# 0.00396f
C1802 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.vout 0.399f
C1803 X1.X2.X2.X2.X3.vin1 a_23126_20264# 1.52e-19
C1804 a_25326_13640# X1.X2.X2.X1.X2.X1.X3.vin2 0.567f
C1805 X1.X1.X2.X1.X1.X1.X1.vin2 a_10686_4110# 0.273f
C1806 a_31476_8010# X2.X1.X1.X2.X2.X2.X1.vin1 1.64e-19
C1807 a_31862_8010# a_31862_6104# 0.00198f
C1808 X2.X2.X1.X2.X2.X2.vout a_48702_5198# 0.418f
C1809 a_49002_7064# X2.X2.X1.X2.X2.X2.X3.vin2 3.85e-19
C1810 X2.X1.X1.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X1.X2.X1.vin1 5.19e-19
C1811 X1.X2.X2.X1.X3.vin1 a_23126_5016# 1.52e-19
C1812 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X3.vin1 0.587f
C1813 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X3.vin1 0.0321f
C1814 a_8572_6962# a_8872_5016# 6.1e-19
C1815 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X1.vin2 3.94e-19
C1816 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.vout 0.335f
C1817 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X1.vin1 0.0689f
C1818 X1.X2.X2.X1.X1.X1.X3.vin2 a_25326_4110# 7.84e-19
C1819 a_8186_10734# X1.X1.X2.X1.X1.X2.X3.vin2 0.00846f
C1820 X2.X2.X1.X2.X2.X2.X3.vin2 a_46116_4198# 0.354f
C1821 a_46116_23258# a_46116_21352# 0.00396f
C1822 a_48702_5198# a_46502_4198# 4.77e-21
C1823 X2.X2.X1.X2.X2.X2.X3.vin2 X2.X2.X2.vrefh 0.172f
C1824 X1.X1.X2.X1.X1.X2.vout X1.X1.X2.X1.X1.X1.vout 0.507f
C1825 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 0.587f
C1826 X1.X1.X1.X1.X2.vrefh a_2196_27070# 0.118f
C1827 a_10686_15546# a_8572_14586# 2.68e-20
C1828 a_49002_26164# X2.X2.X1.X1.X2.X1.X3.vin1 0.00837f
C1829 X2.X2.X1.X1.X2.vrefh a_46502_27070# 0.3f
C1830 a_46502_19446# X2.X2.X1.X2.X1.X1.X1.vin1 8.22e-20
C1831 a_48616_14688# X2.X2.X1.X2.X1.X2.vout 0.0929f
C1832 a_54606_26982# a_52492_25982# 5.36e-21
C1833 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin2 7.84e-19
C1834 a_52492_22210# a_52792_20264# 6.1e-19
C1835 X1.X1.X1.X1.X1.X1.X3.vin1 a_2582_30882# 0.00207f
C1836 X1.X2.X2.X2.X1.X1.vout a_23212_22210# 0.169f
C1837 a_31476_32788# a_31862_32788# 0.419f
C1838 X2.X1.X1.X2.X2.X1.X3.vin2 a_33976_7064# 0.00546f
C1839 a_25326_28888# a_23126_27888# 4.77e-21
C1840 a_10686_30794# a_10686_28888# 0.00198f
C1841 a_52406_27888# X2.X2.X2.X3.vin2 7.93e-20
C1842 X2.X2.X2.X2.X2.X1.X2.vin1 a_54992_28888# 0.197f
C1843 X2.X1.X1.X3.vin1 a_34362_22312# 7.98e-19
C1844 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X2.vrefh 0.00118f
C1845 X1.X1.X1.X1.X1.X2.vrefh a_2582_28976# 8.22e-20
C1846 a_34062_5198# a_31862_4198# 4.77e-21
C1847 X2.X1.X1.X2.X2.X2.X3.vin2 a_31476_4198# 0.354f
C1848 X2.X2.X1.X1.X2.X1.vout a_49002_22312# 0.383f
C1849 X2.X1.X1.X1.X2.X1.X3.vin2 a_31862_21352# 8.07e-19
C1850 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X3.vin1 0.0131f
C1851 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin1 0.195f
C1852 a_46502_28976# X2.X2.X1.X1.X1.X2.X3.vin1 0.52f
C1853 X2.X2.X1.X1.X1.X1.X1.vin2 a_46116_30882# 1.78e-19
C1854 X2.X1.X1.X2.X2.X2.X3.vin2 X2.X1.X2.vrefh 0.172f
C1855 a_31476_27070# a_31862_27070# 0.419f
C1856 a_4396_20446# X1.X1.X1.X1.X2.X2.X3.vin2 0.101f
C1857 X2.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.vrefh 0.117f
C1858 a_39966_25076# a_37766_24076# 4.77e-21
C1859 X2.X2.X3.vin2 a_49952_892# 0.239f
C1860 X2.X2.X1.X1.X1.X1.X3.vin1 a_48702_31882# 0.428f
C1861 a_48702_20446# X2.X2.X3.vin1 1.64e-19
C1862 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.X1.X3.vin1 1.22e-19
C1863 X2.X2.X1.X1.X2.X2.X3.vin2 a_49002_18540# 0.00846f
C1864 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X2.vout 0.0866f
C1865 X2.X3.vin1 X2.X3.vin2 0.514f
C1866 X1.X2.X2.X2.X1.X1.X1.vin1 a_25326_17452# 8.22e-20
C1867 X1.X2.X2.X2.X1.X1.X1.vin2 X1.X2.X2.X1.X2.X2.X3.vin2 3.94e-19
C1868 X1.X1.X3.vin2 a_5082_10916# 3.68e-19
C1869 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.vout 0.326f
C1870 a_2196_9916# X1.X1.X1.X2.X2.X1.X2.vin1 1.78e-19
C1871 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X1.vin2 0.1f
C1872 X1.X2.X1.X2.X2.X2.X3.vin2 a_17222_4198# 0.567f
C1873 a_8872_8828# a_10686_7922# 1.06e-19
C1874 X1.X1.X1.X2.X2.X2.vrefh a_2582_8010# 0.3f
C1875 a_38152_16452# a_37852_14586# 6.71e-19
C1876 X2.X1.X2.X1.X1.X2.vrefh a_40352_6016# 0.118f
C1877 a_10686_15546# X1.X1.X2.X1.X2.X2.X1.vin1 0.417f
C1878 a_46116_6104# X2.X2.X1.X2.X2.X2.X2.vin1 1.78e-19
C1879 X1.X1.X2.X1.X2.X2.X1.vin2 a_11072_15546# 0.12f
C1880 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X3.vin1 0.0174f
C1881 a_54606_30794# X2.X2.X2.X2.X2.X2.vrefh 8.22e-20
C1882 X2.X2.X1.X2.X1.X2.vrefh a_46116_15634# 0.118f
C1883 a_5082_29936# a_4396_28070# 3.31e-19
C1884 a_4696_29936# a_4782_28070# 3.38e-19
C1885 X1.X1.X3.vin1 a_5082_14688# 3.28e-19
C1886 a_31862_32788# a_34062_31882# 4.2e-20
C1887 X1.X1.X1.X1.X2.X2.vrefh a_2196_21352# 1.64e-19
C1888 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.X2.vin1 0.00117f
C1889 X2.X2.X3.vin2 a_52406_5016# 2.33e-19
C1890 a_11072_15546# a_11072_13640# 0.00396f
C1891 a_22826_6962# X1.X2.X2.X1.X1.X1.vout 0.386f
C1892 X1.X1.X2.X1.X2.X2.vout a_8872_16452# 0.36f
C1893 X1.X1.X2.X2.X1.X1.X3.vin2 a_11072_21264# 0.354f
C1894 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.vrefh 0.267f
C1895 a_8486_31700# a_10686_30794# 4.2e-20
C1896 X1.X2.X2.X1.X2.X1.X1.vin2 X2.X1.X1.X2.X2.vrefh 0.0128f
C1897 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 0.22f
C1898 X2.X2.X3.vin1 X2.X2.X2.X1.X1.X2.vout 1.71e-19
C1899 X1.X1.X2.X2.X2.X1.X3.vin1 a_8572_25982# 0.00251f
C1900 X1.X2.X1.X1.X1.X1.X1.vin2 a_17222_30882# 8.88e-20
C1901 a_16836_13728# a_17222_13728# 0.419f
C1902 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X2.X1.X2.X1.X2.X1.vin2 0.00232f
C1903 X1.X1.X2.X2.X1.X2.vout a_8572_22210# 0.0929f
C1904 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X3.vin1 0.206f
C1905 a_25712_30794# a_25712_28888# 0.00396f
C1906 X1.X1.X3.vin1 a_5082_7064# 9.8e-19
C1907 X1.X1.X2.X2.X2.X1.X1.vin2 a_10686_26982# 0.273f
C1908 X2.X1.X1.X1.X1.X2.X3.vin1 X2.X1.X1.X1.X1.X2.X3.vin2 0.587f
C1909 X1.X1.X2.X1.X2.X2.X3.vin2 a_10686_15546# 7.84e-19
C1910 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X1.vin1 0.0689f
C1911 a_8486_8828# a_8572_6962# 3.38e-19
C1912 a_52406_5016# a_52792_5016# 0.419f
C1913 X2.X1.X3.vin1 a_34062_5198# 2.12e-19
C1914 X1.X1.X2.X1.X1.X2.X1.vin2 a_11072_7922# 0.12f
C1915 a_10686_7922# X1.X1.X2.X1.X1.X2.X1.vin1 0.417f
C1916 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X2.vrefh 0.00118f
C1917 X2.X2.X1.X2.X2.X2.vrefh a_46116_8010# 0.118f
C1918 X2.X1.X2.X2.X2.X1.X1.vin1 a_40352_25076# 1.64e-19
C1919 a_31476_11822# a_31476_9916# 0.00396f
C1920 a_8186_25982# a_8486_24076# 4.41e-20
C1921 X1.X1.X2.X2.X2.X1.X3.vin2 a_8186_25982# 3.49e-19
C1922 X2.X1.X1.X2.X2.vrefh a_31862_9916# 8.22e-20
C1923 a_2582_25164# X1.X1.X1.X1.X2.X1.X1.vin2 0.273f
C1924 X1.X2.X1.X1.X2.X1.X3.vin2 a_17222_23258# 0.567f
C1925 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin2 7.84e-19
C1926 a_25326_7922# a_23212_6962# 2.68e-20
C1927 a_8186_22210# X1.X1.X2.X2.X1.X1.vout 0.387f
C1928 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X3.vin1 2.33e-19
C1929 a_33976_14688# X2.X1.X1.X2.X3.vin1 0.363f
C1930 a_25326_30794# X1.X2.X2.X2.X2.X2.vrefh 8.22e-20
C1931 a_52106_14586# a_52792_12640# 2.86e-19
C1932 a_17222_30882# a_19336_29936# 2.95e-20
C1933 X2.X2.X1.X3.vin1 X2.X2.X2.X3.vin2 1.22e-19
C1934 a_17222_17540# X1.X2.X1.X2.X1.X1.X1.vin2 0.273f
C1935 X1.X1.X2.X1.X3.vin2 a_8186_10734# 0.241f
C1936 X2.X2.X2.X1.X2.X1.X1.vin2 a_54606_11734# 0.273f
C1937 a_34062_31882# X2.X1.X1.X1.X1.X1.vout 0.422f
C1938 X1.X2.X1.X1.X2.X2.X1.vin2 a_17222_19446# 8.88e-20
C1939 X1.X2.X2.X1.X1.X1.X3.vin2 a_25712_6016# 0.354f
C1940 a_52492_6962# X2.X2.X2.X1.X1.X1.X3.vin2 0.00546f
C1941 X2.X1.X2.X1.X1.X1.X3.vin1 a_38152_5016# 0.199f
C1942 X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.vout 4.93e-20
C1943 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 0.234f
C1944 X2.X1.X2.X1.X2.X1.X3.vin1 a_37852_10734# 0.00251f
C1945 a_31476_19446# a_31476_17540# 0.00396f
C1946 X1.X2.X1.X1.X3.vin2 a_19336_22312# 0.363f
C1947 X1.X2.X2.X2.X1.X2.X1.vin1 a_25712_21264# 1.64e-19
C1948 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X3.vin1 0.206f
C1949 a_19036_9010# a_19336_7064# 6.1e-19
C1950 a_39966_28888# X2.X1.X2.X2.X2.X1.X2.vin1 0.402f
C1951 X2.X2.X2.X2.X3.vin1 a_52406_24076# 9.54e-19
C1952 a_34362_22312# a_34062_20446# 5.55e-20
C1953 X2.X1.X1.X1.X2.X2.vout a_33676_20446# 0.36f
C1954 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X3.vin2 0.0523f
C1955 a_19422_16634# a_17222_15634# 4.77e-21
C1956 X2.X2.X1.X1.X1.X1.X1.vin2 X2.X2.X1.X1.X1.X1.X2.vin1 0.242f
C1957 X1.X1.X2.X2.X1.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin2 0.0128f
C1958 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.X2.vin1 0.00117f
C1959 a_46502_17540# a_48702_16634# 4.2e-20
C1960 X2.X1.X1.X1.X1.X2.X2.vin1 a_31476_27070# 0.197f
C1961 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 0.139f
C1962 X2.X1.X2.X3.vin2 a_37466_18358# 0.263f
C1963 a_10686_11734# X1.X1.X2.X1.X1.X2.X3.vin2 8.07e-19
C1964 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.vout 0.398f
C1965 X2.X2.X3.vin1 a_52106_18358# 5.87e-20
C1966 a_25326_25076# X1.X2.X2.X2.X1.X2.X1.vin2 8.88e-20
C1967 X1.X1.X1.X1.X2.X2.X3.vin1 a_2582_19446# 0.00207f
C1968 X1.X2.X1.X1.X1.X1.X3.vin2 X1.X2.X1.X1.X1.X2.vrefh 0.165f
C1969 a_22826_22210# a_23512_20264# 2.86e-19
C1970 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X1.X2.X1.X2.X1.X1.vin1 0.668f
C1971 a_54992_28888# a_54992_26982# 0.00396f
C1972 a_37766_20264# a_37852_18358# 3.21e-19
C1973 X2.X1.X2.X2.X2.X1.vout X2.X1.X2.X2.X2.X1.X3.vin2 0.326f
C1974 X2.X1.X2.X2.X2.X2.X3.vin2 a_37766_31700# 0.277f
C1975 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X3.vin1 0.00117f
C1976 X1.X1.X1.X1.X1.X2.X3.vin2 X1.X1.X1.X1.X2.X1.X1.vin1 5.19e-19
C1977 a_5082_7064# X1.X1.X1.X2.X2.X2.X3.vin1 0.00874f
C1978 X1.X1.X1.X2.X1.X2.vrefh a_2196_15634# 0.118f
C1979 X1.X2.X1.X1.X1.X2.X3.vin2 a_16836_27070# 0.354f
C1980 a_19722_14688# a_19422_12822# 5.55e-20
C1981 a_19422_28070# a_17222_27070# 4.77e-21
C1982 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 0.581f
C1983 X2.X2.X1.X2.X1.X1.X2.vin1 X2.X2.X1.X2.X1.X2.vrefh 0.564f
C1984 X2.X2.X1.X2.X1.X2.vout X2.X2.X1.X2.X1.X2.X3.vin1 0.326f
C1985 a_19422_9010# a_17222_8010# 4.77e-21
C1986 a_2582_15634# X1.X1.X1.X2.X1.X2.X1.vin1 8.22e-20
C1987 X2.X1.X1.X1.X2.X2.vout X2.X1.X1.X1.X2.X2.X3.vin1 0.335f
C1988 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin2 0.12f
C1989 X1.X2.X2.X1.X2.X1.X1.vin1 a_25712_11734# 0.195f
C1990 X1.X2.X2.X1.X2.X2.vout a_22826_14586# 0.263f
C1991 a_22826_22210# X1.X2.X2.X2.X1.X1.X3.vin2 0.00815f
C1992 a_54992_26982# X2.X2.X2.X2.X2.vrefh 1.64e-19
C1993 a_39966_15546# a_40352_15546# 0.419f
C1994 X1.X2.X1.X1.X1.X1.X1.vin2 a_19422_31882# 0.00743f
C1995 a_17222_30882# X1.X2.X1.X1.X1.X2.X1.vin1 8.22e-20
C1996 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 0.0565f
C1997 a_10686_17452# a_8872_16452# 1.15e-20
C1998 a_19336_29936# X1.X2.X1.X1.X1.X2.vout 0.0929f
C1999 a_2582_19446# a_4696_18540# 4.72e-20
C2000 X2.X1.X2.X2.X3.vin2 a_37852_25982# 0.0927f
C2001 a_31862_27070# a_31862_25164# 0.00198f
C2002 X1.X2.X2.vrefh X3.vin1 0.0274f
C2003 a_8486_16452# a_8186_14586# 5.55e-20
C2004 a_31476_27070# X2.X1.X1.X1.X2.X1.X1.vin1 1.64e-19
C2005 X2.X1.X2.X2.vrefh a_40352_17452# 0.118f
C2006 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X3.vin1 2.33e-19
C2007 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X1.vout 0.038f
C2008 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 1.22e-19
C2009 X2.X2.X1.X2.X2.X1.X2.vin1 X2.X2.X1.X2.X2.X2.vrefh 0.564f
C2010 X2.X2.X1.X2.X1.X1.X3.vin2 a_46502_13728# 8.07e-19
C2011 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X3.vin2 0.552f
C2012 X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin2 6.26e-19
C2013 X2.X2.X3.vin2 X2.X2.X1.X2.X3.vin1 4.41e-19
C2014 a_19422_24258# X1.X2.X1.X1.X2.X1.X3.vin2 0.267f
C2015 a_39966_7922# a_40352_7922# 0.419f
C2016 a_52406_20264# X2.X2.X2.X2.X1.X1.X3.vin1 0.428f
C2017 X1.X1.X2.X1.X2.vrefh a_11072_9828# 0.118f
C2018 X2.X2.X2.X1.X2.X2.X3.vin2 a_52406_16452# 0.277f
C2019 a_19036_31882# a_19722_29936# 2.86e-19
C2020 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X3.vin1 0.00117f
C2021 a_19422_31882# a_19336_29936# 3.14e-19
C2022 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X2.vrefh 0.183f
C2023 X1.X2.X1.X2.X1.X2.X1.vin2 a_17222_11822# 8.88e-20
C2024 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X2.vin1 0.564f
C2025 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin2 0.12f
C2026 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin1 0.195f
C2027 X2.X2.X2.X1.X2.X2.X3.vin1 a_52106_14586# 0.00874f
C2028 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X3.vin1 0.00118f
C2029 a_16836_23258# X1.X2.X1.X1.X2.X2.X1.vin1 1.64e-19
C2030 a_17222_23258# a_17222_21352# 0.00198f
C2031 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X1.X2.vin1 0.564f
C2032 a_38152_24076# a_37852_22210# 6.71e-19
C2033 a_10686_6016# X1.X1.X2.X1.X1.X1.X3.vin2 0.567f
C2034 X2.X2.X3.vin1 a_49566_892# 0.17f
C2035 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 2.23e-19
C2036 X1.X2.X1.X2.X1.X2.X3.vin1 a_19422_12822# 0.42f
C2037 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X1.X2.X1.X2.X2.vrefh 0.1f
C2038 X1.X1.X2.X2.X2.X2.vout X1.X1.X2.X2.X3.vin2 0.0866f
C2039 a_34362_14688# X2.X1.X1.X2.X1.X2.X3.vin2 3.85e-19
C2040 X2.X1.X1.X2.X3.vin1 a_34062_12822# 9.54e-19
C2041 a_19036_16634# X1.X2.X1.X2.X1.X1.vout 0.359f
C2042 X1.X2.X2.X2.X2.X2.X3.vin1 a_23512_31700# 0.199f
C2043 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X2.vin1 0.0689f
C2044 a_31862_9916# a_33676_9010# 1.06e-19
C2045 X1.X1.X2.X3.vin2 a_8572_25982# 0.355f
C2046 X1.X1.X2.X2.X2.X1.vout X1.X1.X2.X2.X2.X1.X3.vin1 0.118f
C2047 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X2.X1.X1.X1.X2.vrefh 0.0128f
C2048 X1.X1.X2.X1.X2.X2.vrefh a_11072_13640# 0.118f
C2049 X2.X1.X3.vin1 X2.X1.X1.X3.vin2 1.04f
C2050 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.vrefh 2.33e-19
C2051 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.X3.vin1 1.22e-19
C2052 X1.X2.X2.X2.X1.X2.X3.vin1 a_23212_22210# 0.00329f
C2053 a_37766_20264# X2.X1.X2.X2.X1.X1.X3.vin1 0.428f
C2054 X2.X1.X1.X1.X2.X2.X2.vin1 X2.X1.X1.X2.vrefh 0.564f
C2055 X2.X2.X2.X2.X2.X1.X3.vin2 X2.X2.X2.X2.X2.X1.X3.vin1 0.581f
C2056 X2.X2.X2.X2.X2.X1.vout a_52492_29834# 0.169f
C2057 a_31476_23258# a_31862_23258# 0.419f
C2058 a_52492_6962# a_52792_5016# 6.1e-19
C2059 a_54606_7922# a_52492_6962# 2.68e-20
C2060 X1.X2.X2.X2.X2.X2.vrefh a_25712_28888# 0.118f
C2061 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X1.vin2 0.668f
C2062 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 0.587f
C2063 a_5082_22312# a_4396_20446# 3.31e-19
C2064 a_4696_22312# a_4782_20446# 3.38e-19
C2065 a_8186_18358# a_8572_18358# 0.416f
C2066 X2.X2.X2.X2.X2.X1.X1.vin1 a_54606_25076# 8.22e-20
C2067 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X1.X2.X3.vin2 3.94e-19
C2068 a_8572_29834# a_10686_28888# 2.95e-20
C2069 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X2.vrefh 0.076f
C2070 X2.vrefh X1.X2.X2.X2.X2.X2.X3.vin1 0.00118f
C2071 X2.X2.X2.X2.X1.X2.vrefh a_54606_21264# 0.3f
C2072 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X1.X2.X1.X1.X2.vrefh 0.1f
C2073 a_8572_14586# a_8486_12640# 3.14e-19
C2074 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X1.vout 0.399f
C2075 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 0.0903f
C2076 X1.X1.X1.X1.X1.X1.vout X1.X1.X1.X1.X1.X1.X3.vin2 0.342f
C2077 a_19036_9010# X1.X2.X1.X2.X2.X1.vout 0.359f
C2078 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin2 7.84e-19
C2079 a_46502_21352# a_48316_20446# 1.06e-19
C2080 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X2.vin1 0.0689f
C2081 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X1.X3.vin1 0.00789f
C2082 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 0.0903f
C2083 X1.X2.X2.X1.X1.X2.X1.vin1 a_25326_6016# 8.22e-20
C2084 X1.X2.X2.X1.X1.X2.X1.vin2 X1.X2.X2.X1.X1.X1.X3.vin2 3.94e-19
C2085 a_23126_20264# X1.X2.X2.X2.X1.X1.X3.vin1 0.428f
C2086 X1.X2.X1.X1.X2.X2.X2.vin1 X1.X2.X1.X2.vrefh 0.564f
C2087 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.vrefh 2.33e-19
C2088 X1.X2.X2.X2.X1.X2.X1.vin2 X1.X2.X2.X2.X1.X2.X1.vin1 0.668f
C2089 a_8486_20264# a_8572_18358# 3.21e-19
C2090 a_38152_8828# a_37466_6962# 3.31e-19
C2091 X2.X1.X2.vrefh X2.X2.X2.vrefh 0.0959f
C2092 X2.X1.X1.X2.X3.vin1 a_33976_10916# 0.17f
C2093 X2.X1.X1.X1.X1.X2.vrefh a_31476_30882# 0.118f
C2094 X2.X1.X2.X2.X1.X1.X3.vin2 a_37766_20264# 0.267f
C2095 a_54606_25076# a_52792_24076# 1.15e-20
C2096 a_33676_31882# a_33976_29936# 6.1e-19
C2097 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X3.vin1 0.00117f
C2098 a_14082_892# X1.X3.vin2 0.255f
C2099 a_4396_28070# X1.X1.X1.X1.X1.X2.X3.vin2 0.101f
C2100 X1.X2.X3.vin1 a_19422_16634# 2.92e-19
C2101 X1.X1.X1.X2.X1.X1.vout X1.X1.X1.X2.X3.vin1 0.131f
C2102 a_23212_25982# a_25326_25076# 4.72e-20
C2103 a_4696_29936# X1.X1.X1.X1.X3.vin1 0.363f
C2104 X1.X2.X2.X2.X2.X1.vout a_23212_25982# 1.64e-19
C2105 X2.X2.X2.X2.X1.X2.vout X2.X2.X2.X2.X1.X1.vout 0.507f
C2106 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X2.X1.X1.X1.vin1 0.206f
C2107 X1.X2.X2.X2.X3.vin2 X1.X2.X2.X3.vin2 0.17f
C2108 a_19336_7064# a_19036_5198# 6.71e-19
C2109 X1.X2.X2.X2.X2.X2.vout a_23212_29834# 0.0929f
C2110 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 0.0565f
C2111 X2.X1.X2.X1.X2.X2.X1.vin1 a_40352_13640# 1.64e-19
C2112 a_49002_26164# X2.X2.X1.X3.vin1 0.509f
C2113 X1.X1.X1.X1.X1.X2.X1.vin2 a_2582_27070# 8.88e-20
C2114 X1.X2.X2.X1.X1.X2.X3.vin1 a_22826_6962# 0.00874f
C2115 X2.X1.X1.X2.X3.vin2 a_34362_7064# 0.422f
C2116 a_31862_25164# a_31862_23258# 0.00198f
C2117 X1.X2.X2.X1.X2.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin2 0.0128f
C2118 X1.X2.X3.vin1 a_19422_9010# 2.12e-19
C2119 a_33976_18540# X2.X1.X1.X2.X1.X1.X3.vin1 0.00232f
C2120 X1.X2.X2.vrefh X2.X1.X2.vrefh 0.0959f
C2121 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.X1.X1.X1.vin1 5.19e-19
C2122 a_54992_30794# a_54992_28888# 0.00396f
C2123 a_2582_32788# X1.X1.X1.X1.X1.X1.X1.vin2 0.273f
C2124 a_52492_10734# a_52792_8828# 6.48e-19
C2125 X2.X2.X1.X2.X1.X2.X2.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 0.234f
C2126 a_48316_12822# a_48702_12822# 0.419f
C2127 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X2.vin1 0.242f
C2128 a_8486_31700# a_8572_29834# 3.38e-19
C2129 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.X1.vin2 8.93e-19
C2130 a_46502_21352# X2.X2.X1.X1.X2.X2.X1.vin2 0.273f
C2131 a_39966_9828# X2.X1.X2.X1.X1.X2.X3.vin1 0.00207f
C2132 X2.X1.X2.X1.X2.X2.X2.vin1 a_39966_15546# 8.88e-20
C2133 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X1.vin2 0.668f
C2134 a_2196_6104# a_2582_6104# 0.419f
C2135 a_48616_29936# X2.X2.X1.X1.X1.X2.X3.vin1 0.00329f
C2136 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X2.vrefh 2.33e-19
C2137 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X3.vin2 0.234f
C2138 X2.X2.X1.X1.X2.X1.vout X2.X2.X1.X1.X2.X1.X3.vin2 0.326f
C2139 a_10686_21264# X1.X1.X2.X2.X1.X1.X3.vin1 0.00207f
C2140 X1.X1.X2.X2.X2.X1.X3.vin2 a_11072_28888# 0.354f
C2141 a_8572_6962# X1.X1.X2.X1.X1.X1.X3.vin2 0.00546f
C2142 a_23126_27888# X1.X2.X2.X3.vin2 7.93e-20
C2143 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X3.vin1 0.206f
C2144 X1.X1.X2.X1.X1.X1.X3.vin2 a_8872_5016# 0.1f
C2145 X2.X1.X1.X1.X3.vin2 a_34062_24258# 0.00101f
C2146 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X2.vrefh 0.076f
C2147 a_34362_26164# X2.X1.X1.X1.X2.X1.X3.vin2 3.49e-19
C2148 a_54606_28888# a_52792_27888# 1.15e-20
C2149 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin2 7.84e-19
C2150 X1.X1.X1.X2.X1.X2.X3.vin1 a_4396_12822# 0.199f
C2151 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.vout 0.399f
C2152 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X2.vrefh 0.076f
C2153 X1.X2.X2.X1.X1.X2.X3.vin2 a_23512_8828# 0.101f
C2154 a_2582_6104# a_4782_5198# 4.2e-20
C2155 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.X2.vin1 0.00117f
C2156 a_46502_28976# X2.X2.X1.X1.X1.X2.X2.vin1 8.88e-20
C2157 X1.X1.X1.X3.vin1 X1.X1.X3.vin2 7.53e-21
C2158 X1.X2.X1.X2.X1.X1.X1.vin2 a_16836_15634# 1.78e-19
C2159 X2.X2.X2.X2.X1.X1.X3.vin2 X2.X2.X2.X2.X1.X1.X1.vin1 2.23e-19
C2160 X2.X2.X2.X2.X2.X2.X3.vin1 a_52492_29834# 0.00329f
C2161 X2.X1.X2.X2.X1.X2.X3.vin1 a_40352_23170# 0.354f
C2162 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X2.vrefh 0.267f
C2163 X2.X2.X2.X2.X1.X1.X2.vin1 a_54992_19358# 1.78e-19
C2164 a_48702_16634# X2.X2.X1.X2.X1.X1.vout 0.422f
C2165 X2.X2.X2.X1.X1.X1.X1.vin2 X2.X2.X2.X1.X1.X1.X1.vin1 0.668f
C2166 a_39966_25076# a_40352_25076# 0.419f
C2167 a_33676_24258# a_31862_23258# 1.15e-20
C2168 X2.X1.X2.X2.X2.X1.vout X2.X1.X2.X2.X3.vin2 0.399f
C2169 X1.X1.X1.X1.X2.X2.X3.vin2 a_2582_17540# 8.07e-19
C2170 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X2.vrefh 0.00118f
C2171 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.vout 0.118f
C2172 X2.X2.X2.X2.X1.X2.X1.vin1 a_54992_21264# 1.64e-19
C2173 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X2.X1.X1.X1.X2.vrefh 0.00437f
C2174 a_34362_18540# a_34062_16634# 5.25e-20
C2175 a_33976_18540# X2.X1.X1.X2.X1.X1.vout 1.64e-19
C2176 a_31862_25164# X2.X1.X1.X1.X2.X1.X1.vin1 0.417f
C2177 X1.X2.X1.X2.X1.X1.vout X1.X2.X1.X2.X1.X2.vout 0.507f
C2178 X1.X1.X1.X2.X2.X1.X3.vin1 a_2582_8010# 0.00207f
C2179 a_2196_25164# X1.X1.X1.X1.X2.X1.X2.vin1 1.78e-19
C2180 a_31476_25164# X2.X1.X1.X1.X2.X1.X3.vin1 0.354f
C2181 a_19036_20446# a_19336_18540# 6.48e-19
C2182 a_54606_17452# a_54992_17452# 0.419f
C2183 X2.X1.X2.X2.X1.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin2 0.0128f
C2184 a_4782_5198# X1.X1.X1.X2.X2.X2.X3.vin2 0.277f
C2185 a_48616_22312# a_49002_22312# 0.419f
C2186 X1.X2.X2.X1.X2.X1.X3.vin1 a_25326_11734# 0.52f
C2187 a_46502_17540# X2.X2.X1.X2.X1.X1.X1.vin1 0.417f
C2188 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X1.X3.vin2 1.22e-19
C2189 a_46116_17540# X2.X2.X1.X2.X1.X1.X3.vin1 0.354f
C2190 a_54606_11734# a_52492_10734# 5.36e-21
C2191 a_54606_25076# X2.X2.X2.X2.X1.X2.X1.vin2 8.88e-20
C2192 X1.X1.X1.X2.X2.X1.X3.vin2 a_4696_7064# 0.00546f
C2193 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X3.vin2 0.234f
C2194 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.vrefh 0.161f
C2195 X2.X2.X2.X2.X3.vin1 a_52106_22210# 0.436f
C2196 X2.X1.X2.X1.X1.X1.X1.vin2 a_39966_4110# 0.273f
C2197 X2.X2.X2.X1.X2.X1.X3.vin1 a_52106_10734# 0.00837f
C2198 a_10686_32700# a_8486_31700# 4.77e-21
C2199 X1.X2.X2.X1.X1.X1.vout a_23512_5016# 0.359f
C2200 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X2.vrefh 0.267f
C2201 a_31476_21352# X2.X1.X1.X1.X2.X2.X2.vin1 1.78e-19
C2202 a_48702_9010# X2.X2.X1.X2.X2.X1.vout 0.422f
C2203 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X3.vin1 0.00117f
C2204 X2.X1.X2.X1.X2.X1.X3.vin2 a_37766_12640# 0.267f
C2205 X1.X1.X1.X2.vrefh a_2196_19446# 0.118f
C2206 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 0.216f
C2207 a_52406_24076# a_52492_22210# 3.38e-19
C2208 a_52406_20264# a_54606_19358# 4.2e-20
C2209 a_4782_9010# X1.X1.X1.X2.X2.X1.vout 0.422f
C2210 X2.X2.X3.vin1 a_49002_14688# 3.28e-19
C2211 a_39966_26982# a_37852_25982# 5.36e-21
C2212 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 2.23e-19
C2213 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X1.vout 0.0524f
C2214 X1.X1.X1.X1.X1.X1.X3.vin2 a_2582_28976# 8.07e-19
C2215 X1.X2.X2.X2.X3.vin1 a_23212_22210# 0.363f
C2216 a_31862_15634# a_31862_13728# 0.00198f
C2217 X2.X2.X2.X2.X1.X2.X1.vin1 a_54992_23170# 0.195f
C2218 a_31476_15634# X2.X1.X1.X2.X1.X2.X1.vin1 1.64e-19
C2219 X1.X1.X2.X2.X3.vin2 X1.X1.X2.X2.X3.vin1 0.552f
C2220 a_25326_21264# a_23126_20264# 4.77e-21
C2221 a_52406_20264# X2.X2.X3.vin2 7.93e-20
C2222 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X3.vin1 1.22e-19
C2223 X2.X1.X1.X2.X1.X2.X3.vin2 a_34362_10916# 0.00846f
C2224 a_4696_18540# a_4396_16634# 6.2e-19
C2225 X2.X1.X2.X1.X1.X1.vout X2.X1.X2.X1.X1.X1.X3.vin2 0.342f
C2226 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X2.vin1 0.00117f
C2227 a_31862_25164# a_34062_24258# 4.2e-20
C2228 X1.X2.X2.X1.X1.X1.X1.vin2 X1.X2.X2.X1.X1.X1.X1.vin1 0.668f
C2229 a_33976_7064# a_31862_6104# 2.68e-20
C2230 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.vrefh 0.161f
C2231 a_46502_30882# X2.X2.X1.X1.X1.X2.X1.vin1 8.22e-20
C2232 X1.X1.X2.X1.X2.X1.X2.vin1 a_11072_11734# 1.78e-19
C2233 X1.X1.X2.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X1.vin1 2.23e-19
C2234 X1.X1.X3.vin2 X1.X1.X2.X1.X2.X2.X3.vin2 0.0011f
C2235 X2.X1.X1.X1.X1.X1.X3.vin1 a_31862_30882# 0.00207f
C2236 a_25326_9828# a_25712_9828# 0.419f
C2237 a_52492_10734# a_54606_9828# 4.72e-20
C2238 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin2 0.1f
C2239 X1.X1.X1.X2.X2.X1.X3.vin2 a_2582_8010# 0.567f
C2240 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin1 0.195f
C2241 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 0.242f
C2242 a_25326_9828# a_25326_7922# 0.00198f
C2243 a_17222_9916# X1.X2.X1.X2.X2.X1.X1.vin1 0.417f
C2244 a_16836_9916# X1.X2.X1.X2.X2.X1.X3.vin1 0.354f
C2245 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin2 0.12f
C2246 a_49002_18540# a_48316_16634# 2.97e-19
C2247 X2.X1.X1.X2.X1.X1.X3.vin2 a_34362_14688# 0.00815f
C2248 a_48616_18540# a_48702_16634# 3.21e-19
C2249 a_22826_14586# a_23512_12640# 2.86e-19
C2250 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X1.vin2 0.668f
C2251 X1.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X1.X3.vin2 0.0533f
C2252 X1.X2.X3.vin2 X1.X2.X1.X2.X2.X2.vout 1.5e-19
C2253 a_10686_4110# X1.X1.X2.X1.X1.X1.X1.vin1 0.417f
C2254 X1.X1.X2.X1.X1.X1.X1.vin2 a_11072_4110# 0.12f
C2255 X1.X1.X2.X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X1.vin2 0.076f
C2256 X2.X2.X2.X2.X2.X2.X3.vin1 a_54606_30794# 0.52f
C2257 a_54992_21264# X2.X2.X2.X2.X1.X1.X1.vin2 1.78e-19
C2258 X1.X1.X3.vin1 a_6032_892# 0.371f
C2259 X2.X2.X1.X1.X1.X1.X2.vin1 a_46116_30882# 0.197f
C2260 a_52406_8828# a_52106_6962# 5.55e-20
C2261 a_25326_32700# a_23512_31700# 1.15e-20
C2262 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 0.242f
C2263 a_54606_13640# a_54606_11734# 0.00198f
C2264 a_46116_23258# X2.X2.X1.X1.X2.X2.X1.vin1 1.64e-19
C2265 a_22826_10734# a_23126_8828# 4.41e-20
C2266 a_46502_23258# a_46502_21352# 0.00198f
C2267 a_33676_24258# a_34062_24258# 0.419f
C2268 X2.X1.X3.vin2 a_37766_5016# 2.33e-19
C2269 a_33976_10916# X2.X1.X1.X2.X3.vin2 0.0927f
C2270 X2.X1.X2.X1.X2.X1.X1.vin1 a_40352_9828# 1.64e-19
C2271 a_39966_21264# a_39966_19358# 0.00198f
C2272 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 0.242f
C2273 a_39966_32700# a_40352_32700# 0.419f
C2274 a_8572_25982# a_8872_24076# 6.48e-19
C2275 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.vout 0.398f
C2276 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X3.vin2 0.102f
C2277 a_31862_32788# X2.X1.X1.X1.X1.X1.X1.vin1 0.42f
C2278 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 0.581f
C2279 X2.X1.X2.X1.X2.X2.X3.vin1 a_38152_16452# 0.199f
C2280 a_31476_32788# X2.X1.X1.X1.X1.X1.X3.vin1 0.354f
C2281 a_19336_14688# a_17222_13728# 2.68e-20
C2282 X2.X1.X2.X1.X2.X2.vrefh a_40352_13640# 0.118f
C2283 a_37852_29834# a_38152_27888# 6.1e-19
C2284 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin1 0.195f
C2285 X1.X1.X1.X2.X2.X2.X1.vin2 a_2196_4198# 1.78e-19
C2286 X1.X2.X2.X2.X2.X1.X3.vin2 a_23126_27888# 0.267f
C2287 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X1.X3.vin1 0.00117f
C2288 X1.X2.X2.X1.X2.X2.X1.vin2 X2.X1.X1.X2.X1.X2.vrefh 0.0128f
C2289 a_10686_30794# X1.X1.X2.X2.X2.X1.X3.vin2 8.07e-19
C2290 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X2.vin1 0.564f
C2291 a_23212_6962# a_23126_5016# 3.14e-19
C2292 a_25326_32700# X2.vrefh 0.3f
C2293 X1.X2.X2.X2.X2.X2.X2.vin1 a_25712_32700# 0.197f
C2294 X1.X2.X3.vin1 a_19422_5198# 2.12e-19
C2295 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X2.X3.vin1 2.33e-19
C2296 X2.X1.X2.X2.X1.X1.X1.vin1 a_40352_17452# 1.64e-19
C2297 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin1 0.52f
C2298 a_22826_14586# a_23212_14586# 0.419f
C2299 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X3.vin1 1.22e-19
C2300 X2.X1.X2.X3.vin1 X2.X1.X1.X2.X3.vin2 7.46e-20
C2301 a_2196_11822# a_2582_11822# 0.419f
C2302 a_31476_13728# X2.X1.X1.X2.X1.X2.X2.vin1 1.78e-19
C2303 a_37466_18358# X2.X1.X2.X1.X2.X2.X3.vin2 0.00846f
C2304 a_40352_9828# a_40352_7922# 0.00396f
C2305 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X3.vin1 0.00117f
C2306 X2.X1.X2.X2.X1.X2.X3.vin2 a_37766_24076# 0.277f
C2307 X2.X2.X1.X2.X1.X1.X3.vin2 a_48616_14688# 0.00546f
C2308 X2.X1.X2.X1.X2.X1.vout a_38152_12640# 0.359f
C2309 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X3.vin1 0.199f
C2310 X1.X2.X1.X2.X1.X1.X2.vin1 X1.X2.X1.X2.X1.X2.vrefh 0.564f
C2311 a_23126_16452# X1.X2.X2.X1.X2.X2.X3.vin1 0.42f
C2312 a_52106_29834# X2.X2.X2.X2.X2.X1.X3.vin2 0.00815f
C2313 a_25326_26982# X1.X2.X2.X2.X2.vrefh 8.22e-20
C2314 X2.X2.X1.X2.X2.X2.X1.vin2 a_46116_4198# 1.78e-19
C2315 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X2.X1.X2.X2.vrefh 0.0128f
C2316 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 5.19e-19
C2317 X2.X1.X2.X1.X1.X2.X3.vin1 a_38152_8828# 0.199f
C2318 a_2582_9916# a_4396_9010# 1.06e-19
C2319 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X2.vrefh 0.076f
C2320 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X2.vin1 0.0689f
C2321 X2.X2.X2.X1.X1.X2.X1.vin2 X2.X2.X2.X1.X1.X1.X3.vin2 3.94e-19
C2322 X2.X2.X2.X1.X1.X2.X1.vin1 a_54606_6016# 8.22e-20
C2323 a_11072_13640# X1.X1.X2.X1.X2.X1.X1.vin2 1.78e-19
C2324 X1.X2.X2.X1.X1.X2.X1.vin2 X2.X1.X1.X2.X2.X2.vrefh 0.0128f
C2325 a_52492_18358# X2.X2.X2.X1.X2.X2.vout 7.93e-20
C2326 X1.X2.X2.vrefh a_20286_892# 7.23e-19
C2327 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X1.vin1 5.19e-19
C2328 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X2.vin1 0.0689f
C2329 a_46502_6104# a_48316_5198# 1.06e-19
C2330 X1.X1.X2.X2.X1.X2.X1.vin1 a_10686_21264# 8.22e-20
C2331 a_19722_22312# a_19036_20446# 3.31e-19
C2332 X1.X1.X2.X1.X2.X2.X1.vin1 a_11072_15546# 0.195f
C2333 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X1.X2.X2.X1.X1.X3.vin2 3.94e-19
C2334 a_19336_22312# a_19422_20446# 3.38e-19
C2335 a_54992_30794# X2.X2.X2.X2.X2.X2.vrefh 1.64e-19
C2336 a_52792_16452# a_54606_15546# 1.06e-19
C2337 X2.X2.X2.vrefh a_49952_892# 7.3e-19
C2338 a_5082_29936# X1.X1.X1.X1.X1.X2.X3.vin2 3.85e-19
C2339 X1.X1.X1.X1.X3.vin1 a_4782_28070# 9.54e-19
C2340 X2.X1.X1.X1.X1.X1.X3.vin1 a_34062_31882# 0.428f
C2341 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X1.vin1 0.267f
C2342 X1.X2.X1.X1.X2.X1.X3.vin2 a_19722_22312# 0.00815f
C2343 X1.X1.X1.X2.X1.X1.X3.vin2 a_2196_15634# 0.354f
C2344 a_52492_14586# a_54606_13640# 2.95e-20
C2345 a_25326_13640# a_25712_13640# 0.419f
C2346 X2.X2.X1.X1.X1.X2.vrefh X2.X1.X2.X2.X2.X2.vrefh 0.117f
C2347 X1.X2.X2.X1.X2.X1.X1.vin1 X2.X1.X1.X2.X2.vrefh 0.00437f
C2348 X1.X1.X1.X3.vin1 a_5082_18540# 0.389f
C2349 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.X1.vin1 0.206f
C2350 a_17222_13728# X1.X2.X1.X2.X1.X2.X1.vin1 0.417f
C2351 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.vout 0.08f
C2352 a_16836_13728# X1.X2.X1.X2.X1.X2.X3.vin1 0.354f
C2353 a_39966_28888# X2.X1.X2.X2.X2.X1.X1.vin2 8.88e-20
C2354 a_46116_21352# a_46116_19446# 0.00396f
C2355 a_2582_23258# a_4696_22312# 2.95e-20
C2356 X1.X2.X1.X2.X2.X1.X2.vin1 X1.X2.X1.X2.X2.X2.vrefh 0.564f
C2357 a_23126_8828# X1.X2.X2.X1.X1.X2.X3.vin1 0.42f
C2358 X1.X2.X2.X2.X1.X1.X3.vin1 a_22826_18358# 0.00837f
C2359 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X3.vin1 0.00118f
C2360 X1.X1.X2.X2.X2.X1.X1.vin2 a_11072_26982# 0.12f
C2361 a_10686_26982# X1.X1.X2.X2.X2.X1.X1.vin1 0.417f
C2362 X1.X1.X2.X1.X1.X2.X1.vin1 a_11072_7922# 0.195f
C2363 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X3.vin2 8.93e-19
C2364 X1.X2.X1.X1.X1.X2.vrefh a_16836_28976# 1.64e-19
C2365 X1.X1.X3.vin2 X1.X1.X1.X2.X2.X1.vout 4.93e-20
C2366 a_52792_8828# a_54606_7922# 1.06e-19
C2367 X2.X1.X2.X1.X1.X2.X3.vin2 a_37466_6962# 3.85e-19
C2368 a_8872_16452# a_8572_14586# 6.71e-19
C2369 a_31862_11822# a_31862_9916# 0.00198f
C2370 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X3.vin1 0.0174f
C2371 X1.X1.X1.X1.X1.X2.X2.vin1 a_2196_27070# 0.197f
C2372 a_31476_11822# X2.X1.X1.X2.X2.X1.X1.vin1 1.64e-19
C2373 X1.X1.X1.X1.X1.X1.X1.vin2 a_2582_30882# 8.88e-20
C2374 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X3.vin1 2.33e-19
C2375 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X1.vin2 0.216f
C2376 X2.X2.X1.X3.vin1 a_49002_22312# 7.98e-19
C2377 X2.X2.X1.X1.X1.X2.X2.vin1 a_46116_27070# 0.197f
C2378 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 1.22e-19
C2379 X2.X2.X2.X2.X1.X1.X1.vin2 a_54606_19358# 0.273f
C2380 a_52406_27888# X2.X2.X2.X2.X2.X1.X3.vin1 0.428f
C2381 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 0.581f
C2382 X2.X1.X1.X1.X1.X2.vout a_33976_26164# 7.93e-20
C2383 X2.X2.X2.X3.vin2 a_52492_25982# 0.355f
C2384 a_5082_14688# X1.X1.X1.X2.X1.X2.X3.vin1 0.00874f
C2385 a_25712_30794# X1.X2.X2.X2.X2.X2.vrefh 1.64e-19
C2386 a_16836_28976# X1.X2.X1.X1.X1.X2.X2.vin1 1.78e-19
C2387 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.X1.vin2 0.216f
C2388 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X2.vrefh 0.076f
C2389 X2.X2.X2.X1.X2.X1.X1.vin2 a_54992_11734# 0.12f
C2390 a_54606_11734# X2.X2.X2.X1.X2.X1.X1.vin1 0.417f
C2391 a_46502_28976# X2.X2.X1.X1.X1.X2.X1.vin2 0.273f
C2392 X2.X2.X1.X2.X1.X1.X1.vin2 a_46116_15634# 1.78e-19
C2393 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X2.vout 0.0866f
C2394 a_31476_19446# X2.X1.X1.X2.X1.X1.X1.vin1 1.64e-19
C2395 a_31862_19446# a_31862_17540# 0.00198f
C2396 a_19422_9010# a_19722_7064# 4.19e-20
C2397 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X1.X3.vin2 0.234f
C2398 a_10686_28888# X1.X1.X2.X2.X2.X1.X3.vin1 0.00207f
C2399 a_33676_5198# a_34062_5198# 0.419f
C2400 X2.X1.X1.X2.X2.X2.X2.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 0.234f
C2401 X1.X2.X1.X2.X2.X1.vout a_19336_7064# 0.169f
C2402 X1.X2.X3.vin2 a_19722_10916# 3.68e-19
C2403 X2.X1.X1.X1.X2.X2.vout X2.X1.X1.X1.X2.X2.X3.vin2 0.08f
C2404 a_8486_12640# X1.X1.X2.X1.X2.X1.X3.vin1 0.428f
C2405 X1.X1.X1.X2.X1.X2.X2.vin1 X1.X1.X1.X2.X2.vrefh 0.564f
C2406 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.X1.X1.vin2 3.94e-19
C2407 X2.X2.X1.X1.X1.X1.X1.vin2 a_48702_31882# 0.00743f
C2408 a_8186_14586# X1.X1.X2.X1.X3.vin2 0.423f
C2409 X2.X2.X1.X2.X1.X1.X3.vin1 a_48702_16634# 0.428f
C2410 a_33676_28070# a_31862_27070# 1.15e-20
C2411 X2.X1.X2.X1.X3.vin2 a_37766_12640# 0.00101f
C2412 a_52106_18358# a_52492_18358# 0.416f
C2413 X2.X2.X2.X3.vin1 a_52406_12640# 5.28e-19
C2414 a_10686_9828# X1.X1.X2.X1.X1.X2.X3.vin1 0.00207f
C2415 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.vrefh 0.161f
C2416 X1.X2.X2.X2.X1.X2.X2.vin1 a_25326_23170# 8.88e-20
C2417 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X1.vin2 8.93e-19
C2418 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.vrefh 0.161f
C2419 a_39966_15546# a_37852_14586# 2.68e-20
C2420 a_39966_11734# a_40352_11734# 0.419f
C2421 X2.X2.X2.X1.X2.X2.X1.vin2 a_54606_15546# 0.273f
C2422 a_4396_24258# X1.X1.X1.X1.X2.X1.X3.vin2 0.1f
C2423 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X2.vout 0.398f
C2424 a_2196_13728# a_2196_11822# 0.00396f
C2425 a_19036_5198# X1.X2.X1.X2.X2.X2.X3.vin2 0.101f
C2426 a_4696_26164# X1.X1.X1.X1.X3.vin2 0.0927f
C2427 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X2.vin1 0.242f
C2428 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 0.0565f
C2429 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X1.X2.X1.X2.X2.X3.vin2 3.94e-19
C2430 X1.X1.X2.X2.X1.X1.X1.vin1 a_10686_17452# 8.22e-20
C2431 a_34362_10916# X2.X1.X1.X2.X2.X1.X3.vin2 3.49e-19
C2432 X1.X1.X1.X1.X2.X1.X1.vin2 a_2196_23258# 1.78e-19
C2433 X1.X2.X3.vin1 a_19722_7064# 9.8e-19
C2434 X2.X2.X2.X1.X2.X1.X1.vin2 X2.X2.X2.X1.X1.X2.X3.vin2 3.94e-19
C2435 X2.X2.X2.X1.X2.X1.X1.vin1 a_54606_9828# 8.22e-20
C2436 a_48616_29936# X2.X2.X1.X1.X3.vin1 0.363f
C2437 a_8872_27888# a_8572_25982# 6.2e-19
C2438 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X3.vin1 0.0131f
C2439 a_4396_16634# a_4782_16634# 0.419f
C2440 a_54606_32700# X2.X2.X2.X2.X2.X2.X3.vin2 0.567f
C2441 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X1.vin2 0.668f
C2442 a_8486_31700# a_8872_31700# 0.419f
C2443 X1.X2.X2.X1.X2.X1.X1.vin2 X2.X1.X1.X2.X1.X2.X2.vin1 0.00232f
C2444 X2.X1.X2.X2.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin2 0.0128f
C2445 a_8572_10734# a_10686_9828# 4.72e-20
C2446 a_4696_18540# a_5082_18540# 0.413f
C2447 a_52106_22210# a_52492_22210# 0.419f
C2448 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X2.X3.vin2 8.93e-19
C2449 X3.vin2 a_43362_892# 0.472f
C2450 a_25326_6016# X1.X2.X2.X1.X1.X1.X3.vin1 0.00207f
C2451 X2.X2.X2.X1.X1.X2.X1.vin2 a_54606_7922# 0.273f
C2452 a_8872_8828# a_8186_6962# 3.31e-19
C2453 X1.X1.X2.X2.X2.X2.vrefh a_10686_28888# 0.3f
C2454 X1.X1.X2.X1.X2.X2.X3.vin2 a_8872_16452# 0.101f
C2455 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X2.vrefh 0.076f
C2456 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X2.vout 0.398f
C2457 X1.X2.X2.X3.vin1 a_23126_16452# 5.31e-19
C2458 X1.X2.X2.X1.X3.vin2 a_22826_10734# 0.241f
C2459 X2.X1.X1.X1.X1.X1.X3.vin2 a_31476_30882# 0.354f
C2460 a_54606_9828# a_54606_7922# 0.00198f
C2461 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 0.242f
C2462 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X3.vin1 1.22e-19
C2463 X2.X2.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X3.vin1 0.0321f
C2464 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin2 0.1f
C2465 X2.X1.X1.X1.X3.vin2 a_33976_22312# 0.363f
C2466 a_54606_15546# a_52492_14586# 2.68e-20
C2467 X2.X2.X1.X1.X2.X1.X3.vin2 a_48616_22312# 0.00546f
C2468 X1.X2.X2.X3.vin1 a_23126_8828# 1.64e-19
C2469 X1.X1.X2.X1.X2.X2.X2.vin1 a_11072_17452# 0.197f
C2470 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.vrefh 0.161f
C2471 X1.X2.X1.X1.X3.vin1 a_19336_26164# 0.169f
C2472 X2.X1.X2.X2.X3.vin1 a_37852_25982# 0.17f
C2473 a_38152_12640# a_37852_10734# 6.2e-19
C2474 vrefl X2.X2.X2.X2.X2.X2.X3.vin1 0.00118f
C2475 X1.X2.X1.X1.X1.X1.vout a_19722_29936# 0.386f
C2476 a_19422_31882# X1.X2.X1.X1.X3.vin1 1.52e-19
C2477 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X1.vin2 0.668f
C2478 a_54606_9828# X2.X2.X2.X1.X1.X2.X2.vin1 0.402f
C2479 X2.X2.X1.X3.vin1 X2.X2.X3.vin2 7.53e-21
C2480 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X1.vout 0.13f
C2481 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin1 0.52f
C2482 X2.X3.vin2 a_49952_892# 0.684f
C2483 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X2.vin1 0.242f
C2484 a_46502_32788# X2.X2.X1.X1.X1.X1.X3.vin2 7.84e-19
C2485 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin1 0.195f
C2486 X2.X1.X2.X2.X2.X1.X3.vin1 a_38152_27888# 0.199f
C2487 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X2.vrefh 0.267f
C2488 X1.X1.X3.vin1 X1.X1.X1.X2.X3.vin2 0.0816f
C2489 X1.X2.X2.X1.X2.X2.X1.vin2 X1.X2.X2.X1.X2.X1.X3.vin2 3.94e-19
C2490 X1.X2.X2.X1.X2.X2.X1.vin1 a_25326_13640# 8.22e-20
C2491 a_52406_24076# a_52792_24076# 0.419f
C2492 X1.X1.X1.X1.X2.X2.X1.vin2 a_2582_19446# 8.88e-20
C2493 X2.X1.X1.X2.X2.X1.X3.vin1 a_33676_9010# 0.199f
C2494 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X2.X1.X1.X2.X2.vrefh 0.0128f
C2495 a_16836_19446# a_16836_17540# 0.00396f
C2496 a_23126_12640# a_22826_10734# 5.25e-20
C2497 a_37466_18358# X2.X1.X3.vin2 0.451f
C2498 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X2.X1.X1.X1.X2.vrefh 0.00437f
C2499 X2.X1.X2.X3.vin2 a_37766_24076# 6.03e-19
C2500 X2.X1.X2.X1.X2.X2.vout X2.X1.X2.X1.X2.X1.vout 0.514f
C2501 a_49002_10916# X2.X2.X1.X2.X2.X1.X3.vin1 0.00837f
C2502 a_39966_6016# a_39966_4110# 0.00198f
C2503 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 0.242f
C2504 X2.X1.X2.X2.X2.X2.X1.vin1 a_39966_28888# 8.22e-20
C2505 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X1.X2.X2.X2.X1.X3.vin2 3.94e-19
C2506 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X3.vin2 8.93e-19
C2507 a_10686_26982# a_8572_25982# 5.36e-21
C2508 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 0.139f
C2509 X1.X1.X1.X1.X2.X2.vout a_4782_20446# 0.418f
C2510 a_5082_22312# X1.X1.X1.X1.X2.X2.X3.vin2 3.85e-19
C2511 X2.X2.X3.vin2 X2.X2.X1.X2.X2.X1.vout 4.93e-20
C2512 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 5.19e-19
C2513 a_8572_29834# X1.X1.X2.X2.X2.X1.X3.vin2 0.00546f
C2514 a_19036_28070# X1.X2.X1.X1.X1.X2.X3.vin2 0.101f
C2515 a_37466_18358# a_37766_16452# 4.41e-20
C2516 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X3.vin2 0.161f
C2517 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X3.vin2 1.42e-20
C2518 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X1.X2.X1.X1.X2.vrefh 0.267f
C2519 a_48316_9010# a_49002_7064# 2.86e-19
C2520 a_48702_9010# a_48616_7064# 3.14e-19
C2521 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 0.581f
C2522 X2.X1.X2.X1.X3.vin1 a_37852_10734# 0.169f
C2523 X2.X2.X1.X1.X2.X2.X3.vin1 a_48316_20446# 0.199f
C2524 a_46116_32788# a_46502_32788# 0.419f
C2525 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin2 7.84e-19
C2526 X1.X1.X3.vin1 a_4782_5198# 2.12e-19
C2527 X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X3.vin1 0.552f
C2528 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X1.X3.vin2 5.19e-19
C2529 X2.X1.X2.X1.X1.X1.vout a_37766_5016# 0.422f
C2530 a_19336_10916# a_19422_9010# 3.21e-19
C2531 a_19722_10916# a_19036_9010# 2.97e-19
C2532 a_25326_23170# a_25712_23170# 0.419f
C2533 a_40352_13640# a_40352_11734# 0.00396f
C2534 X1.X1.X3.vin1 a_4782_9010# 2.12e-19
C2535 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X3.vin2 0.552f
C2536 X2.X2.X2.X2.X1.X2.X3.vin2 a_52792_24076# 0.101f
C2537 X2.X1.X1.X1.X1.X1.vout a_33976_29936# 0.169f
C2538 a_34062_31882# a_34362_29936# 4.19e-20
C2539 a_39966_23170# a_39966_21264# 0.00198f
C2540 X1.X1.X2.X1.X2.X1.vout X1.X1.X2.X1.X2.X1.X3.vin2 0.326f
C2541 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin2 0.1f
C2542 a_2582_32788# a_4782_31882# 4.2e-20
C2543 a_23212_25982# X1.X2.X2.X2.X1.X2.X3.vin2 0.00535f
C2544 a_19722_7064# a_19422_5198# 5.55e-20
C2545 X1.X2.X1.X2.X2.X2.vout a_19036_5198# 0.36f
C2546 a_33676_31882# X2.X1.X1.X1.X1.X1.X3.vin2 0.1f
C2547 X2.X1.X1.X1.X2.X1.X3.vin1 a_31862_23258# 0.00207f
C2548 a_52406_20264# a_52792_20264# 0.419f
C2549 a_39966_23170# a_37852_22210# 2.68e-20
C2550 a_11072_32700# X1.X2.vrefh 0.118f
C2551 X2.X1.X3.vin2 X2.X1.X2.X1.X3.vin2 0.039f
C2552 X2.X2.X2.X1.X2.X2.vout a_52106_14586# 0.263f
C2553 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.X1.vin2 0.23f
C2554 a_10686_6016# a_11072_6016# 0.419f
C2555 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X3.vin2 0.449f
C2556 a_34926_892# X2.X3.vin1 0.354f
C2557 X1.X2.X2.X2.X2.X2.X3.vin1 a_25326_30794# 0.52f
C2558 a_48702_12822# X2.X2.X1.X2.X1.X2.X3.vin2 0.277f
C2559 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X1.X2.X2.X1.vin2 0.216f
C2560 X2.X1.X2.X1.X2.X2.X2.vin1 a_40352_15546# 1.78e-19
C2561 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.X1.vin1 2.23e-19
C2562 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.X3.vin1 0.587f
C2563 a_11072_26982# a_11072_25076# 0.00396f
C2564 a_33676_24258# a_33976_22312# 6.1e-19
C2565 a_2196_6104# X1.X1.X1.X2.X2.X2.X3.vin1 0.354f
C2566 a_2582_6104# X1.X1.X1.X2.X2.X2.X1.vin1 0.417f
C2567 a_39966_19358# a_37852_18358# 5.36e-21
C2568 a_54606_13640# X2.X2.X2.X1.X2.X1.X2.vin1 0.402f
C2569 X1.X2.X1.X1.X1.X1.X2.vin1 a_16836_30882# 0.197f
C2570 X1.X2.X2.X2.X2.X2.vout a_23512_31700# 0.36f
C2571 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X2.X3.vin1 0.0174f
C2572 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.vout 0.326f
C2573 X1.X1.X2.X2.X1.X1.X3.vin2 X1.X1.X2.X2.X1.X1.X3.vin1 0.581f
C2574 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X2.vrefh 0.00118f
C2575 X2.X2.X1.X1.X1.X2.vrefh a_46116_28976# 1.64e-19
C2576 a_4396_31882# a_4696_29936# 6.1e-19
C2577 X1.X1.X2.X2.X2.X1.vout a_8872_27888# 0.359f
C2578 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X2.vin1 0.564f
C2579 a_37766_16452# X2.X1.X2.X1.X3.vin2 9.7e-20
C2580 X2.X2.X1.X1.X1.X2.X1.vin2 a_46116_27070# 1.78e-19
C2581 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.X1.vin2 3.94e-19
C2582 X1.X2.X2.X2.X1.X2.vout a_23212_22210# 0.0929f
C2583 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 0.216f
C2584 a_37766_12640# a_39966_11734# 4.2e-20
C2585 a_37766_20264# a_38152_20264# 0.419f
C2586 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 0.587f
C2587 X1.X1.X2.X1.X1.X1.X1.vin2 X1.X2.X2.vrefh 0.0128f
C2588 X2.X2.X2.X2.X2.X1.X3.vin2 a_52792_27888# 0.1f
C2589 X1.X1.X2.X3.vin2 a_8572_18358# 0.0927f
C2590 X1.X2.X1.X3.vin2 X1.X2.X3.vin2 3.82e-19
C2591 X1.X1.X1.X2.X2.X2.X3.vin1 a_4782_5198# 0.42f
C2592 a_22826_18358# X1.X2.X2.X3.vin1 0.374f
C2593 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 2.23e-19
C2594 X2.X2.X1.X1.X1.X2.X3.vin1 X2.X2.X1.X1.X1.X2.X2.vin1 0.00117f
C2595 a_46502_28976# a_48702_28070# 4.2e-20
C2596 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X3.vin2 8.93e-19
C2597 X2.X1.X2.X2.X1.X2.X3.vin2 a_40352_25076# 0.354f
C2598 a_54606_4110# a_54992_4110# 0.419f
C2599 X2.X2.X1.X2.X3.vin2 X2.X2.X2.X1.X3.vin1 0.0604f
C2600 X2.X1.X1.X2.X2.X2.vrefh a_31862_6104# 8.22e-20
C2601 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.X1.X1.X3.vin1 1.22e-19
C2602 a_48316_31882# a_49002_29936# 2.86e-19
C2603 a_48702_31882# a_48616_29936# 3.14e-19
C2604 a_2582_25164# a_4396_24258# 1.06e-19
C2605 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X2.vin1 0.0689f
C2606 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X3.vin1 0.206f
C2607 a_23212_22210# a_25326_21264# 2.95e-20
C2608 X2.X1.X3.vin1 X2.X1.X1.X2.X1.X1.vout 2.91e-19
C2609 X1.X2.X1.X1.X2.X2.X3.vin2 a_19336_18540# 0.00504f
C2610 a_19422_20446# a_19722_18540# 4.41e-20
C2611 X2.X2.X2.X1.X2.X2.X3.vin2 a_54992_17452# 0.354f
C2612 X2.X2.vrefh X2.X2.X1.X1.X1.X1.X1.vin2 0.109f
C2613 a_52106_29834# a_52406_27888# 4.19e-20
C2614 X1.X2.X2.X1.X2.X1.X3.vin1 a_25712_11734# 0.354f
C2615 X2.X2.X1.X2.X3.vin1 a_48616_10916# 0.17f
C2616 a_49002_22312# X2.X2.X1.X1.X2.X2.vout 0.263f
C2617 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X3.vin1 0.206f
C2618 a_23126_20264# a_23512_20264# 0.419f
C2619 X2.X2.X2.X2.X1.X2.X2.vin1 a_54606_23170# 8.88e-20
C2620 a_22826_10734# X1.X2.X2.X1.X3.vin1 0.385f
C2621 a_25712_28888# a_25712_26982# 0.00396f
C2622 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X1.vin2 8.93e-19
C2623 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.vrefh 2.33e-19
C2624 X2.X1.X2.X2.X2.X2.X1.vin2 a_39966_30794# 0.273f
C2625 X3.vin1 a_28482_892# 0.426f
C2626 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.vout 0.0215f
C2627 X1.X1.X1.X1.X3.vin2 a_4782_24258# 0.00101f
C2628 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.X3.vin1 0.0131f
C2629 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X2.vin1 0.564f
C2630 X1.X1.X2.X2.X2.X2.X3.vin2 a_8486_31700# 0.277f
C2631 a_39966_4110# X2.X1.X2.X1.X1.X1.X1.vin1 0.417f
C2632 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X3.vin1 0.00117f
C2633 a_5082_26164# X1.X1.X1.X1.X2.X1.X3.vin2 3.49e-19
C2634 X2.X1.X2.X1.X1.X1.X1.vin2 a_40352_4110# 0.12f
C2635 X1.X1.X3.vin1 a_8486_12640# 8.66e-20
C2636 X1.X2.X3.vin2 a_23126_5016# 2.33e-19
C2637 a_31862_21352# a_33676_20446# 1.06e-19
C2638 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X2.vin1 0.0689f
C2639 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.X1.X1.X1.vin1 0.206f
C2640 X1.X1.X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X1.X2.X3.vin1 1.22e-19
C2641 a_54606_23170# X2.X2.X2.X2.X1.X2.vrefh 8.22e-20
C2642 X1.X2.X2.X1.X1.X2.vout a_22826_6962# 0.254f
C2643 a_54606_32700# a_52792_31700# 1.15e-20
C2644 a_23512_16452# a_25326_15546# 1.06e-19
C2645 X1.X2.X2.X2.X1.X1.X3.vin2 a_23126_20264# 0.267f
C2646 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X3.vin1 0.00117f
C2647 X1.X2.X1.X2.X1.X2.vrefh a_17222_15634# 0.3f
C2648 a_19336_14688# a_19722_14688# 0.419f
C2649 a_4696_18540# X1.X1.X1.X2.X1.X1.vout 1.64e-19
C2650 X2.X2.X1.X3.vin1 a_49002_18540# 0.389f
C2651 a_5082_18540# a_4782_16634# 5.25e-20
C2652 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X1.vout 0.399f
C2653 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 0.0903f
C2654 X2.X1.X1.X1.X2.X1.X3.vin1 a_34062_24258# 0.428f
C2655 a_25326_4110# a_25712_4110# 0.419f
C2656 a_8486_24076# a_10686_23170# 4.2e-20
C2657 a_33976_7064# X2.X1.X1.X2.X2.X2.X3.vin1 0.00329f
C2658 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 0.216f
C2659 X1.X2.X3.vin2 X1.X2.X2.X1.X2.X1.vout 3.2e-19
C2660 a_40352_17452# X2.X1.X2.X1.X2.X2.X1.vin2 1.78e-19
C2661 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X3.vin2 0.418f
C2662 X2.X1.X1.X2.X1.X2.vout a_33676_12822# 0.36f
C2663 X1.X2.X1.X2.X1.X1.X2.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 0.234f
C2664 a_10686_21264# a_8872_20264# 1.15e-20
C2665 X2.X1.X2.X2.X2.X2.vrefh a_39966_28888# 0.3f
C2666 X2.X1.X2.X2.X1.X1.X3.vin1 a_39966_19358# 0.52f
C2667 X2.X1.X2.X2.X1.X1.X2.vin1 a_40352_21264# 0.197f
C2668 a_48616_10916# a_48316_9010# 6.2e-19
C2669 a_2582_27070# X1.X1.X1.X1.X2.X1.X1.vin1 8.22e-20
C2670 X1.X2.X2.X1.X1.X2.X3.vin2 a_25712_9828# 0.354f
C2671 a_52492_10734# X2.X2.X2.X1.X1.X2.X3.vin2 0.00535f
C2672 X1.X1.X2.X2.X3.vin2 a_8486_27888# 0.00101f
C2673 a_2582_21352# X1.X1.X1.X1.X2.X2.X2.vin1 8.88e-20
C2674 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X1.vin1 0.0689f
C2675 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin1 0.52f
C2676 X1.X2.X2.X1.X1.X2.X3.vin2 a_25326_7922# 7.84e-19
C2677 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X1.vin2 0.668f
C2678 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.X1.X1.X1.vin1 5.19e-19
C2679 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X3.vin1 0.206f
C2680 X2.X2.X3.vin1 a_48702_16634# 2.92e-19
C2681 a_37852_10734# X2.X1.X2.X1.X1.X2.vout 7.93e-20
C2682 X2.X2.X1.X2.X1.X1.X3.vin2 a_46502_15634# 0.567f
C2683 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X1.vin1 5.19e-19
C2684 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X2.vin1 0.242f
C2685 X1.X2.X1.X2.X2.X2.vrefh a_17222_8010# 0.3f
C2686 a_23512_8828# a_25326_7922# 1.06e-19
C2687 X1.X1.X1.X1.X1.X1.X2.vin1 X1.X1.X1.X1.X1.X2.vrefh 0.564f
C2688 X2.X2.X2.X2.X2.X2.X3.vin1 a_54992_30794# 0.354f
C2689 X1.X1.X2.X1.X1.X1.X1.vin1 a_11072_4110# 0.195f
C2690 X2.X2.X2.X2.X2.X2.vout a_52492_29834# 0.0929f
C2691 a_19336_7064# X1.X2.X1.X2.X2.X2.vout 0.0929f
C2692 a_48316_31882# a_46502_30882# 1.15e-20
C2693 a_10686_25076# X1.X1.X2.X2.X1.X2.X3.vin1 0.00207f
C2694 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X2.X1.X1.X2.vrefh 0.0128f
C2695 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X2.vin1 0.564f
C2696 X1.X2.X2.X2.X2.X2.X3.vin2 a_23512_31700# 0.101f
C2697 X2.X2.X3.vin1 a_48702_9010# 2.12e-19
C2698 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X2.vrefh 0.076f
C2699 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X1.vin1 0.0689f
C2700 X1.X1.X1.X3.vin2 X1.X1.X2.X3.vin1 1.22e-19
C2701 X2.X2.X2.X1.X2.X1.X3.vin2 a_54606_11734# 7.84e-19
C2702 X1.X1.X3.vin1 X1.X1.X3.vin2 3.25f
C2703 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin2 0.12f
C2704 a_25326_23170# X1.X2.X2.X2.X1.X2.vrefh 8.22e-20
C2705 X1.X1.X1.X2.X2.X1.X1.vin2 a_2582_8010# 8.88e-20
C2706 X1.X2.X2.X2.X1.X1.X3.vin1 a_25326_19358# 0.52f
C2707 a_46116_27070# a_46116_25164# 0.00396f
C2708 X1.X2.X2.X3.vin1 a_23126_12640# 5.28e-19
C2709 X1.X2.X1.X2.X2.X1.X2.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 0.234f
C2710 a_34062_24258# X2.X1.X1.X1.X2.X1.vout 0.422f
C2711 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.X3.vin1 0.0174f
C2712 X2.X2.X1.X1.X2.vrefh a_46502_25164# 8.22e-20
C2713 a_25326_25076# X1.X2.X2.X2.X1.X2.X3.vin2 0.567f
C2714 a_5082_10916# X1.X1.X1.X2.X2.X1.X3.vin1 0.00837f
C2715 a_23512_12640# a_25326_11734# 1.06e-19
C2716 X1.X2.X1.X2.X2.vrefh a_17222_11822# 0.3f
C2717 a_52106_14586# X2.X2.X2.X1.X3.vin2 0.423f
C2718 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X1.vin1 0.0689f
C2719 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin2 0.12f
C2720 X2.X1.X2.X2.X1.X1.X3.vin2 a_39966_19358# 7.84e-19
C2721 X2.X1.X2.X2.X2.X2.X3.vin2 a_40352_32700# 0.354f
C2722 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X2.vrefh 0.597f
C2723 X2.X2.X2.X1.X2.X2.X1.vin2 X2.X2.X2.X1.X2.X1.X3.vin2 3.94e-19
C2724 X2.X2.X2.X1.X2.X2.X1.vin1 a_54606_13640# 8.22e-20
C2725 a_16836_8010# a_16836_6104# 0.00396f
C2726 X2.X2.X2.X1.X1.X1.X2.vin1 a_54992_6016# 0.197f
C2727 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X3.vin1 0.206f
C2728 a_19336_14688# X1.X2.X1.X2.X1.X2.X3.vin1 0.00329f
C2729 a_39966_17452# X2.X1.X2.X1.X2.X2.X3.vin2 0.567f
C2730 X2.X2.X1.X2.X2.X1.X3.vin2 a_46502_8010# 0.567f
C2731 a_52792_12640# a_52106_10734# 2.97e-19
C2732 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin1 0.52f
C2733 X1.X1.X1.X2.X1.X1.X3.vin2 a_5082_14688# 0.00815f
C2734 X1.X1.X1.X3.vin2 a_4782_12822# 6.03e-19
C2735 X1.X2.X2.X1.X2.X2.X1.vin1 X2.X1.X1.X2.X1.X2.vrefh 0.00437f
C2736 X2.X1.X2.X2.X3.vin1 a_37852_22210# 0.363f
C2737 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X1.vout 0.0524f
C2738 a_39966_26982# X2.X1.X2.X2.X2.vrefh 8.22e-20
C2739 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.vout 0.335f
C2740 X1.X2.X2.X2.X2.X2.X3.vin2 X2.vrefh 0.183f
C2741 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.vrefh 0.161f
C2742 a_52792_24076# a_52106_22210# 3.31e-19
C2743 X2.X2.X1.X2.vrefh a_46502_19446# 0.3f
C2744 a_4696_22312# X1.X1.X1.X1.X2.X2.vout 0.0929f
C2745 X2.X2.X1.X2.X1.X2.vout a_48702_12822# 0.418f
C2746 a_31862_13728# a_33676_12822# 1.06e-19
C2747 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X2.vin1 0.0689f
C2748 a_48616_26164# X2.X2.X1.X1.X3.vin2 0.0927f
C2749 a_54606_32700# X2.X2.X2.X2.X2.X2.X1.vin2 8.88e-20
C2750 X1.X1.X1.X1.X2.X2.X2.vin1 a_2196_19446# 0.197f
C2751 X1.X2.X2.X2.X2.X1.X1.vin1 a_25326_25076# 8.22e-20
C2752 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X1.X2.X3.vin2 3.94e-19
C2753 a_8486_5016# a_10686_4110# 4.2e-20
C2754 X1.X1.X2.X1.X1.X1.X3.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 0.22f
C2755 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X1.vin2 3.94e-19
C2756 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X3.vin1 0.00118f
C2757 X2.X1.X3.vin2 a_34362_14688# 2.04e-19
C2758 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X2.vin1 0.242f
C2759 X2.X2.X1.X2.X1.X1.vout X2.X2.X1.X2.X1.X2.vout 0.507f
C2760 a_16836_21352# X1.X2.X1.X1.X2.X2.X2.vin1 1.78e-19
C2761 X2.X1.X2.X2.X1.X2.X3.vin1 a_37466_22210# 0.00874f
C2762 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X2.X1.X2.X2.vrefh 0.00437f
C2763 a_25712_26982# X1.X2.X2.X2.X2.vrefh 1.64e-19
C2764 X1.X1.X1.X2.X2.X1.X3.vin1 a_4396_9010# 0.199f
C2765 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X1.X3.vin2 5.19e-19
C2766 a_48616_18540# a_49002_18540# 0.413f
C2767 X1.X2.X2.X1.X1.X2.X1.vin1 X2.X1.X1.X2.X2.X2.vrefh 0.00437f
C2768 X2.X1.X1.X1.X1.X1.X1.vin2 a_31862_30882# 8.88e-20
C2769 X1.X2.X2.vrefh d7 3.76e-19
C2770 a_31476_17540# a_31476_15634# 0.00396f
C2771 X2.X2.X1.X2.X2.X2.X3.vin1 a_48316_5198# 0.199f
C2772 X1.X2.X1.X1.X2.X2.vout a_19422_20446# 0.418f
C2773 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin2 7.84e-19
C2774 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X1.X3.vin2 5.19e-19
C2775 a_19722_22312# X1.X2.X1.X1.X2.X2.X3.vin2 3.85e-19
C2776 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X2.X1.X2.X1.X1.X2.vin1 0.00232f
C2777 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X2.X1.X1.vin1 0.668f
C2778 X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.vout 1.5e-19
C2779 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X1.vout 0.038f
C2780 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin2 0.12f
C2781 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X1.X3.vin1 0.0131f
C2782 X1.X2.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X3.vin1 0.0321f
C2783 a_25326_21264# X1.X2.X2.X2.X1.X1.X2.vin1 0.402f
C2784 a_5082_10916# X1.X1.X1.X2.X2.X1.X3.vin2 3.49e-19
C2785 a_8572_22210# a_8872_20264# 6.1e-19
C2786 a_10686_9828# X1.X1.X2.X1.X1.X2.X3.vin2 0.567f
C2787 a_52492_14586# X2.X2.X2.X1.X2.X1.X3.vin2 0.00546f
C2788 X1.X2.X2.X1.X2.X1.X3.vin2 a_25712_13640# 0.354f
C2789 a_19722_18540# X1.X2.X1.X3.vin2 0.233f
C2790 X2.X1.X2.X1.X2.X1.X3.vin2 a_37466_10734# 3.49e-19
C2791 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 0.242f
C2792 a_25326_32700# a_25326_30794# 0.00198f
C2793 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X3.vin1 0.206f
C2794 a_48316_16634# X2.X2.X1.X2.X1.X1.X3.vin2 0.1f
C2795 X2.X1.X2.X2.X2.X1.X3.vin2 X2.X1.X2.X2.X2.X1.X1.vin2 8.93e-19
C2796 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.vout 0.033f
C2797 X2.X1.X2.X2.X2.X1.X2.vin1 a_39966_26982# 8.88e-20
C2798 a_46502_21352# a_46502_19446# 0.00198f
C2799 a_4782_31882# a_2582_30882# 4.77e-21
C2800 X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin2 0.0128f
C2801 a_37466_29834# a_37852_29834# 0.419f
C2802 a_25712_6016# a_25712_4110# 0.00396f
C2803 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 2.23e-19
C2804 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X1.X3.vin1 0.00118f
C2805 X1.X1.X2.X2.X2.X1.X1.vin1 a_11072_26982# 0.195f
C2806 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X2.X1.X2.X2.X1.X2.vin1 0.00232f
C2807 X2.X1.X2.X1.X2.X2.X3.vin1 a_39966_15546# 0.52f
C2808 X1.X2.X1.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X1.vin1 0.267f
C2809 a_48316_5198# X2.X2.X1.X2.X2.X2.X3.vin2 0.101f
C2810 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X2.X1.X1.X2.X1.X1.vin2 0.00232f
C2811 a_16836_25164# a_17222_25164# 0.419f
C2812 a_4396_28070# a_2582_27070# 1.15e-20
C2813 X1.X2.X1.X2.X1.X2.X2.vin1 X1.X2.X1.X2.X2.vrefh 0.564f
C2814 X2.X1.X2.X1.X2.X2.vout a_38152_16452# 0.36f
C2815 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin2 0.12f
C2816 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X3.vin2 8.93e-19
C2817 a_23126_12640# X1.X2.X2.X1.X2.X1.X3.vin1 0.428f
C2818 X2.X1.X1.X2.X1.X1.X2.vin1 a_31476_15634# 0.197f
C2819 a_48316_28070# a_46502_27070# 1.15e-20
C2820 X2.X2.X2.X2.X1.X1.X1.vin2 a_54992_19358# 0.12f
C2821 a_54606_19358# X2.X2.X2.X2.X1.X1.X1.vin1 0.417f
C2822 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.vrefh 0.161f
C2823 a_31476_17540# a_31862_17540# 0.419f
C2824 X2.X2.X2.X3.vin1 X2.X2.X1.X2.X3.vin2 7.46e-20
C2825 X1.X2.X2.X1.X2.X2.X2.vin1 X2.X1.X1.X2.X1.X1.X1.vin2 0.00232f
C2826 a_37466_14586# X2.X1.X2.X1.X2.X1.vout 0.383f
C2827 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X3.vin2 0.546f
C2828 a_17222_28976# a_19036_28070# 1.06e-19
C2829 X1.X2.X2.X2.X1.X2.X3.vin1 a_23512_24076# 0.199f
C2830 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X2.X2.vin1 0.0689f
C2831 a_39966_6016# X2.X1.X2.X1.X1.X1.X2.vin1 0.402f
C2832 a_48316_9010# X2.X2.X1.X2.X2.X1.X3.vin2 0.1f
C2833 X2.X2.X2.X1.X2.X1.X1.vin1 a_54992_11734# 0.195f
C2834 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X2.X1.vin2 0.1f
C2835 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X1.vin2 3.94e-19
C2836 a_4396_9010# X1.X1.X1.X2.X2.X1.X3.vin2 0.1f
C2837 a_33976_29936# a_33676_28070# 6.71e-19
C2838 a_25326_21264# a_25326_19358# 0.00198f
C2839 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 0.242f
C2840 a_17222_32788# X1.X2.X1.X1.X1.X1.X1.vin2 0.273f
C2841 X1.X2.X2.X2.X2.X2.X3.vin1 a_22826_29834# 0.00874f
C2842 X2.X2.X1.X1.X1.X2.X3.vin1 X2.X2.X1.X1.X1.X2.X1.vin2 0.216f
C2843 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X2.X1.X1.X2.X2.vrefh 0.0128f
C2844 X1.X1.X3.vin1 X1.X3.vin1 0.273f
C2845 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X2.vrefh 0.00118f
C2846 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X1.X3.vin1 0.581f
C2847 a_34062_5198# X2.X1.X1.X2.X2.X2.X3.vin2 0.277f
C2848 X1.X2.X1.X2.X2.X1.vout X1.X2.X1.X2.X2.X2.vout 0.514f
C2849 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X3.vin1 0.199f
C2850 a_37766_27888# a_37852_25982# 3.21e-19
C2851 X2.X1.X1.X1.X1.X2.X3.vin2 a_31862_27070# 0.567f
C2852 a_33976_26164# X2.X1.X1.X3.vin1 0.356f
C2853 X2.X1.X2.X1.X1.X2.X3.vin1 a_39966_7922# 0.52f
C2854 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.X3.vin1 0.587f
C2855 X1.X2.X1.X1.X2.X2.vrefh a_17222_21352# 8.22e-20
C2856 a_23126_16452# X1.X2.X2.X1.X2.X2.vout 0.418f
C2857 X2.X1.X2.X2.X1.X1.X1.vin2 a_39966_19358# 0.273f
C2858 X2.X1.X1.X2.X2.X1.X2.vin1 a_31476_8010# 0.197f
C2859 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X1.vin1 2.23e-19
C2860 X1.X2.X2.X2.X1.X1.X1.vin1 a_25712_17452# 1.64e-19
C2861 X2.X1.X2.X1.X1.X2.vout a_38152_8828# 0.36f
C2862 X1.X2.X2.X2.X1.X2.X2.vin1 a_25712_23170# 1.78e-19
C2863 X2.X2.X2.X1.X3.vin1 a_52406_8828# 9.54e-19
C2864 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X1.X3.vin1 0.0425f
C2865 X2.X1.X3.vin2 a_34926_892# 0.0927f
C2866 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X2.vout 0.197f
C2867 X1.X2.X3.vin1 a_22826_14586# 2.24e-19
C2868 a_54606_15546# X2.X2.X2.X1.X2.X2.X1.vin1 0.417f
C2869 X2.X2.X2.X1.X2.X2.X1.vin2 a_54992_15546# 0.12f
C2870 X1.X1.X1.X1.X2.X1.vout X1.X1.X1.X1.X2.X1.X3.vin2 0.326f
C2871 X1.X3.vin2 a_20672_892# 0.684f
C2872 a_2582_13728# a_2582_11822# 0.00198f
C2873 X2.X1.X1.X1.X1.X2.vout X2.X1.X1.X1.X1.X2.X3.vin1 0.326f
C2874 X2.X1.X1.X1.X1.X1.X1.vin2 a_34062_31882# 0.00743f
C2875 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X3.vin2 0.418f
C2876 a_31862_17540# X2.X1.X1.X2.X1.X1.X2.vin1 8.88e-20
C2877 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 5.19e-19
C2878 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X1.X3.vin1 0.0425f
C2879 a_8486_12640# a_8186_10734# 5.25e-20
C2880 X2.X1.X1.X1.X2.X2.vrefh a_31476_23258# 0.118f
C2881 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 5.19e-19
C2882 a_2196_9916# a_2582_9916# 0.419f
C2883 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X2.vrefh 2.33e-19
C2884 X1.X2.X2.X2.X1.X1.X1.vin2 a_25326_19358# 0.273f
C2885 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin2 0.12f
C2886 a_37852_18358# a_38152_16452# 6.48e-19
C2887 X1.X1.X1.X2.X2.X2.vrefh a_2582_6104# 8.22e-20
C2888 a_4782_16634# X1.X1.X1.X2.X1.X1.vout 0.422f
C2889 a_23512_20264# a_22826_18358# 2.97e-19
C2890 a_23126_8828# X1.X2.X2.X1.X1.X2.vout 0.418f
C2891 a_8572_10734# X1.X1.X2.X1.X1.X2.X3.vin2 0.00535f
C2892 X1.X1.X3.vin2 a_8486_5016# 2.33e-19
C2893 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X3.vin2 0.0523f
C2894 a_10686_13640# X1.X1.X2.X1.X2.X1.X3.vin2 0.567f
C2895 a_5082_18540# X1.X1.X3.vin1 0.47f
C2896 a_19722_22312# X1.X2.X1.X1.X2.X2.X3.vin1 0.00874f
C2897 a_11072_17452# a_11072_15546# 0.00396f
C2898 a_54606_7922# X2.X2.X2.X1.X1.X2.X1.vin1 0.417f
C2899 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X2.vrefh 0.00118f
C2900 X2.X2.X2.X1.X1.X2.X1.vin2 a_54992_7922# 0.12f
C2901 X1.X2.X2.X1.X1.X1.X3.vin2 X1.X2.X2.X1.X1.X1.X3.vin1 0.581f
C2902 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X1.X3.vin2 1.22e-19
C2903 X1.X1.X2.X2.X2.X2.vrefh X1.X1.X2.X2.X2.X1.X3.vin2 0.161f
C2904 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X1.X3.vin1 0.0321f
C2905 a_49002_29936# a_48316_28070# 3.31e-19
C2906 a_22826_29834# X1.X2.X2.X2.X3.vin2 0.422f
C2907 a_48616_29936# a_48702_28070# 3.38e-19
C2908 a_22826_14586# X1.X2.X2.X1.X2.X1.X3.vin2 0.00815f
C2909 X1.X1.X2.X3.vin1 a_8486_8828# 1.64e-19
C2910 a_37766_31700# a_37466_29834# 5.55e-20
C2911 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X2.vout 0.398f
C2912 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin2 0.1f
C2913 X1.X1.X2.X2.X1.X1.X1.vin2 a_10686_19358# 0.273f
C2914 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X3.vin2 8.93e-19
C2915 a_52406_27888# a_52792_27888# 0.419f
C2916 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X1.vin1 0.0689f
C2917 X2.X2.X2.X1.X1.X2.X3.vin2 a_54606_7922# 7.84e-19
C2918 X2.X2.X2.X2.X2.X1.X3.vin1 a_52492_25982# 0.00251f
C2919 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X2.vout 0.0866f
C2920 X1.X2.X2.X2.X1.X1.X3.vin2 a_22826_18358# 3.49e-19
C2921 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X3.vin1 1.42e-20
C2922 X2.X1.X3.vin2 a_34362_10916# 3.68e-19
C2923 a_49002_18540# X2.X2.X1.X2.X1.X1.X3.vin1 0.00837f
C2924 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X3.vin1 0.199f
C2925 X2.X2.X2.X3.vin2 a_52492_18358# 0.0927f
C2926 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 0.234f
C2927 a_25326_13640# a_25326_11734# 0.00198f
C2928 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 0.242f
C2929 X2.X1.X2.X2.X2.X1.X2.vin1 a_40352_28888# 0.197f
C2930 a_10686_28888# a_8872_27888# 1.15e-20
C2931 a_8486_12640# a_8872_12640# 0.419f
C2932 X2.X2.X1.X1.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X1.X3.vin2 0.581f
C2933 a_16836_30882# a_17222_30882# 0.419f
C2934 a_2582_28976# X1.X1.X1.X1.X1.X2.X2.vin1 8.88e-20
C2935 a_31862_28976# X2.X1.X1.X1.X1.X2.X3.vin1 0.52f
C2936 a_22826_29834# a_23126_27888# 4.19e-20
C2937 a_25326_11734# a_23212_10734# 5.36e-21
C2938 X2.X1.X1.X2.X2.X1.X1.vin2 a_31476_8010# 1.78e-19
C2939 a_11072_11734# a_11072_9828# 0.00396f
C2940 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X2.vin1 0.564f
C2941 X1.X1.X3.vin2 a_8186_10734# 6.66e-19
C2942 a_25712_25076# X1.X2.X2.X2.X1.X2.X1.vin2 1.78e-19
C2943 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 5.19e-19
C2944 a_33676_28070# a_34062_28070# 0.419f
C2945 a_28096_892# X3.vin2 0.0927f
C2946 X2.X1.X1.X1.X1.X2.X2.vin1 X2.X1.X1.X1.X1.X2.X3.vin2 0.234f
C2947 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.vout 0.118f
C2948 a_17222_19446# a_17222_17540# 0.00198f
C2949 a_16836_19446# X1.X2.X1.X2.X1.X1.X1.vin1 1.64e-19
C2950 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X2.X1.X1.X2.X2.vrefh 0.00437f
C2951 a_46116_8010# a_46116_6104# 0.00396f
C2952 X2.X2.vrefh X2.X1.X2.X2.X2.X2.X3.vin1 0.00118f
C2953 a_39966_17452# a_37766_16452# 4.77e-21
C2954 X2.X1.X3.vin1 a_34362_7064# 9.8e-19
C2955 X2.X1.X2.X1.X1.X1.X3.vin2 a_39966_4110# 7.84e-19
C2956 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X1.vin1 0.0689f
C2957 a_2196_23258# a_2196_21352# 0.00396f
C2958 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin2 7.84e-19
C2959 X1.X1.X1.X1.X1.X2.vout a_4396_28070# 0.36f
C2960 X1.X1.X3.vin1 X1.X1.X1.X2.X1.X2.vout 3.08e-19
C2961 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 0.0565f
C2962 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin1 0.449f
C2963 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X1.X3.vin2 5.19e-19
C2964 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X1.X2.X2.X2.X2.X1.vin1 0.668f
C2965 X1.X2.X2.X1.X1.X1.vout a_23212_6962# 0.169f
C2966 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.vout 0.335f
C2967 a_33976_10916# a_31862_9916# 5.36e-21
C2968 a_16836_9916# X1.X2.X1.X2.X2.X1.X2.vin1 1.78e-19
C2969 X2.X2.X2.X2.X2.vrefh a_54606_25076# 0.3f
C2970 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X2.vout 0.197f
C2971 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X3.vin1 0.0131f
C2972 a_54606_32700# a_54992_32700# 0.419f
C2973 X2.X1.X2.vrefh a_34926_892# 7.23e-19
C2974 X1.X1.X3.vin1 a_8186_6962# 6.45e-19
C2975 X2.X1.X1.X2.X2.X1.X3.vin2 a_31862_6104# 8.07e-19
C2976 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 0.587f
C2977 X2.X2.X1.X2.X2.X1.vout a_49002_7064# 0.383f
C2978 a_4396_28070# a_4696_26164# 6.48e-19
C2979 a_46116_32788# X2.X2.X1.X1.X1.X1.X3.vin1 0.354f
C2980 a_46502_32788# X2.X2.X1.X1.X1.X1.X1.vin1 0.42f
C2981 a_2196_13728# a_2582_13728# 0.419f
C2982 a_25326_6016# a_23512_5016# 1.15e-20
C2983 X1.X2.X1.X2.X3.vin2 a_19422_9010# 0.00101f
C2984 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X3.vin1 0.00118f
C2985 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X3.vin1 0.0131f
C2986 X2.X1.X2.X1.X3.vin2 a_37466_10734# 0.241f
C2987 a_17222_6104# X1.X2.X1.X2.X2.X2.X2.vin1 8.88e-20
C2988 X1.X1.X2.X3.vin2 a_8486_24076# 6.03e-19
C2989 X2.X1.X1.X1.X1.X1.vout X2.X1.X1.X1.X3.vin1 0.13f
C2990 X1.X1.X2.X1.X2.X2.vout X1.X1.X2.X1.X2.X1.vout 0.514f
C2991 a_39966_23170# X2.X1.X2.X2.X1.X1.X3.vin2 8.07e-19
C2992 X2.X2.X1.X1.X3.vin2 a_48616_22312# 0.363f
C2993 X1.X2.X3.vin2 a_20672_892# 0.239f
C2994 X2.vrefh X2.X1.X1.X1.X1.X1.X1.vin1 0.108f
C2995 a_8186_29834# X1.X1.X2.X2.X2.X1.vout 0.383f
C2996 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.vout 0.326f
C2997 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.vout 0.326f
C2998 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X1.vin2 3.94e-19
C2999 X1.X1.X2.X2.X1.X1.vout a_8572_22210# 0.169f
C3000 X1.X1.X1.X1.X1.X1.X3.vin1 a_4782_31882# 0.428f
C3001 X1.X2.X2.X2.X1.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin1 0.00437f
C3002 X2.X1.X2.X2.X2.X1.vout a_37766_27888# 0.422f
C3003 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.X1.X1.vin1 5.19e-19
C3004 a_34362_14688# X2.X1.X1.X2.X1.X2.vout 0.254f
C3005 X1.X2.X1.X2.X2.X2.vout X1.X2.X1.X2.X2.X2.X3.vin2 0.08f
C3006 X2.X1.X1.X1.X1.X1.vout X2.X1.X1.X1.X1.X1.X3.vin2 0.342f
C3007 X1.X1.X2.X1.X3.vin2 a_8572_10734# 0.0927f
C3008 a_10686_28888# a_10686_26982# 0.00198f
C3009 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X3.vin1 0.00118f
C3010 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X1.vin2 0.242f
C3011 a_8486_12640# a_10686_11734# 4.2e-20
C3012 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 0.216f
C3013 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 0.216f
C3014 a_8186_18358# a_8486_16452# 4.41e-20
C3015 a_39966_19358# X2.X1.X2.X2.vrefh 8.22e-20
C3016 a_52406_12640# a_54606_11734# 4.2e-20
C3017 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X3.vin1 0.0131f
C3018 X2.X1.X1.X2.X1.X2.vrefh a_31862_13728# 8.22e-20
C3019 a_2582_17540# X1.X1.X1.X2.X1.X1.X1.vin2 0.273f
C3020 X1.X2.X1.X2.X1.X1.X3.vin2 a_17222_15634# 0.567f
C3021 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin1 0.195f
C3022 X1.X2.X3.vin1 X1.X2.X1.X2.X3.vin2 0.0816f
C3023 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin2 7.84e-19
C3024 X2.X2.X2.X2.X1.X2.X3.vin1 a_54606_23170# 0.52f
C3025 X1.X1.X2.X1.X1.X1.X3.vin2 a_11072_6016# 0.354f
C3026 X1.X2.X2.X2.X2.X2.X3.vin1 a_25712_30794# 0.354f
C3027 X2.X1.X2.X3.vin2 X2.X1.X3.vin2 0.171f
C3028 X2.X2.X3.vin1 X2.X2.X3.vin2 3.25f
C3029 X2.X2.X1.X3.vin2 X2.X2.X2.X3.vin1 1.22e-19
C3030 a_25326_28888# X1.X2.X2.X2.X2.X1.X2.vin1 0.402f
C3031 X2.X1.X1.X1.X2.X1.vout a_33976_22312# 0.169f
C3032 a_34062_24258# a_34362_22312# 4.19e-20
C3033 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X3.vin1 0.206f
C3034 X2.X2.X1.X1.X2.X1.X2.vin1 a_46116_23258# 0.197f
C3035 a_2582_11822# X1.X1.X1.X2.X2.X1.X1.vin1 8.22e-20
C3036 a_19036_31882# a_17222_30882# 1.15e-20
C3037 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 0.234f
C3038 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X1.vin1 0.267f
C3039 a_23212_22210# a_23512_20264# 6.1e-19
C3040 a_4782_31882# a_5082_29936# 4.19e-20
C3041 X1.X1.X1.X1.X1.X1.vout a_4696_29936# 0.169f
C3042 a_16836_25164# a_16836_23258# 0.00396f
C3043 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X2.vrefh 0.00118f
C3044 a_37466_25982# a_38152_24076# 3.08e-19
C3045 a_8572_10734# X1.X1.X2.X1.X1.X2.vout 7.93e-20
C3046 X2.X2.X2.X3.vin1 a_52406_16452# 5.31e-19
C3047 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X2.X1.X1.vin1 0.206f
C3048 X1.X2.X2.X2.X1.X1.X1.vin2 X1.X2.X2.X2.vrefh 0.1f
C3049 X1.X1.X2.X1.X1.X1.X1.vin1 X1.X2.X2.vrefh 0.00437f
C3050 X1.X2.X1.X2.X1.X2.vout a_19422_12822# 0.418f
C3051 X2.X1.X3.vin1 a_34062_12822# 2.12e-19
C3052 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X2.X3.vin2 2.23e-19
C3053 X2.X2.X1.X1.X1.X2.X3.vin1 a_48702_28070# 0.42f
C3054 a_25326_17452# X1.X2.X2.X1.X2.X2.X1.vin2 8.88e-20
C3055 X1.X2.X1.X2.X2.X1.X3.vin2 a_17222_8010# 0.567f
C3056 a_2196_19446# a_2196_17540# 0.00396f
C3057 X1.X1.X1.X1.X1.X1.X2.vin1 X1.X1.X1.X1.X1.X1.X3.vin2 0.234f
C3058 X2.X2.X2.X3.vin1 a_52406_8828# 1.64e-19
C3059 X2.X2.X2.X2.X2.X1.X1.vin1 a_54992_25076# 1.64e-19
C3060 a_23212_25982# a_23126_24076# 3.3e-19
C3061 X2.X2.X2.X2.X1.X2.vrefh a_54992_21264# 0.118f
C3062 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X3.vin1 2.33e-19
C3063 a_8186_6962# X1.X1.X2.X1.X1.X1.vout 0.386f
C3064 X2.X2.X1.X1.X1.X1.vout a_49002_29936# 0.386f
C3065 a_48702_31882# X2.X2.X1.X1.X3.vin1 1.52e-19
C3066 a_46116_11822# a_46116_9916# 0.00396f
C3067 X1.X2.X2.X1.X2.X2.vout X1.X2.X2.X1.X3.vin2 0.0866f
C3068 X2.X1.X2.X2.X2.X1.X3.vin2 a_37466_25982# 3.49e-19
C3069 a_23212_22210# X1.X2.X2.X2.X1.X1.X3.vin2 0.00546f
C3070 X1.X1.X1.X1.X2.X1.X3.vin1 a_4396_24258# 0.199f
C3071 X2.X2.X1.X2.X2.vrefh a_46502_9916# 8.22e-20
C3072 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X3.vin2 8.93e-19
C3073 X2.X2.X2.X2.X2.X1.vout X2.X2.X2.X2.X2.X1.X3.vin1 0.118f
C3074 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X3.vin2 0.552f
C3075 a_37466_6962# a_38152_5016# 2.86e-19
C3076 X2.X2.X1.X1.X2.X2.vrefh a_46502_21352# 8.22e-20
C3077 X1.X2.X2.X1.X1.X2.X1.vin1 a_25712_6016# 1.64e-19
C3078 X2.X1.X2.X2.X2.X2.X1.vin2 a_40352_30794# 0.12f
C3079 a_39966_30794# X2.X1.X2.X2.X2.X2.X1.vin1 0.417f
C3080 X2.X2.X2.X2.X1.X2.X2.vin1 a_54992_23170# 1.78e-19
C3081 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X1.X2.X2.vrefh 0.1f
C3082 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X1.vin1 2.23e-19
C3083 X1.X1.X2.X1.X1.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin2 0.0128f
C3084 a_8486_16452# X1.X1.X2.X1.X3.vin2 9.7e-20
C3085 X2.X1.X2.X1.X1.X1.X1.vin1 a_40352_4110# 0.195f
C3086 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin2 7.84e-19
C3087 X2.X1.X1.X1.X2.X2.X3.vin1 a_33676_20446# 0.199f
C3088 X2.X2.X1.X2.vrefh a_46502_17540# 8.22e-20
C3089 a_48316_12822# a_49002_10916# 3.08e-19
C3090 a_48702_12822# a_48616_10916# 3.3e-19
C3091 X2.X2.X2.X1.X3.vin1 a_52106_6962# 0.436f
C3092 a_52492_14586# a_52406_12640# 3.14e-19
C3093 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 0.139f
C3094 X1.X2.X2.X1.X2.X1.X1.vin1 a_25326_9828# 8.22e-20
C3095 X1.X2.X2.X1.X2.X1.X1.vin2 X1.X2.X2.X1.X1.X2.X3.vin2 3.94e-19
C3096 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.vout 0.038f
C3097 a_54992_23170# X2.X2.X2.X2.X1.X2.vrefh 1.64e-19
C3098 X2.X1.X1.X1.X2.X1.X1.vin2 a_31862_23258# 8.88e-20
C3099 X1.X2.X1.X1.X1.X1.X3.vin2 a_19336_29936# 0.00546f
C3100 X2.X2.X2.X2.X2.X2.X3.vin2 a_52792_31700# 0.101f
C3101 X1.X1.X2.X2.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin2 0.0128f
C3102 a_19722_14688# X1.X2.X1.X2.X3.vin1 0.436f
C3103 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin2 1.42e-20
C3104 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X2.vin1 0.564f
C3105 X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.vout 2.91e-19
C3106 X2.X1.X1.X1.X2.vrefh X1.X2.X2.X2.X2.vrefh 0.117f
C3107 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X1.vin2 0.076f
C3108 X2.X2.X1.X1.X2.X2.vrefh X2.X1.X2.X2.X1.X2.vrefh 0.117f
C3109 X2.X1.X2.X2.X2.X2.X3.vin2 a_37466_29834# 3.85e-19
C3110 X2.X1.X1.X2.X2.X2.vout X2.X1.X1.X2.X2.X2.X3.vin1 0.335f
C3111 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X1.vin1 0.206f
C3112 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.vout 0.075f
C3113 X2.X1.X1.X2.X1.X2.vout X2.X1.X1.X2.X1.X2.X3.vin2 0.075f
C3114 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin2 0.12f
C3115 X1.X1.X1.X3.vin2 a_5082_10916# 0.452f
C3116 a_19422_16634# X1.X2.X1.X2.X1.X1.X3.vin2 0.267f
C3117 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X2.vrefh 0.076f
C3118 a_48616_10916# X2.X2.X1.X2.X2.X1.vout 1.64e-19
C3119 a_49002_10916# a_48702_9010# 5.25e-20
C3120 X2.X1.X2.X2.X2.X2.vrefh X2.X1.X2.X2.X2.X1.X3.vin2 0.161f
C3121 X2.X1.X2.X2.X1.X1.X3.vin1 a_40352_19358# 0.354f
C3122 a_22826_6962# X1.X2.X2.X1.X1.X1.X3.vin2 0.00815f
C3123 X1.X1.X1.X1.X2.X1.X2.vin1 a_2582_23258# 0.402f
C3124 X1.X1.X2.X2.X1.X1.X3.vin2 a_8872_20264# 0.1f
C3125 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin1 0.195f
C3126 X1.X2.X2.X3.vin2 X1.X2.X2.X3.vin1 0.559f
C3127 a_16836_15634# a_16836_13728# 0.00396f
C3128 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X1.X2.X2.X2.vin1 0.00117f
C3129 a_39966_32700# a_38152_31700# 1.15e-20
C3130 a_2582_21352# a_4782_20446# 4.2e-20
C3131 a_38152_16452# a_37466_14586# 3.31e-19
C3132 a_19036_31882# a_19422_31882# 0.419f
C3133 X2.X1.X3.vin1 X2.X1.X2.X3.vin1 3.45e-19
C3134 a_13696_892# X3.vin1 0.369f
C3135 X2.X1.X1.X2.X2.vrefh a_31476_11822# 0.118f
C3136 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X3.vin2 8.93e-19
C3137 X2.X2.X2.X2.X1.X1.vout X2.X2.X2.X2.X1.X1.X3.vin2 0.342f
C3138 a_17222_25164# X1.X2.X1.X1.X2.X1.X2.vin1 8.88e-20
C3139 a_48616_22312# a_46502_21352# 2.68e-20
C3140 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X2.X2.vin1 0.242f
C3141 a_31476_30882# a_31476_28976# 0.00396f
C3142 X1.X1.X2.X1.X1.X1.X1.vin2 X1.X2.X1.X2.X2.X2.X2.vin1 0.00232f
C3143 X1.X2.X1.X1.X3.vin2 a_19422_20446# 9.7e-20
C3144 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X3.vin1 0.587f
C3145 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.X1.X1.X1.vin2 3.94e-19
C3146 X1.X1.X3.vin2 a_8572_18358# 0.355f
C3147 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X2.X1.X1.X2.vrefh 0.00437f
C3148 X1.X2.X1.X2.X3.vin2 a_19422_5198# 9.7e-20
C3149 a_23126_16452# a_23212_14586# 3.38e-19
C3150 X1.X1.X2.X2.X2.X1.X3.vin1 a_8186_25982# 0.00837f
C3151 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X1.vin2 0.668f
C3152 X1.X2.X2.X2.X1.X1.X3.vin1 a_25712_19358# 0.354f
C3153 a_25712_23170# X1.X2.X2.X2.X1.X2.vrefh 1.64e-19
C3154 a_8186_6962# a_8486_5016# 4.19e-20
C3155 a_46502_27070# a_46502_25164# 0.00198f
C3156 a_19422_9010# X1.X2.X1.X2.X2.X1.X3.vin2 0.267f
C3157 a_46116_27070# X2.X2.X1.X1.X2.X1.X1.vin1 1.64e-19
C3158 a_33976_29936# a_34362_29936# 0.419f
C3159 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X3.vin1 2.33e-19
C3160 a_4696_29936# a_2582_28976# 2.68e-20
C3161 a_31476_15634# a_31862_15634# 0.419f
C3162 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X2.vin1 0.564f
C3163 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X1.vin2 0.668f
C3164 a_54992_25076# X2.X2.X2.X2.X1.X2.X1.vin2 1.78e-19
C3165 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 5.19e-19
C3166 a_17222_8010# a_17222_6104# 0.00198f
C3167 X1.X2.X1.X1.X1.X1.X3.vin2 X1.X2.X1.X1.X1.X2.X1.vin1 5.19e-19
C3168 a_38152_8828# a_37852_6962# 6.71e-19
C3169 a_16836_8010# X1.X2.X1.X2.X2.X2.X1.vin1 1.64e-19
C3170 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X3.vin1 0.0174f
C3171 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X1.X2.X1.X2.vrefh 0.1f
C3172 a_52106_22210# a_52406_20264# 4.19e-20
C3173 a_10686_6016# X1.X1.X2.X1.X1.X1.X1.vin2 8.88e-20
C3174 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X1.vout 0.0524f
C3175 X1.X2.X3.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 8.36e-19
C3176 X2.X1.X1.X2.X1.X2.X1.vin2 a_31476_11822# 1.78e-19
C3177 a_40352_26982# X2.X1.X2.X2.X2.vrefh 1.64e-19
C3178 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X1.vin2 0.076f
C3179 a_5082_29936# X1.X1.X1.X1.X1.X2.vout 0.254f
C3180 X1.X2.X3.vin1 a_20286_892# 0.17f
C3181 X2.X1.X1.X2.X1.X2.X3.vin1 a_33676_12822# 0.199f
C3182 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin2 7.84e-19
C3183 X1.X1.X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X1.X2.X1.vin2 3.94e-19
C3184 X2.X2.X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X2.X1.vin2 8.93e-19
C3185 a_4396_20446# a_2582_19446# 1.15e-20
C3186 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X3.vin2 0.418f
C3187 X2.X2.X2.X2.X2.X2.X2.vin1 a_54606_30794# 8.88e-20
C3188 X1.X2.X2.X1.X1.X2.X3.vin1 a_23212_6962# 0.00329f
C3189 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 5.19e-19
C3190 X1.X2.X2.X1.X2.X2.X1.vin2 X1.X2.X2.X1.X2.X2.X1.vin1 0.668f
C3191 a_19336_26164# a_17222_25164# 5.36e-21
C3192 X2.X1.X2.X2.X2.X1.X1.vin2 a_39966_26982# 0.273f
C3193 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.vrefh 2.33e-19
C3194 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 0.049f
C3195 a_54606_17452# a_52792_16452# 1.15e-20
C3196 X1.X1.X2.X1.X1.X1.X3.vin1 X1.X1.X2.X1.X1.X1.X1.vin1 0.206f
C3197 a_31476_8010# a_31862_8010# 0.419f
C3198 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X2.vin1 0.0689f
C3199 a_17222_21352# a_19036_20446# 1.06e-19
C3200 a_10686_30794# a_8572_29834# 2.68e-20
C3201 a_42976_892# a_43362_892# 0.419f
C3202 a_19722_29936# a_19036_28070# 3.31e-19
C3203 a_23212_18358# a_25326_17452# 4.72e-20
C3204 a_19336_29936# a_19422_28070# 3.38e-19
C3205 a_22826_25982# a_23212_25982# 0.414f
C3206 a_54606_6016# X2.X2.X2.X1.X1.X1.X1.vin2 8.88e-20
C3207 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.vout 0.118f
C3208 X2.X2.X2.X1.X1.X2.vrefh a_54606_6016# 0.3f
C3209 X1.X2.X1.X1.X2.X1.X3.vin2 a_17222_21352# 8.07e-19
C3210 a_49002_18540# X2.X2.X3.vin1 0.47f
C3211 a_8486_24076# a_8872_24076# 0.419f
C3212 X2.X1.X1.X2.vrefh a_31862_19446# 0.3f
C3213 a_38152_20264# a_39966_19358# 1.06e-19
C3214 a_31862_17540# a_31862_15634# 0.00198f
C3215 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 0.587f
C3216 a_37852_29834# a_39966_28888# 2.95e-20
C3217 a_25326_26982# a_25712_26982# 0.419f
C3218 a_31862_21352# X2.X1.X1.X1.X2.X2.X1.vin2 0.273f
C3219 a_25326_25076# a_23126_24076# 4.77e-21
C3220 a_37766_20264# a_37466_18358# 5.25e-20
C3221 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X1.vin2 0.668f
C3222 X1.X2.X2.X2.X2.X1.X3.vin1 a_23212_25982# 0.00251f
C3223 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X1.X3.vin2 0.0533f
C3224 X1.X2.X2.X1.X1.X2.X1.vin2 X1.X2.X2.X1.X1.X2.X1.vin1 0.668f
C3225 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X3.vin2 0.234f
C3226 X1.X2.X2.X2.X2.X2.X3.vin2 a_25326_30794# 7.84e-19
C3227 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X1.vin1 0.0689f
C3228 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X3.vin1 0.00118f
C3229 X2.X2.X1.X2.X1.X1.vout X2.X2.X1.X2.X1.X1.X3.vin2 0.342f
C3230 X2.X1.X1.X1.X2.X1.X3.vin2 a_31476_23258# 0.354f
C3231 X2.X2.X1.X1.X2.X2.X3.vin1 a_46502_19446# 0.00207f
C3232 X2.X1.X2.X2.X2.X1.X3.vin2 X2.X1.X2.X2.X2.X1.X1.vin1 2.23e-19
C3233 X2.X1.X2.X2.X2.X1.X2.vin1 a_40352_26982# 1.78e-19
C3234 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 1.22e-19
C3235 X2.X2.X2.X1.X1.X2.vout X2.X2.X2.X1.X1.X1.vout 0.507f
C3236 X1.X1.X1.X2.X2.X1.X3.vin2 a_2582_6104# 8.07e-19
C3237 a_39966_30794# X2.X1.X2.X2.X2.X2.vrefh 8.22e-20
C3238 a_8486_24076# a_8186_22210# 5.55e-20
C3239 a_23512_20264# a_25326_19358# 1.06e-19
C3240 X1.X2.X1.X2.vrefh a_17222_19446# 0.3f
C3241 a_48316_31882# X2.X2.X1.X1.X1.X1.vout 0.359f
C3242 a_34362_18540# X2.X1.X1.X2.X1.X1.X3.vin2 3.49e-19
C3243 X2.X1.X1.X3.vin2 a_34062_16634# 5.21e-19
C3244 X2.X2.X2.X1.X1.X1.X3.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 0.22f
C3245 a_52406_5016# a_54606_4110# 4.2e-20
C3246 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X2.X1.X1.X1.X2.X2.vin1 0.00232f
C3247 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.vout 0.398f
C3248 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X3.vin1 0.00118f
C3249 a_25326_25076# a_25712_25076# 0.419f
C3250 a_52492_25982# a_54606_25076# 4.72e-20
C3251 a_38152_31700# a_37852_29834# 6.71e-19
C3252 X2.X1.X2.X1.X2.X2.X3.vin1 a_40352_15546# 0.354f
C3253 a_16836_25164# X1.X2.X1.X1.X2.X1.X3.vin1 0.354f
C3254 a_17222_25164# X1.X2.X1.X1.X2.X1.X1.vin1 0.417f
C3255 X1.X2.X1.X2.X1.X2.X2.vin1 a_17222_11822# 0.402f
C3256 X1.X1.X1.X1.X1.X2.X3.vin2 a_2582_27070# 0.567f
C3257 X2.X2.X2.X2.X3.vin1 a_52492_22210# 0.363f
C3258 a_10686_32700# a_10686_30794# 0.00198f
C3259 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X1.vout 0.0524f
C3260 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 0.242f
C3261 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X1.vin2 0.696f
C3262 a_39966_17452# a_40352_17452# 0.419f
C3263 a_33676_16634# a_31862_15634# 1.15e-20
C3264 X1.X2.X1.X1.X1.X2.X1.vin2 a_16836_27070# 1.78e-19
C3265 X2.X1.X1.X3.vin2 a_34062_9010# 7.93e-20
C3266 X2.X2.X2.X2.X1.X1.X1.vin1 a_54992_19358# 0.195f
C3267 a_46116_25164# a_46116_23258# 0.00396f
C3268 X2.X2.X1.X1.X1.X2.X3.vin2 a_46502_27070# 0.567f
C3269 X2.X1.X2.X2.X3.vin2 a_37466_25982# 0.263f
C3270 X2.X2.X2.X1.X2.X1.X3.vin1 a_52492_10734# 0.00251f
C3271 a_46502_6104# X2.X2.X1.X2.X2.X2.X1.vin2 0.273f
C3272 a_11072_30794# a_11072_28888# 0.00396f
C3273 a_31476_17540# X2.X1.X1.X2.X1.X1.X3.vin1 0.354f
C3274 a_2196_17540# X1.X1.X1.X2.X1.X1.X2.vin1 1.78e-19
C3275 a_31862_17540# X2.X1.X1.X2.X1.X1.X1.vin1 0.417f
C3276 a_17222_28976# X1.X2.X1.X1.X1.X2.X3.vin2 7.84e-19
C3277 X1.X2.X1.X1.X1.X2.X3.vin1 a_19036_28070# 0.199f
C3278 a_25712_32700# X2.vrefh 0.118f
C3279 X2.X2.X1.X2.X2.X1.vout X2.X2.X1.X2.X2.X1.X3.vin2 0.326f
C3280 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X3.vin2 0.234f
C3281 X1.X1.X1.X2.X2.X1.vout X1.X1.X1.X2.X2.X1.X3.vin2 0.326f
C3282 a_54606_11734# X2.X2.X2.X1.X2.vrefh 8.22e-20
C3283 a_34362_29936# a_34062_28070# 5.55e-20
C3284 a_37766_5016# a_39966_4110# 4.2e-20
C3285 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X1.vin1 0.0689f
C3286 X2.X1.X2.X1.X1.X1.X3.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 0.22f
C3287 X1.X2.X2.X2.X1.X1.X3.vin2 a_25326_19358# 7.84e-19
C3288 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.X1.vin2 0.23f
C3289 X2.X2.X1.X1.X2.X2.X2.vin1 a_46116_19446# 0.197f
C3290 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X2.X1.X1.X2.X2.vrefh 0.00437f
C3291 X2.X2.X3.vin1 X2.X2.X1.X2.X1.X2.vout 3.08e-19
C3292 a_54606_17452# X2.X2.X2.X1.X2.X2.X1.vin2 8.88e-20
C3293 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X3.vin1 0.449f
C3294 X1.X1.X2.vrefh a_5646_892# 7.23e-19
C3295 X2.X2.X2.X2.X1.X1.X3.vin1 a_52492_18358# 0.00255f
C3296 X1.X1.X2.vrefh a_2196_4198# 0.119f
C3297 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X1.vin2 0.076f
C3298 X2.X1.X2.X1.X1.X2.X3.vin1 a_40352_7922# 0.354f
C3299 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin2 7.84e-19
C3300 X1.X2.X1.X2.X3.vin2 a_19722_7064# 0.422f
C3301 a_5082_26164# X1.X1.X1.X1.X2.X1.X3.vin1 0.00837f
C3302 X2.X1.X2.X2.X1.X1.X1.vin2 a_40352_19358# 0.12f
C3303 X2.X1.X2.X2.X1.X2.vout a_37466_22210# 0.254f
C3304 a_39966_19358# X2.X1.X2.X2.X1.X1.X1.vin1 0.417f
C3305 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X3.vin1 2.33e-19
C3306 a_33676_9010# a_31862_8010# 1.15e-20
C3307 X2.X1.X3.vin2 X2.X3.vin1 0.238f
C3308 X2.X2.X3.vin2 X2.X2.X1.X2.X2.X2.vout 1.5e-19
C3309 X2.X2.X2.X1.X1.X2.X1.vin1 a_54992_6016# 1.64e-19
C3310 X1.X2.X2.X1.X1.X1.X3.vin1 a_25326_4110# 0.52f
C3311 X2.X2.X2.X1.X2.X2.X1.vin1 a_54992_15546# 0.195f
C3312 X1.X1.X2.X2.X1.X2.X1.vin1 a_11072_21264# 1.64e-19
C3313 X2.X1.X2.X1.X1.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin2 0.0128f
C3314 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X1.vin2 0.076f
C3315 X1.X1.X1.X2.X1.X2.X3.vin1 a_2582_11822# 0.00207f
C3316 a_48616_7064# a_49002_7064# 0.419f
C3317 a_8186_25982# X1.X1.X2.X3.vin2 0.452f
C3318 X1.X1.X1.X1.X1.X1.X1.vin1 vrefh 0.103f
C3319 a_31862_17540# a_34062_16634# 4.2e-20
C3320 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X2.vin1 0.00117f
C3321 a_10686_9828# a_11072_9828# 0.419f
C3322 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X1.vout 0.033f
C3323 a_52106_29834# X2.X2.X2.X2.X2.X1.vout 0.383f
C3324 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin1 0.195f
C3325 a_10686_25076# X1.X1.X2.X2.X1.X2.X1.vin2 8.88e-20
C3326 a_2196_9916# X1.X1.X1.X2.X2.X1.X3.vin1 0.354f
C3327 X2.X2.X2.X1.X2.vrefh a_54606_9828# 0.3f
C3328 a_2582_9916# X1.X1.X1.X2.X2.X1.X1.vin1 0.417f
C3329 a_25326_19358# X1.X2.X2.X2.X1.X1.X1.vin1 0.417f
C3330 X1.X2.X2.X2.X1.X1.X1.vin2 a_25712_19358# 0.12f
C3331 X1.X1.X1.X2.X2.X2.vrefh X1.X1.X1.X2.X2.X2.X3.vin1 2.33e-19
C3332 a_40352_28888# X2.X1.X2.X2.X2.X1.X1.vin2 1.78e-19
C3333 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X1.vin2 0.668f
C3334 a_52406_8828# a_52492_6962# 3.38e-19
C3335 a_8186_14586# a_8486_12640# 4.19e-20
C3336 a_23212_10734# a_23126_8828# 3.3e-19
C3337 a_33676_24258# X2.X1.X1.X1.X2.X1.X3.vin2 0.1f
C3338 X2.X2.X2.X1.X1.X2.X1.vin1 a_54992_7922# 0.195f
C3339 a_49002_29936# X2.X2.X1.X1.X1.X2.X3.vin2 3.85e-19
C3340 X2.X2.X1.X1.X3.vin1 a_48702_28070# 9.54e-19
C3341 a_54606_13640# X2.X2.X2.X1.X2.X1.X3.vin1 0.00207f
C3342 X1.X1.X2.X2.X1.X1.vout X1.X1.X2.X2.X1.X1.X3.vin2 0.342f
C3343 a_33976_22312# a_34362_22312# 0.419f
C3344 a_4696_22312# a_2582_21352# 2.68e-20
C3345 a_23126_12640# a_23512_12640# 0.419f
C3346 a_8486_20264# a_8186_18358# 5.25e-20
C3347 a_46116_15634# a_46116_13728# 0.00396f
C3348 X1.X1.X2.X2.X1.X1.X1.vin2 a_11072_19358# 0.12f
C3349 X1.X2.X2.X2.X1.X2.X3.vin1 a_25326_23170# 0.52f
C3350 a_10686_19358# X1.X1.X2.X2.X1.X1.X1.vin1 0.417f
C3351 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X1.vin1 5.19e-19
C3352 a_37766_31700# a_38152_31700# 0.419f
C3353 a_33676_16634# a_34062_16634# 0.419f
C3354 a_2582_30882# X1.X1.X1.X1.X1.X2.X1.vin1 8.22e-20
C3355 a_46116_25164# X2.X2.X1.X1.X2.X1.X2.vin1 1.78e-19
C3356 X1.X2.X2.X2.X1.X2.vout a_23512_24076# 0.36f
C3357 X1.X2.X1.X1.X2.X1.X2.vin1 a_16836_23258# 0.197f
C3358 X1.X2.X2.X1.X3.vin2 a_23212_14586# 0.363f
C3359 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X3.vin1 0.199f
C3360 X1.X2.X2.X2.X2.X2.vout a_22826_29834# 0.263f
C3361 a_8572_18358# a_8872_16452# 6.48e-19
C3362 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin1 0.195f
C3363 X2.X1.X3.vin2 X2.X1.X2.X1.X2.X2.X3.vin2 0.0011f
C3364 X1.X2.X2.X1.X2.X1.X3.vin2 a_25326_11734# 7.84e-19
C3365 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X1.vin1 0.0689f
C3366 X1.X1.X2.X2.X2.X1.X3.vin2 a_8872_27888# 0.1f
C3367 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X2.vrefh 0.076f
C3368 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X2.vrefh 0.00118f
C3369 a_16836_27070# a_16836_25164# 0.00396f
C3370 X1.X2.X1.X1.X2.vrefh a_17222_25164# 8.22e-20
C3371 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X2.X2.vin1 0.00117f
C3372 a_2582_28976# a_4782_28070# 4.2e-20
C3373 X1.X2.X2.X2.X2.X1.vout X1.X2.X2.X2.X2.X1.X3.vin1 0.118f
C3374 X2.X1.X1.X2.X1.X1.X3.vin2 a_31862_13728# 8.07e-19
C3375 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.vout 0.075f
C3376 X2.X1.X3.vin1 X2.X1.X1.X2.X3.vin1 7.18e-19
C3377 X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X1.X3.vin2 0.0533f
C3378 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 0.242f
C3379 a_10686_21264# a_10686_19358# 0.00198f
C3380 a_34062_28070# X2.X1.X1.X1.X1.X2.X3.vin2 0.277f
C3381 a_8486_31700# a_8186_29834# 5.55e-20
C3382 vout X3.vin2 0.0726f
C3383 X2.X1.X1.X3.vin1 a_33976_18540# 0.17f
C3384 X2.X1.X1.X3.vin1 a_34062_20446# 5.31e-19
C3385 d7 a_28482_892# 0.00777f
C3386 a_46502_8010# a_46502_6104# 0.00198f
C3387 a_33676_9010# a_34062_9010# 0.419f
C3388 a_46116_8010# X2.X2.X1.X2.X2.X2.X1.vin1 1.64e-19
C3389 X2.X2.X1.X1.X1.X1.X3.vin2 a_46502_28976# 8.07e-19
C3390 a_19036_12822# a_19336_10916# 6.48e-19
C3391 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X3.vin1 0.00117f
C3392 X2.X1.X2.X1.X2.X2.X3.vin2 a_37766_16452# 0.277f
C3393 X1.X1.X1.X1.X1.X2.vout X1.X1.X1.X1.X1.X2.X3.vin2 0.075f
C3394 X1.X1.X3.vin2 a_8186_14586# 3.67e-19
C3395 a_2196_23258# X1.X1.X1.X1.X2.X2.X1.vin1 1.64e-19
C3396 X1.X3.vin1 X1.X3.vin2 0.514f
C3397 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 0.581f
C3398 a_2582_23258# a_2582_21352# 0.00198f
C3399 a_23212_14586# a_23126_12640# 3.14e-19
C3400 X2.X1.X3.vin2 a_37766_12640# 2.33e-19
C3401 X2.X1.X2.X2.X1.X2.X1.vin2 a_39966_23170# 0.273f
C3402 a_10686_30794# a_11072_30794# 0.419f
C3403 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X1.X1.vin2 0.216f
C3404 a_23126_27888# a_25326_26982# 4.2e-20
C3405 X1.X1.X2.X2.X1.X1.X1.vin1 a_11072_17452# 1.64e-19
C3406 a_33976_10916# X2.X1.X1.X2.X2.X1.X3.vin1 0.00251f
C3407 X2.X2.X1.X1.X1.X2.vrefh a_46502_30882# 0.3f
C3408 X2.X2.X2.X1.X2.X1.X1.vin1 a_54992_9828# 1.64e-19
C3409 X1.X1.X1.X3.vin1 X1.X1.X1.X3.vin2 0.552f
C3410 X2.X2.X2.X2.X2.X2.X3.vin1 a_52106_29834# 0.00874f
C3411 a_17222_9916# a_19036_9010# 1.06e-19
C3412 a_52106_6962# a_52406_5016# 4.19e-20
C3413 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X2.vin1 0.0689f
C3414 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X3.vin2 0.161f
C3415 X2.X2.X2.X2.X2.X2.X2.vin1 vrefl 0.597f
C3416 X2.X2.X2.X2.X2.X2.X3.vin2 a_54992_32700# 0.354f
C3417 X1.X1.X1.X2.X1.X2.vrefh a_2196_13728# 1.64e-19
C3418 a_48616_14688# a_46502_13728# 2.68e-20
C3419 X2.X1.X2.vrefh X2.X3.vin1 0.0451f
C3420 a_10686_13640# a_11072_13640# 0.419f
C3421 X2.X1.X1.X1.X3.vin1 X2.X1.X2.X2.X3.vin2 0.0604f
C3422 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.X3.vin1 1.22e-19
C3423 a_31476_28976# a_31476_27070# 0.00396f
C3424 a_4782_28070# a_5082_26164# 4.41e-20
C3425 X1.X1.X1.X1.X1.X2.X3.vin2 a_4696_26164# 0.00535f
C3426 X2.X2.X1.X1.X1.X1.X1.vin1 X2.X2.X1.X1.X1.X1.X3.vin1 0.206f
C3427 a_39966_28888# X2.X1.X2.X2.X2.X1.X3.vin1 0.00207f
C3428 X1.X2.X1.X2.X2.X2.X1.vin2 a_16836_4198# 1.78e-19
C3429 a_2196_13728# X1.X1.X1.X2.X1.X2.X3.vin1 0.354f
C3430 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X2.vin1 0.564f
C3431 a_2582_13728# X1.X1.X1.X2.X1.X2.X1.vin1 0.417f
C3432 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X2.vrefh 0.076f
C3433 X1.X2.X2.X1.X1.X1.X3.vin2 a_23512_5016# 0.1f
C3434 X1.X1.X2.X2.X2.X2.vrefh a_11072_28888# 0.118f
C3435 a_34362_7064# a_33676_5198# 3.31e-19
C3436 X1.X2.X2.X2.X1.X2.X3.vin2 a_22826_22210# 3.85e-19
C3437 a_17222_6104# a_19422_5198# 4.2e-20
C3438 a_33976_7064# a_34062_5198# 3.38e-19
C3439 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X2.vin1 0.00117f
C3440 a_19336_10916# X1.X2.X1.X2.X3.vin2 0.0927f
C3441 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X1.X3.vin2 0.0943f
C3442 X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin2 0.0128f
C3443 a_2582_15634# a_4696_14688# 2.95e-20
C3444 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X2.vout 0.0866f
C3445 a_46502_27070# a_48616_26164# 4.72e-20
C3446 X2.X2.X3.vin2 a_49002_10916# 3.68e-19
C3447 a_52792_27888# a_52492_25982# 6.2e-19
C3448 X1.X1.X1.X2.X1.X2.vout X1.X1.X1.X2.X1.X2.X3.vin1 0.326f
C3449 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X1.X2.X1.X1.X1.X3.vin2 3.94e-19
C3450 X1.X1.X2.X1.X1.X2.X1.vin1 a_10686_6016# 8.22e-20
C3451 a_54606_19358# a_52492_18358# 5.36e-21
C3452 X1.X1.X2.X2.X2.X1.X3.vin2 a_10686_26982# 7.84e-19
C3453 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X1.vin1 0.0689f
C3454 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X2.X1.X1.vin1 0.206f
C3455 X1.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin2 0.0128f
C3456 a_40352_19358# X2.X1.X2.X2.vrefh 1.64e-19
C3457 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X3.vin1 0.0131f
C3458 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X2.X1.X1.vin1 0.206f
C3459 X2.X2.X2.X1.X1.X2.X2.vin1 a_54992_9828# 0.197f
C3460 X1.X2.X1.X2.X2.X1.X3.vin2 a_19722_7064# 0.00815f
C3461 X1.X2.X2.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin1 0.00437f
C3462 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X3.vin2 0.0565f
C3463 a_39966_25076# a_38152_24076# 1.15e-20
C3464 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X1.vin2 0.216f
C3465 a_48316_20446# X2.X2.X1.X1.X2.X2.X3.vin2 0.101f
C3466 X1.X2.X3.vin2 a_22826_10734# 6.66e-19
C3467 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X3.vin1 2.33e-19
C3468 X2.X2.X1.X1.X1.X1.X1.vin2 X2.X2.X1.X1.X1.X1.X3.vin2 8.93e-19
C3469 X1.X1.X2.X2.X3.vin2 X1.X1.X1.X3.vin1 7.46e-20
C3470 a_31862_28976# X2.X1.X1.X1.X1.X2.X1.vin2 0.273f
C3471 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin1 0.52f
C3472 X1.X1.X2.X1.X2.X1.vout a_8572_14586# 0.169f
C3473 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 0.581f
C3474 X2.X2.X2.X2.X1.X2.X3.vin1 a_54992_23170# 0.354f
C3475 X2.X2.X3.vin2 a_52492_18358# 0.355f
C3476 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X1.X3.vin2 0.234f
C3477 a_2582_8010# a_4696_7064# 2.95e-20
C3478 a_48316_24258# a_46502_23258# 1.15e-20
C3479 X2.X1.X1.X1.X2.X1.vout X2.X1.X1.X1.X2.X2.vout 0.514f
C3480 X1.X2.X2.X1.X2.X2.X1.vin1 a_25712_13640# 1.64e-19
C3481 a_17222_25164# a_17222_23258# 0.00198f
C3482 X2.X1.X3.vin1 a_35312_892# 0.371f
C3483 X1.X1.X1.X1.X1.X1.vout X1.X1.X1.X1.X3.vin1 0.13f
C3484 X2.X2.X3.vin1 a_49002_7064# 9.8e-19
C3485 X1.X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin2 0.0128f
C3486 X1.X1.X1.X1.X2.vrefh a_2196_25164# 1.64e-19
C3487 X1.X2.X2.X2.X2.X2.X3.vin2 a_22826_29834# 3.85e-19
C3488 a_54606_28888# X2.X2.X2.X2.X2.X1.X1.vin2 8.88e-20
C3489 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X2.vrefh 0.267f
C3490 X2.X1.X2.X2.X2.X2.X1.vin1 a_40352_28888# 1.64e-19
C3491 a_34062_20446# a_33976_18540# 3.3e-19
C3492 a_33676_20446# a_34362_18540# 3.08e-19
C3493 X2.X2.X2.vrefh a_43362_892# 2.22e-19
C3494 a_33676_20446# X2.X1.X1.X1.X2.X2.X3.vin2 0.101f
C3495 X1.X2.X2.X1.X2.X2.X2.vin1 a_25326_15546# 8.88e-20
C3496 a_25326_9828# X1.X2.X2.X1.X1.X2.X3.vin1 0.00207f
C3497 X2.X2.X3.vin1 X2.X2.X2.vrefh 0.178f
C3498 a_54606_25076# X2.X2.X2.X2.X1.X2.X2.vin1 0.402f
C3499 X1.X2.X2.X2.X2.X2.vrefh X2.X1.X1.X1.X1.X2.X1.vin2 0.0128f
C3500 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X1.vin2 8.93e-19
C3501 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.vrefh 0.161f
C3502 X1.X2.X3.vin1 a_22826_6962# 6.45e-19
C3503 X1.X1.X1.X1.X1.X2.vrefh a_2582_30882# 0.3f
C3504 a_49002_29936# X2.X2.X1.X1.X1.X2.vout 0.254f
C3505 a_2582_19446# a_2582_17540# 0.00198f
C3506 a_8872_31700# a_10686_30794# 1.06e-19
C3507 a_2196_19446# X1.X1.X1.X2.X1.X1.X1.vin1 1.64e-19
C3508 a_4396_16634# X1.X1.X1.X2.X1.X1.X3.vin2 0.1f
C3509 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X2.vout 0.2f
C3510 a_46116_11822# X2.X2.X1.X2.X2.X1.X1.vin1 1.64e-19
C3511 a_52406_31700# X2.X2.X2.X2.X2.X2.X3.vin1 0.42f
C3512 a_46502_11822# a_46502_9916# 0.00198f
C3513 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.vout 0.326f
C3514 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.vout 0.118f
C3515 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X3.vin1 2.33e-19
C3516 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X3.vin2 8.93e-19
C3517 a_4696_18540# X1.X1.X1.X3.vin2 0.0927f
C3518 X2.X2.X2.X1.X3.vin2 a_52106_10734# 0.241f
C3519 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin2 0.12f
C3520 a_4396_24258# a_5082_22312# 2.86e-19
C3521 a_4782_24258# a_4696_22312# 3.14e-19
C3522 a_19336_26164# a_19036_24258# 6.2e-19
C3523 a_34362_14688# X2.X1.X1.X2.X1.X2.X3.vin1 0.00874f
C3524 a_16836_32788# X1.X2.X1.X1.X1.X1.X2.vin1 1.78e-19
C3525 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X3.vin1 2.33e-19
C3526 a_8872_8828# a_8572_6962# 6.71e-19
C3527 X2.X1.X2.X2.X2.X2.X1.vin1 a_40352_30794# 0.195f
C3528 X1.X1.X1.X3.vin1 a_4782_20446# 5.31e-19
C3529 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X2.vrefh 0.267f
C3530 X1.X1.X1.X2.X1.X1.X1.vin2 a_2196_15634# 1.78e-19
C3531 a_19036_20446# X1.X2.X1.X1.X2.X2.X3.vin2 0.101f
C3532 a_8186_25982# a_8872_24076# 3.08e-19
C3533 a_2196_32788# X1.X1.X1.X1.X1.X1.X2.vin1 1.78e-19
C3534 X2.X1.X2.X1.X1.X1.X1.vin2 X2.X2.X1.X2.X2.X2.X2.vin1 0.00232f
C3535 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.vrefh 0.161f
C3536 X1.X2.X2.X1.X3.vin2 a_23212_10734# 0.0927f
C3537 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X3.vin1 2.33e-19
C3538 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 0.587f
C3539 a_37466_29834# a_38152_27888# 2.86e-19
C3540 X2.X2.X1.X2.X1.X2.X3.vin2 a_49002_10916# 0.00846f
C3541 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.vrefh 2.33e-19
C3542 X1.X1.X1.X1.X1.X1.X1.vin2 a_4782_31882# 0.00743f
C3543 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 5.19e-19
C3544 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X3.vin1 0.00836f
C3545 X2.X1.X3.vin1 X2.X1.X1.X2.X3.vin2 0.0816f
C3546 X1.X1.X1.X2.X2.vrefh a_2196_11822# 0.118f
C3547 X1.X2.X1.X1.X1.X1.vout X1.X2.X1.X1.X1.X2.vout 0.507f
C3548 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X3.vin1 0.00789f
C3549 X2.X2.X1.X2.X2.vrefh a_46502_11822# 0.3f
C3550 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X2.vout 0.197f
C3551 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 0.0903f
C3552 a_25326_13640# a_23126_12640# 4.77e-21
C3553 a_39966_9828# X2.X1.X2.X1.X1.X2.X2.vin1 0.402f
C3554 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X1.vin2 0.668f
C3555 X2.X2.X2.X1.X2.X1.X2.vin1 a_54992_13640# 0.197f
C3556 X1.X1.X3.vin1 X1.X1.X2.X1.X3.vin1 0.00304f
C3557 a_4782_24258# a_2582_23258# 4.77e-21
C3558 X2.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.vout 0.399f
C3559 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 2.23e-19
C3560 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin1 0.195f
C3561 a_52106_6962# a_52492_6962# 0.419f
C3562 a_23126_12640# a_23212_10734# 3.21e-19
C3563 X2.X1.X2.X3.vin1 a_37852_18358# 0.17f
C3564 a_19336_26164# a_19722_26164# 0.414f
C3565 a_17222_15634# a_17222_13728# 0.00198f
C3566 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin1 0.52f
C3567 a_16836_15634# X1.X2.X1.X2.X1.X2.X1.vin1 1.64e-19
C3568 a_10686_30794# X1.X1.X2.X2.X2.X2.vrefh 8.22e-20
C3569 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X2.vrefh 0.076f
C3570 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 2.23e-19
C3571 X2.X1.X2.X2.X2.X2.X3.vin2 a_38152_31700# 0.101f
C3572 X1.X1.X1.X1.X2.X2.X3.vin1 a_4782_20446# 0.42f
C3573 a_19422_31882# X1.X2.X1.X1.X1.X1.vout 0.422f
C3574 a_31476_11822# a_31862_11822# 0.419f
C3575 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X2.vin1 0.00117f
C3576 a_17222_25164# a_19422_24258# 4.2e-20
C3577 a_31862_30882# a_31862_28976# 0.00198f
C3578 a_31476_30882# X2.X1.X1.X1.X1.X2.X1.vin1 1.64e-19
C3579 a_48616_22312# X2.X2.X1.X1.X2.X2.X3.vin1 0.00329f
C3580 a_52406_16452# a_52792_16452# 0.419f
C3581 a_39966_6016# X2.X1.X2.X1.X1.X1.X3.vin1 0.00207f
C3582 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X2.X1.X2.X1.X2.vrefh 0.0128f
C3583 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin2 0.1f
C3584 X2.X1.X3.vin2 a_37766_16452# 3.98e-19
C3585 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 0.242f
C3586 X1.X1.X2.X1.X1.X1.vout X1.X1.X2.X1.X1.X1.X3.vin1 0.118f
C3587 a_10686_9828# a_10686_7922# 0.00198f
C3588 X2.X2.X1.X2.X2.X1.X3.vin2 a_48616_7064# 0.00546f
C3589 X2.X2.X2.X2.X2.X1.vout a_52792_27888# 0.359f
C3590 a_4696_29936# X1.X1.X1.X1.X1.X2.X3.vin1 0.00329f
C3591 a_34362_29936# X2.X1.X1.X1.X3.vin1 0.434f
C3592 a_5082_14688# a_4396_12822# 3.31e-19
C3593 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X2.X1.X1.vin1 0.668f
C3594 a_4696_14688# a_4782_12822# 3.38e-19
C3595 a_19036_16634# a_19336_14688# 6.1e-19
C3596 X3.vin2 a_35312_892# 5.64e-19
C3597 a_37466_22210# a_37852_22210# 0.419f
C3598 X2.X2.X2.X1.X2.X2.vrefh a_54606_13640# 0.3f
C3599 X2.X1.X3.vin2 a_37766_8828# 2.33e-19
C3600 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 0.049f
C3601 X2.X1.X1.X1.X1.X1.X3.vin2 a_34362_29936# 0.00815f
C3602 a_8872_16452# a_8186_14586# 3.31e-19
C3603 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X2.vrefh 0.267f
C3604 X1.X1.X2.X1.X1.X1.X2.vin1 a_10686_4110# 8.88e-20
C3605 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X1.vin2 8.93e-19
C3606 X1.X2.vrefh X1.X1.X2.X2.X2.X2.X3.vin1 0.00118f
C3607 X2.X2.X2.X2.X1.X1.vout X2.X2.X2.X2.X1.X1.X3.vin1 0.118f
C3608 a_52406_8828# a_52792_8828# 0.419f
C3609 a_4782_20446# a_4696_18540# 3.3e-19
C3610 a_4396_20446# a_5082_18540# 3.08e-19
C3611 a_8486_8828# a_8872_8828# 0.419f
C3612 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin2 7.84e-19
C3613 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X2.X1.X2.X2.X2.vrefh 0.0128f
C3614 a_52106_25982# X2.X2.X2.X3.vin2 0.452f
C3615 X1.X1.X2.X1.X2.X1.X1.vin2 a_10686_11734# 0.273f
C3616 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 0.587f
C3617 X1.X1.X1.X1.X2.X2.X3.vin2 a_2582_19446# 0.567f
C3618 X2.X2.X2.X2.X2.X2.X2.vin1 a_54992_30794# 1.78e-19
C3619 a_25326_15546# a_25712_15546# 0.419f
C3620 X2.X2.X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X2.X1.vin1 2.23e-19
C3621 a_39966_26982# X2.X1.X2.X2.X2.X1.X1.vin1 0.417f
C3622 X2.X1.X2.X2.X2.X1.X1.vin2 a_40352_26982# 0.12f
C3623 a_19336_26164# X1.X2.X1.X1.X2.X1.X3.vin1 0.00251f
C3624 a_46502_9916# X2.X2.X1.X2.X2.X1.X2.vin1 8.88e-20
C3625 X2.X2.X2.X1.X2.X2.X3.vin2 a_52792_16452# 0.101f
C3626 a_52492_25982# a_52406_24076# 3.3e-19
C3627 X2.X1.X1.X2.vrefh a_31476_17540# 1.64e-19
C3628 X2.X2.X2.X1.X2.X2.vout X2.X2.X2.X1.X3.vin2 0.0866f
C3629 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin2 7.84e-19
C3630 X1.X2.X1.X1.X2.X2.X3.vin1 a_19036_20446# 0.199f
C3631 X1.X2.X1.X3.vin2 a_19722_10916# 0.452f
C3632 a_43362_892# X2.X3.vin2 0.255f
C3633 a_23212_18358# X1.X2.X2.X1.X2.X2.X3.vin2 0.00517f
C3634 X1.X1.X1.X1.X3.vin1 a_5082_26164# 0.385f
C3635 X2.X2.X2.X1.X1.X1.X2.vin1 a_54606_4110# 8.88e-20
C3636 a_19722_29936# X1.X2.X1.X1.X1.X2.X3.vin2 3.85e-19
C3637 X1.X2.X1.X1.X3.vin1 a_19422_28070# 9.54e-19
C3638 X2.X2.X2.X1.X1.X1.X3.vin2 X2.X2.X2.X1.X1.X1.X1.vin2 8.93e-19
C3639 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X1.vout 0.13f
C3640 X2.X2.X3.vin1 X2.X3.vin2 0.12f
C3641 X2.X2.X3.vin1 a_52406_12640# 8.66e-20
C3642 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X3.vin2 0.165f
C3643 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X3.vin1 1.22e-19
C3644 X2.X1.X2.X2.X2.X2.vrefh a_40352_28888# 0.118f
C3645 a_39966_32700# a_39966_30794# 0.00198f
C3646 X2.X1.X1.X2.X1.X1.X3.vin1 a_31862_15634# 0.00207f
C3647 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 0.242f
C3648 a_37852_29834# X2.X1.X2.X2.X2.X1.X3.vin2 0.00546f
C3649 X1.X2.X2.X2.X1.X2.X3.vin2 a_23126_24076# 0.277f
C3650 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X1.X2.X2.X1.vin2 0.216f
C3651 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X2.vin1 0.242f
C3652 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X3.vin1 0.00117f
C3653 X1.X1.X2.X1.X1.X2.X3.vin1 a_10686_7922# 0.52f
C3654 a_25712_9828# a_25712_7922# 0.00396f
C3655 X2.X1.X2.X1.X2.X2.X3.vin1 a_37852_14586# 0.00329f
C3656 a_39966_13640# X2.X1.X2.X1.X2.X1.X2.vin1 0.402f
C3657 a_25326_7922# a_25712_7922# 0.419f
C3658 X1.X1.X1.X2.X2.X1.X2.vin1 a_2196_8010# 0.197f
C3659 X1.X2.X2.X3.vin1 X1.X2.X3.vin2 1.16f
C3660 X1.X2.X2.X2.X1.X1.X1.vin2 X2.X1.X1.X2.vrefh 0.0128f
C3661 X2.X1.X1.X2.X1.X2.X2.vin1 a_31476_11822# 0.197f
C3662 a_39966_7922# a_39966_6016# 0.00198f
C3663 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.vout 0.335f
C3664 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.vout 0.075f
C3665 X1.X1.X1.X2.X2.X1.X3.vin2 X1.X1.X1.X2.X2.X2.X3.vin1 1.22e-19
C3666 X2.X2.X1.X1.X1.X1.X3.vin2 a_48616_29936# 0.00546f
C3667 a_8872_27888# a_8186_25982# 2.97e-19
C3668 a_54992_13640# a_54992_11734# 0.00396f
C3669 a_40352_30794# X2.X1.X2.X2.X2.X2.vrefh 1.64e-19
C3670 X2.X1.X2.X1.X2.X1.vout X2.X1.X2.X1.X2.X1.X3.vin2 0.326f
C3671 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin2 0.1f
C3672 X2.X1.X3.vin2 X2.X1.X2.vrefh 0.15f
C3673 X2.X2.X2.X1.X1.X1.X3.vin1 X2.X2.X2.X1.X1.X1.X1.vin1 0.206f
C3674 X2.X2.X2.X2.X3.vin2 a_52406_27888# 0.00101f
C3675 a_8486_5016# X1.X1.X2.X1.X1.X1.X3.vin1 0.428f
C3676 X1.X1.X1.X2.X2.X2.X2.vin1 X1.X1.X2.vrefh 0.564f
C3677 X1.X2.X2.X2.X1.X2.X3.vin2 a_25712_25076# 0.354f
C3678 a_52492_25982# X2.X2.X2.X2.X1.X2.X3.vin2 0.00535f
C3679 a_39966_7922# a_37852_6962# 2.68e-20
C3680 a_40352_21264# a_40352_19358# 0.00396f
C3681 X1.X2.X2.X1.X3.vin1 a_23212_10734# 0.169f
C3682 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X3.vin1 0.206f
C3683 X1.X2.X1.X2.X1.X2.X3.vin2 a_16836_11822# 0.354f
C3684 X2.X2.X2.X2.X1.X1.X1.vin1 a_54606_17452# 8.22e-20
C3685 a_19422_12822# a_17222_11822# 4.77e-21
C3686 X2.X2.X2.X1.X2.X2.X1.vin1 a_54992_13640# 1.64e-19
C3687 X2.X2.X2.X2.X1.X1.X1.vin2 X2.X2.X2.X1.X2.X2.X3.vin2 3.94e-19
C3688 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X1.vin1 0.0689f
C3689 X1.X1.X2.X2.X2.X2.X3.vin2 a_10686_30794# 7.84e-19
C3690 X2.X1.X2.X1.X2.X2.X3.vin2 a_40352_17452# 0.354f
C3691 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X2.X1.X2.vrefh 0.0128f
C3692 a_54606_19358# X2.X2.X2.X2.vrefh 8.22e-20
C3693 a_16836_23258# a_17222_23258# 0.419f
C3694 a_46502_25164# a_46502_23258# 0.00198f
C3695 X2.X1.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin2 0.0128f
C3696 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X1.vin2 0.22f
C3697 a_2582_17540# a_4396_16634# 1.06e-19
C3698 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.vrefh 0.00118f
C3699 X1.X2.X3.vin1 a_23126_16452# 8.66e-20
C3700 X1.X2.X2.X2.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin1 0.00437f
C3701 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X2.vin1 0.0689f
C3702 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X1.X3.vin2 0.0533f
C3703 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X3.vin1 0.206f
C3704 a_33676_9010# a_33976_7064# 6.1e-19
C3705 X1.X2.X1.X1.X1.X2.X3.vin1 X1.X2.X1.X1.X1.X2.X3.vin2 0.587f
C3706 X2.X1.X2.X1.X1.X1.X3.vin1 X2.X1.X2.X1.X1.X1.X1.vin1 0.206f
C3707 a_54992_11734# X2.X2.X2.X1.X2.vrefh 1.64e-19
C3708 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X2.X3.vin2 0.0565f
C3709 X2.X2.X3.vin2 a_52106_14586# 3.67e-19
C3710 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X1.vin2 8.93e-19
C3711 a_54992_32700# X2.X2.X2.X2.X2.X2.X1.vin2 1.78e-19
C3712 X1.X2.X2.X2.X2.X1.X1.vin1 a_25712_25076# 1.64e-19
C3713 X2.X2.X2.X1.X2.X2.X2.vin1 a_54606_15546# 8.88e-20
C3714 a_48316_20446# a_46502_19446# 1.15e-20
C3715 a_54606_9828# a_52406_8828# 4.77e-21
C3716 X1.X2.X2.X1.X1.X2.vout a_23212_6962# 0.0929f
C3717 a_16836_11822# a_16836_9916# 0.00396f
C3718 X1.X2.X3.vin1 a_23126_8828# 8.66e-20
C3719 a_19336_14688# X1.X2.X1.X2.X1.X2.vout 0.0929f
C3720 X1.X2.X1.X2.X2.vrefh a_17222_9916# 8.22e-20
C3721 a_37466_25982# X2.X1.X2.X2.X3.vin1 0.372f
C3722 X2.X1.X1.X1.X3.vin2 X2.X1.X2.X3.vin2 7.46e-20
C3723 X1.X1.X1.X3.vin2 a_4782_16634# 5.21e-19
C3724 a_5082_18540# X1.X1.X1.X2.X1.X1.X3.vin2 3.49e-19
C3725 X2.X2.X1.X3.vin1 X2.X2.X1.X3.vin2 0.552f
C3726 a_52406_16452# a_52492_14586# 3.38e-19
C3727 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X1.X2.X2.X1.X2.X1.vin1 0.668f
C3728 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 0.581f
C3729 X2.X1.X2.X2.X1.X1.X1.vin1 a_40352_19358# 0.195f
C3730 X1.X2.X1.X1.X1.X2.vrefh a_16836_30882# 0.118f
C3731 a_8872_31700# a_8572_29834# 6.71e-19
C3732 X2.X2.X1.X3.vin2 a_48702_12822# 6.03e-19
C3733 X2.X1.X2.X3.vin2 a_37766_20264# 5.21e-19
C3734 X1.X2.X2.X1.X1.X1.X3.vin1 a_25712_4110# 0.354f
C3735 a_23212_6962# a_25326_6016# 2.95e-20
C3736 X1.X1.X2.X1.X3.vin1 a_8486_5016# 1.52e-19
C3737 a_54606_15546# X2.X2.X2.X1.X2.X2.vrefh 8.22e-20
C3738 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X3.vin2 8.93e-19
C3739 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X3.vin1 0.00789f
C3740 a_49002_7064# X2.X2.X1.X2.X2.X2.vout 0.263f
C3741 X2.X1.X1.X1.X2.X2.X2.vin1 a_31862_19446# 0.402f
C3742 a_34362_18540# X2.X1.X3.vin2 6.58e-20
C3743 a_23512_27888# a_23212_25982# 6.2e-19
C3744 X2.X2.X3.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 8.36e-19
C3745 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X1.vout 0.0524f
C3746 X2.X1.X1.X2.X1.X1.X3.vin1 a_34062_16634# 0.428f
C3747 X1.X2.X2.X2.X1.X1.X2.vin1 a_25712_21264# 0.197f
C3748 X1.X1.X2.X1.X1.X2.X3.vin2 a_11072_9828# 0.354f
C3749 a_8486_16452# a_10686_15546# 4.2e-20
C3750 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 0.216f
C3751 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X1.vin2 8.93e-19
C3752 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin1 0.52f
C3753 X1.X1.X1.X1.X1.X1.X2.vin1 a_2196_30882# 0.197f
C3754 X1.X1.X2.X2.X1.X2.X2.vin1 a_10686_23170# 8.88e-20
C3755 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X3.vin2 0.161f
C3756 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X3.vin1 0.206f
C3757 X1.X2.X2.X2.X1.X1.X1.vin1 a_25712_19358# 0.195f
C3758 X2.vrefh X1.X2.X2.X2.X2.X2.X1.vin2 0.0763f
C3759 a_4396_12822# a_4696_10916# 6.48e-19
C3760 X2.X2.X1.X1.X1.X1.X3.vin2 a_46116_30882# 0.354f
C3761 X2.X2.X1.X1.X2.X2.X1.vin2 a_46502_19446# 8.88e-20
C3762 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 0.049f
C3763 a_46116_4198# a_46502_4198# 0.419f
C3764 a_8186_29834# X1.X1.X2.X2.X2.X1.X3.vin2 0.00815f
C3765 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.X3.vin1 0.0131f
C3766 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X2.vin1 0.564f
C3767 X2.X2.X2.vrefh a_46502_4198# 0.301f
C3768 X1.X1.X2.X1.X2.X1.vout X1.X1.X2.X1.X2.X1.X3.vin1 0.118f
C3769 X2.X1.X1.X1.X2.X1.vout X2.X1.X1.X1.X2.X1.X3.vin2 0.326f
C3770 a_39966_30794# a_37852_29834# 2.68e-20
C3771 X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X3.vin1 0.0604f
C3772 a_54606_7922# X2.X2.X2.X1.X1.X2.vrefh 8.22e-20
C3773 X1.X2.X1.X1.X2.X2.X2.vin1 a_17222_19446# 0.402f
C3774 X2.X2.X2.X1.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X3.vin1 0.581f
C3775 X2.X2.X2.X2.X3.vin2 X2.X2.X1.X3.vin1 7.46e-20
C3776 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin2 0.12f
C3777 X2.X2.X2.X1.X2.X1.vout a_52492_14586# 0.169f
C3778 a_34362_22312# X2.X1.X1.X1.X2.X2.vout 0.263f
C3779 a_4696_22312# X1.X1.X1.X1.X2.X2.X3.vin1 0.00329f
C3780 a_10686_17452# X1.X1.X2.X1.X2.X2.X3.vin1 0.00207f
C3781 a_10686_25076# X1.X1.X2.X2.X1.X2.X3.vin2 0.567f
C3782 a_52792_12640# a_52492_10734# 6.2e-19
C3783 a_46502_15634# a_46502_13728# 0.00198f
C3784 a_46116_15634# X2.X2.X1.X2.X1.X2.X1.vin1 1.64e-19
C3785 a_8186_10734# X1.X1.X2.X1.X3.vin1 0.385f
C3786 X1.X1.X2.X2.X1.X1.X1.vin1 a_11072_19358# 0.195f
C3787 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin2 0.12f
C3788 a_10686_32700# a_8872_31700# 1.15e-20
C3789 X1.X2.X2.X2.X1.X2.X3.vin1 a_25712_23170# 0.354f
C3790 a_25326_15546# X1.X2.X2.X1.X2.X2.vrefh 8.22e-20
C3791 a_8572_14586# a_10686_13640# 2.95e-20
C3792 a_34062_16634# X2.X1.X1.X2.X1.X1.vout 0.422f
C3793 a_48316_28070# X2.X2.X1.X1.X1.X2.X3.vin2 0.101f
C3794 X2.X1.X2.X1.X1.X1.X2.vin1 a_40352_6016# 0.197f
C3795 a_52792_24076# a_52492_22210# 6.71e-19
C3796 a_46502_25164# a_48316_24258# 1.06e-19
C3797 a_19036_24258# a_17222_23258# 1.15e-20
C3798 a_25326_17452# X1.X2.X2.X1.X2.X2.X3.vin2 0.567f
C3799 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X2.vin1 0.0689f
C3800 X2.X1.X2.vrefh a_31476_4198# 0.119f
C3801 a_22826_25982# X1.X2.X2.X2.X1.X2.X3.vin2 0.00846f
C3802 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin1 0.52f
C3803 a_16836_27070# X1.X2.X1.X1.X2.X1.X1.vin1 1.64e-19
C3804 a_17222_27070# a_17222_25164# 0.00198f
C3805 a_46116_32788# a_46116_30882# 0.00396f
C3806 a_37766_12640# a_37466_10734# 5.25e-20
C3807 a_52792_20264# a_52492_18358# 6.2e-19
C3808 a_31862_27070# a_33976_26164# 4.72e-20
C3809 X2.X1.X1.X3.vin2 X2.X1.X2.X1.X3.vin2 7.46e-20
C3810 X2.X1.X2.X3.vin1 a_37466_14586# 7.98e-19
C3811 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 1.22e-19
C3812 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X3.vin1 2.33e-19
C3813 X1.X1.X1.X1.X1.X2.X3.vin1 a_4782_28070# 0.42f
C3814 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 2.23e-19
C3815 X1.X1.X1.X2.X2.X2.X2.vin1 a_2196_4198# 0.197f
C3816 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X3.vin1 1.22e-19
C3817 a_39966_9828# X2.X1.X2.X1.X1.X2.X1.vin2 8.88e-20
C3818 a_4396_12822# X1.X1.X1.X2.X1.X2.X3.vin2 0.101f
C3819 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin2 0.1f
C3820 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.vrefh 0.161f
C3821 X2.X1.X2.X2.X1.X2.X3.vin1 a_37852_22210# 0.00329f
C3822 X1.X1.X2.X2.X1.X1.X3.vin2 a_10686_19358# 7.84e-19
C3823 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X1.vin1 0.0689f
C3824 a_4696_14688# X1.X1.X1.X2.X3.vin1 0.363f
C3825 a_16836_4198# a_17222_4198# 0.419f
C3826 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 2.23e-19
C3827 X1.X2.X1.X3.vin1 X1.X2.X2.X3.vin2 1.22e-19
C3828 a_48616_18540# X2.X2.X1.X3.vin2 0.0927f
C3829 X1.X2.X2.vrefh a_17222_4198# 0.301f
C3830 a_23512_5016# a_25326_4110# 1.06e-19
C3831 a_25326_7922# X1.X2.X2.X1.X1.X2.vrefh 8.22e-20
C3832 X2.X1.X1.X3.vin1 X2.X1.X3.vin1 0.188f
C3833 a_34062_9010# X2.X1.X1.X2.X2.X1.vout 0.422f
C3834 X1.X1.X1.X2.X2.vrefh a_2196_9916# 1.64e-19
C3835 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X2.X3.vin1 1.22e-19
C3836 X1.X2.X1.X2.X1.X2.X3.vin2 a_19336_10916# 0.00535f
C3837 X1.X1.X1.X2.X1.X2.X1.vin2 a_2582_11822# 8.88e-20
C3838 a_19422_12822# a_19722_10916# 4.41e-20
C3839 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X1.vout 0.033f
C3840 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X2.vin1 0.242f
C3841 X2.X1.X2.X2.X1.X2.X1.vin2 a_40352_23170# 0.12f
C3842 a_39966_23170# X2.X1.X2.X2.X1.X2.X1.vin1 0.417f
C3843 a_54606_30794# a_52492_29834# 2.68e-20
C3844 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X1.X1.vin1 0.206f
C3845 X1.X1.X2.X3.vin2 a_8186_18358# 0.263f
C3846 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X3.vin1 0.0321f
C3847 X1.X1.X2.X1.X2.X2.X1.vin1 a_10686_13640# 8.22e-20
C3848 X1.X2.X3.vin1 a_22826_18358# 5.87e-20
C3849 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X1.X2.X1.X2.X1.X3.vin2 3.94e-19
C3850 X2.X2.X2.X1.X1.X1.vout X2.X2.X2.X1.X1.X1.X3.vin1 0.118f
C3851 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin2 0.12f
C3852 X1.X2.X1.X2.X2.X1.X3.vin1 a_19036_9010# 0.199f
C3853 X1.X1.X2.vrefh a_6032_892# 7.3e-19
C3854 X1.X1.X1.X2.X2.X2.vrefh X1.X1.X1.X2.X2.X2.X1.vin2 0.1f
C3855 a_22826_10734# X1.X2.X2.X1.X1.X2.X3.vin2 0.00846f
C3856 a_10686_21264# X1.X1.X2.X2.X1.X1.X2.vin1 0.402f
C3857 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X1.vin1 0.267f
C3858 X1.X1.X1.X1.X1.X1.X3.vin2 a_2582_30882# 0.567f
C3859 X1.X2.X1.X2.X2.X1.X3.vin2 X1.X2.X1.X2.X2.X2.vrefh 0.161f
C3860 a_52792_8828# a_52106_6962# 3.31e-19
C3861 a_48616_14688# X2.X2.X1.X2.X1.X2.X3.vin1 0.00329f
C3862 X2.X1.X2.X2.X3.vin2 a_37852_29834# 0.363f
C3863 X1.X1.X2.X1.X2.X1.X3.vin2 a_11072_13640# 0.354f
C3864 a_4696_7064# X1.X1.X1.X2.X2.X2.vout 0.0929f
C3865 a_31862_28976# a_31862_27070# 0.00198f
C3866 X2.X2.X1.X1.X1.X1.X2.vin1 X2.X2.X1.X1.X1.X1.X3.vin2 0.234f
C3867 X2.X1.X1.X1.X1.X2.X3.vin1 X2.X1.X1.X1.X2.vrefh 0.00118f
C3868 X2.X1.X2.X2.X2.X1.X3.vin2 X2.X1.X2.X2.X2.X1.X3.vin1 0.581f
C3869 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X3.vin1 0.206f
C3870 X1.X2.X2.X2.X2.X2.X1.vin1 a_25326_28888# 8.22e-20
C3871 X1.X2.X2.X2.X2.X2.X1.vin2 X1.X2.X2.X2.X2.X1.X3.vin2 3.94e-19
C3872 a_22826_10734# a_23512_8828# 3.08e-19
C3873 X1.X1.X2.X3.vin2 a_8486_20264# 5.21e-19
C3874 a_54606_13640# a_52792_12640# 1.15e-20
C3875 a_34362_7064# X2.X1.X1.X2.X2.X2.X3.vin2 3.85e-19
C3876 X1.X2.X1.X2.X2.X2.X3.vin1 a_19422_5198# 0.42f
C3877 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 2.23e-19
C3878 X2.X1.X1.X2.X2.X2.vout a_34062_5198# 0.418f
C3879 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X1.vin1 5.19e-19
C3880 X2.X1.X2.X2.X2.X2.vout X2.X1.X2.X2.X2.X1.vout 0.514f
C3881 a_46502_13728# X2.X2.X1.X2.X1.X2.X2.vin1 8.88e-20
C3882 a_39966_26982# a_39966_25076# 0.00198f
C3883 X2.X1.X2.X1.X1.X2.X3.vin1 a_37466_6962# 0.00874f
C3884 X3.vin1 a_20286_892# 5.17e-19
C3885 a_37766_31700# a_39966_30794# 4.2e-20
C3886 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 0.22f
C3887 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin1 0.199f
C3888 X2.X1.X2.X1.X2.X1.vout X2.X1.X2.X1.X3.vin2 0.399f
C3889 a_54606_25076# X2.X2.X2.X2.X1.X2.X3.vin1 0.00207f
C3890 a_54992_9828# a_54992_7922# 0.00396f
C3891 a_2196_25164# a_2582_25164# 0.419f
C3892 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X1.X2.X1.X1.X1.X3.vin2 5.19e-19
C3893 X2.X2.X1.X2.X3.vin2 a_48616_7064# 0.363f
C3894 X1.X2.X2.X1.X2.X2.X3.vin2 a_22826_14586# 3.85e-19
C3895 a_16836_17540# a_17222_17540# 0.419f
C3896 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X2.X1.X2.X1.X1.X1.vin2 0.00232f
C3897 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X2.X1.X1.X1.X1.X1.vin2 0.00232f
C3898 a_19036_24258# a_19422_24258# 0.419f
C3899 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X2.vrefh 0.076f
C3900 a_25326_6016# X1.X2.X2.X1.X1.X1.X2.vin1 0.402f
C3901 X2.X1.X2.X2.X1.X2.X3.vin2 a_38152_24076# 0.101f
C3902 X1.X1.X2.X2.X3.vin2 a_8572_25982# 0.0927f
C3903 a_25326_23170# a_25326_21264# 0.00198f
C3904 X2.X1.X1.X1.X1.X2.X3.vin1 X2.X1.X1.X1.X1.X2.X1.vin2 0.216f
C3905 a_34362_26164# X2.X1.X1.X1.X3.vin2 0.241f
C3906 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X2.vin1 0.242f
C3907 X1.X2.X2.X2.X2.X1.vout a_23512_27888# 0.359f
C3908 X1.X2.X2.X1.X2.X2.X3.vin1 a_23512_16452# 0.199f
C3909 a_46116_32788# X2.X2.X1.X1.X1.X1.X2.vin1 1.78e-19
C3910 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X2.X1.X2.X1.X2.vrefh 0.0128f
C3911 X1.X2.X3.vin2 X1.X2.X1.X2.X3.vin1 4.41e-19
C3912 X1.X2.X3.vin1 X1.X2.X2.X1.X3.vin2 6.26e-19
C3913 X1.X2.X1.X1.X2.X1.X3.vin1 a_17222_23258# 0.00207f
C3914 X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X2.X1.X1.vin1 0.267f
C3915 X1.X2.X2.vrefh X1.X3.vin2 4.75e-20
C3916 X2.X2.X2.X2.X2.X1.X2.vin1 a_54606_26982# 8.88e-20
C3917 X2.X2.X2.X2.X2.X1.X3.vin2 X2.X2.X2.X2.X2.X1.X1.vin2 8.93e-19
C3918 a_40352_6016# a_40352_4110# 0.00396f
C3919 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X3.vin2 8.93e-19
C3920 a_33976_18540# X2.X1.X3.vin1 0.354f
C3921 X2.X1.X1.X1.X2.X2.X3.vin2 a_34362_18540# 0.00846f
C3922 X2.X2.X2.X2.X2.X2.X1.vin2 X2.X2.X2.X2.X2.X2.X1.vin1 0.668f
C3923 a_34062_20446# X2.X1.X3.vin1 1.64e-19
C3924 a_23126_24076# a_22826_22210# 5.55e-20
C3925 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 0.234f
C3926 X1.X2.X1.X1.X2.vrefh a_16836_27070# 0.118f
C3927 X1.X2.X2.X1.X2.X2.X2.vin1 a_25712_15546# 1.78e-19
C3928 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X3.vin1 0.587f
C3929 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X1.vin1 2.23e-19
C3930 a_8486_12640# a_8572_10734# 3.21e-19
C3931 X2.X2.X2.X2.X2.X2.vout a_52106_29834# 0.263f
C3932 X2.X2.X2.X2.X2.vrefh a_54992_25076# 0.118f
C3933 X1.X1.X1.X2.X1.X1.vout X1.X1.X1.X2.X1.X1.X3.vin2 0.342f
C3934 X1.X2.X2.X1.X1.X2.X3.vin1 a_23512_8828# 0.199f
C3935 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.X1.vin2 3.94e-19
C3936 X2.X2.X1.X1.X1.X1.X1.vin1 X2.X2.X1.X1.X1.X1.X1.vin2 0.696f
C3937 X1.X1.X3.vin1 X1.X1.X1.X3.vin2 1.04f
C3938 a_19722_26164# a_19422_24258# 5.25e-20
C3939 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X2.X1.X2.X2.X2.vrefh 0.0128f
C3940 a_19336_26164# X1.X2.X1.X1.X2.X1.vout 1.64e-19
C3941 a_39966_28888# a_38152_27888# 1.15e-20
C3942 X1.X2.X3.vin1 a_23126_12640# 8.66e-20
C3943 X1.X1.X1.X1.X2.X1.vout a_5082_22312# 0.383f
C3944 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin2 0.12f
C3945 a_4396_31882# X1.X1.X1.X1.X1.X1.vout 0.359f
C3946 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X2.vin1 0.0689f
C3947 a_17222_32788# a_19036_31882# 1.06e-19
C3948 X2.X2.X1.X1.X1.X2.vout a_48316_28070# 0.36f
C3949 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X2.X1.X1.X1.X1.X2.vin1 0.00232f
C3950 a_31862_28976# X2.X1.X1.X1.X1.X2.X2.vin1 8.88e-20
C3951 X1.X2.X2.X2.X2.X1.vout a_23212_29834# 0.169f
C3952 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.vrefh 2.33e-19
C3953 X1.X2.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X3.vin2 0.0533f
C3954 X2.X1.X1.X2.X1.X2.vrefh a_31476_15634# 0.118f
C3955 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.X3.vin1 0.00836f
C3956 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X2.vin1 0.242f
C3957 X2.X2.X1.X1.X3.vin1 a_49002_26164# 0.385f
C3958 a_37766_31700# X2.X1.X2.X2.X3.vin2 9.7e-20
C3959 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X2.vin1 0.0689f
C3960 X1.X2.X1.X2.X2.X2.vrefh a_17222_6104# 8.22e-20
C3961 a_40352_23170# a_40352_21264# 0.00396f
C3962 a_5646_892# a_6032_892# 0.419f
C3963 X2.X1.X3.vin2 a_37466_10734# 6.66e-19
C3964 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X1.X3.vin1 0.0425f
C3965 a_48316_28070# a_48616_26164# 6.48e-19
C3966 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 0.242f
C3967 a_39966_25076# a_39966_23170# 0.00198f
C3968 X2.X2.X2.X2.X3.vin1 a_52406_20264# 1.52e-19
C3969 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X2.vout 0.2f
C3970 X2.X1.X2.X2.X1.X1.vout a_37766_20264# 0.422f
C3971 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin2 0.1f
C3972 a_10686_32700# X1.X1.X2.X2.X2.X2.X3.vin2 0.567f
C3973 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X3.vin2 8.93e-19
C3974 X2.X1.X1.X2.X2.X2.vrefh a_31476_8010# 0.118f
C3975 a_46502_9916# X2.X2.X1.X2.X2.X1.X1.vin2 0.273f
C3976 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X1.vout 0.131f
C3977 X1.X2.X2.X2.X3.vin2 a_23126_27888# 0.00101f
C3978 a_37852_14586# a_38152_12640# 6.1e-19
C3979 X2.X2.X2.X1.X3.vin1 a_52406_5016# 1.52e-19
C3980 X2.X1.X1.X3.vin2 a_34362_14688# 0.00292f
C3981 X1.X2.X2.X1.X2.X1.X3.vin2 a_23126_12640# 0.267f
C3982 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X3.vin1 0.00117f
C3983 a_54606_21264# X2.X2.X2.X2.X1.X1.X3.vin2 0.567f
C3984 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 0.234f
C3985 X1.X2.X2.X2.X2.X1.X2.vin1 a_25712_28888# 0.197f
C3986 a_19722_26164# X1.X2.X1.X3.vin1 0.509f
C3987 a_17222_28976# X1.X2.X1.X1.X1.X2.X3.vin1 0.52f
C3988 X1.X2.X2.vrefh a_28096_892# 4.63e-19
C3989 a_39966_23170# X2.X1.X2.X2.X1.X2.vrefh 8.22e-20
C3990 X1.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin1 0.00437f
C3991 a_11072_30794# X1.X1.X2.X2.X2.X2.vrefh 1.64e-19
C3992 a_19722_7064# X1.X2.X1.X2.X2.X2.X3.vin1 0.00874f
C3993 a_48316_24258# X2.X2.X1.X1.X2.X1.vout 0.359f
C3994 a_31862_15634# a_33976_14688# 2.95e-20
C3995 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X1.X3.vin2 1.22e-19
C3996 X1.X2.X1.X1.X2.X1.X3.vin1 a_19422_24258# 0.428f
C3997 X2.X1.X3.vin1 a_37466_6962# 6.45e-19
C3998 a_33976_26164# a_34062_24258# 3.21e-19
C3999 a_34362_26164# a_33676_24258# 2.97e-19
C4000 a_37466_10734# a_37766_8828# 4.41e-20
C4001 X2.X2.X1.X1.X2.X2.vout X2.X2.X1.X1.X2.X2.X3.vin1 0.335f
C4002 a_25712_17452# X1.X2.X2.X1.X2.X2.X1.vin2 1.78e-19
C4003 X2.X1.X2.X1.X1.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X3.vin1 0.581f
C4004 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X2.vrefh 0.00118f
C4005 a_52106_14586# X2.X2.X2.X1.X2.X1.X3.vin2 0.00815f
C4006 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin1 0.195f
C4007 a_25326_11734# X1.X2.X2.X1.X2.vrefh 8.22e-20
C4008 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X2.X1.X2.X1.X2.vrefh 0.00437f
C4009 a_37466_22210# X2.X1.X2.X2.X1.X1.X3.vin2 0.00815f
C4010 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X1.vin2 0.076f
C4011 a_52406_31700# X2.X2.X2.X2.X2.X2.vout 0.418f
C4012 a_23126_20264# a_23212_18358# 3.21e-19
C4013 X1.X1.X2.X1.X1.X2.X3.vin2 a_10686_7922# 7.84e-19
C4014 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X1.vin1 0.0689f
C4015 X1.X2.X2.X2.X2.X2.X2.vin1 a_23126_31700# 0.00351f
C4016 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin2 0.1f
C4017 a_25326_32700# X1.X2.X2.X2.X2.X2.X3.vin1 0.00207f
C4018 a_48616_10916# a_49002_10916# 0.414f
C4019 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.X3.vin1 0.0174f
C4020 X1.X2.X1.X2.X1.X1.vout a_19336_14688# 0.169f
C4021 X1.X1.X1.X2.X3.vin1 a_4782_12822# 9.54e-19
C4022 X1.X2.X1.X3.vin2 a_19422_12822# 6.03e-19
C4023 a_19422_16634# a_19722_14688# 4.19e-20
C4024 a_4696_7064# a_4396_5198# 6.71e-19
C4025 a_5082_14688# X1.X1.X1.X2.X1.X2.X3.vin2 3.85e-19
C4026 X2.X2.X2.X2.X1.X1.X3.vin2 a_52106_18358# 3.49e-19
C4027 a_54606_26982# a_54992_26982# 0.419f
C4028 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin2 0.1f
C4029 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X3.vin2 0.0533f
C4030 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X3.vin1 1.42e-20
C4031 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X3.vin2 0.161f
C4032 X2.X1.X2.X1.X3.vin2 a_37852_10734# 0.0927f
C4033 X1.X2.X3.vin2 X1.X2.X2.X1.X2.X2.vout 3.38e-19
C4034 a_4396_9010# a_4696_7064# 6.1e-19
C4035 X1.X1.X2.X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X2.vin1 0.564f
C4036 X1.X2.X2.X1.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin1 0.00437f
C4037 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X1.vin1 2.23e-19
C4038 X1.X1.X2.X1.X1.X1.X2.vin1 a_11072_4110# 1.78e-19
C4039 a_39966_13640# X2.X1.X2.X1.X2.X1.X1.vin2 8.88e-20
C4040 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin2 0.1f
C4041 X1.X1.X2.X2.X2.X1.vout X1.X1.X2.X2.X3.vin2 0.399f
C4042 X1.X1.X1.X1.X2.X2.X3.vin2 a_5082_18540# 0.00846f
C4043 a_4782_20446# X1.X1.X3.vin1 1.64e-19
C4044 X1.X2.X3.vin2 X1.X2.X2.vrefh 0.15f
C4045 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X3.vin2 8.93e-19
C4046 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.X3.vin2 0.581f
C4047 X2.X1.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X1.X3.vin1 0.0321f
C4048 X2.X2.X3.vin1 X2.X2.X1.X2.X3.vin2 0.0816f
C4049 a_31862_23258# X2.X1.X1.X1.X2.X2.X1.vin1 8.22e-20
C4050 a_48616_22312# a_48316_20446# 6.71e-19
C4051 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X2.X1.X2.X2.X2.vrefh 0.00437f
C4052 a_10686_11734# X1.X1.X2.X1.X2.X1.X1.vin1 0.417f
C4053 X1.X1.X2.X1.X2.X1.X1.vin2 a_11072_11734# 0.12f
C4054 X1.X2.X2.X1.X2.X1.X1.vin1 a_25712_9828# 1.64e-19
C4055 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.vout 0.0898f
C4056 X2.X1.X2.X2.X2.X1.X1.vin1 a_40352_26982# 0.195f
C4057 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X3.vin1 0.0131f
C4058 a_39966_15546# a_39966_13640# 0.00198f
C4059 a_2196_8010# a_2196_6104# 0.00396f
C4060 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.X2.vin1 0.00117f
C4061 a_46502_9916# a_48702_9010# 4.2e-20
C4062 X1.X1.X3.vin2 a_8486_16452# 3.98e-19
C4063 a_46502_15634# a_48616_14688# 2.95e-20
C4064 X1.X1.X1.X2.X1.X2.X2.vin1 a_2196_11822# 0.197f
C4065 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin1 0.267f
C4066 X1.X2.X3.vin1 X1.X2.X2.X1.X3.vin1 0.00304f
C4067 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 0.587f
C4068 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X2.vin1 0.564f
C4069 X2.X2.X1.X2.X1.X2.X2.vin1 a_46116_11822# 0.197f
C4070 a_37766_27888# a_37466_25982# 5.25e-20
C4071 X2.X2.X2.X1.X1.X1.X3.vin2 X2.X2.X2.X1.X1.X1.X1.vin1 2.23e-19
C4072 X2.X2.X2.X1.X1.X1.X2.vin1 a_54992_4110# 1.78e-19
C4073 a_52406_12640# X2.X2.X2.X1.X2.X1.X3.vin1 0.428f
C4074 a_48616_26164# a_48316_24258# 6.2e-19
C4075 a_2196_32788# a_2582_32788# 0.419f
C4076 X2.X2.X2.X2.X2.X2.X1.vin1 a_54606_28888# 8.22e-20
C4077 X2.X2.X2.X2.X2.X2.X1.vin2 X2.X2.X2.X2.X2.X1.X3.vin2 3.94e-19
C4078 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X3.vin1 0.00118f
C4079 a_16836_13728# X1.X2.X1.X2.X1.X2.X2.vin1 1.78e-19
C4080 X2.X1.X1.X1.X2.X1.X3.vin2 a_34362_22312# 0.00815f
C4081 X1.X2.X1.X1.X1.X1.X3.vin2 a_16836_30882# 0.354f
C4082 a_46116_21352# a_46502_21352# 0.419f
C4083 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X1.vin1 0.0689f
C4084 X2.X1.X2.X2.X2.X2.X3.vin2 a_39966_30794# 7.84e-19
C4085 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X2.X1.X1.X2.X2.X1.vin2 0.00232f
C4086 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin1 0.195f
C4087 X1.X1.X1.X1.X1.X1.X3.vin2 a_5082_29936# 0.00815f
C4088 a_46502_13728# X2.X2.X1.X2.X1.X2.X1.vin2 0.273f
C4089 X1.X2.X3.vin1 a_19722_14688# 3.28e-19
C4090 a_37852_25982# X2.X1.X2.X2.X1.X2.vout 7.93e-20
C4091 X1.X1.X2.X1.X1.X2.X3.vin1 a_11072_7922# 0.354f
C4092 a_17222_23258# a_19336_22312# 2.95e-20
C4093 a_10686_28888# X1.X1.X2.X2.X2.X1.X2.vin1 0.402f
C4094 a_10686_13640# X1.X1.X2.X1.X2.X1.X3.vin1 0.00207f
C4095 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 0.234f
C4096 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X2.vin1 0.242f
C4097 X2.X2.X2.X1.X2.X2.X3.vin1 a_54606_15546# 0.52f
C4098 a_4396_9010# a_2582_8010# 1.15e-20
C4099 a_34062_16634# a_33976_14688# 3.14e-19
C4100 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X3.vin2 0.102f
C4101 a_10686_6016# a_8486_5016# 4.77e-21
C4102 X1.X2.X2.X2.X1.X1.X1.vin1 X2.X1.X1.X2.vrefh 0.00437f
C4103 a_33676_16634# a_34362_14688# 2.86e-19
C4104 a_33676_12822# a_31862_11822# 1.15e-20
C4105 X2.X2.X1.X2.X1.X1.X2.vin1 a_46116_15634# 0.197f
C4106 a_39966_7922# X2.X1.X2.X1.X1.X1.X3.vin2 8.07e-19
C4107 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.vrefh 0.161f
C4108 a_39966_6016# a_38152_5016# 1.15e-20
C4109 X1.X1.X2.X2.X2.X2.vrefh X1.X1.X2.X2.X2.X1.X3.vin1 0.00118f
C4110 a_8186_22210# a_8486_20264# 4.19e-20
C4111 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X3.vin1 0.00836f
C4112 a_16836_17540# a_16836_15634# 0.00396f
C4113 X1.X1.X1.X2.vrefh a_2582_17540# 8.22e-20
C4114 a_31862_6104# X2.X1.X1.X2.X2.X2.X2.vin1 8.88e-20
C4115 X1.X2.X2.X1.X1.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin1 0.00437f
C4116 X1.X1.X2.X1.X1.X1.vout a_8572_6962# 0.169f
C4117 a_37466_18358# a_38152_16452# 3.08e-19
C4118 a_2582_27070# a_4696_26164# 4.72e-20
C4119 X2.X2.X1.X1.X1.X1.vout X2.X2.X1.X1.X1.X2.vout 0.507f
C4120 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 2.23e-19
C4121 a_37766_24076# a_38152_24076# 0.419f
C4122 X1.X1.X2.X1.X1.X1.vout a_8872_5016# 0.359f
C4123 a_54606_23170# a_54606_21264# 0.00198f
C4124 a_37852_6962# a_38152_5016# 6.1e-19
C4125 X2.X2.X1.X1.X1.X2.X3.vin2 a_46502_25164# 8.07e-19
C4126 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 5.19e-19
C4127 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X2.X1.X2.vrefh 0.00437f
C4128 X1.X1.X3.vin1 a_8486_8828# 8.66e-20
C4129 X2.X2.X2.X1.X1.X2.X3.vin1 a_54606_7922# 0.52f
C4130 X2.X2.X1.X1.X2.X1.X3.vin1 a_46502_23258# 0.00207f
C4131 a_25326_28888# X1.X2.X2.X2.X2.X1.X1.vin2 8.88e-20
C4132 a_23212_18358# a_23126_16452# 3.3e-19
C4133 a_48616_14688# X2.X2.X1.X2.X3.vin1 0.363f
C4134 a_54992_19358# X2.X2.X2.X2.vrefh 1.64e-19
C4135 X1.X1.X2.X1.X2.X2.X3.vin1 a_8572_14586# 0.00329f
C4136 a_11072_6016# X1.X1.X2.X1.X1.X1.X1.vin2 1.78e-19
C4137 X1.X1.X1.X2.X1.X1.X3.vin1 a_4396_16634# 0.199f
C4138 X2.X2.X2.X2.X1.X1.vout a_52792_20264# 0.359f
C4139 X2.X2.X1.X2.X2.X1.X2.vin1 a_46116_8010# 0.197f
C4140 X2.X1.X1.X2.X2.X1.vout a_33976_7064# 0.169f
C4141 a_34062_9010# a_34362_7064# 4.19e-20
C4142 X2.X2.X2.X1.X3.vin1 a_52492_6962# 0.363f
C4143 X2.X2.X2.X2.X2.X1.X3.vin1 a_52106_25982# 0.00837f
C4144 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X3.vin2 8.93e-19
C4145 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X3.vin1 0.00117f
C4146 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X1.vin1 2.23e-19
C4147 X2.X2.X2.X1.X1.X2.X3.vin2 a_52406_8828# 0.277f
C4148 X2.X2.X2.X1.X2.X2.X2.vin1 a_54992_15546# 1.78e-19
C4149 X2.X2.X1.X1.X2.X2.X3.vin2 a_46502_19446# 0.567f
C4150 X2.X1.X1.X3.vin2 a_34362_10916# 0.452f
C4151 a_17222_11822# a_17222_9916# 0.00198f
C4152 a_16836_11822# X1.X2.X1.X2.X2.X1.X1.vin1 1.64e-19
C4153 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.vout 0.398f
C4154 X1.X1.X2.vrefh a_10686_4110# 4.89e-19
C4155 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X3.vin1 2.33e-19
C4156 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 1.22e-19
C4157 X2.X2.X2.X3.vin2 a_52106_18358# 0.263f
C4158 a_10686_23170# a_11072_23170# 0.419f
C4159 X2.X2.X1.X1.X2.X2.vrefh a_46502_23258# 0.3f
C4160 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X2.X1.X1.X2.X2.X2.vin1 0.00232f
C4161 a_54992_6016# X2.X2.X2.X1.X1.X1.X1.vin2 1.78e-19
C4162 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X2.vout 0.2f
C4163 a_48316_16634# a_48616_14688# 6.1e-19
C4164 X2.X2.X2.X1.X1.X2.vrefh a_54992_6016# 0.118f
C4165 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X1.vin2 3.94e-19
C4166 a_23212_6962# X1.X2.X2.X1.X1.X1.X3.vin2 0.00546f
C4167 a_49002_10916# X2.X2.X1.X2.X2.X1.X3.vin2 3.49e-19
C4168 X2.X1.X1.X2.X1.X1.X1.vin2 a_31862_15634# 8.88e-20
C4169 a_54992_15546# X2.X2.X2.X1.X2.X2.vrefh 1.64e-19
C4170 a_31862_19446# a_33976_18540# 4.72e-20
C4171 X2.X1.X1.X1.X2.X2.X3.vin2 a_31476_19446# 0.354f
C4172 X2.X1.X2.X1.X2.X2.vout a_37852_14586# 0.0929f
C4173 a_34062_20446# a_31862_19446# 4.77e-21
C4174 X2.X2.X1.X2.X2.X2.vrefh a_46502_6104# 8.22e-20
C4175 a_19036_31882# X1.X2.X1.X1.X1.X1.X3.vin2 0.1f
C4176 X1.X2.X1.X2.vrefh a_16836_17540# 1.64e-19
C4177 X2.X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X2.X2.vrefh 0.117f
C4178 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin1 0.195f
C4179 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X1.vin1 0.206f
C4180 X1.X1.X2.X2.X1.X2.X2.vin1 a_11072_23170# 1.78e-19
C4181 a_19036_24258# a_19722_22312# 2.86e-19
C4182 a_19422_24258# a_19336_22312# 3.14e-19
C4183 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X1.vin1 2.23e-19
C4184 X2.X1.X2.X1.X2.X1.X3.vin1 a_38152_12640# 0.199f
C4185 a_25712_32700# a_25712_30794# 0.00396f
C4186 X1.X1.X1.X2.X1.X1.X2.vin1 a_2582_15634# 0.402f
C4187 a_4782_12822# a_5082_10916# 4.41e-20
C4188 X1.X1.X1.X2.X1.X2.X3.vin2 a_4696_10916# 0.00535f
C4189 X1.X2.X2.X2.X1.X1.X1.vin2 X2.X1.X1.X1.X2.X2.X2.vin1 0.00232f
C4190 X1.X1.X1.X2.X2.X1.X3.vin2 X1.X1.X1.X2.X2.X2.X1.vin2 3.94e-19
C4191 X1.X1.X2.X2.X1.X2.vout X1.X1.X2.X2.X1.X1.vout 0.507f
C4192 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X1.vin1 5.19e-19
C4193 a_8572_6962# a_8486_5016# 3.14e-19
C4194 a_8486_31700# X1.X1.X2.X2.X2.X2.X3.vin1 0.42f
C4195 X2.X2.X2.vrefh X2.X2.X2.X1.X1.X1.X1.vin2 0.096f
C4196 X1.X1.X2.X2.X2.X1.X3.vin1 X1.X1.X2.X2.X2.vrefh 2.33e-19
C4197 a_17222_17540# X1.X2.X1.X2.X1.X1.X2.vin1 8.88e-20
C4198 a_54992_7922# X2.X2.X2.X1.X1.X2.vrefh 1.64e-19
C4199 a_8486_5016# a_8872_5016# 0.419f
C4200 a_33976_29936# X2.X1.X1.X1.X1.X2.vout 0.0929f
C4201 a_19422_20446# a_17222_19446# 4.77e-21
C4202 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X1.vin2 0.076f
C4203 X1.X2.X1.X1.X2.X2.X3.vin2 a_16836_19446# 0.354f
C4204 X2.X2.X2.X2.X3.vin2 a_52492_25982# 0.0927f
C4205 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X1.vin2 0.668f
C4206 X1.X1.X2.X1.X1.X2.X3.vin1 a_8186_6962# 0.00874f
C4207 X1.X2.vrefh X1.X1.X2.X2.X2.X2.X1.vin2 0.0763f
C4208 X1.X1.X1.X1.X2.X2.vout X1.X1.X1.X1.X2.X2.X3.vin1 0.335f
C4209 a_39966_11734# a_39966_9828# 0.00198f
C4210 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.X3.vin1 0.587f
C4211 X2.X2.X1.X2.X2.X2.vrefh X2.X1.X2.X1.X1.X2.vrefh 0.117f
C4212 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X2.vrefh 0.076f
C4213 X1.X1.X2.X2.X2.X2.X3.vin2 a_8872_31700# 0.101f
C4214 a_52492_22210# a_52406_20264# 3.14e-19
C4215 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X1.vin2 0.668f
C4216 a_8572_14586# X1.X1.X2.X1.X2.X1.X3.vin2 0.00546f
C4217 a_25712_15546# X1.X2.X2.X1.X2.X2.vrefh 1.64e-19
C4218 a_19036_12822# X1.X2.X1.X2.X1.X2.X3.vin2 0.101f
C4219 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X2.X1.X1.X2.X2.X2.vin1 0.00232f
C4220 a_46502_23258# a_48616_22312# 2.95e-20
C4221 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X2.X3.vin2 8.93e-19
C4222 a_2196_6104# a_2196_4198# 0.00396f
C4223 X2.X2.X1.X1.X2.X1.X3.vin1 a_48316_24258# 0.199f
C4224 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X1.X3.vin2 1.22e-19
C4225 a_25712_21264# a_25712_19358# 0.00396f
C4226 a_39966_11734# a_37852_10734# 5.36e-21
C4227 a_54606_28888# X2.X2.X2.X2.X2.X1.X3.vin2 0.567f
C4228 a_54992_17452# X2.X2.X2.X1.X2.X2.X1.vin2 1.78e-19
C4229 a_39966_19358# a_39966_17452# 0.00198f
C4230 X2.X1.X2.X1.X3.vin1 a_37466_6962# 0.436f
C4231 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.vrefh 0.161f
C4232 a_46502_32788# a_46502_30882# 0.00198f
C4233 X2.X2.X2.X1.X1.X1.vout X2.X2.X2.X1.X1.X1.X3.vin2 0.342f
C4234 X1.X2.X2.X2.X2.X2.X1.vin2 a_25326_30794# 0.273f
C4235 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X3.vin2 8.93e-19
C4236 a_48616_7064# a_46502_6104# 2.68e-20
C4237 X2.X1.X2.X2.X2.X1.X3.vin1 a_39966_26982# 0.52f
C4238 X2.X1.X2.X1.X1.X2.X2.vin1 a_39966_7922# 8.88e-20
C4239 a_4396_5198# a_2582_4198# 1.15e-20
C4240 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.X1.vin2 8.93e-19
C4241 X1.X1.X1.X1.X1.X2.vout a_4696_26164# 7.93e-20
C4242 X1.X2.X1.X1.X1.X2.vout a_19036_28070# 0.36f
C4243 a_8872_24076# a_10686_23170# 1.06e-19
C4244 X1.X2.X2.X3.vin2 a_23212_25982# 0.355f
C4245 X1.X1.X1.X1.X2.X2.vrefh a_2582_23258# 0.3f
C4246 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.vrefh 2.33e-19
C4247 X2.X2.X3.vin1 X2.X2.X1.X3.vin2 1.04f
C4248 a_46116_6104# a_46116_4198# 0.00396f
C4249 a_25712_7922# X1.X2.X2.X1.X1.X2.vrefh 1.64e-19
C4250 a_52406_24076# X2.X2.X2.X2.X1.X2.X3.vin1 0.42f
C4251 X1.X2.X2.vrefh X1.X2.X2.X1.X1.X1.X1.vin2 0.096f
C4252 a_19336_18540# a_17222_17540# 5.36e-21
C4253 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X1.vin1 0.267f
C4254 X1.X1.X1.X1.X2.X2.vout a_4696_18540# 7.93e-20
C4255 a_8572_29834# a_8872_27888# 6.1e-19
C4256 a_37766_20264# X2.X1.X3.vin2 7.93e-20
C4257 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X2.vin1 0.564f
C4258 X2.X2.X3.vin1 a_52406_16452# 8.66e-20
C4259 X2.X1.X2.X2.X1.X2.X1.vin1 a_40352_23170# 0.195f
C4260 X1.X2.X1.X2.X2.X1.X1.vin2 a_16836_8010# 1.78e-19
C4261 a_33976_29936# a_31862_28976# 2.68e-20
C4262 a_22826_18358# a_23212_18358# 0.416f
C4263 a_19036_28070# a_19336_26164# 6.48e-19
C4264 a_11072_25076# X1.X1.X2.X2.X1.X2.X1.vin2 1.78e-19
C4265 a_17222_21352# X1.X2.X1.X1.X2.X2.X1.vin2 0.273f
C4266 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 5.19e-19
C4267 X2.X2.X2.X1.X2.vrefh a_54992_9828# 0.118f
C4268 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X1.vin2 0.668f
C4269 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.vout 0.118f
C4270 a_34362_10916# a_33676_9010# 2.97e-19
C4271 a_33976_10916# a_34062_9010# 3.21e-19
C4272 a_8486_16452# a_8872_16452# 0.419f
C4273 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X3.vin2 0.234f
C4274 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X3.vin1 0.0174f
C4275 a_48616_7064# a_48316_5198# 6.71e-19
C4276 X2.X2.X3.vin1 a_52406_8828# 8.66e-20
C4277 a_52106_10734# a_52492_10734# 0.414f
C4278 X1.X1.X3.vin2 X1.X1.X2.vrefh 0.15f
C4279 a_25326_17452# a_23126_16452# 4.77e-21
C4280 X2.X1.X1.X1.X1.X2.X3.vin1 a_31862_27070# 0.00207f
C4281 a_22826_25982# a_23126_24076# 4.41e-20
C4282 a_8486_24076# a_8572_22210# 3.38e-19
C4283 X1.X1.X2.X1.X2.X1.vout a_8872_12640# 0.359f
C4284 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X1.X3.vin2 0.0943f
C4285 a_48702_31882# X2.X2.X1.X1.X1.X1.X3.vin2 0.267f
C4286 a_25326_6016# X1.X2.X2.X1.X1.X1.X1.vin2 8.88e-20
C4287 X2.X2.X1.X2.X1.X2.X1.vin2 a_46116_11822# 1.78e-19
C4288 X1.X2.X2.X2.X2.X2.X1.vin1 X1.X2.X2.X2.X2.X1.X3.vin2 5.19e-19
C4289 X2.X2.X2.X1.X2.X1.X3.vin2 a_52792_12640# 0.1f
C4290 X2.X2.X1.X2.X2.X2.X2.vin1 a_46116_4198# 0.197f
C4291 X2.X2.X1.X2.X2.X2.X2.vin1 X2.X2.X2.vrefh 0.564f
C4292 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X2.vin1 0.00117f
C4293 a_46502_13728# a_48702_12822# 4.2e-20
C4294 a_48616_26164# a_46502_25164# 5.36e-21
C4295 a_39966_26982# X2.X1.X2.X2.X1.X2.X3.vin2 8.07e-19
C4296 X2.X1.X1.X2.X1.X1.X3.vin2 a_31476_15634# 0.354f
C4297 X2.X1.X1.X1.X2.X2.X1.vin2 a_31476_19446# 1.78e-19
C4298 a_19336_29936# X1.X2.X1.X1.X3.vin1 0.363f
C4299 a_10686_25076# a_11072_25076# 0.419f
C4300 X3.vin1 d7 0.0163f
C4301 X2.X1.X2.X2.X3.vin2 X2.X1.X2.X3.vin2 0.17f
C4302 X2.X1.X2.X2.X2.X1.vout a_37852_25982# 1.64e-19
C4303 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.X1.vin1 0.206f
C4304 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X3.vin1 0.587f
C4305 a_46116_19446# a_46116_17540# 0.00396f
C4306 a_2582_25164# X1.X1.X1.X1.X2.X1.X1.vin1 0.417f
C4307 a_2196_25164# X1.X1.X1.X1.X2.X1.X3.vin1 0.354f
C4308 X1.X2.X1.X2.X2.X1.X3.vin2 a_17222_6104# 8.07e-19
C4309 X2.X1.X1.X1.X1.X1.X2.vin1 a_31862_30882# 0.402f
C4310 a_52492_18358# a_54606_17452# 4.72e-20
C4311 a_25326_17452# a_25712_17452# 0.419f
C4312 X2.X1.X1.X1.X1.X2.vout a_34062_28070# 0.418f
C4313 a_52106_14586# a_52406_12640# 4.19e-20
C4314 X2.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X2.vout 0.0866f
C4315 a_31862_6104# X2.X1.X1.X2.X2.X2.X1.vin2 0.273f
C4316 a_10686_23170# X1.X1.X2.X2.X1.X2.vrefh 8.22e-20
C4317 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.X3.vin2 0.0523f
C4318 a_17222_17540# X1.X2.X1.X2.X1.X1.X1.vin1 0.417f
C4319 a_16836_17540# X1.X2.X1.X2.X1.X1.X3.vin1 0.354f
C4320 a_48316_24258# a_48616_22312# 6.1e-19
C4321 X2.X1.X1.X2.X2.X2.X2.vin1 a_31476_4198# 0.197f
C4322 a_19422_24258# X1.X2.X1.X1.X2.X1.vout 0.422f
C4323 a_25712_13640# a_25712_11734# 0.00396f
C4324 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X2.vrefh 2.33e-19
C4325 X1.X1.X2.X2.X1.X1.X3.vin1 a_8872_20264# 0.199f
C4326 a_46116_28976# a_46502_28976# 0.419f
C4327 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X2.X1.X1.X1.X2.X1.vin2 0.00232f
C4328 a_37766_5016# X2.X1.X2.X1.X1.X1.X3.vin1 0.428f
C4329 X2.X1.X1.X2.X2.X2.X2.vin1 X2.X1.X2.vrefh 0.564f
C4330 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X3.vin2 0.234f
C4331 a_46116_17540# a_46116_15634# 0.00396f
C4332 a_25326_23170# X1.X2.X2.X2.X1.X1.X3.vin2 8.07e-19
C4333 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin2 0.1f
C4334 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X1.X3.vin1 0.0321f
C4335 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X1.vin2 3.94e-19
C4336 a_46502_32788# a_48316_31882# 1.06e-19
C4337 X1.X1.X2.X2.X1.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin1 0.00437f
C4338 X2.X2.X1.X1.X1.X1.X1.vin1 X2.X2.X1.X1.X1.X1.X2.vin1 0.0689f
C4339 X2.X1.X2.X2.X1.X2.vout a_37852_22210# 0.0929f
C4340 a_48316_20446# a_48616_18540# 6.48e-19
C4341 X2.X1.X1.X2.X2.X1.X3.vin2 a_31476_8010# 0.354f
C4342 a_33676_28070# a_34362_26164# 3.08e-19
C4343 a_34062_28070# a_33976_26164# 3.3e-19
C4344 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X1.vout 0.033f
C4345 X1.X1.X2.X2.X2.X2.vout X1.X1.X2.X2.X2.X1.vout 0.514f
C4346 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X2.X1.X2.X1.X2.vrefh 0.00437f
C4347 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.vout 0.335f
C4348 a_22826_22210# a_23126_20264# 4.19e-20
C4349 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X2.X1.vin2 3.94e-19
C4350 X1.X1.X2.X2.X3.vin1 a_8572_25982# 0.17f
C4351 X2.X2.X2.X2.X2.X1.X3.vin2 X2.X2.X2.X2.X2.X1.X1.vin1 2.23e-19
C4352 X2.X2.X2.X2.X2.X1.X2.vin1 a_54992_26982# 1.78e-19
C4353 X1.X2.X1.X2.X2.X2.X2.vin1 a_17222_4198# 0.402f
C4354 X1.X2.X1.X3.vin1 X1.X2.X3.vin2 7.53e-21
C4355 X1.X2.X1.X2.X1.X2.vrefh a_17222_13728# 8.22e-20
C4356 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin2 7.84e-19
C4357 a_5082_18540# X1.X1.X1.X2.X1.X1.X3.vin1 0.00837f
C4358 a_54606_30794# a_54992_30794# 0.419f
C4359 a_8186_10734# a_8486_8828# 4.41e-20
C4360 a_16836_27070# a_17222_27070# 0.419f
C4361 a_31476_32788# X2.X1.X1.X1.X1.X1.X2.vin1 1.78e-19
C4362 X2.X2.X2.X2.X2.X1.vout X2.X2.X2.X2.X3.vin2 0.399f
C4363 X2.X2.X2.X1.X1.X1.vout a_52792_5016# 0.359f
C4364 X2.X1.X1.X1.X1.X2.vrefh a_31862_28976# 8.22e-20
C4365 a_2196_25164# a_2196_23258# 0.00396f
C4366 a_19722_29936# X1.X2.X1.X1.X1.X2.X3.vin1 0.00874f
C4367 a_8186_18358# X1.X1.X3.vin2 0.451f
C4368 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin1 0.195f
C4369 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X3.vin1 0.00118f
C4370 X1.X1.X2.X1.X3.vin2 a_8486_12640# 0.00101f
C4371 a_23126_16452# a_22826_14586# 5.55e-20
C4372 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.vout 0.038f
C4373 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X2.X1.X2.X2.X2.vrefh 0.00437f
C4374 X2.X1.X2.X2.X2.X1.X3.vin2 a_38152_27888# 0.1f
C4375 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X2.vrefh 0.076f
C4376 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X1.vin2 0.668f
C4377 X1.X2.X1.X1.X1.X1.X3.vin1 a_19036_31882# 0.199f
C4378 X2.X2.X2.X1.X1.X2.X3.vin2 a_52106_6962# 3.85e-19
C4379 X2.X1.X1.X1.X1.X2.X3.vin1 X2.X1.X1.X1.X1.X2.X2.vin1 0.00117f
C4380 X2.X2.X1.X1.X1.X2.vout X2.X2.X1.X1.X1.X2.X3.vin2 0.075f
C4381 a_31862_28976# a_34062_28070# 4.2e-20
C4382 a_10686_17452# X1.X1.X2.X1.X2.X2.X1.vin2 8.88e-20
C4383 a_8486_20264# X1.X1.X3.vin2 7.93e-20
C4384 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X2.X3.vin1 2.33e-19
C4385 X2.X1.X2.X1.X1.X2.vout a_37466_6962# 0.254f
C4386 X2.X1.X1.X1.X1.X2.vrefh X1.X2.X2.X2.X2.X2.vrefh 0.117f
C4387 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 1.22e-19
C4388 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X2.X1.X2.X2.vrefh 0.0128f
C4389 a_34362_26164# X2.X1.X1.X1.X2.X1.X3.vin1 0.00837f
C4390 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X2.vin1 0.564f
C4391 a_33676_16634# X2.X1.X1.X2.X1.X1.X3.vin2 0.1f
C4392 X1.X3.vin1 a_14082_892# 0.413f
C4393 X2.X1.X1.X1.X2.X2.vrefh a_31476_21352# 1.64e-19
C4394 X1.X1.X2.X1.X1.X2.X1.vin1 a_11072_6016# 1.64e-19
C4395 X1.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X3.vin1 0.552f
C4396 X2.X2.X1.X1.X1.X2.X3.vin2 a_48616_26164# 0.00535f
C4397 a_48702_28070# a_49002_26164# 4.41e-20
C4398 X1.X2.X2.X2.X2.X2.vout X1.X2.X2.X2.X3.vin2 0.0866f
C4399 a_11072_28888# a_11072_26982# 0.00396f
C4400 X2.X1.X2.X2.X1.X2.X3.vin2 a_39966_23170# 7.84e-19
C4401 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X1.vin1 0.0689f
C4402 X1.X1.X3.vin2 a_5646_892# 0.0927f
C4403 X1.X1.X2.vrefh X1.X3.vin1 0.0451f
C4404 X1.X1.X1.X2.X3.vin1 a_5082_10916# 0.372f
C4405 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X2.vin1 0.564f
C4406 a_54606_32700# X2.X2.X2.X2.X2.X2.X3.vin1 0.00207f
C4407 X2.X2.X2.X2.X2.X2.X2.vin1 a_52406_31700# 0.00351f
C4408 X1.X2.X2.X1.X2.X2.X3.vin1 a_25326_15546# 0.52f
C4409 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.X1.vin2 0.216f
C4410 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin1 0.195f
C4411 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X3.vin1 0.0131f
C4412 a_46116_17540# X2.X2.X1.X2.X1.X1.X2.vin1 1.78e-19
C4413 a_39966_11734# X2.X1.X2.X1.X2.vrefh 8.22e-20
C4414 X1.X2.X2.X1.X2.X2.vout a_23512_16452# 0.36f
C4415 X1.X2.X1.X2.X1.X1.X2.vin1 a_16836_15634# 0.197f
C4416 a_52492_10734# X2.X2.X2.X1.X1.X2.vout 7.93e-20
C4417 a_8486_31700# X1.X1.X2.X2.X3.vin2 9.7e-20
C4418 X1.X1.X1.X2.X3.vin2 a_5082_7064# 0.422f
C4419 a_40352_23170# X2.X1.X2.X2.X1.X2.vrefh 1.64e-19
C4420 X1.X2.X1.X1.X2.X1.X1.vin2 a_17222_23258# 8.88e-20
C4421 a_33676_9010# X2.X1.X1.X2.X2.X1.X3.vin2 0.1f
C4422 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X2.vrefh 0.00118f
C4423 a_54992_28888# X2.X2.X2.X2.X2.X1.X1.vin2 1.78e-19
C4424 X1.X1.X3.vin2 X1.X1.X2.X1.X3.vin2 0.039f
C4425 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X2.vin1 0.564f
C4426 X1.X1.X2.X1.X1.X1.vout X1.X1.X2.X1.X1.X1.X3.vin2 0.342f
C4427 X1.X2.X2.X2.X2.X1.X3.vin1 a_22826_25982# 0.00837f
C4428 X2.X1.X1.X3.vin1 a_34062_24258# 5.28e-19
C4429 a_33976_7064# a_34362_7064# 0.419f
C4430 a_4696_7064# a_2582_6104# 2.68e-20
C4431 X2.X2.X2.X2.X1.X2.X2.vin1 a_54992_25076# 0.197f
C4432 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.X3.vin1 0.0174f
C4433 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.vout 0.075f
C4434 a_25712_11734# X1.X2.X2.X1.X2.vrefh 1.64e-19
C4435 a_52492_6962# a_52406_5016# 3.14e-19
C4436 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin1 0.52f
C4437 X1.X2.X2.X1.X1.X2.X3.vin1 a_25326_7922# 0.52f
C4438 X1.X2.X1.X1.X1.X2.X2.vin1 a_16836_27070# 0.197f
C4439 X1.X2.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X2.X1.X2.vin1 0.564f
C4440 a_23212_10734# a_25326_9828# 4.72e-20
C4441 a_2196_15634# a_2196_13728# 0.00396f
C4442 X1.X2.X1.X2.X2.X1.X2.vin1 a_16836_8010# 0.197f
C4443 X1.X2.X2.X1.X1.X2.vout a_23512_8828# 0.36f
C4444 a_49002_10916# X2.X2.X1.X2.X3.vin2 0.263f
C4445 a_54606_21264# X2.X2.X2.X2.X1.X1.X3.vin1 0.00207f
C4446 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.X3.vin1 0.587f
C4447 X1.X2.X2.X1.X2.X1.X1.vin2 X1.X2.X2.X1.X2.X1.X1.vin1 0.668f
C4448 X1.X1.X1.X2.X2.X2.vout a_4396_5198# 0.36f
C4449 X1.X2.X1.X2.X1.X1.vout X1.X2.X1.X2.X3.vin1 0.131f
C4450 X2.X2.X1.X2.X1.X2.X3.vin2 a_46502_9916# 8.07e-19
C4451 a_5082_7064# a_4782_5198# 5.55e-20
C4452 X2.X1.X2.X1.X2.X2.X1.vin2 a_39966_15546# 0.273f
C4453 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X2.vrefh 0.1f
C4454 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.vrefh 2.33e-19
C4455 a_16836_30882# a_16836_28976# 0.00396f
C4456 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.vout 0.0898f
C4457 a_38152_31700# a_37466_29834# 3.31e-19
C4458 a_4782_9010# a_5082_7064# 4.19e-20
C4459 X1.X1.X1.X2.X2.X1.vout a_4696_7064# 0.169f
C4460 X1.X1.X1.X1.X1.X2.X3.vin2 X1.X1.X1.X1.X2.vrefh 0.161f
C4461 X2.X1.X2.X1.X2.X1.X2.vin1 a_39966_11734# 8.88e-20
C4462 X2.X1.X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X1.vin2 8.93e-19
C4463 X1.X2.X1.X1.X2.X2.vrefh a_16836_23258# 0.118f
C4464 a_37466_14586# a_37852_14586# 0.419f
C4465 X2.X2.X3.vin2 a_52106_10734# 6.66e-19
C4466 a_4696_26164# a_4782_24258# 3.21e-19
C4467 a_49002_22312# a_48702_20446# 5.55e-20
C4468 a_19336_22312# a_19722_22312# 0.419f
C4469 a_5082_26164# a_4396_24258# 2.97e-19
C4470 X2.X2.X1.X1.X2.X2.vout a_48316_20446# 0.36f
C4471 X2.X1.X1.X1.X2.vrefh a_31476_25164# 1.64e-19
C4472 X2.X2.X1.X1.X2.X2.X3.vin2 a_46502_17540# 8.07e-19
C4473 X1.X1.X2.X1.X2.X1.X1.vin1 a_11072_11734# 0.195f
C4474 X2.X2.X1.X2.X2.X1.X1.vin2 a_46116_8010# 1.78e-19
C4475 X1.X2.X2.X2.X1.X2.vrefh a_25326_21264# 0.3f
C4476 X2.X2.X2.X2.X1.X2.X3.vin1 a_52106_22210# 0.00874f
C4477 a_23126_31700# a_23212_29834# 3.38e-19
C4478 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X2.X1.X1.X1.X2.X2.vin1 0.00232f
C4479 a_39966_15546# X2.X1.X2.X1.X2.X1.X3.vin2 8.07e-19
C4480 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X1.vout 0.131f
C4481 a_2582_8010# a_2582_6104# 0.00198f
C4482 a_2196_8010# X1.X1.X1.X2.X2.X2.X1.vin1 1.64e-19
C4483 X2.X2.X1.X2.X2.X1.X3.vin1 a_48702_9010# 0.428f
C4484 X2.X1.X2.X1.X1.X2.X1.vin2 a_39966_7922# 0.273f
C4485 a_37466_22210# a_38152_20264# 2.86e-19
C4486 X1.X2.X2.X1.X2.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin1 0.00437f
C4487 a_4396_12822# a_2582_11822# 1.15e-20
C4488 a_10686_32700# a_11072_32700# 0.419f
C4489 a_48316_12822# a_46502_11822# 1.15e-20
C4490 X2.X2.X2.X2.X1.X1.X3.vin1 a_52106_18358# 0.00837f
C4491 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.vrefh 0.161f
C4492 a_54606_21264# a_54992_21264# 0.419f
C4493 a_48616_26164# X2.X2.X1.X1.X2.X1.vout 1.64e-19
C4494 a_49002_26164# a_48702_24258# 5.25e-20
C4495 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X1.X3.vin2 5.19e-19
C4496 a_2196_32788# X1.X1.X1.X1.X1.X1.X3.vin1 0.354f
C4497 a_2582_32788# X1.X1.X1.X1.X1.X1.X1.vin1 0.42f
C4498 X2.X1.X2.X1.X1.X2.X2.vin1 a_40352_9828# 0.197f
C4499 X2.X2.X1.X1.X2.X1.X3.vin2 a_46116_23258# 0.354f
C4500 a_17222_13728# a_19036_12822# 1.06e-19
C4501 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X2.vin1 0.0689f
C4502 a_46116_21352# X2.X2.X1.X1.X2.X2.X3.vin1 0.354f
C4503 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X1.X3.vin2 0.0523f
C4504 a_46502_21352# X2.X2.X1.X1.X2.X2.X1.vin1 0.417f
C4505 a_33976_14688# a_33676_12822# 6.71e-19
C4506 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X1.X2.X3.vin2 3.94e-19
C4507 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin1 0.52f
C4508 X1.X1.X2.X2.X2.X1.X1.vin1 a_10686_25076# 8.22e-20
C4509 a_17222_28976# X1.X2.X1.X1.X1.X2.X1.vin2 0.273f
C4510 X2.X2.X3.vin1 a_52106_6962# 6.45e-19
C4511 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X1.vin2 0.216f
C4512 a_39966_17452# a_38152_16452# 1.15e-20
C4513 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 0.139f
C4514 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X3.vin2 0.234f
C4515 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X2.vrefh 0.00118f
C4516 X1.X1.X2.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X3.vin1 0.581f
C4517 X2.X2.X2.X1.X2.X2.X3.vin1 a_54992_15546# 0.354f
C4518 X1.X2.X1.X3.vin1 a_19722_18540# 0.389f
C4519 a_46116_28976# a_46116_27070# 0.00396f
C4520 X2.X1.X1.X2.X1.X1.vout a_34362_14688# 0.387f
C4521 a_34062_16634# X2.X1.X1.X2.X3.vin1 1.52e-19
C4522 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X3.vin1 0.00117f
C4523 X1.X1.X2.X1.X1.X1.X3.vin2 a_8486_5016# 0.267f
C4524 X2.X1.X1.X2.X1.X2.X3.vin2 a_31862_11822# 0.567f
C4525 X2.X1.X1.X2.X2.X2.X1.vin2 a_31476_4198# 1.78e-19
C4526 a_54606_28888# a_52406_27888# 4.77e-21
C4527 a_5646_892# X1.X3.vin1 0.354f
C4528 a_48316_16634# a_46502_15634# 1.15e-20
C4529 X2.X1.X2.X1.X1.X1.X3.vin2 a_38152_5016# 0.1f
C4530 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X2.vrefh 0.076f
C4531 X1.X1.X2.X2.X1.X1.vout X1.X1.X2.X2.X1.X1.X3.vin1 0.118f
C4532 X1.X2.X2.X2.X2.X1.vout X1.X2.X2.X2.X2.X1.X3.vin2 0.326f
C4533 a_2196_30882# a_2582_30882# 0.419f
C4534 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X1.vin2 0.076f
C4535 a_17222_17540# a_17222_15634# 0.00198f
C4536 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X3.vin1 2.33e-19
C4537 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 1.22e-19
C4538 a_31862_6104# a_34062_5198# 4.2e-20
C4539 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X1.X3.vin2 0.0943f
C4540 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X1.X2.X2.X2.X2.vin1 0.00117f
C4541 a_39966_25076# X2.X1.X2.X2.X1.X2.X2.vin1 0.402f
C4542 a_54606_23170# X2.X2.X2.X2.X1.X1.X3.vin2 8.07e-19
C4543 X2.X2.X2.X1.X3.vin2 a_52492_10734# 0.0927f
C4544 X1.X1.X1.X1.X2.X1.X3.vin2 a_4696_22312# 0.00546f
C4545 X2.X1.X1.X2.X1.X2.vout X2.X1.X1.X2.X1.X2.X3.vin1 0.326f
C4546 X2.X1.X2.X2.X1.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin1 0.00437f
C4547 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.X1.X3.vin1 1.22e-19
C4548 a_54606_17452# X2.X2.X2.X1.X2.X2.X2.vin1 0.402f
C4549 X2.X2.X2.X1.X2.X2.vrefh a_54992_13640# 0.118f
C4550 X2.X2.X2.X2.vrefh a_54606_17452# 0.3f
C4551 X2.X2.X1.X1.X1.X2.vout a_48616_26164# 7.93e-20
C4552 X1.X2.X2.X2.X2.X1.X3.vin2 X1.X2.X2.X2.X2.X1.X1.vin2 8.93e-19
C4553 X1.X2.X2.X2.X2.X1.X2.vin1 a_25326_26982# 8.88e-20
C4554 a_8572_25982# X1.X1.X2.X2.X1.X2.vout 7.93e-20
C4555 X2.X2.X2.X1.X1.X2.X3.vin1 a_54992_7922# 0.354f
C4556 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 0.0565f
C4557 X1.X1.X2.X2.X2.X1.X3.vin1 a_8872_27888# 0.199f
C4558 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.vout 0.335f
C4559 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.vout 0.118f
C4560 a_48316_9010# a_46502_8010# 1.15e-20
C4561 X2.X1.X1.X2.X2.X1.vout X2.X1.X1.X2.X2.X2.vout 0.514f
C4562 a_4696_10916# X1.X1.X1.X2.X3.vin2 0.0927f
C4563 X2.X2.X1.X2.X1.X2.vrefh a_46502_13728# 8.22e-20
C4564 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X3.vin2 8.93e-19
C4565 a_4396_16634# a_5082_14688# 2.86e-19
C4566 a_4782_16634# a_4696_14688# 3.14e-19
C4567 a_19336_18540# a_19036_16634# 6.2e-19
C4568 X1.X2.X2.X1.X1.X1.vout a_23126_5016# 0.422f
C4569 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X1.X3.vin2 1.22e-19
C4570 X1.X1.X2.X1.X1.X2.X3.vin2 a_8186_6962# 3.85e-19
C4571 a_48616_14688# a_48702_12822# 3.38e-19
C4572 X2.X1.X3.vin1 X2.X1.X2.X1.X3.vin1 0.00304f
C4573 a_49002_14688# a_48316_12822# 3.31e-19
C4574 a_22826_14586# X1.X2.X2.X1.X3.vin2 0.423f
C4575 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X2.vin1 0.242f
C4576 a_8186_18358# a_8872_16452# 3.08e-19
C4577 X1.X1.X2.vrefh a_11072_4110# 9.79e-19
C4578 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X3.vin2 8.93e-19
C4579 X1.X1.X2.X3.vin2 a_8186_22210# 0.00292f
C4580 a_52406_12640# a_52792_12640# 0.419f
C4581 X2.X2.X1.X2.X1.X1.vout a_48616_14688# 0.169f
C4582 a_48702_16634# a_49002_14688# 4.19e-20
C4583 X2.X2.vrefh X2.X1.X2.X2.X2.X2.X1.vin2 0.0763f
C4584 X1.X1.X1.X1.X2.X1.X3.vin2 a_2582_23258# 0.567f
C4585 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.vout 0.326f
C4586 a_19336_26164# X1.X2.X1.X1.X3.vin2 0.0927f
C4587 a_28096_892# a_28482_892# 0.419f
C4588 X2.X2.X1.X1.X2.X1.X2.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 0.234f
C4589 a_25326_9828# X1.X2.X2.X1.X1.X2.X2.vin1 0.402f
C4590 X1.X2.X1.X1.X1.X1.vout X1.X2.X1.X1.X1.X1.X3.vin2 0.342f
C4591 X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.vout 3.38e-19
C4592 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin1 0.267f
C4593 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X3.vin1 2.33e-19
C4594 a_10686_13640# a_8872_12640# 1.15e-20
C4595 X2.X1.X2.X1.X2.X1.X2.vin1 a_40352_13640# 0.197f
C4596 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin2 7.84e-19
C4597 X1.X1.X3.vin2 a_5082_14688# 2.04e-19
C4598 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin1 0.195f
C4599 a_2582_13728# X1.X1.X1.X2.X1.X2.X2.vin1 8.88e-20
C4600 a_22826_14586# a_23126_12640# 4.19e-20
C4601 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin1 0.52f
C4602 a_5082_10916# a_4396_9010# 2.97e-19
C4603 a_4696_10916# a_4782_9010# 3.21e-19
C4604 X1.X2.X1.X1.X2.X1.vout a_19722_22312# 0.383f
C4605 a_25326_19358# a_23212_18358# 5.36e-21
C4606 a_2196_6104# X1.X1.X1.X2.X2.X2.X2.vin1 1.78e-19
C4607 a_4782_16634# a_2582_15634# 4.77e-21
C4608 a_37766_24076# a_39966_23170# 4.2e-20
C4609 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X2.vout 0.0898f
C4610 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 0.242f
C4611 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 0.216f
C4612 a_37852_22210# a_39966_21264# 2.95e-20
C4613 a_54606_21264# a_54606_19358# 0.00198f
C4614 a_19336_18540# a_19722_18540# 0.413f
C4615 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X1.X1.vin2 0.076f
C4616 a_33676_12822# a_34062_12822# 0.419f
C4617 X2.X1.X1.X2.X1.X2.X2.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 0.234f
C4618 a_23212_25982# a_23512_24076# 6.48e-19
C4619 X1.X1.X3.vin2 a_5082_7064# 5.84e-19
C4620 X2.X2.X2.vrefh X2.X2.X2.X1.X1.X1.X1.vin1 0.142f
C4621 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X2.vout 0.398f
C4622 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.X2.vin1 0.00117f
C4623 a_17222_17540# a_19422_16634# 4.2e-20
C4624 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X1.vin2 0.076f
C4625 X1.X1.X1.X2.X1.X2.vout a_4396_12822# 0.36f
C4626 a_39966_11734# X2.X1.X2.X1.X1.X2.X3.vin2 8.07e-19
C4627 X1.X1.X2.X2.X2.X1.X3.vin1 a_10686_26982# 0.52f
C4628 X2.X2.X2.X2.X1.X1.X1.vin1 a_54992_17452# 1.64e-19
C4629 a_11072_32700# a_11072_30794# 0.00396f
C4630 a_39966_32700# X2.X1.X2.X2.X2.X2.X2.vin1 0.402f
C4631 X2.X2.X1.X1.X2.X1.X1.vin2 a_46502_23258# 8.88e-20
C4632 X2.X2.X2.X2.X2.X1.X3.vin1 a_54606_26982# 0.52f
C4633 X1.X1.X2.X1.X2.X2.vout a_8572_14586# 0.0929f
C4634 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X3.vin1 0.00789f
C4635 a_8186_29834# a_8572_29834# 0.419f
C4636 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 0.0903f
C4637 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X2.vin1 0.564f
C4638 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.vout 0.118f
C4639 a_37852_29834# a_37766_27888# 3.14e-19
C4640 a_2582_6104# a_2582_4198# 0.00198f
C4641 X2.X2.X1.X3.vin2 a_49002_10916# 0.452f
C4642 a_52792_27888# a_52106_25982# 2.97e-19
C4643 X2.X1.X1.X1.X3.vin1 a_33976_26164# 0.169f
C4644 X2.X1.X2.vrefh a_39966_4110# 4.89e-19
C4645 X2.X2.X2.X2.X3.vin1 a_52492_25982# 0.17f
C4646 a_25326_32700# X1.X2.X2.X2.X2.X2.X3.vin2 0.567f
C4647 a_39966_19358# X2.X1.X2.X1.X2.X2.X3.vin2 8.07e-19
C4648 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 0.139f
C4649 X2.X2.X1.X1.X1.X1.X3.vin1 a_46502_30882# 0.00207f
C4650 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin2 0.1f
C4651 a_8572_25982# a_10686_25076# 4.72e-20
C4652 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.vout 0.2f
C4653 X2.X2.X2.X2.X1.X2.X1.vin2 X2.X2.X2.X2.X1.X2.X1.vin1 0.668f
C4654 a_25326_30794# X1.X2.X2.X2.X2.X2.X1.vin1 0.417f
C4655 X1.X2.X2.X2.X2.X2.X1.vin2 a_25712_30794# 0.12f
C4656 X2.X1.X2.X1.X1.X2.X2.vin1 a_40352_7922# 1.78e-19
C4657 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.X1.vin1 2.23e-19
C4658 X2.X1.X2.X2.X2.X1.X3.vin1 a_40352_26982# 0.354f
C4659 a_48616_7064# X2.X2.X1.X2.X2.X2.X3.vin1 0.00329f
C4660 X1.X1.X1.X2.X2.X2.X3.vin2 a_2582_4198# 0.567f
C4661 a_33676_12822# a_33976_10916# 6.48e-19
C4662 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X3.vin2 0.546f
C4663 a_8186_14586# X1.X1.X2.X1.X2.X1.vout 0.383f
C4664 X1.X2.X1.X1.X1.X2.vout X1.X2.X1.X1.X1.X2.X3.vin2 0.075f
C4665 a_31476_25164# X2.X1.X1.X1.X2.X1.X2.vin1 1.78e-19
C4666 X2.X1.X2.X1.X2.X1.vout a_37766_12640# 0.422f
C4667 a_52106_18358# X2.X2.X3.vin2 0.451f
C4668 a_46116_30882# a_46116_28976# 0.00396f
C4669 X1.X2.X2.vrefh X1.X2.X2.X1.X1.X1.X1.vin1 0.142f
C4670 a_46502_6104# a_46502_4198# 0.00198f
C4671 a_19336_18540# X1.X2.X1.X2.X1.X1.X3.vin1 0.00232f
C4672 a_54606_6016# X2.X2.X2.X1.X1.X1.X3.vin1 0.00207f
C4673 a_10686_13640# a_10686_11734# 0.00198f
C4674 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 0.242f
C4675 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.vrefh 0.00118f
C4676 a_52492_18358# a_52406_16452# 3.3e-19
C4677 a_4396_24258# X1.X1.X1.X1.X2.X1.vout 0.359f
C4678 a_37466_6962# a_37852_6962# 0.419f
C4679 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X2.X1.X1.X2.X1.X2.vin1 0.00232f
C4680 a_33976_29936# X2.X1.X1.X1.X1.X2.X3.vin1 0.00329f
C4681 X1.X2.X1.X2.X1.X1.X3.vin2 a_17222_13728# 8.07e-19
C4682 a_4696_26164# X1.X1.X1.X3.vin1 0.356f
C4683 a_19422_28070# a_19722_26164# 4.41e-20
C4684 X1.X2.X1.X1.X1.X2.X3.vin2 a_19336_26164# 0.00535f
C4685 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X1.X2.X2.X1.vin2 0.216f
C4686 X2.X1.X1.X2.X3.vin2 a_34062_9010# 0.00101f
C4687 a_25326_13640# X1.X2.X2.X1.X2.X1.X2.vin1 0.402f
C4688 X2.X1.X1.X1.X1.X1.X3.vin2 a_31862_28976# 8.07e-19
C4689 a_49002_7064# a_48702_5198# 5.55e-20
C4690 X2.X2.X1.X2.X2.X2.vout a_48316_5198# 0.36f
C4691 X1.X2.X2.X1.X2.X2.X3.vin2 a_23126_16452# 0.277f
C4692 a_19722_10916# X1.X2.X1.X2.X2.X1.X3.vin1 0.00837f
C4693 a_23512_16452# a_23212_14586# 6.71e-19
C4694 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X3.vin1 0.00117f
C4695 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X3.vin1 0.0174f
C4696 a_8486_31700# X1.X1.X2.X2.X2.X2.vout 0.418f
C4697 X1.X2.X2.X1.X1.X1.X3.vin2 X1.X2.X2.X1.X1.X1.X1.vin2 8.93e-19
C4698 X1.X2.X2.X1.X1.X1.X2.vin1 a_25326_4110# 8.88e-20
C4699 a_52106_22210# X2.X2.X2.X2.X1.X1.vout 0.387f
C4700 a_48316_5198# a_46502_4198# 1.15e-20
C4701 X1.X1.X2.X1.X1.X2.vout a_8186_6962# 0.254f
C4702 X2.X2.X1.X2.X1.X2.X3.vin1 a_48702_12822# 0.42f
C4703 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 2.23e-19
C4704 a_48616_26164# X2.X2.X1.X1.X2.X1.X3.vin1 0.00251f
C4705 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.vout 0.08f
C4706 X1.X1.X2.X2.X1.X2.X3.vin2 a_11072_25076# 0.354f
C4707 X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.vout 1.71e-19
C4708 X2.X2.X1.X1.X2.vrefh a_46116_27070# 0.118f
C4709 a_22826_22210# a_23212_22210# 0.419f
C4710 a_46116_19446# X2.X2.X1.X2.X1.X1.X1.vin1 1.64e-19
C4711 a_46502_19446# a_46502_17540# 0.00198f
C4712 X1.X2.X1.X2.X2.X1.X3.vin2 X1.X2.X1.X2.X2.X2.X3.vin1 1.22e-19
C4713 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X1.X3.vin1 0.0131f
C4714 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X3.vin1 0.206f
C4715 a_34062_31882# a_31862_30882# 4.77e-21
C4716 X1.X2.X2.X1.X2.X2.X3.vin2 a_25712_17452# 0.354f
C4717 X1.X2.X3.vin1 X1.X3.vin2 0.12f
C4718 a_52492_18358# X2.X2.X2.X1.X2.X2.X3.vin2 0.00517f
C4719 X2.X2.X2.X1.X2.X1.vout X2.X2.X2.X1.X2.X1.X3.vin1 0.118f
C4720 X2.X2.X3.vin2 X2.X2.X2.X1.X3.vin2 0.039f
C4721 a_54606_28888# a_54992_28888# 0.419f
C4722 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X1.X2.X2.X2.X1.vin2 0.22f
C4723 X1.X1.X1.X1.X1.X2.vrefh a_2196_28976# 1.64e-19
C4724 a_11072_23170# X1.X1.X2.X2.X1.X2.vrefh 1.64e-19
C4725 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X3.vin1 0.206f
C4726 X2.X2.X1.X1.X2.X1.vout a_48616_22312# 0.169f
C4727 a_33676_5198# a_31862_4198# 1.15e-20
C4728 a_48702_24258# a_49002_22312# 4.19e-20
C4729 a_46116_28976# X2.X2.X1.X1.X1.X2.X3.vin1 0.354f
C4730 a_16836_32788# a_17222_32788# 0.419f
C4731 a_46502_28976# X2.X2.X1.X1.X1.X2.X1.vin1 0.417f
C4732 a_46502_17540# a_46502_15634# 0.00198f
C4733 a_16836_15634# a_17222_15634# 0.419f
C4734 a_4396_20446# a_4782_20446# 0.419f
C4735 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X3.vin2 0.449f
C4736 X1.X1.X1.X1.X2.X2.X2.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 0.234f
C4737 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X1.X3.vin2 0.0943f
C4738 X2.X1.X1.X1.X2.vrefh a_31862_27070# 0.3f
C4739 a_38152_27888# a_39966_26982# 1.06e-19
C4740 a_40352_9828# X2.X1.X2.X1.X1.X2.X1.vin2 1.78e-19
C4741 X2.X2.X1.X1.X1.X1.X3.vin1 a_48316_31882# 0.199f
C4742 X2.X2.X3.vin2 a_49566_892# 0.0912f
C4743 a_48702_20446# a_49002_18540# 4.41e-20
C4744 X2.X2.X1.X1.X2.X2.X3.vin2 a_48616_18540# 0.00504f
C4745 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.X1.X1.vin1 5.19e-19
C4746 X2.X3.vin1 a_43362_892# 0.413f
C4747 a_11072_21264# a_11072_19358# 0.00396f
C4748 X1.X1.X1.X1.X3.vin2 a_5082_22312# 0.423f
C4749 X1.X2.X1.X1.X2.X2.vout a_19336_18540# 7.93e-20
C4750 X2.X1.X1.X1.X1.X2.X3.vin2 a_34362_26164# 0.00846f
C4751 a_34062_28070# X2.X1.X1.X3.vin1 1.64e-19
C4752 a_2582_30882# a_4696_29936# 2.95e-20
C4753 a_25326_19358# a_25326_17452# 0.00198f
C4754 a_52406_24076# X2.X2.X2.X2.X1.X2.vout 0.418f
C4755 X1.X2.X2.X2.X1.X1.vout X1.X2.X2.X2.X1.X1.X3.vin1 0.118f
C4756 X1.X2.X2.X3.vin2 a_23212_18358# 0.0927f
C4757 a_25326_25076# a_23512_24076# 1.15e-20
C4758 X1.X2.X1.X2.X2.X2.X3.vin2 a_16836_4198# 0.354f
C4759 a_19422_5198# a_17222_4198# 4.77e-21
C4760 a_37466_18358# X2.X1.X2.X3.vin1 0.374f
C4761 X2.X1.X1.X3.vin2 X2.X1.X3.vin2 3.82e-19
C4762 X1.X1.X1.X2.X2.X2.vrefh a_2196_8010# 0.118f
C4763 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X3.vin1 2.33e-19
C4764 X2.X1.X2.X2.X3.vin1 a_37766_24076# 9.54e-19
C4765 X1.X2.X1.X2.X2.X2.X3.vin2 X1.X2.X2.vrefh 0.172f
C4766 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.X3.vin1 0.0174f
C4767 X2.X2.X2.X2.X2.X2.X1.vin2 X2.X2.X2.X2.X2.X2.vrefh 0.1f
C4768 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X1.X2.X1.X2.X2.X1.vin1 0.668f
C4769 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 0.581f
C4770 X2.X2.X2.X1.X2.X1.X3.vin2 a_52106_10734# 3.49e-19
C4771 X2.X1.X1.X2.X2.vrefh X1.X2.X2.X1.X2.vrefh 0.117f
C4772 a_4696_29936# a_4396_28070# 6.71e-19
C4773 a_31862_32788# a_33676_31882# 1.06e-19
C4774 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X2.vin1 0.0689f
C4775 a_16836_8010# a_17222_8010# 0.419f
C4776 X1.X1.X2.X1.X2.X2.X1.vin1 a_11072_13640# 1.64e-19
C4777 X2.X1.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X3.vin1 2.33e-19
C4778 X1.X1.X2.X2.X1.X1.X2.vin1 a_11072_21264# 0.197f
C4779 a_2582_25164# a_2582_23258# 0.00198f
C4780 X1.X2.X1.X1.X1.X1.X1.vin2 a_16836_30882# 1.78e-19
C4781 a_10686_26982# X1.X1.X2.X2.X2.vrefh 8.22e-20
C4782 X1.X1.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X1.X3.vin2 0.0533f
C4783 a_8486_27888# a_8572_25982# 3.21e-19
C4784 a_8872_24076# a_8186_22210# 3.31e-19
C4785 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin1 0.52f
C4786 X2.X1.X1.X1.X1.X2.X1.vin2 a_31862_27070# 8.88e-20
C4787 X1.X2.X2.X2.X2.X2.X1.vin1 a_25712_28888# 1.64e-19
C4788 X2.X1.X2.X2.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin1 0.00437f
C4789 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.vout 0.118f
C4790 X2.X1.X1.X1.X1.X2.X3.vin1 a_34062_28070# 0.42f
C4791 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X2.X3.vin2 2.23e-19
C4792 X1.X1.X2.X2.X2.X2.vrefh X1.X2.X1.X1.X1.X2.X1.vin2 0.0128f
C4793 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.X1.vin2 8.93e-19
C4794 X1.X1.X2.X1.X2.X2.X2.vin1 a_10686_15546# 8.88e-20
C4795 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X1.X2.X1.X1.X2.X1.vin1 0.668f
C4796 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X2.vin1 0.242f
C4797 X1.X1.X2.X1.X3.vin1 a_8572_10734# 0.169f
C4798 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.vout 0.075f
C4799 X2.X1.X1.X2.X2.vrefh a_31476_9916# 1.64e-19
C4800 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X2.X1.X2.X2.vrefh 0.00437f
C4801 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin2 0.12f
C4802 X2.X1.X1.X2.X1.X1.vout X2.X1.X1.X2.X1.X1.X3.vin2 0.342f
C4803 X1.X2.X1.X1.X2.X1.X3.vin2 a_16836_23258# 0.354f
C4804 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X3.vin2 0.102f
C4805 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin1 0.267f
C4806 a_4696_14688# a_2582_13728# 2.68e-20
C4807 a_33976_14688# a_34362_14688# 0.419f
C4808 X1.X2.X2.X2.X2.X2.X1.vin2 X1.X2.X2.X2.X2.X2.vrefh 0.1f
C4809 a_33676_31882# X2.X1.X1.X1.X1.X1.vout 0.359f
C4810 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin2 0.12f
C4811 X1.X2.X1.X1.X2.X2.X1.vin2 a_16836_19446# 1.78e-19
C4812 X1.X2.vrefh X1.X2.X1.X1.X1.X1.X1.vin2 0.109f
C4813 a_37766_5016# a_38152_5016# 0.419f
C4814 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X3.vin1 0.00789f
C4815 a_10686_17452# X1.X1.X2.X1.X2.X2.X3.vin2 0.567f
C4816 X1.X2.X2.X1.X1.X1.X2.vin1 a_25712_6016# 0.197f
C4817 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X3.vin1 0.00118f
C4818 a_37766_12640# a_37852_10734# 3.21e-19
C4819 X2.X2.X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X2.X3.vin1 0.587f
C4820 X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.vout 3.2e-19
C4821 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X3.vin2 0.418f
C4822 X1.X2.X2.X1.X2.X2.X3.vin1 a_25712_15546# 0.354f
C4823 a_52106_25982# a_52406_24076# 4.41e-20
C4824 a_34362_22312# a_33676_20446# 3.31e-19
C4825 a_33976_22312# a_34062_20446# 3.38e-19
C4826 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin1 0.52f
C4827 a_19036_16634# a_17222_15634# 1.15e-20
C4828 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X2.vin1 0.0689f
C4829 a_40352_11734# X2.X1.X2.X1.X2.vrefh 1.64e-19
C4830 a_46502_17540# a_48316_16634# 1.06e-19
C4831 a_22826_18358# X1.X2.X2.X1.X2.X2.X3.vin2 0.00846f
C4832 a_31476_9916# a_31476_8010# 0.00396f
C4833 a_5082_14688# X1.X1.X1.X2.X1.X2.vout 0.254f
C4834 X1.X1.X2.X1.X2.X1.X1.vin1 a_10686_9828# 8.22e-20
C4835 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X1.X2.X1.X1.X2.X3.vin2 3.94e-19
C4836 X2.X1.X1.X1.X1.X2.X2.vin1 X2.X1.X1.X1.X2.vrefh 0.564f
C4837 a_37766_27888# X2.X1.X2.X2.X2.X1.X3.vin1 0.428f
C4838 X2.X1.X1.X2.X2.X1.vout X2.X1.X1.X2.X2.X1.X3.vin2 0.326f
C4839 X2.X1.X2.X1.X2.X1.X1.vin2 a_39966_11734# 0.273f
C4840 a_37466_29834# X2.X1.X2.X2.X2.X1.X3.vin2 0.00815f
C4841 X2.X1.X2.X2.X2.X2.X2.vin1 a_37766_31700# 0.00351f
C4842 X1.X2.X2.X1.X1.X1.X3.vin1 a_23512_5016# 0.199f
C4843 a_39966_32700# X2.X1.X2.X2.X2.X2.X3.vin1 0.00207f
C4844 X2.X1.X2.X1.X2.X2.X3.vin1 a_37466_14586# 0.00874f
C4845 X1.X1.X1.X1.X1.X2.X3.vin2 a_2582_25164# 8.07e-19
C4846 X1.X2.X2.X2.X1.X2.vout X1.X2.X2.X2.X1.X1.vout 0.507f
C4847 a_34362_7064# X2.X1.X1.X2.X2.X2.vout 0.263f
C4848 a_4696_7064# X1.X1.X1.X2.X2.X2.X3.vin1 0.00329f
C4849 a_2582_11822# a_4696_10916# 4.72e-20
C4850 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X1.vin2 0.076f
C4851 X1.X1.X2.X3.vin2 X1.X1.X3.vin2 0.171f
C4852 X1.X2.X1.X3.vin2 X1.X2.X2.X3.vin1 1.22e-19
C4853 X1.X2.X3.vin1 X1.X2.X3.vin2 3.25f
C4854 a_19722_14688# a_19036_12822# 3.31e-19
C4855 a_19036_28070# a_17222_27070# 1.15e-20
C4856 X1.X2.X2.X1.X1.X2.X3.vin1 a_25712_7922# 0.354f
C4857 a_19336_14688# a_19422_12822# 3.38e-19
C4858 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 2.23e-19
C4859 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 0.049f
C4860 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.vrefh 0.161f
C4861 a_23212_10734# X1.X2.X2.X1.X1.X2.X3.vin2 0.00535f
C4862 a_19036_9010# a_17222_8010# 1.15e-20
C4863 a_52792_8828# a_52492_6962# 6.71e-19
C4864 a_2196_15634# X1.X1.X1.X2.X1.X2.X1.vin1 1.64e-19
C4865 a_2582_15634# a_2582_13728# 0.00198f
C4866 a_34362_22312# X2.X1.X1.X1.X2.X2.X3.vin1 0.00874f
C4867 X2.X2.X2.X2.X1.X1.X3.vin2 X2.X2.X2.X2.X1.X1.X3.vin1 0.581f
C4868 a_37852_14586# a_39966_13640# 2.95e-20
C4869 a_25326_11734# a_25712_11734# 0.419f
C4870 a_23212_10734# a_23512_8828# 6.48e-19
C4871 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X3.vin1 1.22e-19
C4872 a_39966_15546# X2.X1.X2.X1.X2.X2.X1.vin1 0.417f
C4873 X1.X1.X1.X2.X2.X2.vout X1.X1.X1.X2.X2.X2.X3.vin2 0.08f
C4874 X2.X1.X2.X1.X2.X2.X1.vin2 a_40352_15546# 0.12f
C4875 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.vrefh 0.267f
C4876 X1.X2.X1.X1.X1.X1.X1.vin2 a_19036_31882# 0.00113f
C4877 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X2.X2.vin1 0.242f
C4878 a_17222_30882# a_17222_28976# 0.00198f
C4879 a_52106_25982# X2.X2.X2.X2.X1.X2.X3.vin2 0.00846f
C4880 a_16836_30882# X1.X2.X1.X1.X1.X2.X1.vin1 1.64e-19
C4881 X1.X2.X1.X2.X3.vin2 X1.X2.X2.X1.X3.vin1 0.0604f
C4882 X1.X1.X1.X2.X2.X1.vout X1.X1.X1.X2.X2.X2.vout 0.514f
C4883 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin2 0.1f
C4884 X2.X1.X2.X1.X1.X2.X3.vin1 a_37852_6962# 0.00329f
C4885 X2.X1.X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X1.vin1 2.23e-19
C4886 X2.X1.X2.X1.X2.X1.X2.vin1 a_40352_11734# 1.78e-19
C4887 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.vrefh 0.00118f
C4888 X1.X2.X2.vrefh a_14082_892# 2.22e-19
C4889 X1.X1.X1.X3.vin1 a_4782_24258# 5.28e-19
C4890 X2.X2.X1.X1.X2.X2.vout X2.X2.X1.X1.X2.X2.X3.vin2 0.08f
C4891 a_19722_22312# X1.X2.X1.X1.X2.X2.vout 0.263f
C4892 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin1 0.267f
C4893 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.X1.X1.X3.vin1 1.22e-19
C4894 X1.X2.X1.X2.X3.vin1 a_19722_10916# 0.372f
C4895 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X2.X1.X2.X1.X2.X2.vin1 0.00232f
C4896 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X3.vin2 0.161f
C4897 X1.X1.X2.vrefh X1.X2.X2.vrefh 0.0959f
C4898 X2.X2.X3.vin2 a_49002_14688# 2.04e-19
C4899 a_19036_24258# X1.X2.X1.X1.X2.X1.X3.vin2 0.1f
C4900 a_39966_7922# X2.X1.X2.X1.X1.X2.X1.vin1 0.417f
C4901 X2.X1.X2.X1.X1.X2.X1.vin2 a_40352_7922# 0.12f
C4902 X2.X2.X1.X1.X2.X2.X2.vin1 X2.X2.X1.X2.vrefh 0.564f
C4903 X1.X1.X1.X2.X1.X2.X3.vin2 a_2582_11822# 0.567f
C4904 a_19036_31882# a_19336_29936# 6.1e-19
C4905 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X2.vrefh 0.597f
C4906 X1.X1.X2.X2.X2.X2.X3.vin2 a_11072_32700# 0.354f
C4907 X2.X2.X1.X2.X1.X2.X3.vin2 a_46502_11822# 0.567f
C4908 X1.X2.X2.X2.vrefh a_25326_17452# 0.3f
C4909 a_54606_17452# X2.X2.X2.X1.X2.X2.X3.vin1 0.00207f
C4910 X1.X2.X1.X2.X1.X2.X1.vin2 a_16836_11822# 1.78e-19
C4911 a_2196_17540# a_2582_17540# 0.419f
C4912 a_52406_16452# a_52106_14586# 5.55e-20
C4913 X2.X2.X2.X2.X1.X1.X3.vin2 a_54992_21264# 0.354f
C4914 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.vout 0.038f
C4915 X2.X2.X2.X2.X2.X2.vrefh a_54606_28888# 0.3f
C4916 a_10686_6016# X1.X1.X2.X1.X1.X1.X2.vin1 0.402f
C4917 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X3.vin1 0.206f
C4918 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin2 7.84e-19
C4919 X1.X2.X1.X2.X1.X2.X3.vin1 a_19036_12822# 0.199f
C4920 a_8872_31700# a_8186_29834# 3.31e-19
C4921 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X3.vin1 0.206f
C4922 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.vout 0.038f
C4923 a_34362_14688# a_34062_12822# 5.55e-20
C4924 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X1.X2.X3.vin2 5.19e-19
C4925 X1.X2.X1.X1.X1.X2.X3.vin1 X1.X2.X1.X1.X1.X2.X1.vin2 0.216f
C4926 a_23126_31700# a_23512_31700# 0.419f
C4927 a_19036_16634# a_19422_16634# 0.419f
C4928 a_8486_24076# X1.X1.X2.X2.X1.X2.X3.vin1 0.42f
C4929 X1.X1.X1.X1.X2.X1.X2.vin1 X1.X1.X1.X1.X2.X2.vrefh 0.564f
C4930 a_31862_9916# X2.X1.X1.X2.X2.X1.X2.vin1 8.88e-20
C4931 X2.X2.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 0.0565f
C4932 X2.X1.X2.X1.X2.X2.X3.vin2 a_38152_16452# 0.101f
C4933 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X2.vrefh 0.076f
C4934 X1.X1.X2.X2.X2.X1.vout a_8486_27888# 0.422f
C4935 a_34362_18540# X2.X1.X1.X3.vin2 0.233f
C4936 a_48616_10916# a_46502_9916# 5.36e-21
C4937 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.X1.vin1 5.19e-19
C4938 a_46502_28976# a_46502_27070# 0.00198f
C4939 a_23512_27888# a_22826_25982# 2.97e-19
C4940 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X3.vin1 0.00118f
C4941 a_23126_24076# a_23212_22210# 3.38e-19
C4942 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X1.X3.vin1 0.00117f
C4943 X2.X2.X1.X1.X1.X2.X3.vin1 X2.X2.X1.X1.X2.vrefh 0.00118f
C4944 X2.X2.X2.X2.X2.X1.X3.vin2 a_52406_27888# 0.267f
C4945 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.vout 0.398f
C4946 a_52106_29834# a_52492_29834# 0.419f
C4947 X1.X2.X1.X2.X1.X1.X3.vin1 a_17222_15634# 0.00207f
C4948 a_46502_25164# X2.X2.X1.X1.X2.X1.X1.vin2 0.273f
C4949 X2.X2.X2.X2.X2.X2.vout X2.X2.X2.X2.X3.vin2 0.0866f
C4950 X1.X1.X3.vin2 a_6032_892# 0.268f
C4951 X1.X2.X2.X2.X2.X1.X3.vin1 a_23512_27888# 0.199f
C4952 a_4696_22312# a_4396_20446# 6.71e-19
C4953 X2.X1.X1.X2.X2.X2.X3.vin1 a_34062_5198# 0.42f
C4954 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 2.23e-19
C4955 a_11072_9828# a_11072_7922# 0.00396f
C4956 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 0.234f
C4957 a_54606_26982# a_54606_25076# 0.00198f
C4958 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.vout 0.08f
C4959 a_54606_21264# a_52792_20264# 1.15e-20
C4960 X1.X1.X3.vin1 X1.X1.X2.X3.vin1 3.45e-19
C4961 X1.X2.X1.X1.X3.vin2 a_19422_24258# 0.00101f
C4962 a_19722_26164# X1.X2.X1.X1.X2.X1.X3.vin2 3.49e-19
C4963 a_4782_31882# X1.X1.X1.X1.X1.X1.X3.vin2 0.267f
C4964 a_19036_9010# a_19422_9010# 0.419f
C4965 a_46502_21352# X2.X2.X1.X1.X2.X2.X2.vin1 8.88e-20
C4966 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 0.234f
C4967 X2.X2.vrefh X2.X2.X1.X1.X1.X1.X1.vin1 0.108f
C4968 X2.X2.X2.X1.X2.X2.X3.vin2 a_52106_14586# 3.85e-19
C4969 X1.X1.X2.X1.X2.X1.X3.vin2 a_8186_10734# 3.49e-19
C4970 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X3.vin2 0.161f
C4971 a_25326_7922# a_25326_6016# 0.00198f
C4972 X2.X1.X2.X2.X2.X2.X3.vin1 a_37852_29834# 0.00329f
C4973 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X1.X3.vin2 0.546f
C4974 X1.X2.X2.X2.X2.X1.X2.vin1 a_25712_26982# 1.78e-19
C4975 a_52106_14586# X2.X2.X2.X1.X2.X1.vout 0.383f
C4976 X1.X2.X2.X2.X2.X1.X3.vin2 X1.X2.X2.X2.X2.X1.X1.vin1 2.23e-19
C4977 X1.X2.X2.X2.X1.X2.X1.vin2 a_25326_23170# 0.273f
C4978 a_40352_13640# X2.X1.X2.X1.X2.X1.X1.vin2 1.78e-19
C4979 a_39966_21264# X2.X1.X2.X2.X1.X1.X3.vin1 0.00207f
C4980 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X1.vin2 0.076f
C4981 a_13696_892# X1.X3.vin2 0.0927f
C4982 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X3.vin1 2.33e-19
C4983 a_4396_28070# a_4782_28070# 0.419f
C4984 X1.X1.X1.X1.X1.X2.X2.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 0.234f
C4985 a_19336_18540# X1.X2.X1.X2.X1.X1.vout 1.64e-19
C4986 a_19722_18540# a_19422_16634# 5.25e-20
C4987 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X3.vin1 0.00118f
C4988 X1.X1.X3.vin1 a_4782_12822# 2.12e-19
C4989 a_4782_16634# X1.X1.X1.X2.X3.vin1 1.52e-19
C4990 X1.X1.X1.X2.X1.X1.vout a_5082_14688# 0.387f
C4991 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X1.vout 0.131f
C4992 a_4696_29936# a_5082_29936# 0.419f
C4993 X1.X1.X2.X2.X1.X1.X3.vin1 a_10686_19358# 0.52f
C4994 X2.X2.X2.X2.X1.X2.vout a_52106_22210# 0.254f
C4995 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.vrefh 2.33e-19
C4996 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X1.X3.vin1 0.0425f
C4997 X2.X2.X1.X2.X3.vin1 a_48702_12822# 9.54e-19
C4998 a_49002_14688# X2.X2.X1.X2.X1.X2.X3.vin2 3.85e-19
C4999 a_48616_26164# X2.X2.X1.X3.vin1 0.356f
C5000 a_23126_8828# a_22826_6962# 5.55e-20
C5001 X1.X1.X1.X2.X1.X2.vout a_4696_10916# 7.93e-20
C5002 X1.X1.X1.X1.X1.X2.X1.vin2 a_2196_27070# 1.78e-19
C5003 X2.X1.X1.X2.X3.vin2 a_33976_7064# 0.363f
C5004 a_46502_19446# a_48616_18540# 4.72e-20
C5005 a_52792_20264# a_52106_18358# 2.97e-19
C5006 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.vout 0.197f
C5007 X2.X1.X3.vin1 a_37466_14586# 2.24e-19
C5008 X2.X1.X1.X1.X2.X2.X3.vin2 a_31862_17540# 8.07e-19
C5009 X2.X2.X2.X2.X2.X2.X1.vin1 a_54992_28888# 1.64e-19
C5010 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin2 0.12f
C5011 X2.X2.X1.X2.X1.X1.vout X2.X2.X1.X2.X3.vin1 0.131f
C5012 a_40352_32700# a_40352_30794# 0.00396f
C5013 X2.X1.X2.X2.X2.X2.vrefh X2.X2.X1.X1.X1.X2.X1.vin2 0.0128f
C5014 a_39966_9828# a_37766_8828# 4.77e-21
C5015 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 0.242f
C5016 a_39966_17452# a_39966_15546# 0.00198f
C5017 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin2 0.12f
C5018 a_31862_9916# X2.X1.X1.X2.X2.X1.X1.vin2 0.273f
C5019 a_28482_892# vout 0.399f
C5020 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X3.vin2 0.418f
C5021 X1.X1.X1.X2.X3.vin2 a_4782_5198# 9.7e-20
C5022 a_39966_21264# X2.X1.X2.X2.X1.X1.X3.vin2 0.567f
C5023 a_10686_21264# a_8486_20264# 4.77e-21
C5024 a_48702_24258# X2.X2.X1.X1.X2.X1.X3.vin2 0.267f
C5025 X1.X1.X2.X2.X2.X1.X2.vin1 a_11072_28888# 0.197f
C5026 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 0.234f
C5027 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X1.vin2 0.076f
C5028 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X2.vrefh 0.076f
C5029 X1.X1.X2.X1.X2.X1.X3.vin2 a_8872_12640# 0.1f
C5030 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.vrefh 2.33e-19
C5031 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 0.581f
C5032 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X3.vin1 0.00118f
C5033 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin1 0.52f
C5034 X1.X2.X2.X1.X2.X1.vout X1.X2.X2.X1.X2.X1.X3.vin1 0.118f
C5035 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X2.vin1 0.00117f
C5036 X1.X1.X1.X2.X3.vin2 a_4782_9010# 0.00101f
C5037 a_2582_13728# a_4782_12822# 4.2e-20
C5038 a_37852_10734# a_37766_8828# 3.3e-19
C5039 a_40352_7922# a_40352_6016# 0.00396f
C5040 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X2.vin1 0.0689f
C5041 a_2582_6104# a_4396_5198# 1.06e-19
C5042 X1.X1.X2.X2.X1.X1.vout a_8872_20264# 0.359f
C5043 a_46116_28976# X2.X2.X1.X1.X1.X2.X2.vin1 1.78e-19
C5044 X2.X2.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X3.vin2 0.0533f
C5045 a_37852_22210# X2.X1.X2.X2.X1.X1.X3.vin2 0.00546f
C5046 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X1.vin1 0.206f
C5047 X2.X2.X2.X2.X1.X1.X3.vin2 a_54606_19358# 7.84e-19
C5048 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X1.vin1 0.0689f
C5049 a_19722_18540# X1.X2.X3.vin1 0.47f
C5050 a_52406_31700# a_52492_29834# 3.38e-19
C5051 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X2.vin1 0.242f
C5052 a_39966_15546# X2.X1.X2.X1.X2.X2.vrefh 8.22e-20
C5053 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X1.vin2 0.1f
C5054 a_34062_12822# X2.X1.X1.X2.X1.X2.X3.vin2 0.277f
C5055 X2.X2.X2.X2.X2.X2.X3.vin1 a_52792_31700# 0.199f
C5056 a_48316_16634# X2.X2.X1.X2.X1.X1.vout 0.359f
C5057 X2.X1.X1.X1.X2.X1.X2.vin1 a_31862_23258# 0.402f
C5058 X2.X2.X2.X1.X1.X1.X1.vin2 a_54606_4110# 0.273f
C5059 a_37466_29834# X2.X1.X2.X2.X3.vin2 0.422f
C5060 X1.X2.X1.X2.X1.X1.X3.vin1 a_19422_16634# 0.428f
C5061 a_33976_18540# a_34062_16634# 3.21e-19
C5062 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin1 0.195f
C5063 a_34362_18540# a_33676_16634# 2.97e-19
C5064 X1.X1.X1.X2.X1.X2.vout X1.X1.X1.X2.X1.X2.X3.vin2 0.075f
C5065 X1.X2.X1.X2.X1.X1.X3.vin2 a_19722_14688# 0.00815f
C5066 a_4396_5198# X1.X1.X1.X2.X2.X2.X3.vin2 0.101f
C5067 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.X1.X1.vin2 3.94e-19
C5068 X1.X1.X2.X2.X2.X1.X3.vin1 a_11072_26982# 0.354f
C5069 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 0.216f
C5070 a_23126_12640# a_25326_11734# 4.2e-20
C5071 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin1 0.195f
C5072 X2.X2.X2.X2.X2.X1.X3.vin1 a_54992_26982# 0.354f
C5073 a_25712_28888# X1.X2.X2.X2.X2.X1.X1.vin2 1.78e-19
C5074 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X3.vin2 0.237f
C5075 a_54606_6016# X2.X2.X2.X1.X1.X1.X3.vin2 0.567f
C5076 X1.X1.X1.X2.X2.X2.X3.vin1 a_2582_4198# 0.00207f
C5077 a_52406_12640# a_52106_10734# 5.25e-20
C5078 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X3.vin1 0.199f
C5079 a_31476_13728# a_31476_11822# 0.00396f
C5080 a_22826_6962# a_23512_5016# 2.86e-19
C5081 a_39966_7922# X2.X1.X2.X1.X1.X2.vrefh 8.22e-20
C5082 X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin1 0.00304f
C5083 X2.X1.X2.vrefh a_40352_4110# 9.79e-19
C5084 a_39966_13640# X2.X1.X2.X1.X2.X1.X3.vin1 0.00207f
C5085 X2.X1.X1.X1.X1.X1.X2.vin1 X2.X1.X1.X1.X1.X2.vrefh 0.564f
C5086 a_6032_892# X1.X3.vin1 0.461f
C5087 a_48316_9010# X2.X2.X1.X2.X2.X1.vout 0.359f
C5088 a_37766_31700# X2.X1.X2.X2.X2.X2.X3.vin1 0.42f
C5089 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.vout 0.326f
C5090 a_4396_9010# X1.X1.X1.X2.X2.X1.vout 0.359f
C5091 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin2 7.84e-19
C5092 X1.X2.X2.X3.vin2 a_22826_22210# 0.00292f
C5093 a_8572_25982# X1.X1.X2.X2.X1.X2.X3.vin2 0.00535f
C5094 a_54606_23170# a_54992_23170# 0.419f
C5095 X2.X2.X1.X2.X2.X2.vout X2.X2.X1.X2.X2.X2.X3.vin1 0.335f
C5096 X1.X2.X2.X2.X2.X2.X1.vin1 a_25712_30794# 0.195f
C5097 X1.X1.X2.X2.X3.vin2 a_8186_25982# 0.263f
C5098 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X1.vin1 5.19e-19
C5099 X2.X1.X1.X2.X1.X2.X3.vin2 a_33976_10916# 0.00535f
C5100 a_34062_12822# a_34362_10916# 4.41e-20
C5101 a_37766_27888# X2.X1.X2.X3.vin2 7.93e-20
C5102 a_37466_6962# X2.X1.X2.X1.X1.X1.X3.vin2 0.00815f
C5103 a_31862_25164# a_33676_24258# 1.06e-19
C5104 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X2.vin1 0.0689f
C5105 X1.X2.X2.X1.X1.X1.X1.vin2 a_25326_4110# 0.273f
C5106 X2.X2.X1.X2.X2.X2.X3.vin1 a_46502_4198# 0.00207f
C5107 a_46116_30882# X2.X2.X1.X1.X1.X2.X1.vin1 1.64e-19
C5108 a_46502_30882# a_46502_28976# 0.00198f
C5109 X2.X2.X2.X1.X1.X1.X3.vin2 X2.X2.X2.X1.X1.X1.X3.vin1 0.581f
C5110 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X3.vin1 0.449f
C5111 X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.vout 3.08e-19
C5112 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X1.vin1 0.0689f
C5113 X1.X1.X2.X1.X2.X1.X3.vin2 a_10686_11734# 7.84e-19
C5114 a_2196_27070# a_2196_25164# 0.00396f
C5115 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin2 0.1f
C5116 a_31476_21352# a_31862_21352# 0.419f
C5117 X1.X1.X1.X2.X2.X1.X3.vin2 a_2196_8010# 0.354f
C5118 X1.X2.X2.X2.X1.X1.X2.vin1 X2.X1.X1.X1.X2.X2.X1.vin2 0.00232f
C5119 a_25326_9828# X1.X2.X2.X1.X1.X2.X1.vin2 8.88e-20
C5120 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X2.X3.vin1 0.0174f
C5121 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin1 0.195f
C5122 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X3.vin1 1.22e-19
C5123 a_48616_18540# a_48316_16634# 6.2e-19
C5124 X2.X1.X1.X2.X1.X1.X3.vin2 a_33976_14688# 0.00546f
C5125 a_31862_13728# X2.X1.X1.X2.X1.X2.X1.vin2 0.273f
C5126 X1.X2.X3.vin2 a_19722_7064# 5.84e-19
C5127 a_8572_22210# a_8486_20264# 3.14e-19
C5128 X1.X1.X2.X2.X2.X2.X3.vin2 a_8186_29834# 3.85e-19
C5129 X1.X1.X2.X1.X1.X1.X1.vin2 X1.X1.X2.X1.X1.X1.X1.vin1 0.668f
C5130 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.X1.vin2 0.22f
C5131 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 0.234f
C5132 a_52406_31700# a_54606_30794# 4.2e-20
C5133 X2.X1.X1.X1.X2.X2.vrefh X1.X2.X2.X2.X1.X2.vrefh 0.117f
C5134 X2.X2.X1.X2.X2.X2.vout X2.X2.X1.X2.X2.X2.X3.vin2 0.08f
C5135 a_31862_8010# X2.X1.X1.X2.X2.X2.X1.vin1 8.22e-20
C5136 X2.X1.X1.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X1.X2.X3.vin1 1.22e-19
C5137 a_37852_18358# X2.X1.X2.X1.X2.X2.vout 7.93e-20
C5138 X1.X2.X2.X1.X1.X1.X3.vin2 X1.X2.X2.X1.X1.X1.X1.vin1 2.23e-19
C5139 X1.X2.X2.X1.X1.X1.X2.vin1 a_25712_4110# 1.78e-19
C5140 X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin1 0.00437f
C5141 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X2.vin1 0.242f
C5142 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 0.0565f
C5143 a_54606_13640# X2.X2.X2.X1.X2.X1.X1.vin2 8.88e-20
C5144 X2.X2.X1.X2.X2.X2.X3.vin2 a_46502_4198# 0.567f
C5145 a_4696_10916# a_2582_9916# 5.36e-21
C5146 a_33976_10916# a_34362_10916# 0.414f
C5147 X1.X1.X1.X1.X2.vrefh a_2582_27070# 0.3f
C5148 a_22826_29834# X1.X2.X2.X2.X2.X1.vout 0.383f
C5149 a_8872_27888# a_10686_26982# 1.06e-19
C5150 a_46116_27070# a_46502_27070# 0.419f
C5151 a_39966_21264# X2.X1.X2.X2.X1.X1.X1.vin2 8.88e-20
C5152 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X3.vin1 0.0131f
C5153 a_52792_27888# a_54606_26982# 1.06e-19
C5154 a_49002_14688# X2.X2.X1.X2.X1.X2.vout 0.254f
C5155 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X2.vrefh 2.33e-19
C5156 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 2.23e-19
C5157 a_37766_16452# a_38152_16452# 0.419f
C5158 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin1 0.195f
C5159 a_16836_28976# a_16836_27070# 0.00396f
C5160 X2.X1.X1.X2.X2.X1.X3.vin2 a_34362_7064# 0.00815f
C5161 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X2.X1.X2.X2.X2.X1.vin2 0.00232f
C5162 a_25326_28888# X1.X2.X2.X2.X2.X1.X3.vin1 0.00207f
C5163 a_46116_6104# a_46502_6104# 0.419f
C5164 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X1.X2.X2.X2.X1.X3.vin2 3.94e-19
C5165 X1.X2.X2.X2.X2.vrefh a_25326_25076# 0.3f
C5166 X1.X1.X2.X2.X2.X2.X1.vin1 a_10686_28888# 8.22e-20
C5167 a_25326_32700# a_25712_32700# 0.419f
C5168 X2.X2.X2.X2.X2.X1.X3.vin2 a_54992_28888# 0.354f
C5169 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X2.X1.vin1 0.267f
C5170 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X2.vout 0.2f
C5171 a_17222_8010# a_19336_7064# 2.95e-20
C5172 X2.X1.X1.X2.X2.X2.X3.vin2 a_31862_4198# 0.567f
C5173 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X1.vin1 5.19e-19
C5174 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X2.X3.vin1 0.0131f
C5175 X2.X2.X1.X1.X2.X1.vout X2.X2.X1.X1.X2.X2.vout 0.514f
C5176 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X2.X3.vin1 0.206f
C5177 a_16836_32788# X1.X2.X1.X1.X1.X1.X3.vin1 0.354f
C5178 a_17222_32788# X1.X2.X1.X1.X1.X1.X1.vin1 0.42f
C5179 X2.X2.X1.X1.X1.X1.X1.vin2 a_46502_30882# 8.88e-20
C5180 X2.X2.X1.X2.X1.X1.X3.vin1 a_46502_15634# 0.00207f
C5181 X2.X2.X2.X3.vin2 X2.X2.X3.vin2 0.171f
C5182 a_4782_20446# X1.X1.X1.X1.X2.X2.X3.vin2 0.277f
C5183 a_52492_25982# a_52792_24076# 6.48e-19
C5184 a_39966_25076# X2.X1.X2.X2.X1.X2.X3.vin1 0.00207f
C5185 X2.X2.X1.X1.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X1.vout 0.118f
C5186 a_37466_14586# a_38152_12640# 2.86e-19
C5187 X1.X1.X2.X3.vin1 a_8186_10734# 0.509f
C5188 a_25326_19358# X1.X2.X2.X1.X2.X2.X3.vin2 8.07e-19
C5189 a_37766_8828# a_38152_8828# 0.419f
C5190 X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin2 0.00254f
C5191 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X2.vrefh 0.1f
C5192 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X1.vin2 0.076f
C5193 a_2582_9916# X1.X1.X1.X2.X2.X1.X2.vin1 8.88e-20
C5194 a_54606_7922# a_54606_6016# 0.00198f
C5195 a_54606_6016# a_52792_5016# 1.15e-20
C5196 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X2.vrefh 0.076f
C5197 X1.X2.X2.X2.X1.X2.X3.vin2 a_23512_24076# 0.101f
C5198 a_46502_6104# X2.X2.X1.X2.X2.X2.X2.vin1 8.88e-20
C5199 X1.X1.X1.X2.X1.X2.X3.vin2 a_2582_9916# 8.07e-19
C5200 a_19336_22312# a_19036_20446# 6.71e-19
C5201 a_10686_23170# a_10686_21264# 0.00198f
C5202 a_10686_15546# a_11072_15546# 0.419f
C5203 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X2.vrefh 0.267f
C5204 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.vrefh 2.33e-19
C5205 X2.X2.X1.X2.X1.X2.vrefh a_46502_15634# 0.3f
C5206 a_5082_29936# a_4782_28070# 5.55e-20
C5207 X1.X1.X1.X1.X2.X2.vrefh a_2582_21352# 8.22e-20
C5208 X1.X1.X3.vin1 X1.X1.X1.X2.X3.vin1 7.18e-19
C5209 X2.X1.X1.X1.X1.X1.X3.vin1 a_33676_31882# 0.199f
C5210 X2.X2.X2.vrefh a_49566_892# 7.23e-19
C5211 X1.X2.X1.X1.X2.X1.X3.vin2 a_19336_22312# 0.00546f
C5212 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X1.X3.vin1 0.00836f
C5213 a_25326_15546# a_23212_14586# 2.68e-20
C5214 X1.X1.X1.X1.X2.X1.X3.vin1 a_2582_23258# 0.00207f
C5215 X1.X1.X2.X2.X2.X2.X3.vin1 a_10686_30794# 0.52f
C5216 a_11072_26982# X1.X1.X2.X2.X2.vrefh 1.64e-19
C5217 X1.X1.X1.X3.vin1 a_4696_18540# 0.17f
C5218 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin1 0.195f
C5219 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X2.vout 0.398f
C5220 a_25712_6016# X1.X2.X2.X1.X1.X1.X1.vin2 1.78e-19
C5221 a_23126_20264# a_22826_18358# 5.25e-20
C5222 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X2.vout 0.0857f
C5223 a_52492_29834# a_52792_27888# 6.1e-19
C5224 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.X1.X1.vin1 0.668f
C5225 X1.X1.X2.X1.X2.X2.X2.vin1 a_11072_15546# 1.78e-19
C5226 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.X1.vin1 2.23e-19
C5227 X2.X2.X2.X1.X1.X1.X3.vin1 a_52792_5016# 0.199f
C5228 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 0.049f
C5229 X1.X1.X2.X1.X1.X2.X3.vin1 a_8572_6962# 0.00329f
C5230 a_10686_7922# a_11072_7922# 0.419f
C5231 a_40352_26982# a_40352_25076# 0.00396f
C5232 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X3.vin1 0.00118f
C5233 X2.X2.X1.X2.X2.X2.vrefh a_46502_8010# 0.3f
C5234 X1.X1.X2.X2.X3.vin1 a_8486_24076# 9.54e-19
C5235 X1.X1.X1.X1.X1.X1.X1.vin2 a_2196_30882# 1.78e-19
C5236 X1.X2.X1.X2.X2.X1.X3.vin2 X1.X2.X1.X2.X2.X2.X1.vin2 3.94e-19
C5237 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X1.vin2 0.668f
C5238 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin1 0.267f
C5239 X2.X2.X1.X1.X1.X2.X2.vin1 X2.X2.X1.X1.X2.vrefh 0.564f
C5240 X1.X1.X1.X1.X3.vin1 X1.X1.X2.X2.X3.vin2 0.0604f
C5241 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 2.23e-19
C5242 X2.X2.X2.X1.X2.X1.vout a_52792_12640# 0.359f
C5243 X1.X2.X2.X2.X2.X2.X1.vin1 X1.X2.X2.X2.X2.X2.vrefh 0.267f
C5244 a_4696_14688# X1.X1.X1.X2.X1.X2.X3.vin1 0.00329f
C5245 a_34362_14688# X2.X1.X1.X2.X3.vin1 0.436f
C5246 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X1.vin2 0.668f
C5247 a_54606_9828# a_52792_8828# 1.15e-20
C5248 X1.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X3.vin1 0.546f
C5249 X1.X1.X2.X1.X2.X1.vout a_8572_10734# 1.64e-19
C5250 X2.X2.X2.X1.X2.X1.X1.vin2 X2.X2.X2.X1.X2.X1.X1.vin1 0.668f
C5251 X2.X1.X2.X1.X3.vin1 a_37852_6962# 0.363f
C5252 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin2 0.12f
C5253 X2.X2.X1.X1.X3.vin2 a_48702_20446# 9.7e-20
C5254 a_25712_23170# a_25712_21264# 0.00396f
C5255 X1.X2.X1.X1.X3.vin2 a_19722_22312# 0.423f
C5256 X2.X1.X1.X1.X2.X2.vout a_33976_18540# 7.93e-20
C5257 a_10686_28888# a_8486_27888# 4.77e-21
C5258 a_52792_16452# a_52492_14586# 6.71e-19
C5259 a_19422_9010# a_19336_7064# 3.14e-19
C5260 a_19036_9010# a_19722_7064# 2.86e-19
C5261 a_39966_28888# X2.X1.X2.X2.X2.X1.X3.vin2 0.567f
C5262 a_34362_22312# X2.X1.X1.X1.X2.X2.X3.vin2 3.85e-19
C5263 X2.X1.X1.X1.X2.X2.vout a_34062_20446# 0.418f
C5264 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X3.vin1 0.0174f
C5265 X2.X2.X1.X2.X1.X1.X3.vin1 a_48316_16634# 0.199f
C5266 X2.X2.X1.X1.X1.X1.X1.vin2 a_48316_31882# 0.00113f
C5267 X2.X1.X1.X1.X1.X2.X2.vin1 a_31862_27070# 0.402f
C5268 X2.X2.X1.X2.X3.vin2 a_48702_5198# 9.7e-20
C5269 a_2196_23258# a_2582_23258# 0.419f
C5270 a_31862_9916# a_31862_8010# 0.00198f
C5271 a_10686_9828# a_8486_8828# 4.77e-21
C5272 X2.X1.X2.X3.vin2 X2.X1.X2.X3.vin1 0.559f
C5273 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 5.19e-19
C5274 X2.X2.X3.vin1 X2.X2.X2.X3.vin1 3.45e-19
C5275 a_25326_25076# a_25326_23170# 0.00198f
C5276 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 0.242f
C5277 X1.X2.X2.X2.X1.X1.vout a_23512_20264# 0.359f
C5278 X2.X1.X2.X1.X2.X1.X1.vin2 a_40352_11734# 0.12f
C5279 a_39966_11734# X2.X1.X2.X1.X2.X1.X1.vin1 0.417f
C5280 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin2 0.1f
C5281 X2.X1.X2.X2.X1.X1.X3.vin1 a_37852_18358# 0.00255f
C5282 X2.X1.X2.X2.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X2.X3.vin1 0.587f
C5283 X1.X1.X1.X1.X2.X1.X2.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 0.234f
C5284 X1.X1.X1.X1.X1.X2.X3.vin2 X1.X1.X1.X1.X2.X1.X3.vin1 1.22e-19
C5285 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X3.vin2 8.93e-19
C5286 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.vout 0.398f
C5287 X1.X1.X1.X2.X2.X2.vout X1.X1.X1.X2.X2.X2.X3.vin1 0.335f
C5288 a_19036_5198# a_19422_5198# 0.419f
C5289 X1.X2.X1.X2.X2.X2.X2.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 0.234f
C5290 X1.X1.X1.X2.X1.X2.vrefh a_2582_15634# 0.3f
C5291 a_8872_16452# a_10686_15546# 1.06e-19
C5292 X1.X2.X3.vin2 a_23212_18358# 0.355f
C5293 a_10686_19358# a_10686_17452# 0.00198f
C5294 X1.X2.X1.X1.X1.X2.X3.vin2 a_17222_27070# 0.567f
C5295 a_19722_14688# X1.X2.X1.X2.X1.X2.X3.vin2 3.85e-19
C5296 X1.X2.X1.X2.X3.vin1 a_19422_12822# 9.54e-19
C5297 a_52406_16452# X2.X2.X2.X1.X2.X2.X3.vin1 0.42f
C5298 X2.X1.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X1.vin2 0.1f
C5299 a_10686_23170# a_8572_22210# 2.68e-20
C5300 a_48616_29936# a_49002_29936# 0.419f
C5301 a_54606_11734# a_54606_9828# 0.00198f
C5302 a_46502_8010# a_48616_7064# 2.95e-20
C5303 X1.X2.X2.X3.vin2 a_23126_24076# 6.03e-19
C5304 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X1.X3.vin2 1.22e-19
C5305 a_2582_21352# X1.X1.X1.X1.X2.X2.X1.vin2 0.273f
C5306 X1.X2.X2.X1.X2.X2.vout X1.X2.X2.X1.X2.X1.vout 0.514f
C5307 a_54606_32700# X2.X2.X2.X2.X2.X2.X2.vin1 0.402f
C5308 a_37852_14586# X2.X1.X2.X1.X2.X1.X3.vin2 0.00546f
C5309 X1.X2.X2.X2.X1.X1.vout X1.X2.X2.X2.X1.X1.X3.vin2 0.342f
C5310 X2.X1.X2.X1.X2.X2.X1.vin1 a_40352_15546# 0.195f
C5311 a_16836_6104# a_16836_4198# 0.00396f
C5312 a_11072_17452# X1.X1.X2.X1.X2.X2.X1.vin2 1.78e-19
C5313 a_19336_22312# a_17222_21352# 2.68e-20
C5314 X3.vin2 a_42976_892# 0.37f
C5315 a_25326_6016# a_23126_5016# 4.77e-21
C5316 a_31862_30882# a_33976_29936# 2.95e-20
C5317 a_19722_29936# X1.X2.X1.X1.X1.X2.vout 0.254f
C5318 X2.X1.X3.vin2 X2.X1.X1.X2.X2.X1.vout 4.93e-20
C5319 X1.X1.X2.X1.X2.X2.X3.vin1 a_8186_14586# 0.00874f
C5320 a_22826_18358# a_23126_16452# 4.41e-20
C5321 X1.X1.X3.vin2 a_8486_12640# 2.33e-19
C5322 a_31862_27070# X2.X1.X1.X1.X2.X1.X1.vin1 8.22e-20
C5323 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X1.vin2 0.076f
C5324 a_52406_8828# X2.X2.X2.X1.X1.X2.X3.vin1 0.42f
C5325 a_54606_9828# X2.X2.X2.X1.X1.X2.X1.vin2 8.88e-20
C5326 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X1.vin1 5.19e-19
C5327 X1.X1.X1.X2.X2.X1.X2.vin1 X1.X1.X1.X2.X2.X2.vrefh 0.564f
C5328 a_8486_8828# X1.X1.X2.X1.X1.X2.X3.vin1 0.42f
C5329 X2.X2.X2.X1.X3.vin2 a_52406_12640# 0.00101f
C5330 a_40352_25076# a_40352_23170# 0.00396f
C5331 X1.X2.X1.X1.X2.X1.vout X1.X2.X1.X1.X2.X1.X3.vin2 0.326f
C5332 a_48616_18540# a_46502_17540# 5.36e-21
C5333 X2.X1.X2.X1.X1.X2.X1.vin1 a_40352_7922# 0.195f
C5334 a_10686_17452# a_11072_17452# 0.419f
C5335 a_37466_25982# a_37852_25982# 0.414f
C5336 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X3.vin1 0.587f
C5337 X1.X2.X1.X1.X1.X1.vout a_19336_29936# 0.169f
C5338 a_19422_31882# a_19722_29936# 4.19e-20
C5339 X2.X2.X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X2.vout 0.08f
C5340 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X3.vin2 0.161f
C5341 a_17222_6104# X1.X2.X1.X2.X2.X2.X1.vin2 0.273f
C5342 X1.X2.X2.X1.X3.vin1 a_22826_6962# 0.436f
C5343 a_2582_17540# X1.X1.X1.X2.X1.X1.X1.vin1 0.417f
C5344 a_2196_17540# X1.X1.X1.X2.X1.X1.X3.vin1 0.354f
C5345 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X1.X3.vin2 0.161f
C5346 X2.X3.vin2 a_49566_892# 0.51f
C5347 a_17222_23258# X1.X2.X1.X1.X2.X2.X1.vin1 8.22e-20
C5348 a_31476_28976# a_31862_28976# 0.419f
C5349 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X3.vin2 0.234f
C5350 X1.X2.X2.X2.X2.X1.X2.vin1 X2.X1.X1.X1.X1.X2.X1.vin2 0.00232f
C5351 X2.X2.X3.vin1 a_49952_892# 0.386f
C5352 a_37766_27888# a_38152_27888# 0.419f
C5353 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 0.587f
C5354 a_10686_15546# X1.X1.X2.X1.X2.X2.vrefh 8.22e-20
C5355 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 0.0565f
C5356 a_19422_16634# X1.X2.X1.X2.X1.X1.vout 0.422f
C5357 X1.X1.X1.X1.X2.X2.X1.vin2 a_2196_19446# 1.78e-19
C5358 a_25326_15546# a_25326_13640# 0.00198f
C5359 X1.X1.X3.vin1 a_5082_10916# 6.09e-19
C5360 a_31862_9916# a_34062_9010# 4.2e-20
C5361 a_23212_22210# a_23126_20264# 3.14e-19
C5362 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X2.vin1 0.00117f
C5363 X2.X1.X2.X1.X2.X2.vout a_37466_14586# 0.263f
C5364 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X1.X3.vin1 0.0425f
C5365 a_8572_10734# a_8486_8828# 3.3e-19
C5366 a_48616_10916# X2.X2.X1.X2.X2.X1.X3.vin1 0.00251f
C5367 X2.X2.X1.X1.X1.X2.X3.vin1 a_46502_27070# 0.00207f
C5368 a_39966_6016# X2.X1.X2.X1.X1.X1.X1.vin2 8.88e-20
C5369 a_39966_30794# a_39966_28888# 0.00198f
C5370 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X1.vin2 0.216f
C5371 X2.X2.X3.vin1 a_52406_5016# 8.66e-20
C5372 a_46502_30882# a_48616_29936# 2.95e-20
C5373 X1.X2.X1.X1.X1.X2.vout X1.X2.X1.X1.X1.X2.X3.vin1 0.326f
C5374 X1.X2.X1.X3.vin1 a_19422_20446# 5.31e-19
C5375 X1.X1.X1.X1.X2.X2.vout a_4396_20446# 0.36f
C5376 a_5082_22312# a_4782_20446# 5.55e-20
C5377 X1.X1.X2.X3.vin1 a_8572_18358# 0.17f
C5378 a_54606_26982# X2.X2.X2.X2.X1.X2.X3.vin2 8.07e-19
C5379 a_19036_28070# a_19422_28070# 0.419f
C5380 X1.X2.X1.X1.X1.X2.X2.vin1 X1.X2.X1.X1.X1.X2.X3.vin2 0.234f
C5381 X2.X2.X2.X2.X1.X1.X3.vin2 a_52792_20264# 0.1f
C5382 a_23126_16452# X1.X2.X2.X1.X3.vin2 9.7e-20
C5383 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X2.vin1 0.564f
C5384 a_10686_7922# X1.X1.X2.X1.X1.X2.vrefh 8.22e-20
C5385 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X1.vin2 3.94e-19
C5386 a_48316_9010# a_48616_7064# 6.1e-19
C5387 a_19422_9010# X1.X2.X1.X2.X2.X1.vout 0.422f
C5388 a_37466_10734# a_37852_10734# 0.414f
C5389 X2.X1.X2.X2.X1.X2.X3.vin2 a_37466_22210# 3.85e-19
C5390 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 2.23e-19
C5391 a_46502_21352# a_48702_20446# 4.2e-20
C5392 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X1.X2.X2.X2.vin1 0.00117f
C5393 X2.X2.X2.X2.X3.vin2 a_52106_25982# 0.263f
C5394 a_37466_6962# a_37766_5016# 4.19e-20
C5395 a_25326_7922# X1.X2.X2.X1.X1.X1.X3.vin2 8.07e-19
C5396 a_19336_10916# a_19036_9010# 6.2e-19
C5397 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X2.X3.vin2 0.0523f
C5398 a_25326_23170# X1.X2.X2.X2.X1.X2.X1.vin1 0.417f
C5399 X1.X2.X2.X2.X1.X2.X1.vin2 a_25712_23170# 0.12f
C5400 a_2196_17540# a_2196_15634# 0.00396f
C5401 X1.X1.X2.X2.X1.X1.X3.vin1 a_8572_18358# 0.00255f
C5402 X2.X1.X2.X1.X1.X2.vout a_37852_6962# 0.0929f
C5403 X1.X1.X2.X1.X1.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin1 0.00437f
C5404 a_38152_31700# a_39966_30794# 1.06e-19
C5405 X2.X1.X1.X1.X1.X2.vrefh a_31862_30882# 0.3f
C5406 a_46502_11822# a_48616_10916# 4.72e-20
C5407 X2.X1.X1.X2.X3.vin1 a_34362_10916# 0.372f
C5408 a_33676_31882# a_34362_29936# 2.86e-19
C5409 a_34062_31882# a_33976_29936# 3.14e-19
C5410 X2.X1.X2.X2.X1.X1.X3.vin2 X2.X1.X2.X2.X1.X1.X3.vin1 0.581f
C5411 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X2.vrefh 0.076f
C5412 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X2.vrefh 0.00118f
C5413 X3.vin1 X1.X3.vin2 0.246f
C5414 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X1.X3.vin1 0.0321f
C5415 a_4782_28070# X1.X1.X1.X1.X1.X2.X3.vin2 0.277f
C5416 a_8186_14586# X1.X1.X2.X1.X2.X1.X3.vin2 0.00815f
C5417 X1.X2.X3.vin1 X1.X2.X1.X2.X1.X1.vout 2.91e-19
C5418 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.X1.X1.X1.vin2 3.94e-19
C5419 a_5082_29936# X1.X1.X1.X1.X3.vin1 0.434f
C5420 X1.X2.X2.X2.X1.X2.vrefh a_25712_21264# 0.118f
C5421 X1.X1.X2.X2.X1.X1.X3.vin1 a_11072_19358# 0.354f
C5422 a_2582_32788# a_4396_31882# 1.06e-19
C5423 a_19722_7064# a_19036_5198# 3.31e-19
C5424 a_19336_7064# a_19422_5198# 3.38e-19
C5425 a_40352_15546# a_40352_13640# 0.00396f
C5426 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X1.vin2 0.076f
C5427 X2.X1.X1.X1.X1.X1.X2.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 0.234f
C5428 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X2.vout 0.0866f
C5429 X1.X1.X2.X2.X1.X1.X3.vin2 a_8186_18358# 3.49e-19
C5430 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X1.vout 0.0215f
C5431 X2.X2.X1.X1.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X2.vrefh 0.00118f
C5432 X1.X1.X2.X2.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin1 0.00437f
C5433 a_34362_18540# X2.X1.X1.X2.X1.X1.X3.vin1 0.00837f
C5434 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.X1.X1.X3.vin1 1.22e-19
C5435 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X1.vin2 0.696f
C5436 a_48316_12822# X2.X2.X1.X2.X1.X2.X3.vin2 0.101f
C5437 a_22826_25982# X1.X2.X2.X3.vin2 0.452f
C5438 a_34926_892# a_35312_892# 0.419f
C5439 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 0.22f
C5440 a_23126_31700# a_25326_30794# 4.2e-20
C5441 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X1.vin1 0.0689f
C5442 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X1.vin2 0.668f
C5443 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X3.vin1 0.00117f
C5444 X1.X1.X2.X2.X2.X2.X3.vin1 a_8572_29834# 0.00329f
C5445 X1.X1.X2.X2.X2.X1.X1.vin1 a_11072_25076# 1.64e-19
C5446 X2.X1.X2.X1.X2.X2.X3.vin2 a_39966_15546# 7.84e-19
C5447 X2.X1.X2.X1.X1.X2.X3.vin2 a_37766_8828# 0.277f
C5448 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin1 0.195f
C5449 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X1.vin2 0.216f
C5450 a_25326_26982# a_23212_25982# 5.36e-21
C5451 a_49002_29936# X2.X2.X1.X1.X1.X2.X3.vin1 0.00874f
C5452 a_8486_24076# X1.X1.X2.X2.X1.X2.vout 0.418f
C5453 a_2196_11822# a_2196_9916# 0.00396f
C5454 X1.X1.X2.X2.X1.X1.X3.vin2 a_8486_20264# 0.267f
C5455 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X3.vin1 0.00117f
C5456 a_8186_29834# a_8872_27888# 2.86e-19
C5457 X1.X1.X2.X2.vrefh a_10686_17452# 0.3f
C5458 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 0.0903f
C5459 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X1.vout 0.399f
C5460 X1.X1.X1.X2.X1.X2.X3.vin1 a_4782_12822# 0.42f
C5461 a_23512_24076# a_22826_22210# 3.31e-19
C5462 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 2.23e-19
C5463 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X2.vrefh 0.076f
C5464 a_46116_30882# a_46502_30882# 0.419f
C5465 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin2 7.84e-19
C5466 X1.X1.X1.X2.X2.X2.X3.vin1 a_4396_5198# 0.199f
C5467 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X2.X2.vin1 0.0689f
C5468 a_46502_28976# a_48316_28070# 1.06e-19
C5469 a_40352_15546# X2.X1.X2.X1.X2.X2.vrefh 1.64e-19
C5470 X1.X2.X1.X2.X1.X1.X1.vin2 a_17222_15634# 8.88e-20
C5471 X2.X2.X2.X1.X1.X1.X1.vin2 a_54992_4110# 0.12f
C5472 a_54606_4110# X2.X2.X2.X1.X1.X1.X1.vin1 0.417f
C5473 X2.X1.X2.X2.X1.X2.X2.vin1 a_40352_25076# 0.197f
C5474 a_34062_24258# a_31862_23258# 4.77e-21
C5475 X2.X1.X1.X2.X2.X2.vrefh a_31476_6104# 1.64e-19
C5476 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.X1.X1.X1.vin1 5.19e-19
C5477 a_48316_31882# a_48616_29936# 6.1e-19
C5478 a_54992_23170# a_54992_21264# 0.00396f
C5479 a_2582_25164# X1.X1.X1.X1.X2.X1.X2.vin1 8.88e-20
C5480 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin1 0.52f
C5481 X2.X1.X3.vin1 a_34062_16634# 2.92e-19
C5482 a_19422_20446# a_19336_18540# 3.3e-19
C5483 a_19036_20446# a_19722_18540# 3.08e-19
C5484 X2.X2.X2.X1.X2.X2.X2.vin1 a_54992_17452# 0.197f
C5485 a_48616_22312# X2.X2.X1.X1.X2.X2.vout 0.0929f
C5486 X2.X2.X2.X2.vrefh a_54992_17452# 0.118f
C5487 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X2.X1.X1.vin1 0.206f
C5488 X2.X1.X2.X2.X2.X2.vout a_37852_29834# 0.0929f
C5489 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin1 0.52f
C5490 a_54606_25076# a_54606_23170# 0.00198f
C5491 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 0.242f
C5492 X1.X1.X1.X2.X2.X1.X3.vin2 a_5082_7064# 0.00815f
C5493 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X1.vout 0.131f
C5494 X3.vin1 a_28096_892# 0.196f
C5495 X2.X1.X3.vin1 a_34062_9010# 2.12e-19
C5496 a_39966_21264# a_38152_20264# 1.15e-20
C5497 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin2 0.1f
C5498 X2.X1.X2.X1.X3.vin2 a_37852_14586# 0.363f
C5499 a_10686_32700# X1.X1.X2.X2.X2.X2.X3.vin1 0.00207f
C5500 X2.X1.X2.X1.X1.X1.X1.vin2 X2.X1.X2.X1.X1.X1.X1.vin1 0.668f
C5501 X1.X1.X2.X2.X2.X2.X2.vin1 a_8486_31700# 0.00351f
C5502 X1.X2.X2.X1.X2.vrefh a_25326_9828# 0.3f
C5503 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X3.vin1 0.0131f
C5504 a_40352_7922# X2.X1.X2.X1.X1.X2.vrefh 1.64e-19
C5505 a_31862_13728# a_31862_11822# 0.00198f
C5506 a_31862_21352# X2.X1.X1.X1.X2.X2.X2.vin1 8.88e-20
C5507 X1.X2.X1.X2.X1.X2.vout a_19336_10916# 7.93e-20
C5508 X2.X1.X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X3.vin1 0.581f
C5509 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X2.vrefh 0.00118f
C5510 X2.X2.X2.X2.X1.X1.X3.vin1 a_54606_19358# 0.52f
C5511 X2.X2.X2.X2.X1.X2.X3.vin1 a_52492_22210# 0.00329f
C5512 a_8872_20264# a_10686_19358# 1.06e-19
C5513 X1.X1.X1.X2.vrefh a_2582_19446# 0.3f
C5514 X1.X1.X3.vin2 X1.X3.vin1 0.238f
C5515 X1.X1.X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X1.X2.X1.vin1 5.19e-19
C5516 X2.X2.X3.vin1 X2.X2.X1.X2.X3.vin1 7.18e-19
C5517 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 0.581f
C5518 X2.X2.X2.X2.X1.X2.X1.vin2 X2.X2.X2.X2.X1.X2.vrefh 0.1f
C5519 a_37852_22210# a_38152_20264# 6.1e-19
C5520 a_31862_15634# X2.X1.X1.X2.X1.X2.X1.vin1 8.22e-20
C5521 X1.X2.X2.X2.X2.X2.X1.vin2 X2.X1.X1.X1.X1.X1.X2.vin1 0.00232f
C5522 X1.X2.X1.X2.X1.X2.vrefh a_16836_15634# 0.118f
C5523 a_25326_21264# X1.X2.X2.X2.X1.X1.X3.vin1 0.00207f
C5524 X1.X2.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X2.X1.X1.vin2 0.076f
C5525 a_23212_29834# a_23512_27888# 6.1e-19
C5526 a_5082_18540# a_4396_16634# 2.97e-19
C5527 a_4696_18540# a_4782_16634# 3.21e-19
C5528 X2.X2.X1.X3.vin1 a_48616_18540# 0.17f
C5529 a_49002_26164# X2.X2.X1.X1.X2.X1.X3.vin2 3.49e-19
C5530 X2.X2.X1.X1.X3.vin2 a_48702_24258# 0.00101f
C5531 X2.X1.X1.X1.X2.X1.X3.vin1 a_33676_24258# 0.199f
C5532 X1.X2.X2.X1.X1.X1.X1.vin2 a_25712_4110# 0.12f
C5533 a_25326_4110# X1.X2.X2.X1.X1.X1.X1.vin1 0.417f
C5534 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X1.X3.vin2 1.22e-19
C5535 X1.X2.X3.vin2 a_22826_14586# 3.67e-19
C5536 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 0.216f
C5537 a_2196_27070# X1.X1.X1.X1.X2.X1.X1.vin1 1.64e-19
C5538 a_39966_21264# a_40352_21264# 0.419f
C5539 a_2582_27070# a_2582_25164# 0.00198f
C5540 a_37766_20264# a_39966_19358# 4.2e-20
C5541 X1.X2.X2.X1.X1.X2.X2.vin1 a_25712_9828# 0.197f
C5542 a_8186_25982# X1.X1.X2.X2.X3.vin1 0.372f
C5543 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X3.vin2 8.93e-19
C5544 X1.X1.X1.X1.X3.vin2 X1.X1.X2.X3.vin2 7.46e-20
C5545 X1.X2.X2.X1.X1.X2.X2.vin1 a_25326_7922# 8.88e-20
C5546 a_31476_21352# X2.X1.X1.X1.X2.X2.X3.vin1 0.354f
C5547 a_31862_21352# X2.X1.X1.X1.X2.X2.X1.vin1 0.417f
C5548 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X1.vin2 8.93e-19
C5549 a_2196_21352# X1.X1.X1.X1.X2.X2.X2.vin1 1.78e-19
C5550 X1.X2.X1.X1.X2.X2.X3.vin2 a_17222_17540# 8.07e-19
C5551 X1.X2.X1.X3.vin1 X1.X2.X1.X3.vin2 0.552f
C5552 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin1 0.52f
C5553 a_2582_28976# X1.X1.X1.X1.X1.X2.X1.vin2 0.273f
C5554 a_48616_18540# X2.X2.X1.X2.X1.X1.vout 1.64e-19
C5555 X1.X2.X3.vin2 X3.vin1 0.00523f
C5556 a_49002_18540# a_48702_16634# 5.25e-20
C5557 X1.X2.X2.X1.X2.X1.vout a_23512_12640# 0.359f
C5558 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X1.vin2 0.216f
C5559 X2.X1.X1.X2.X1.X1.vout X2.X1.X1.X2.X1.X2.vout 0.507f
C5560 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X2.vin1 0.242f
C5561 X2.X2.X1.X2.X1.X1.X3.vin2 a_46116_15634# 0.354f
C5562 a_37466_10734# a_38152_8828# 3.08e-19
C5563 X1.X1.X1.X1.X2.X1.X3.vin2 a_2582_21352# 8.07e-19
C5564 X1.X2.X1.X1.X2.vrefh X1.X1.X2.X2.X2.vrefh 0.117f
C5565 a_10686_4110# a_11072_4110# 0.419f
C5566 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.X1.vin1 0.206f
C5567 X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.X3.vin2 0.0604f
C5568 X1.X2.X1.X2.X2.X2.vrefh a_16836_8010# 0.118f
C5569 a_19336_7064# a_19722_7064# 0.419f
C5570 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X1.X3.vin2 1.22e-19
C5571 X2.X2.X1.X1.X1.X1.X2.vin1 a_46502_30882# 0.402f
C5572 X2.X2.X2.X2.X2.X2.vout a_52792_31700# 0.36f
C5573 a_10686_25076# a_8486_24076# 4.77e-21
C5574 X2.X2.X2.X1.X1.X2.X3.vin1 a_52106_6962# 0.00874f
C5575 X1.X2.X2.X2.X2.X2.X2.vin1 a_23512_31700# 5.34e-19
C5576 X1.X2.X2.X1.X1.X2.vrefh a_25326_6016# 0.3f
C5577 a_5082_18540# X1.X1.X3.vin2 6.58e-20
C5578 X2.X2.X2.X1.X2.X1.X2.vin1 a_54606_11734# 8.88e-20
C5579 X1.X2.X2.X2.X1.X2.X1.vin2 X1.X2.X2.X2.X1.X2.vrefh 0.1f
C5580 X2.X2.X2.X1.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X1.vin2 8.93e-19
C5581 X1.X1.X1.X2.X2.X1.X1.vin2 a_2196_8010# 1.78e-19
C5582 a_23126_20264# a_25326_19358# 4.2e-20
C5583 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 0.216f
C5584 a_33676_24258# X2.X1.X1.X1.X2.X1.vout 0.359f
C5585 X2.X2.X1.X1.X2.vrefh a_46116_25164# 1.64e-19
C5586 a_46502_23258# X2.X2.X1.X1.X2.X2.X1.vin1 8.22e-20
C5587 X1.X2.X2.X1.X3.vin1 a_23126_8828# 9.54e-19
C5588 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X3.vin1 0.00836f
C5589 a_4696_10916# X1.X1.X1.X2.X2.X1.X3.vin1 0.00251f
C5590 a_34362_10916# X2.X1.X1.X2.X3.vin2 0.263f
C5591 a_25326_25076# X1.X2.X2.X2.X1.X2.X2.vin1 0.402f
C5592 X1.X2.X2.X2.X2.X1.X3.vin2 a_22826_25982# 3.49e-19
C5593 a_40352_11734# a_40352_9828# 0.00396f
C5594 X1.X2.X1.X2.X2.vrefh a_16836_11822# 0.118f
C5595 X2.X1.X2.X2.X1.X1.X2.vin1 a_39966_19358# 8.88e-20
C5596 X2.X1.X2.X2.X1.X1.X3.vin2 X2.X1.X2.X2.X1.X1.X1.vin2 8.93e-19
C5597 a_39966_32700# X2.X2.vrefh 0.3f
C5598 X2.X1.X2.X2.X2.X2.X2.vin1 a_40352_32700# 0.197f
C5599 a_54606_15546# a_54606_13640# 0.00198f
C5600 a_54606_6016# a_54992_6016# 0.419f
C5601 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin1 0.52f
C5602 a_39966_17452# X2.X1.X2.X1.X2.X2.X2.vin1 0.402f
C5603 a_17222_28976# a_17222_27070# 0.00198f
C5604 X2.X2.X1.X2.X2.X1.X3.vin2 a_46116_8010# 0.354f
C5605 X1.X1.X1.X2.X2.X2.X1.vin2 a_2582_4198# 8.88e-20
C5606 a_46502_6104# X2.X2.X1.X2.X2.X2.X1.vin1 0.417f
C5607 a_46116_6104# X2.X2.X1.X2.X2.X2.X3.vin1 0.354f
C5608 X1.X2.X2.X2.X2.X1.X3.vin2 X1.X2.X2.X2.X2.X1.X3.vin1 0.581f
C5609 X1.X2.X1.X1.X1.X2.X3.vin1 X1.X2.X1.X1.X2.vrefh 0.00118f
C5610 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X3.vin2 0.161f
C5611 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X1.X2.X2.X2.X1.X3.vin2 5.19e-19
C5612 X1.X1.X1.X2.X1.X1.X3.vin2 a_4696_14688# 0.00546f
C5613 X2.X1.X2.X3.vin2 a_37466_22210# 0.00292f
C5614 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X2.vrefh 0.1f
C5615 a_39966_13640# a_38152_12640# 1.15e-20
C5616 X1.X2.X2.X2.X2.X2.X3.vin2 a_25712_32700# 0.354f
C5617 X1.X2.X2.X2.X2.X2.X2.vin1 X2.vrefh 0.597f
C5618 a_37766_31700# X2.X1.X2.X2.X2.X2.vout 0.418f
C5619 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 0.049f
C5620 X2.X2.X1.X2.vrefh a_46116_19446# 0.118f
C5621 a_40352_19358# a_40352_17452# 0.00396f
C5622 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X3.vin1 0.206f
C5623 a_4696_22312# a_5082_22312# 0.419f
C5624 X1.X2.X2.X1.X2.X1.vout a_23212_14586# 0.169f
C5625 a_31862_13728# X2.X1.X1.X2.X1.X2.X2.vin1 8.88e-20
C5626 X2.X2.X1.X2.X1.X2.vout a_48316_12822# 0.36f
C5627 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X1.X3.vin2 0.0523f
C5628 X1.X2.X2.X2.X3.vin2 X1.X2.X1.X3.vin1 7.46e-20
C5629 a_25326_26982# a_25326_25076# 0.00198f
C5630 a_8572_18358# X1.X1.X2.X1.X2.X2.vout 7.93e-20
C5631 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 0.139f
C5632 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X3.vin1 0.587f
C5633 X2.X2.X1.X2.X1.X1.X3.vin2 a_49002_14688# 0.00815f
C5634 a_37766_24076# a_37466_22210# 5.55e-20
C5635 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.vrefh 0.267f
C5636 X2.X2.X1.X2.X2.X2.X1.vin2 a_46502_4198# 8.88e-20
C5637 X2.X2.X2.X2.X2.X1.vout X2.X2.X2.X2.X2.X1.X3.vin2 0.326f
C5638 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X2.vin1 0.00117f
C5639 X2.X2.X2.X1.X1.X1.X3.vin2 a_52792_5016# 0.1f
C5640 a_54606_7922# X2.X2.X2.X1.X1.X1.X3.vin2 8.07e-19
C5641 a_2582_9916# a_4782_9010# 4.2e-20
C5642 X2.X1.X1.X1.X1.X1.X1.vin2 a_31476_30882# 1.78e-19
C5643 X1.X2.X2.vrefh a_20672_892# 7.3e-19
C5644 X2.X1.X2.X1.X1.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin1 0.00437f
C5645 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X2.vin1 0.00117f
C5646 a_46502_6104# a_48702_5198# 4.2e-20
C5647 a_10686_23170# X1.X1.X2.X2.X1.X1.X3.vin2 8.07e-19
C5648 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X3.vin1 1.22e-19
C5649 X1.X2.X1.X1.X2.X2.vout a_19036_20446# 0.36f
C5650 a_19722_22312# a_19422_20446# 5.55e-20
C5651 X1.X2.X2.X2.X2.X1.X1.vin2 a_25326_26982# 0.273f
C5652 X2.X1.X3.vin2 a_34362_7064# 5.84e-19
C5653 X1.X1.X2.X3.vin1 a_8186_14586# 7.98e-19
C5654 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X1.vin2 3.94e-19
C5655 X1.X1.X1.X3.vin2 X1.X1.X2.X1.X3.vin2 7.46e-20
C5656 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X3.vin1 2.33e-19
C5657 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.vout 0.118f
C5658 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 0.0565f
C5659 X1.X2.X2.X1.X3.vin2 a_23126_12640# 0.00101f
C5660 X2.X1.X2.X3.vin1 a_37766_12640# 5.28e-19
C5661 a_10686_9828# X1.X1.X2.X1.X1.X2.X2.vin1 0.402f
C5662 X1.X2.X2.X1.X2.X1.X2.vin1 a_25712_13640# 0.197f
C5663 X1.X1.X1.X2.X1.X1.X3.vin2 a_2582_15634# 0.567f
C5664 a_19336_18540# X1.X2.X1.X3.vin2 0.0927f
C5665 X1.X1.X2.X2.X2.X2.X3.vin1 a_11072_30794# 0.354f
C5666 a_25326_32700# X1.X2.X2.X2.X2.X2.X1.vin2 8.88e-20
C5667 X1.X1.X1.X3.vin1 X1.X1.X3.vin1 0.188f
C5668 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin1 0.52f
C5669 X2.X1.X1.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X1.X2.X1.vin2 3.94e-19
C5670 X2.X2.X1.X2.X1.X1.X2.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 0.234f
C5671 a_39966_28888# a_39966_26982# 0.00198f
C5672 X1.X1.X3.vin2 a_8186_6962# 0.00111f
C5673 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X1.X1.vin2 0.242f
C5674 X1.X1.X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X1.X2.vrefh 0.165f
C5675 a_4396_31882# a_2582_30882# 1.15e-20
C5676 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin2 7.84e-19
C5677 a_10686_26982# a_11072_26982# 0.419f
C5678 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 0.216f
C5679 a_37766_16452# a_39966_15546# 4.2e-20
C5680 X1.X2.X1.X1.X1.X2.vrefh a_17222_28976# 8.22e-20
C5681 X2.X2.X1.X2.X2.X2.X2.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 0.234f
C5682 a_48316_5198# a_48702_5198# 0.419f
C5683 a_23212_18358# a_23512_16452# 6.48e-19
C5684 a_31862_11822# X2.X1.X1.X2.X2.X1.X1.vin1 8.22e-20
C5685 X1.X1.X1.X1.X1.X2.X2.vin1 a_2582_27070# 0.402f
C5686 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.vout 0.2f
C5687 X1.X1.X2.X2.X3.vin2 a_8572_29834# 0.363f
C5688 X2.X2.X1.X1.X1.X2.X2.vin1 a_46502_27070# 0.402f
C5689 X2.X2.X2.X2.X1.X1.X1.vin2 X2.X2.X2.X2.X1.X1.X1.vin1 0.668f
C5690 a_25326_28888# a_23512_27888# 1.15e-20
C5691 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X3.vin1 0.0174f
C5692 X2.X2.X1.X2.X2.X1.X2.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 0.234f
C5693 a_23126_24076# a_23512_24076# 0.419f
C5694 a_17222_28976# X1.X2.X1.X1.X1.X2.X2.vin1 8.88e-20
C5695 X2.X2.X2.X1.X1.X2.X3.vin2 a_52792_8828# 0.101f
C5696 X1.X1.X1.X2.X2.X1.X2.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 0.234f
C5697 a_54606_11734# a_54992_11734# 0.419f
C5698 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin2 0.12f
C5699 a_25326_21264# X1.X2.X2.X2.X1.X1.X1.vin2 8.88e-20
C5700 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X2.X1.vin2 0.668f
C5701 a_23126_31700# a_22826_29834# 5.55e-20
C5702 X2.X2.X1.X2.X1.X1.X1.vin2 a_46502_15634# 8.88e-20
C5703 a_31862_19446# X2.X1.X1.X2.X1.X1.X1.vin1 8.22e-20
C5704 a_33676_5198# X2.X1.X1.X2.X2.X2.X3.vin2 0.101f
C5705 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X3.vin1 0.00117f
C5706 X1.X1.X2.X2.X2.X1.X3.vin2 a_8486_27888# 0.267f
C5707 X1.X2.X1.X2.X2.X1.vout a_19722_7064# 0.383f
C5708 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X1.vin2 0.076f
C5709 X1.X2.X3.vin2 X1.X2.X1.X2.X3.vin2 0.00254f
C5710 X1.X2.X2.X3.vin1 a_22826_10734# 0.509f
C5711 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 1.22e-19
C5712 X1.X1.X2.X1.X2.X1.vout X1.X1.X2.X1.X3.vin2 0.399f
C5713 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.vout 0.118f
C5714 a_34062_28070# a_31862_27070# 4.77e-21
C5715 a_37852_6962# a_39966_6016# 2.95e-20
C5716 a_4696_26164# a_2582_25164# 5.36e-21
C5717 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 0.216f
C5718 a_33976_26164# a_34362_26164# 0.414f
C5719 a_37766_8828# a_39966_7922# 4.2e-20
C5720 X2.X1.X1.X1.X1.X2.X3.vin2 a_31476_27070# 0.354f
C5721 X2.X2.X2.X3.vin1 a_52492_18358# 0.17f
C5722 X2.X1.X1.X2.X2.X1.X3.vin1 a_31862_8010# 0.00207f
C5723 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X2.vrefh 2.33e-19
C5724 X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X3.vin1 0.0321f
C5725 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.X3.vin1 0.0131f
C5726 X1.X1.X2.X1.X1.X2.X3.vin2 a_8486_8828# 0.277f
C5727 X1.X2.X1.X1.X2.X2.vrefh a_16836_21352# 1.64e-19
C5728 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X3.vin1 0.00117f
C5729 X1.X2.X2.X2.X1.X2.X3.vin2 a_25326_23170# 7.84e-19
C5730 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X1.vin1 0.0689f
C5731 a_52106_10734# a_52406_8828# 4.41e-20
C5732 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X1.X3.vin2 1.22e-19
C5733 X2.X1.X2.X1.X2.X1.X1.vin1 a_40352_11734# 0.195f
C5734 a_8572_18358# a_10686_17452# 4.72e-20
C5735 X2.X2.X2.X1.X2.X2.X1.vin2 X2.X2.X2.X1.X2.X2.X1.vin1 0.668f
C5736 a_4782_24258# X1.X1.X1.X1.X2.X1.X3.vin2 0.267f
C5737 X1.X3.vin2 a_20286_892# 0.51f
C5738 X2.X1.X1.X1.X1.X1.X1.vin2 a_33676_31882# 0.00113f
C5739 a_5082_26164# X1.X1.X1.X1.X3.vin2 0.241f
C5740 a_19422_5198# X1.X2.X1.X2.X2.X2.X3.vin2 0.277f
C5741 a_31476_17540# X2.X1.X1.X2.X1.X1.X2.vin1 1.78e-19
C5742 a_23212_29834# a_25326_28888# 2.95e-20
C5743 a_10686_19358# X1.X1.X2.X1.X2.X2.X3.vin2 8.07e-19
C5744 X1.X2.X2.X3.vin2 a_23126_20264# 5.21e-19
C5745 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X3.vin2 0.0533f
C5746 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X2.vout 0.0857f
C5747 X1.X1.X1.X1.X2.X1.X1.vin2 a_2582_23258# 8.88e-20
C5748 a_54606_11734# X2.X2.X2.X1.X1.X2.X3.vin2 8.07e-19
C5749 a_49002_29936# X2.X2.X1.X1.X3.vin1 0.434f
C5750 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X2.vrefh 0.00118f
C5751 X1.X1.X1.X2.X2.X2.vrefh a_2196_6104# 1.64e-19
C5752 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X1.X2.X2.X1.vin2 0.216f
C5753 X1.X1.X2.X2.X2.X2.X3.vin1 a_8872_31700# 0.199f
C5754 X2.X2.X2.X2.X2.X2.X2.vin1 X2.X2.X2.X2.X2.X2.X3.vin2 0.237f
C5755 a_4396_16634# X1.X1.X1.X2.X1.X1.vout 0.359f
C5756 a_10686_13640# X1.X1.X2.X1.X2.X1.X2.vin1 0.402f
C5757 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X2.X1.X2.X1.X1.X2.vin1 0.00232f
C5758 X2.X2.X2.X2.X1.X1.vout a_52492_22210# 0.169f
C5759 a_4696_18540# X1.X1.X3.vin1 0.354f
C5760 a_19336_22312# X1.X2.X1.X1.X2.X2.X3.vin1 0.00329f
C5761 a_17222_6104# a_17222_4198# 0.00198f
C5762 X3.vin2 X2.X3.vin2 0.215f
C5763 X2.X1.X3.vin1 a_37766_5016# 8.66e-20
C5764 X1.X2.X2.X1.X1.X1.X3.vin2 a_23126_5016# 0.267f
C5765 X2.X2.X2.X1.X1.X2.X1.vin2 X2.X2.X2.X1.X1.X2.X1.vin1 0.668f
C5766 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X3.vin1 0.00117f
C5767 X1.X1.X2.X1.X1.X2.vout a_8572_6962# 0.0929f
C5768 a_48616_29936# a_48316_28070# 6.71e-19
C5769 X1.X1.X2.X2.X2.X2.vrefh X1.X1.X2.X2.X2.X1.X2.vin1 0.564f
C5770 a_37852_25982# a_39966_25076# 4.72e-20
C5771 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X3.vin1 0.0131f
C5772 X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin1 0.00437f
C5773 X1.X2.X2.X1.X3.vin2 X1.X2.X2.X1.X3.vin1 0.546f
C5774 X1.X2.X2.X1.X2.X1.vout a_23212_10734# 1.64e-19
C5775 X2.X1.X1.X1.X1.X1.X3.vin2 a_31862_30882# 0.567f
C5776 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X1.vin2 8.93e-19
C5777 X2.X2.X2.X1.X1.X2.X2.vin1 a_54606_7922# 8.88e-20
C5778 a_52406_27888# a_52492_25982# 3.21e-19
C5779 X2.X1.X1.X1.X3.vin2 a_34362_22312# 0.423f
C5780 a_2196_30882# a_2196_28976# 0.00396f
C5781 X2.X2.X1.X1.X2.X1.X3.vin2 a_49002_22312# 0.00815f
C5782 X2.X2.X1.X1.X2.X2.vout a_48616_18540# 7.93e-20
C5783 a_48616_18540# X2.X2.X1.X2.X1.X1.X3.vin1 0.00232f
C5784 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X2.X1.X2.X2.X1.X2.vin1 0.00232f
C5785 X1.X2.X1.X1.X3.vin1 a_19722_26164# 0.385f
C5786 X1.X1.X2.X1.X2.X2.X3.vin2 a_11072_17452# 0.354f
C5787 X1.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin1 0.00437f
C5788 a_25326_13640# X1.X2.X2.X1.X2.X1.X1.vin2 8.88e-20
C5789 X1.X2.X1.X1.X1.X1.vout X1.X2.X1.X1.X3.vin1 0.13f
C5790 a_54606_9828# X2.X2.X2.X1.X1.X2.X3.vin2 0.567f
C5791 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X1.vin2 0.22f
C5792 a_39966_28888# a_40352_28888# 0.419f
C5793 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X2.vout 0.398f
C5794 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X3.vin1 0.206f
C5795 a_31862_23258# a_33976_22312# 2.95e-20
C5796 X2.X2.X1.X1.X1.X1.X1.vin1 X2.X2.X1.X1.X1.X1.X3.vin2 2.23e-19
C5797 a_2196_28976# X1.X1.X1.X1.X1.X2.X2.vin1 1.78e-19
C5798 a_31476_28976# X2.X1.X1.X1.X1.X2.X3.vin1 0.354f
C5799 a_31862_28976# X2.X1.X1.X1.X1.X2.X1.vin1 0.417f
C5800 X1.X1.X2.X1.X2.X1.X1.vin1 a_11072_9828# 1.64e-19
C5801 X1.X1.X2.X2.X1.X2.vrefh a_10686_21264# 0.3f
C5802 a_11072_15546# X1.X1.X2.X1.X2.X2.vrefh 1.64e-19
C5803 X2.X2.X2.X2.X1.X2.X3.vin1 a_52792_24076# 0.199f
C5804 a_25326_15546# X1.X2.X2.X1.X2.X1.X3.vin2 8.07e-19
C5805 X1.X2.X2.X1.X2.X1.X3.vin1 a_22826_10734# 0.00837f
C5806 X2.X1.X1.X2.X2.X1.X3.vin1 a_34062_9010# 0.428f
C5807 a_52106_6962# X2.X2.X2.X1.X1.X1.vout 0.386f
C5808 X2.X1.X2.X3.vin1 X2.X1.X3.vin2 1.16f
C5809 X1.X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin1 0.00437f
C5810 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X3.vin1 0.0131f
C5811 a_38152_20264# a_37852_18358# 6.2e-19
C5812 X2.X1.X2.X2.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X2.vout 0.08f
C5813 X1.X1.X1.X1.X1.X2.X3.vin2 X1.X1.X1.X1.X2.X1.X1.vin2 3.94e-19
C5814 X2.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X3.vin1 0.0321f
C5815 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.vrefh 2.33e-19
C5816 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.vrefh 0.161f
C5817 X2.X1.X2.X1.X1.X1.X2.vin1 a_39966_4110# 8.88e-20
C5818 X2.X1.X2.X1.X1.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X1.vin2 8.93e-19
C5819 X1.X1.X1.X3.vin2 a_5082_14688# 0.00292f
C5820 a_39966_30794# X2.X1.X2.X2.X2.X1.X3.vin2 8.07e-19
C5821 a_37466_10734# X2.X1.X2.X1.X1.X2.X3.vin2 0.00846f
C5822 X1.X1.X2.X2.X2.X2.X1.vin2 a_10686_30794# 0.273f
C5823 a_22826_6962# a_23212_6962# 0.419f
C5824 X1.X2.X2.X2.X2.X2.vrefh X2.X1.X1.X1.X1.X2.X1.vin1 0.00437f
C5825 a_52406_16452# X2.X2.X2.X1.X2.X2.vout 0.418f
C5826 X1.X1.X1.X1.X2.X2.vout X1.X1.X1.X1.X2.X2.X3.vin2 0.08f
C5827 a_25326_17452# a_23512_16452# 1.15e-20
C5828 a_22826_25982# a_23512_24076# 3.08e-19
C5829 a_19422_28070# X1.X2.X1.X1.X1.X2.X3.vin2 0.277f
C5830 a_8872_24076# a_8572_22210# 6.71e-19
C5831 X2.X1.X2.X3.vin1 a_37766_16452# 5.31e-19
C5832 a_11072_7922# X1.X1.X2.X1.X1.X2.vrefh 1.64e-19
C5833 a_37766_24076# X2.X1.X2.X2.X1.X2.X3.vin1 0.42f
C5834 X2.X1.X1.X1.X2.X1.X2.vin1 X2.X1.X1.X1.X2.X2.vrefh 0.564f
C5835 a_48702_9010# a_49002_7064# 4.19e-20
C5836 X2.X2.X1.X2.X2.X1.vout a_48616_7064# 0.169f
C5837 X2.X2.X1.X1.X2.X2.X3.vin1 a_48702_20446# 0.42f
C5838 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 2.23e-19
C5839 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin1 0.195f
C5840 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 0.049f
C5841 X2.X1.X2.X1.X1.X1.vout X2.X1.X2.X1.X1.X1.X3.vin1 0.118f
C5842 a_19722_10916# a_19422_9010# 5.25e-20
C5843 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.vrefh 0.161f
C5844 a_19336_10916# X1.X2.X1.X2.X2.X1.vout 1.64e-19
C5845 X1.X2.X2.X2.X1.X2.X1.vin1 a_25712_23170# 0.195f
C5846 a_37466_22210# X2.X1.X2.X2.X1.X1.vout 0.387f
C5847 a_2582_17540# a_2582_15634# 0.00198f
C5848 X2.X1.X2.X3.vin1 a_37766_8828# 1.64e-19
C5849 a_16836_6104# X1.X2.X1.X2.X2.X2.X2.vin1 1.78e-19
C5850 X2.X1.X2.X1.X1.X1.X1.vin2 X2.X2.X2.vrefh 0.0128f
C5851 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X1.vout 0.0215f
C5852 a_34062_31882# X2.X1.X1.X1.X3.vin1 1.52e-19
C5853 X2.X1.X1.X1.X1.X1.vout a_34362_29936# 0.386f
C5854 X1.X1.X2.X1.X2.X2.vout a_8186_14586# 0.263f
C5855 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X1.X2.X2.X1.X1.X3.vin2 3.94e-19
C5856 X2.X1.X2.X2.X1.X2.X1.vin1 a_39966_21264# 8.22e-20
C5857 X1.X2.X3.vin2 a_20286_892# 0.0912f
C5858 X1.X2.X2.X2.X2.X2.X2.vin1 X2.X1.X1.X1.X1.X1.X1.vin2 0.00232f
C5859 a_52406_8828# X2.X2.X2.X1.X1.X2.vout 0.418f
C5860 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X2.vrefh 2.33e-19
C5861 a_8486_8828# X1.X1.X2.X1.X1.X2.vout 0.418f
C5862 a_37466_29834# a_37766_27888# 4.19e-20
C5863 a_8186_22210# a_8572_22210# 0.419f
C5864 X1.X1.X1.X1.X1.X1.X3.vin1 a_4396_31882# 0.199f
C5865 a_33976_14688# X2.X1.X1.X2.X1.X2.vout 0.0929f
C5866 X2.X1.X1.X1.X1.X2.X3.vin2 a_31862_25164# 8.07e-19
C5867 X2.X2.X1.X1.X3.vin2 X2.X2.X2.X3.vin2 7.46e-20
C5868 X1.X2.X1.X2.X2.X2.vout a_19422_5198# 0.418f
C5869 a_19722_7064# X1.X2.X1.X2.X2.X2.X3.vin2 3.85e-19
C5870 a_52106_25982# X2.X2.X2.X2.X3.vin1 0.372f
C5871 a_34062_31882# X2.X1.X1.X1.X1.X1.X3.vin2 0.267f
C5872 a_10686_28888# X1.X1.X2.X2.X2.X1.X1.vin2 8.88e-20
C5873 X2.X2.X2.X2.X1.X1.X3.vin1 a_52792_20264# 0.199f
C5874 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X1.X2.X2.vrefh 0.1f
C5875 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.vout 0.08f
C5876 X1.X2.X2.X2.vrefh a_25712_17452# 0.118f
C5877 X1.X2.X2.X1.X1.X1.X1.vin2 X2.X1.X2.vrefh 0.0128f
C5878 X2.X2.X2.X3.vin2 a_52406_24076# 6.03e-19
C5879 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin2 0.12f
C5880 X2.X1.X1.X2.X1.X2.vrefh a_31476_13728# 1.64e-19
C5881 X2.X2.X2.X1.X2.X2.vout X2.X2.X2.X1.X2.X1.vout 0.514f
C5882 X1.X2.X1.X2.X1.X1.X3.vin2 a_16836_15634# 0.354f
C5883 X2.X2.X2.X2.X2.X2.vrefh a_54992_28888# 0.118f
C5884 X1.X2.X3.vin1 a_19722_10916# 6.09e-19
C5885 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 0.216f
C5886 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X2.X1.X2.X2.X1.X1.vin2 0.00232f
C5887 a_46116_9916# a_46502_9916# 0.419f
C5888 a_52406_24076# a_54606_23170# 4.2e-20
C5889 X1.X1.X2.X1.X1.X1.X2.vin1 a_11072_6016# 0.197f
C5890 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.X1.vin1 0.206f
C5891 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X3.vin2 8.93e-19
C5892 X1.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X3.vin2 0.0011f
C5893 a_35312_892# X2.X3.vin1 0.461f
C5894 a_49002_18540# X2.X2.X3.vin2 6.58e-20
C5895 a_34062_24258# a_33976_22312# 3.14e-19
C5896 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin1 0.52f
C5897 a_33676_24258# a_34362_22312# 2.86e-19
C5898 a_54606_13640# X2.X2.X2.X1.X2.X1.X3.vin2 0.567f
C5899 a_2582_11822# a_2582_9916# 0.00198f
C5900 X1.X2.X1.X1.X1.X1.X2.vin1 a_17222_30882# 0.402f
C5901 a_2196_11822# X1.X1.X1.X2.X2.X1.X1.vin1 1.64e-19
C5902 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X2.vin1 0.242f
C5903 X2.X2.X1.X1.X1.X2.vrefh a_46502_28976# 8.22e-20
C5904 a_4396_31882# a_5082_29936# 2.86e-19
C5905 a_4782_31882# a_4696_29936# 3.14e-19
C5906 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X3.vin2 0.161f
C5907 X2.X1.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X1.X3.vin2 0.0533f
C5908 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X3.vin2 1.42e-20
C5909 a_52106_18358# a_52406_16452# 4.41e-20
C5910 a_8186_10734# a_8872_8828# 3.08e-19
C5911 X2.X2.X1.X1.X1.X2.X1.vin2 a_46502_27070# 8.88e-20
C5912 X2.X1.X2.X2.X1.X1.X3.vin1 a_38152_20264# 0.199f
C5913 X2.X1.X2.X1.X2.X1.X3.vin1 a_39966_11734# 0.52f
C5914 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 0.587f
C5915 X1.X2.X1.X2.X1.X2.vout a_19036_12822# 0.36f
C5916 X2.X2.X1.X1.X1.X2.X3.vin1 a_48316_28070# 0.199f
C5917 a_46502_28976# X2.X2.X1.X1.X1.X2.X3.vin2 7.84e-19
C5918 X2.X2.X2.X1.X1.X1.X1.vin1 a_54992_4110# 0.195f
C5919 X1.X2.X1.X2.X2.X1.X3.vin2 a_16836_8010# 0.354f
C5920 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin1 0.267f
C5921 a_48702_31882# a_49002_29936# 4.19e-20
C5922 a_8572_14586# a_8872_12640# 6.1e-19
C5923 a_23512_16452# a_22826_14586# 3.31e-19
C5924 X2.X2.X1.X1.X1.X1.vout a_48616_29936# 0.169f
C5925 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X2.vin1 0.00117f
C5926 a_2582_25164# a_4782_24258# 4.2e-20
C5927 X2.X2.X1.X2.X2.vrefh a_46116_9916# 1.64e-19
C5928 a_19422_20446# X1.X2.X3.vin1 1.64e-19
C5929 X1.X2.X1.X1.X2.X2.X3.vin2 a_19722_18540# 0.00846f
C5930 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X2.vin1 0.242f
C5931 X2.X2.X2.X2.X2.X1.vout a_52406_27888# 0.422f
C5932 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X3.vin2 0.102f
C5933 a_33976_14688# a_31862_13728# 2.68e-20
C5934 X2.X2.X1.X2.X3.vin1 a_49002_10916# 0.372f
C5935 X2.X2.X1.X1.X2.X2.vrefh a_46116_21352# 1.64e-19
C5936 X1.X2.X2.X2.X1.X1.X3.vin1 a_23512_20264# 0.199f
C5937 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X1.X2.X2.X2.X2.X1.vin1 0.668f
C5938 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X1.vin1 0.0689f
C5939 X2.X2.X2.X2.X1.X2.X3.vin2 a_54606_23170# 7.84e-19
C5940 a_8872_20264# a_8572_18358# 6.2e-19
C5941 X3.vin1 vout 0.104f
C5942 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X2.vrefh 0.076f
C5943 X2.X1.X2.X2.X1.X1.X3.vin2 a_38152_20264# 0.1f
C5944 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X3.vin2 0.161f
C5945 a_39966_4110# a_40352_4110# 0.419f
C5946 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X1.vout 0.399f
C5947 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 0.0903f
C5948 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.X3.vin1 0.587f
C5949 X2.X1.X1.X2.X1.X2.X3.vin1 a_31862_11822# 0.00207f
C5950 X2.X2.X1.X2.vrefh a_46116_17540# 1.64e-19
C5951 a_31862_21352# a_34062_20446# 4.2e-20
C5952 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X1.X3.vin1 0.00836f
C5953 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X1.X2.X2.X2.vin1 0.00117f
C5954 a_48316_12822# a_48616_10916# 6.48e-19
C5955 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X1.X3.vin2 0.0943f
C5956 a_52106_18358# X2.X2.X2.X1.X2.X2.X3.vin2 0.00846f
C5957 X2.X2.X2.X2.X1.X1.X3.vin1 a_54992_19358# 0.354f
C5958 a_25326_11734# a_25326_9828# 0.00198f
C5959 X2.X2.X2.X3.vin1 a_52106_14586# 7.98e-19
C5960 X2.X2.X1.X3.vin2 X2.X2.X2.X1.X3.vin2 7.46e-20
C5961 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X2.vrefh 0.267f
C5962 X2.X1.X1.X1.X2.X1.X1.vin2 a_31476_23258# 1.78e-19
C5963 X1.X2.X2.X1.X1.X2.vout X1.X2.X2.X1.X1.X1.vout 0.507f
C5964 X2.X2.X2.X2.X2.X2.X2.vin1 a_52792_31700# 5.34e-19
C5965 X1.X2.X2.X2.X1.X1.X3.vin2 X1.X2.X2.X2.X1.X1.X3.vin1 0.581f
C5966 X2.X2.X1.X1.X1.X1.X1.vin2 X2.X2.X1.X1.X1.X2.vrefh 0.076f
C5967 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X2.vrefh 0.00118f
C5968 a_19336_14688# X1.X2.X1.X2.X3.vin1 0.363f
C5969 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X2.vrefh 0.00118f
C5970 X2.X1.X1.X3.vin1 X2.X1.X2.X3.vin2 1.22e-19
C5971 X1.X2.X2.X1.X2.X2.vrefh a_25326_13640# 0.3f
C5972 a_52406_16452# X2.X2.X2.X1.X3.vin2 9.7e-20
C5973 X1.X1.X3.vin1 a_4782_16634# 2.92e-19
C5974 X2.X2.X1.X3.vin1 X2.X2.X3.vin1 0.188f
C5975 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.X1.X1.X1.vin2 3.94e-19
C5976 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.vout 0.118f
C5977 X1.X2.X2.X1.X1.X1.X1.vin1 a_25712_4110# 0.195f
C5978 X1.X2.X1.X1.X1.X2.vrefh X1.X1.X2.X2.X2.X2.vrefh 0.117f
C5979 a_34362_7064# X2.X1.X1.X2.X2.X2.X3.vin1 0.00874f
C5980 X1.X1.X2.X2.X2.X2.vout a_8572_29834# 0.0929f
C5981 X1.X1.X2.X2.X1.X2.X3.vin1 a_10686_23170# 0.52f
C5982 X2.X2.X3.vin1 a_48702_12822# 2.12e-19
C5983 X2.X1.X1.X2.X1.X2.vout a_34062_12822# 0.418f
C5984 X2.X1.X2.X2.X3.vin1 a_37766_20264# 1.52e-19
C5985 a_19036_16634# X1.X2.X1.X2.X1.X1.X3.vin2 0.1f
C5986 X1.X1.X1.X3.vin2 a_4696_10916# 0.355f
C5987 X2.X1.X2.X2.X1.X1.X3.vin2 a_40352_21264# 0.354f
C5988 X1.X1.X1.X1.X2.X1.X2.vin1 a_2196_23258# 0.197f
C5989 a_48616_10916# a_48702_9010# 3.21e-19
C5990 a_49002_10916# a_48316_9010# 2.97e-19
C5991 X2.X1.X2.X2.X2.X2.vrefh X2.X1.X2.X2.X2.X1.X2.vin1 0.564f
C5992 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X2.X1.X1.X1.vin1 0.206f
C5993 X1.X2.X2.X3.vin2 a_22826_18358# 0.263f
C5994 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X2.X1.X2.X1.X2.X1.vin2 0.00232f
C5995 a_46116_13728# a_46502_13728# 0.419f
C5996 a_2582_21352# a_4396_20446# 1.06e-19
C5997 X1.X1.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X1.X3.vin1 0.0321f
C5998 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X3.vin1 0.206f
C5999 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X2.vin1 0.0689f
C6000 X2.X1.X3.vin1 a_37466_18358# 5.87e-20
C6001 X1.X2.X2.X1.X1.X2.X2.vin1 a_25712_7922# 1.78e-19
C6002 X2.X1.X2.X1.X3.vin1 a_37766_5016# 1.52e-19
C6003 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X1.vin1 2.23e-19
C6004 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.X1.X1.X3.vin1 1.22e-19
C6005 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X2.X1.vin2 0.216f
C6006 a_13696_892# a_14082_892# 0.419f
C6007 X2.X2.X3.vin1 X2.X2.X1.X2.X1.X1.vout 2.91e-19
C6008 a_16836_25164# X1.X2.X1.X1.X2.X1.X2.vin1 1.78e-19
C6009 a_52106_22210# X2.X2.X2.X2.X1.X1.X3.vin2 0.00815f
C6010 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X3.vin1 1.22e-19
C6011 X2.X2.X2.X2.X3.vin2 a_52492_29834# 0.363f
C6012 a_54992_21264# a_54992_19358# 0.00396f
C6013 a_19722_7064# X1.X2.X1.X2.X2.X2.vout 0.263f
C6014 X1.X1.X1.X2.X1.X1.X2.vin1 X1.X1.X1.X2.X1.X2.vrefh 0.564f
C6015 a_8486_16452# X1.X1.X2.X1.X2.X2.X3.vin1 0.42f
C6016 a_48702_31882# a_46502_30882# 4.77e-21
C6017 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X3.vin1 0.00117f
C6018 X1.X1.X2.X2.X1.X2.X3.vin2 a_8486_24076# 0.277f
C6019 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X3.vin2 0.165f
C6020 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X1.vout 0.0215f
C6021 a_8486_27888# a_8186_25982# 5.25e-20
C6022 X2.X2.X2.X1.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X1.vin1 2.23e-19
C6023 X2.X2.X2.X1.X2.X1.X2.vin1 a_54992_11734# 1.78e-19
C6024 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X1.X3.vin2 0.0533f
C6025 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X2.vrefh 0.267f
C6026 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X2.X1.X1.X1.vin1 0.206f
C6027 a_31862_25164# X2.X1.X1.X1.X2.X1.X1.vin2 0.273f
C6028 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.X3.vin1 0.0131f
C6029 a_19036_9010# X1.X2.X1.X2.X2.X1.X3.vin2 0.1f
C6030 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X3.vin1 0.0321f
C6031 a_16836_11822# a_17222_11822# 0.419f
C6032 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin1 0.267f
C6033 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 0.234f
C6034 X2.X1.X2.X2.X1.X1.X2.vin1 a_40352_19358# 1.78e-19
C6035 X2.X1.X2.X2.X1.X2.vrefh a_39966_21264# 0.3f
C6036 X2.X1.X2.X2.X1.X1.X3.vin2 X2.X1.X2.X2.X1.X1.X1.vin1 2.23e-19
C6037 X2.X2.X2.X1.X2.X1.vout X2.X2.X2.X1.X3.vin2 0.399f
C6038 a_46502_17540# X2.X2.X1.X2.X1.X1.X1.vin2 0.273f
C6039 X2.X1.X2.X2.X2.X2.X3.vin2 X2.X2.vrefh 0.183f
C6040 a_54606_15546# X2.X2.X2.X1.X2.X1.X3.vin2 8.07e-19
C6041 X2.X2.X2.X1.X1.X1.X3.vin2 a_54992_6016# 0.354f
C6042 X1.X2.X1.X1.X1.X1.X3.vin2 a_17222_28976# 8.07e-19
C6043 a_19722_14688# X1.X2.X1.X2.X1.X2.X3.vin1 0.00874f
C6044 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 0.234f
C6045 X2.X1.X1.X2.X1.X2.vout a_33976_10916# 7.93e-20
C6046 X1.X2.X1.X1.X1.X2.X3.vin1 a_17222_27070# 0.00207f
C6047 X1.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X3.vin1 0.0604f
C6048 X2.X1.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin1 0.00437f
C6049 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X3.vin1 0.206f
C6050 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X3.vin2 0.102f
C6051 a_19722_18540# X1.X2.X1.X2.X1.X1.X3.vin2 3.49e-19
C6052 X1.X1.X1.X2.X1.X1.vout X1.X1.X1.X2.X1.X2.vout 0.507f
C6053 X1.X2.X1.X3.vin2 a_19422_16634# 5.21e-19
C6054 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.vrefh 0.267f
C6055 X2.X1.X2.X1.X2.X1.X3.vin2 a_38152_12640# 0.1f
C6056 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X2.vrefh 0.076f
C6057 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X1.vin2 0.076f
C6058 X2.X2.X2.X2.X1.X2.vout a_52492_22210# 0.0929f
C6059 a_4696_29936# X1.X1.X1.X1.X1.X2.vout 0.0929f
C6060 X1.X2.X2.X2.X3.vin2 a_23212_25982# 0.0927f
C6061 a_52792_20264# a_54606_19358# 1.06e-19
C6062 a_5082_22312# X1.X1.X1.X1.X2.X2.vout 0.263f
C6063 a_23512_31700# a_23212_29834# 6.71e-19
C6064 X2.X2.X1.X2.X1.X2.vout X2.X2.X1.X2.X1.X2.X3.vin2 0.075f
C6065 a_31862_13728# a_34062_12822# 4.2e-20
C6066 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X2.vin1 0.00117f
C6067 a_49002_26164# X2.X2.X1.X1.X3.vin2 0.241f
C6068 X1.X1.X1.X1.X2.X2.X2.vin1 a_2582_19446# 0.402f
C6069 a_54606_32700# a_54606_30794# 0.00198f
C6070 X2.X2.X2.X2.X2.X2.X2.vin1 X2.X2.X2.X2.X2.X2.X1.vin2 0.242f
C6071 a_25326_26982# X1.X2.X2.X2.X1.X2.X3.vin2 8.07e-19
C6072 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X3.vin2 8.93e-19
C6073 X1.X2.X2.X1.X2.X2.X1.vin2 a_25326_15546# 0.273f
C6074 a_23126_8828# a_23212_6962# 3.38e-19
C6075 X1.X2.X1.X3.vin2 a_19422_9010# 7.93e-20
C6076 a_25326_21264# a_23512_20264# 1.15e-20
C6077 X1.X1.X2.X1.X1.X1.X3.vin1 a_10686_4110# 0.52f
C6078 X2.X1.X3.vin1 X2.X1.X2.X1.X3.vin2 6.26e-19
C6079 X2.X1.X3.vin2 X2.X1.X1.X2.X3.vin1 4.41e-19
C6080 a_17222_21352# X1.X2.X1.X1.X2.X2.X2.vin1 8.88e-20
C6081 a_19336_29936# a_19036_28070# 6.71e-19
C6082 X1.X1.X1.X2.X2.X1.X3.vin1 a_4782_9010# 0.428f
C6083 a_11072_13640# a_11072_11734# 0.00396f
C6084 a_48616_18540# X2.X2.X3.vin1 0.354f
C6085 X2.X1.X1.X2.vrefh a_31476_19446# 0.118f
C6086 X1.X2.X1.X1.X2.X2.vout X1.X2.X1.X1.X2.X2.X3.vin2 0.08f
C6087 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 2.23e-19
C6088 X2.X2.X1.X2.X2.X2.X3.vin1 a_48702_5198# 0.42f
C6089 a_25712_9828# X1.X2.X2.X1.X1.X2.X1.vin2 1.78e-19
C6090 a_25326_26982# X1.X2.X2.X2.X2.X1.X1.vin1 0.417f
C6091 X1.X2.X2.X2.X2.X1.X1.vin2 a_25712_26982# 0.12f
C6092 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin2 0.12f
C6093 a_17222_9916# X1.X2.X1.X2.X2.X1.X1.vin2 0.273f
C6094 a_23126_27888# a_23212_25982# 3.21e-19
C6095 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X3.vin2 0.0533f
C6096 a_25326_21264# X1.X2.X2.X2.X1.X1.X3.vin2 0.567f
C6097 X1.X2.X2.X1.X1.X2.X1.vin2 a_25326_7922# 0.273f
C6098 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 0.234f
C6099 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X3.vin1 0.00118f
C6100 X1.X2.X3.vin1 X1.X2.X1.X3.vin2 1.04f
C6101 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.X1.vin2 8.93e-19
C6102 X1.X2.X2.X2.X2.X2.X2.vin1 a_25326_30794# 8.88e-20
C6103 a_48702_16634# X2.X2.X1.X2.X1.X1.X3.vin2 0.267f
C6104 X2.X1.X2.X2.X2.X1.X3.vin2 a_39966_26982# 7.84e-19
C6105 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X1.X1.vin1 0.0689f
C6106 X2.X2.X2.X1.X1.X2.vout a_52106_6962# 0.254f
C6107 X2.X1.X2.X2.X2.X1.vout a_37852_29834# 0.169f
C6108 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 0.581f
C6109 a_54992_13640# X2.X2.X2.X1.X2.X1.X1.vin2 1.78e-19
C6110 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X1.X2.X2.X2.X2.vrefh 0.1f
C6111 X1.X2.X1.X2.vrefh a_16836_19446# 0.118f
C6112 a_48316_31882# a_48702_31882# 0.419f
C6113 X1.X1.X2.X2.X3.vin1 a_8486_20264# 1.52e-19
C6114 a_40352_21264# X2.X1.X2.X2.X1.X1.X1.vin2 1.78e-19
C6115 X1.X2.X1.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X3.vin1 2.33e-19
C6116 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X1.vin1 0.206f
C6117 a_48702_5198# X2.X2.X1.X2.X2.X2.X3.vin2 0.277f
C6118 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin1 0.195f
C6119 X1.X2.X1.X2.X1.X2.X2.vin1 a_16836_11822# 0.197f
C6120 a_10686_32700# X1.X1.X2.X2.X2.X2.X1.vin2 8.88e-20
C6121 X1.X1.X1.X1.X1.X2.X3.vin2 a_2196_27070# 0.354f
C6122 a_4782_28070# a_2582_27070# 4.77e-21
C6123 X2.X2.X2.X3.vin2 a_52106_22210# 0.00292f
C6124 X2.X1.X1.X2.X1.X1.X2.vin1 a_31862_15634# 0.402f
C6125 a_31862_32788# X2.X1.X1.X1.X1.X1.X1.vin2 0.273f
C6126 a_48702_28070# a_46502_27070# 4.77e-21
C6127 X2.X2.X1.X1.X1.X2.X3.vin2 a_46116_27070# 0.354f
C6128 a_52406_12640# a_52492_10734# 3.21e-19
C6129 a_54606_19358# a_54992_19358# 0.419f
C6130 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X2.vrefh 0.076f
C6131 X1.X2.X2.X2.X2.X1.X3.vin2 a_23512_27888# 0.1f
C6132 X1.X1.X2.X2.X2.X2.X1.vin1 a_11072_28888# 1.64e-19
C6133 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin2 0.12f
C6134 X1.X2.X2.X2.X2.vrefh a_25712_25076# 0.118f
C6135 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin1 0.195f
C6136 a_23212_6962# a_23512_5016# 6.1e-19
C6137 X1.X2.X1.X1.X1.X2.X3.vin1 X1.X2.X1.X1.X1.X2.X2.vin1 0.00117f
C6138 a_39966_6016# X2.X1.X2.X1.X1.X1.X3.vin2 0.567f
C6139 a_48702_9010# X2.X2.X1.X2.X2.X1.X3.vin2 0.267f
C6140 a_17222_28976# a_19422_28070# 4.2e-20
C6141 X1.X2.X3.vin1 a_23126_5016# 8.66e-20
C6142 X2.X2.X2.X1.X2.X1.X1.vin2 X2.X2.X2.X1.X2.vrefh 0.1f
C6143 a_4782_9010# X1.X1.X1.X2.X2.X1.X3.vin2 0.267f
C6144 X1.X2.X2.X2.X1.X1.X3.vin2 X1.X2.X2.X2.X1.X1.X1.vin2 8.93e-19
C6145 X1.X2.X2.X2.X1.X1.X2.vin1 a_25326_19358# 8.88e-20
C6146 a_33976_29936# a_34062_28070# 3.38e-19
C6147 a_34362_29936# a_33676_28070# 3.31e-19
C6148 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X1.vin2 0.696f
C6149 X2.X2.X1.X3.vin2 a_49002_14688# 0.00292f
C6150 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.vout 0.075f
C6151 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.vrefh 0.161f
C6152 X1.X1.X2.X2.X2.X1.vout a_8572_25982# 1.64e-19
C6153 X1.X1.X2.X2.X3.vin2 X1.X1.X2.X3.vin2 0.17f
C6154 a_52406_20264# a_52492_18358# 3.21e-19
C6155 X2.X1.X2.X2.X2.X1.X3.vin1 a_37852_25982# 0.00251f
C6156 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.X1.vin1 0.206f
C6157 a_4696_26164# X1.X1.X1.X1.X2.X1.X3.vin1 0.00251f
C6158 a_34362_26164# X2.X1.X1.X3.vin1 0.509f
C6159 a_37852_6962# X2.X1.X2.X1.X1.X1.X3.vin2 0.00546f
C6160 X1.X2.X1.X2.X3.vin2 a_19336_7064# 0.363f
C6161 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X1.X2.X2.X1.X1.X1.vin1 0.668f
C6162 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin1 0.267f
C6163 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.vout 0.335f
C6164 X2.X2.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.X3.vin1 0.0174f
C6165 X2.X1.X1.X2.X2.X1.X2.vin1 a_31862_8010# 0.402f
C6166 a_25712_19358# a_25712_17452# 0.00396f
C6167 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X2.vin1 0.242f
C6168 a_17222_11822# a_19336_10916# 4.72e-20
C6169 X1.X1.X2.X2.X1.X1.vout a_8572_18358# 1.64e-19
C6170 X2.X1.X3.vin2 a_35312_892# 0.268f
C6171 X2.X2.X3.vin2 a_49002_7064# 5.84e-19
C6172 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X2.X1.X2.X1.X2.X2.vin1 0.00232f
C6173 X1.X2.X2.X1.X1.X1.X3.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 0.22f
C6174 a_23126_5016# a_25326_4110# 4.2e-20
C6175 a_54606_15546# a_54992_15546# 0.419f
C6176 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X1.vin2 3.94e-19
C6177 a_8572_18358# X1.X1.X2.X1.X2.X2.X3.vin2 0.00517f
C6178 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X2.vin1 0.242f
C6179 X1.X2.X2.vrefh X1.X3.vin1 0.00136f
C6180 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X1.vin2 0.1f
C6181 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X2.vin1 0.0689f
C6182 a_31862_17540# a_33676_16634# 1.06e-19
C6183 a_16836_9916# a_16836_8010# 0.00396f
C6184 X2.X2.X3.vin2 X2.X2.X2.vrefh 0.15f
C6185 a_23212_29834# X1.X2.X2.X2.X2.X1.X3.vin2 0.00546f
C6186 X1.X2.X3.vin2 a_22826_6962# 0.00111f
C6187 X1.X1.X2.X1.X2.X1.X3.vin1 a_8186_10734# 0.00837f
C6188 a_38152_24076# a_39966_23170# 1.06e-19
C6189 X2.X1.X1.X1.X2.X2.vrefh a_31862_23258# 0.3f
C6190 a_16836_21352# a_17222_21352# 0.419f
C6191 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X2.X1.X1.X2.X2.X1.vin2 0.00232f
C6192 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin1 0.195f
C6193 X1.X2.X2.X2.X1.X1.X1.vin2 X1.X2.X2.X2.X1.X1.X1.vin1 0.668f
C6194 a_49952_892# vss 0.973f
C6195 a_49566_892# vss 1.67f
C6196 X2.X3.vin2 vss 3.86f
C6197 a_43362_892# vss 0.997f
C6198 a_42976_892# vss 1.67f
C6199 X2.X3.vin1 vss 2.94f
C6200 a_35312_892# vss 1.01f
C6201 a_34926_892# vss 1.67f
C6202 X3.vin2 vss 7.74f
C6203 vout vss 0.355f
C6204 a_28482_892# vss 1.03f
C6205 a_28096_892# vss 1.67f
C6206 d7 vss 0.864f
C6207 a_20672_892# vss 0.97f
C6208 a_20286_892# vss 1.67f
C6209 X1.X3.vin2 vss 3.74f
C6210 X3.vin1 vss 7.99f
C6211 a_14082_892# vss 0.996f
C6212 a_13696_892# vss 1.67f
C6213 X1.X3.vin1 vss 2.98f
C6214 a_6032_892# vss 1.01f
C6215 a_5646_892# vss 1.67f
C6216 a_54992_4110# vss 1.66f
C6217 X2.X2.X2.X1.X1.X1.X1.vin1 vss 2.17f
C6218 a_54606_4110# vss 0.858f
C6219 X2.X2.X2.X1.X1.X1.X1.vin2 vss 2.21f
C6220 a_46502_4198# vss 0.888f
C6221 a_46116_4198# vss 1.67f
C6222 X2.X2.X2.vrefh vss 16.5f
C6223 a_52792_5016# vss 1.67f
C6224 X2.X2.X2.X1.X1.X1.X3.vin1 vss 0.982f
C6225 a_52406_5016# vss 0.854f
C6226 X2.X2.X1.X2.X2.X2.X3.vin2 vss 1.69f
C6227 a_48702_5198# vss 0.947f
C6228 a_48316_5198# vss 1.67f
C6229 X2.X2.X1.X2.X2.X2.X2.vin1 vss 1.8f
C6230 a_40352_4110# vss 1.66f
C6231 X2.X1.X2.X1.X1.X1.X1.vin1 vss 2.16f
C6232 a_39966_4110# vss 0.858f
C6233 X2.X1.X2.X1.X1.X1.X1.vin2 vss 2.19f
C6234 a_31862_4198# vss 0.888f
C6235 a_31476_4198# vss 1.67f
C6236 X2.X1.X2.vrefh vss 16.4f
C6237 a_38152_5016# vss 1.67f
C6238 X2.X1.X2.X1.X1.X1.X3.vin1 vss 0.982f
C6239 a_37766_5016# vss 0.854f
C6240 X2.X1.X1.X2.X2.X2.X3.vin2 vss 1.69f
C6241 a_34062_5198# vss 0.947f
C6242 a_33676_5198# vss 1.67f
C6243 X2.X1.X1.X2.X2.X2.X2.vin1 vss 1.8f
C6244 a_25712_4110# vss 1.66f
C6245 X1.X2.X2.X1.X1.X1.X1.vin1 vss 2.16f
C6246 a_25326_4110# vss 0.858f
C6247 X1.X2.X2.X1.X1.X1.X1.vin2 vss 2.19f
C6248 a_17222_4198# vss 0.888f
C6249 a_16836_4198# vss 1.67f
C6250 X1.X2.X2.vrefh vss 16.4f
C6251 a_23512_5016# vss 1.67f
C6252 X1.X2.X2.X1.X1.X1.X3.vin1 vss 0.982f
C6253 a_23126_5016# vss 0.854f
C6254 X1.X2.X1.X2.X2.X2.X3.vin2 vss 1.69f
C6255 a_19422_5198# vss 0.947f
C6256 a_19036_5198# vss 1.67f
C6257 X1.X2.X1.X2.X2.X2.X2.vin1 vss 1.8f
C6258 a_11072_4110# vss 1.66f
C6259 X1.X1.X2.X1.X1.X1.X1.vin1 vss 2.16f
C6260 a_10686_4110# vss 0.858f
C6261 X1.X1.X2.X1.X1.X1.X1.vin2 vss 2.19f
C6262 a_2582_4198# vss 0.888f
C6263 a_2196_4198# vss 1.67f
C6264 X1.X1.X2.vrefh vss 16.5f
C6265 a_8872_5016# vss 1.67f
C6266 X1.X1.X2.X1.X1.X1.X3.vin1 vss 0.982f
C6267 a_8486_5016# vss 0.854f
C6268 X1.X1.X1.X2.X2.X2.X3.vin2 vss 1.69f
C6269 a_4782_5198# vss 0.947f
C6270 a_4396_5198# vss 1.67f
C6271 X1.X1.X1.X2.X2.X2.X2.vin1 vss 1.8f
C6272 a_54992_6016# vss 1.66f
C6273 X2.X2.X2.X1.X1.X1.X3.vin2 vss 1.34f
C6274 X2.X2.X2.X1.X1.X1.X2.vin1 vss 1.8f
C6275 a_54606_6016# vss 0.883f
C6276 X2.X2.X1.X2.X2.X2.X1.vin2 vss 2.19f
C6277 X2.X2.X1.X2.X2.X2.X3.vin1 vss 0.896f
C6278 X2.X2.X1.X2.X2.X2.X1.vin1 vss 2.05f
C6279 a_46502_6104# vss 0.856f
C6280 a_46116_6104# vss 1.66f
C6281 a_40352_6016# vss 1.66f
C6282 X2.X1.X2.X1.X1.X1.X3.vin2 vss 1.34f
C6283 X2.X1.X2.X1.X1.X1.X2.vin1 vss 1.8f
C6284 a_39966_6016# vss 0.883f
C6285 X2.X1.X1.X2.X2.X2.X1.vin2 vss 2.19f
C6286 X2.X1.X1.X2.X2.X2.X3.vin1 vss 0.896f
C6287 X2.X1.X1.X2.X2.X2.X1.vin1 vss 2.05f
C6288 a_31862_6104# vss 0.856f
C6289 a_31476_6104# vss 1.66f
C6290 a_25712_6016# vss 1.66f
C6291 X1.X2.X2.X1.X1.X1.X3.vin2 vss 1.34f
C6292 X1.X2.X2.X1.X1.X1.X2.vin1 vss 1.8f
C6293 a_25326_6016# vss 0.883f
C6294 X1.X2.X1.X2.X2.X2.X1.vin2 vss 2.19f
C6295 X1.X2.X1.X2.X2.X2.X3.vin1 vss 0.896f
C6296 X1.X2.X1.X2.X2.X2.X1.vin1 vss 2.05f
C6297 a_17222_6104# vss 0.856f
C6298 a_16836_6104# vss 1.66f
C6299 a_11072_6016# vss 1.66f
C6300 X1.X1.X2.X1.X1.X1.X3.vin2 vss 1.34f
C6301 X1.X1.X2.X1.X1.X1.X2.vin1 vss 1.8f
C6302 a_10686_6016# vss 0.883f
C6303 X1.X1.X1.X2.X2.X2.X1.vin2 vss 2.21f
C6304 X1.X1.X1.X2.X2.X2.X3.vin1 vss 0.896f
C6305 X1.X1.X1.X2.X2.X2.X1.vin1 vss 2.05f
C6306 a_2582_6104# vss 0.856f
C6307 a_2196_6104# vss 1.66f
C6308 a_52492_6962# vss 1.66f
C6309 X2.X2.X2.X1.X1.X1.vout vss 0.861f
C6310 a_52106_6962# vss 0.96f
C6311 X2.X2.X1.X2.X2.X2.vout vss 1.18f
C6312 a_49002_7064# vss 0.962f
C6313 a_48616_7064# vss 1.66f
C6314 a_37852_6962# vss 1.66f
C6315 X2.X1.X2.X1.X1.X1.vout vss 0.861f
C6316 a_37466_6962# vss 0.96f
C6317 X2.X1.X1.X2.X2.X2.vout vss 1.18f
C6318 a_34362_7064# vss 0.962f
C6319 a_33976_7064# vss 1.66f
C6320 a_23212_6962# vss 1.66f
C6321 X1.X2.X2.X1.X1.X1.vout vss 0.861f
C6322 a_22826_6962# vss 0.96f
C6323 X1.X2.X1.X2.X2.X2.vout vss 1.18f
C6324 a_19722_7064# vss 0.962f
C6325 a_19336_7064# vss 1.66f
C6326 a_8572_6962# vss 1.66f
C6327 X1.X1.X2.X1.X1.X1.vout vss 0.861f
C6328 a_8186_6962# vss 0.96f
C6329 X1.X1.X1.X2.X2.X2.vout vss 1.18f
C6330 a_5082_7064# vss 0.962f
C6331 a_4696_7064# vss 1.66f
C6332 X2.X2.X2.X1.X1.X2.vrefh vss 4.22f
C6333 a_54992_7922# vss 1.66f
C6334 X2.X2.X2.X1.X1.X2.X1.vin1 vss 2.05f
C6335 a_54606_7922# vss 0.856f
C6336 X2.X2.X2.X1.X1.X2.X1.vin2 vss 2.19f
C6337 a_46502_8010# vss 0.883f
C6338 a_46116_8010# vss 1.66f
C6339 X2.X1.X2.X1.X1.X2.vrefh vss 4.07f
C6340 X2.X2.X1.X2.X2.X2.vrefh vss 4.05f
C6341 a_52792_8828# vss 1.67f
C6342 X2.X2.X2.X1.X1.X2.vout vss 1.11f
C6343 X2.X2.X2.X1.X1.X2.X3.vin1 vss 0.892f
C6344 a_52406_8828# vss 0.945f
C6345 X2.X2.X1.X2.X2.X1.X3.vin2 vss 1.32f
C6346 X2.X2.X1.X2.X2.X1.vout vss 0.816f
C6347 a_48702_9010# vss 0.854f
C6348 a_48316_9010# vss 1.67f
C6349 X2.X2.X1.X2.X2.X1.X2.vin1 vss 1.79f
C6350 a_40352_7922# vss 1.66f
C6351 X2.X1.X2.X1.X1.X2.X1.vin1 vss 2.05f
C6352 a_39966_7922# vss 0.856f
C6353 X2.X1.X2.X1.X1.X2.X1.vin2 vss 2.17f
C6354 a_31862_8010# vss 0.883f
C6355 a_31476_8010# vss 1.66f
C6356 X1.X2.X2.X1.X1.X2.vrefh vss 4.07f
C6357 X2.X1.X1.X2.X2.X2.vrefh vss 4.05f
C6358 a_38152_8828# vss 1.67f
C6359 X2.X1.X2.X1.X1.X2.vout vss 1.11f
C6360 X2.X1.X2.X1.X1.X2.X3.vin1 vss 0.892f
C6361 a_37766_8828# vss 0.945f
C6362 X2.X1.X1.X2.X2.X1.X3.vin2 vss 1.32f
C6363 X2.X1.X1.X2.X2.X1.vout vss 0.816f
C6364 a_34062_9010# vss 0.854f
C6365 a_33676_9010# vss 1.67f
C6366 X2.X1.X1.X2.X2.X1.X2.vin1 vss 1.79f
C6367 a_25712_7922# vss 1.66f
C6368 X1.X2.X2.X1.X1.X2.X1.vin1 vss 2.05f
C6369 a_25326_7922# vss 0.856f
C6370 X1.X2.X2.X1.X1.X2.X1.vin2 vss 2.17f
C6371 a_17222_8010# vss 0.883f
C6372 a_16836_8010# vss 1.66f
C6373 X1.X1.X2.X1.X1.X2.vrefh vss 4.07f
C6374 X1.X2.X1.X2.X2.X2.vrefh vss 4.05f
C6375 a_23512_8828# vss 1.67f
C6376 X1.X2.X2.X1.X1.X2.vout vss 1.11f
C6377 X1.X2.X2.X1.X1.X2.X3.vin1 vss 0.892f
C6378 a_23126_8828# vss 0.945f
C6379 X1.X2.X1.X2.X2.X1.X3.vin2 vss 1.32f
C6380 X1.X2.X1.X2.X2.X1.vout vss 0.816f
C6381 a_19422_9010# vss 0.854f
C6382 a_19036_9010# vss 1.67f
C6383 X1.X2.X1.X2.X2.X1.X2.vin1 vss 1.79f
C6384 a_11072_7922# vss 1.66f
C6385 X1.X1.X2.X1.X1.X2.X1.vin1 vss 2.05f
C6386 a_10686_7922# vss 0.856f
C6387 X1.X1.X2.X1.X1.X2.X1.vin2 vss 2.17f
C6388 a_2582_8010# vss 0.883f
C6389 a_2196_8010# vss 1.66f
C6390 X1.X1.X1.X2.X2.X2.vrefh vss 4.21f
C6391 a_8872_8828# vss 1.67f
C6392 X1.X1.X2.X1.X1.X2.vout vss 1.11f
C6393 X1.X1.X2.X1.X1.X2.X3.vin1 vss 0.892f
C6394 a_8486_8828# vss 0.945f
C6395 X1.X1.X1.X2.X2.X1.X3.vin2 vss 1.32f
C6396 X1.X1.X1.X2.X2.X1.vout vss 0.816f
C6397 a_4782_9010# vss 0.854f
C6398 a_4396_9010# vss 1.67f
C6399 X1.X1.X1.X2.X2.X1.X2.vin1 vss 1.8f
C6400 a_54992_9828# vss 1.66f
C6401 X2.X2.X2.X1.X1.X2.X3.vin2 vss 1.55f
C6402 X2.X2.X2.X1.X1.X2.X2.vin1 vss 1.8f
C6403 a_54606_9828# vss 0.884f
C6404 X2.X2.X1.X2.X2.X1.X1.vin2 vss 2.17f
C6405 X2.X2.X1.X2.X2.X1.X3.vin1 vss 0.91f
C6406 X2.X2.X1.X2.X2.X1.X1.vin1 vss 2.05f
C6407 a_46502_9916# vss 0.855f
C6408 a_46116_9916# vss 1.66f
C6409 a_40352_9828# vss 1.66f
C6410 X2.X1.X2.X1.X1.X2.X3.vin2 vss 1.55f
C6411 X2.X1.X2.X1.X1.X2.X2.vin1 vss 1.79f
C6412 a_39966_9828# vss 0.884f
C6413 X2.X1.X1.X2.X2.X1.X1.vin2 vss 2.17f
C6414 X2.X1.X1.X2.X2.X1.X3.vin1 vss 0.91f
C6415 X2.X1.X1.X2.X2.X1.X1.vin1 vss 2.05f
C6416 a_31862_9916# vss 0.855f
C6417 a_31476_9916# vss 1.66f
C6418 a_25712_9828# vss 1.66f
C6419 X1.X2.X2.X1.X1.X2.X3.vin2 vss 1.55f
C6420 X1.X2.X2.X1.X1.X2.X2.vin1 vss 1.79f
C6421 a_25326_9828# vss 0.884f
C6422 X1.X2.X1.X2.X2.X1.X1.vin2 vss 2.17f
C6423 X1.X2.X1.X2.X2.X1.X3.vin1 vss 0.91f
C6424 X1.X2.X1.X2.X2.X1.X1.vin1 vss 2.05f
C6425 a_17222_9916# vss 0.855f
C6426 a_16836_9916# vss 1.66f
C6427 a_11072_9828# vss 1.66f
C6428 X1.X1.X2.X1.X1.X2.X3.vin2 vss 1.55f
C6429 X1.X1.X2.X1.X1.X2.X2.vin1 vss 1.79f
C6430 a_10686_9828# vss 0.884f
C6431 X1.X1.X1.X2.X2.X1.X1.vin2 vss 2.18f
C6432 X1.X1.X1.X2.X2.X1.X3.vin1 vss 0.91f
C6433 X1.X1.X1.X2.X2.X1.X1.vin1 vss 2.05f
C6434 a_2582_9916# vss 0.855f
C6435 a_2196_9916# vss 1.66f
C6436 a_52492_10734# vss 1.67f
C6437 X2.X2.X2.X1.X3.vin1 vss 2.32f
C6438 a_52106_10734# vss 0.926f
C6439 X2.X2.X1.X2.X3.vin2 vss 1.96f
C6440 a_49002_10916# vss 0.93f
C6441 a_48616_10916# vss 1.67f
C6442 a_37852_10734# vss 1.67f
C6443 X2.X1.X2.X1.X3.vin1 vss 2.32f
C6444 a_37466_10734# vss 0.926f
C6445 X2.X1.X1.X2.X3.vin2 vss 1.96f
C6446 a_34362_10916# vss 0.93f
C6447 a_33976_10916# vss 1.67f
C6448 a_23212_10734# vss 1.67f
C6449 X1.X2.X2.X1.X3.vin1 vss 2.32f
C6450 a_22826_10734# vss 0.926f
C6451 X1.X2.X1.X2.X3.vin2 vss 1.96f
C6452 a_19722_10916# vss 0.93f
C6453 a_19336_10916# vss 1.67f
C6454 a_8572_10734# vss 1.67f
C6455 X1.X1.X2.X1.X3.vin1 vss 2.32f
C6456 a_8186_10734# vss 0.926f
C6457 X1.X1.X1.X2.X3.vin2 vss 1.96f
C6458 a_5082_10916# vss 0.93f
C6459 a_4696_10916# vss 1.67f
C6460 X2.X2.X2.X1.X2.vrefh vss 4.21f
C6461 a_54992_11734# vss 1.66f
C6462 X2.X2.X2.X1.X2.X1.X1.vin1 vss 2.05f
C6463 a_54606_11734# vss 0.855f
C6464 X2.X2.X2.X1.X2.X1.X1.vin2 vss 2.18f
C6465 a_46502_11822# vss 0.884f
C6466 a_46116_11822# vss 1.66f
C6467 X2.X1.X2.X1.X2.vrefh vss 4.06f
C6468 X2.X2.X1.X2.X2.vrefh vss 4.06f
C6469 a_52792_12640# vss 1.67f
C6470 X2.X2.X2.X1.X2.X1.X3.vin1 vss 0.905f
C6471 a_52406_12640# vss 0.854f
C6472 X2.X2.X1.X2.X1.X2.X3.vin2 vss 1.5f
C6473 a_48702_12822# vss 0.945f
C6474 a_48316_12822# vss 1.67f
C6475 X2.X2.X1.X2.X1.X2.X2.vin1 vss 1.79f
C6476 a_40352_11734# vss 1.66f
C6477 X2.X1.X2.X1.X2.X1.X1.vin1 vss 2.05f
C6478 a_39966_11734# vss 0.855f
C6479 X2.X1.X2.X1.X2.X1.X1.vin2 vss 2.17f
C6480 a_31862_11822# vss 0.884f
C6481 a_31476_11822# vss 1.66f
C6482 X1.X2.X2.X1.X2.vrefh vss 4.06f
C6483 X2.X1.X1.X2.X2.vrefh vss 4.06f
C6484 a_38152_12640# vss 1.67f
C6485 X2.X1.X2.X1.X2.X1.X3.vin1 vss 0.905f
C6486 a_37766_12640# vss 0.854f
C6487 X2.X1.X1.X2.X1.X2.X3.vin2 vss 1.5f
C6488 a_34062_12822# vss 0.945f
C6489 a_33676_12822# vss 1.67f
C6490 X2.X1.X1.X2.X1.X2.X2.vin1 vss 1.79f
C6491 a_25712_11734# vss 1.66f
C6492 X1.X2.X2.X1.X2.X1.X1.vin1 vss 2.05f
C6493 a_25326_11734# vss 0.855f
C6494 X1.X2.X2.X1.X2.X1.X1.vin2 vss 2.17f
C6495 a_17222_11822# vss 0.884f
C6496 a_16836_11822# vss 1.66f
C6497 X1.X1.X2.X1.X2.vrefh vss 4.06f
C6498 X1.X2.X1.X2.X2.vrefh vss 4.06f
C6499 a_23512_12640# vss 1.67f
C6500 X1.X2.X2.X1.X2.X1.X3.vin1 vss 0.905f
C6501 a_23126_12640# vss 0.854f
C6502 X1.X2.X1.X2.X1.X2.X3.vin2 vss 1.5f
C6503 a_19422_12822# vss 0.945f
C6504 a_19036_12822# vss 1.67f
C6505 X1.X2.X1.X2.X1.X2.X2.vin1 vss 1.79f
C6506 a_11072_11734# vss 1.66f
C6507 X1.X1.X2.X1.X2.X1.X1.vin1 vss 2.05f
C6508 a_10686_11734# vss 0.855f
C6509 X1.X1.X2.X1.X2.X1.X1.vin2 vss 2.17f
C6510 a_2582_11822# vss 0.884f
C6511 a_2196_11822# vss 1.66f
C6512 X1.X1.X1.X2.X2.vrefh vss 4.21f
C6513 a_8872_12640# vss 1.67f
C6514 X1.X1.X2.X1.X2.X1.X3.vin1 vss 0.905f
C6515 a_8486_12640# vss 0.854f
C6516 X1.X1.X1.X2.X1.X2.X3.vin2 vss 1.5f
C6517 a_4782_12822# vss 0.945f
C6518 a_4396_12822# vss 1.67f
C6519 X1.X1.X1.X2.X1.X2.X2.vin1 vss 1.8f
C6520 a_54992_13640# vss 1.66f
C6521 X2.X2.X2.X1.X2.X1.X3.vin2 vss 1.28f
C6522 X2.X2.X2.X1.X2.X1.X2.vin1 vss 1.8f
C6523 a_54606_13640# vss 0.883f
C6524 X2.X2.X1.X2.X1.X2.X1.vin2 vss 2.17f
C6525 X2.X2.X1.X2.X1.X2.X3.vin1 vss 0.887f
C6526 X2.X2.X1.X2.X1.X2.X1.vin1 vss 2.05f
C6527 a_46502_13728# vss 0.856f
C6528 a_46116_13728# vss 1.66f
C6529 a_40352_13640# vss 1.66f
C6530 X2.X1.X2.X1.X2.X1.X3.vin2 vss 1.28f
C6531 X2.X1.X2.X1.X2.X1.X2.vin1 vss 1.79f
C6532 a_39966_13640# vss 0.883f
C6533 X2.X1.X1.X2.X1.X2.X1.vin2 vss 2.17f
C6534 X2.X1.X1.X2.X1.X2.X3.vin1 vss 0.887f
C6535 X2.X1.X1.X2.X1.X2.X1.vin1 vss 2.05f
C6536 a_31862_13728# vss 0.856f
C6537 a_31476_13728# vss 1.66f
C6538 a_25712_13640# vss 1.66f
C6539 X1.X2.X2.X1.X2.X1.X3.vin2 vss 1.28f
C6540 X1.X2.X2.X1.X2.X1.X2.vin1 vss 1.79f
C6541 a_25326_13640# vss 0.883f
C6542 X1.X2.X1.X2.X1.X2.X1.vin2 vss 2.17f
C6543 X1.X2.X1.X2.X1.X2.X3.vin1 vss 0.887f
C6544 X1.X2.X1.X2.X1.X2.X1.vin1 vss 2.05f
C6545 a_17222_13728# vss 0.856f
C6546 a_16836_13728# vss 1.66f
C6547 a_11072_13640# vss 1.66f
C6548 X1.X1.X2.X1.X2.X1.X3.vin2 vss 1.28f
C6549 X1.X1.X2.X1.X2.X1.X2.vin1 vss 1.79f
C6550 a_10686_13640# vss 0.883f
C6551 X1.X1.X1.X2.X1.X2.X1.vin2 vss 2.19f
C6552 X1.X1.X1.X2.X1.X2.X3.vin1 vss 0.887f
C6553 X1.X1.X1.X2.X1.X2.X1.vin1 vss 2.05f
C6554 a_2582_13728# vss 0.856f
C6555 a_2196_13728# vss 1.66f
C6556 a_52492_14586# vss 1.66f
C6557 X2.X2.X2.X1.X3.vin2 vss 1.74f
C6558 X2.X2.X2.X1.X2.X1.vout vss 0.788f
C6559 a_52106_14586# vss 0.876f
C6560 X2.X2.X1.X2.X1.X2.vout vss 1.04f
C6561 X2.X2.X1.X2.X3.vin1 vss 2.11f
C6562 a_49002_14688# vss 0.909f
C6563 a_48616_14688# vss 1.66f
C6564 a_37852_14586# vss 1.66f
C6565 X2.X1.X2.X1.X3.vin2 vss 1.74f
C6566 X2.X1.X2.X1.X2.X1.vout vss 0.788f
C6567 a_37466_14586# vss 0.876f
C6568 X2.X1.X1.X2.X1.X2.vout vss 1.04f
C6569 X2.X1.X1.X2.X3.vin1 vss 2.11f
C6570 a_34362_14688# vss 0.909f
C6571 a_33976_14688# vss 1.66f
C6572 a_23212_14586# vss 1.66f
C6573 X1.X2.X2.X1.X3.vin2 vss 1.74f
C6574 X1.X2.X2.X1.X2.X1.vout vss 0.788f
C6575 a_22826_14586# vss 0.876f
C6576 X1.X2.X1.X2.X1.X2.vout vss 1.04f
C6577 X1.X2.X1.X2.X3.vin1 vss 2.11f
C6578 a_19722_14688# vss 0.909f
C6579 a_19336_14688# vss 1.66f
C6580 a_8572_14586# vss 1.66f
C6581 X1.X1.X2.X1.X3.vin2 vss 1.74f
C6582 X1.X1.X2.X1.X2.X1.vout vss 0.788f
C6583 a_8186_14586# vss 0.876f
C6584 X1.X1.X1.X2.X1.X2.vout vss 1.04f
C6585 X1.X1.X1.X2.X3.vin1 vss 2.11f
C6586 a_5082_14688# vss 0.909f
C6587 a_4696_14688# vss 1.66f
C6588 X2.X2.X2.X1.X2.X2.vrefh vss 4.21f
C6589 a_54992_15546# vss 1.66f
C6590 X2.X2.X2.X1.X2.X2.X1.vin1 vss 2.05f
C6591 a_54606_15546# vss 0.856f
C6592 X2.X2.X2.X1.X2.X2.X1.vin2 vss 2.18f
C6593 a_46502_15634# vss 0.883f
C6594 a_46116_15634# vss 1.66f
C6595 X2.X1.X2.X1.X2.X2.vrefh vss 4.05f
C6596 X2.X2.X1.X2.X1.X2.vrefh vss 4.05f
C6597 a_52792_16452# vss 1.67f
C6598 X2.X2.X2.X1.X2.X2.vout vss 1.04f
C6599 X2.X2.X2.X1.X2.X2.X3.vin1 vss 0.888f
C6600 a_52406_16452# vss 0.945f
C6601 X2.X2.X1.X2.X1.X1.X3.vin2 vss 1.3f
C6602 X2.X2.X1.X2.X1.X1.vout vss 0.842f
C6603 a_48702_16634# vss 0.854f
C6604 a_48316_16634# vss 1.67f
C6605 X2.X2.X1.X2.X1.X1.X2.vin1 vss 1.79f
C6606 a_40352_15546# vss 1.66f
C6607 X2.X1.X2.X1.X2.X2.X1.vin1 vss 2.05f
C6608 a_39966_15546# vss 0.856f
C6609 X2.X1.X2.X1.X2.X2.X1.vin2 vss 2.17f
C6610 a_31862_15634# vss 0.883f
C6611 a_31476_15634# vss 1.66f
C6612 X1.X2.X2.X1.X2.X2.vrefh vss 4.05f
C6613 X2.X1.X1.X2.X1.X2.vrefh vss 4.05f
C6614 a_38152_16452# vss 1.67f
C6615 X2.X1.X2.X1.X2.X2.vout vss 1.04f
C6616 X2.X1.X2.X1.X2.X2.X3.vin1 vss 0.888f
C6617 a_37766_16452# vss 0.945f
C6618 X2.X1.X1.X2.X1.X1.X3.vin2 vss 1.3f
C6619 X2.X1.X1.X2.X1.X1.vout vss 0.842f
C6620 a_34062_16634# vss 0.854f
C6621 a_33676_16634# vss 1.67f
C6622 X2.X1.X1.X2.X1.X1.X2.vin1 vss 1.79f
C6623 a_25712_15546# vss 1.66f
C6624 X1.X2.X2.X1.X2.X2.X1.vin1 vss 2.05f
C6625 a_25326_15546# vss 0.856f
C6626 X1.X2.X2.X1.X2.X2.X1.vin2 vss 2.17f
C6627 a_17222_15634# vss 0.883f
C6628 a_16836_15634# vss 1.66f
C6629 X1.X1.X2.X1.X2.X2.vrefh vss 4.05f
C6630 X1.X2.X1.X2.X1.X2.vrefh vss 4.05f
C6631 a_23512_16452# vss 1.67f
C6632 X1.X2.X2.X1.X2.X2.vout vss 1.04f
C6633 X1.X2.X2.X1.X2.X2.X3.vin1 vss 0.888f
C6634 a_23126_16452# vss 0.945f
C6635 X1.X2.X1.X2.X1.X1.X3.vin2 vss 1.3f
C6636 X1.X2.X1.X2.X1.X1.vout vss 0.842f
C6637 a_19422_16634# vss 0.854f
C6638 a_19036_16634# vss 1.67f
C6639 X1.X2.X1.X2.X1.X1.X2.vin1 vss 1.79f
C6640 a_11072_15546# vss 1.66f
C6641 X1.X1.X2.X1.X2.X2.X1.vin1 vss 2.05f
C6642 a_10686_15546# vss 0.856f
C6643 X1.X1.X2.X1.X2.X2.X1.vin2 vss 2.17f
C6644 a_2582_15634# vss 0.883f
C6645 a_2196_15634# vss 1.66f
C6646 X1.X1.X1.X2.X1.X2.vrefh vss 4.21f
C6647 a_8872_16452# vss 1.67f
C6648 X1.X1.X2.X1.X2.X2.vout vss 1.04f
C6649 X1.X1.X2.X1.X2.X2.X3.vin1 vss 0.888f
C6650 a_8486_16452# vss 0.945f
C6651 X1.X1.X1.X2.X1.X1.X3.vin2 vss 1.3f
C6652 X1.X1.X1.X2.X1.X1.vout vss 0.842f
C6653 a_4782_16634# vss 0.854f
C6654 a_4396_16634# vss 1.67f
C6655 X1.X1.X1.X2.X1.X1.X2.vin1 vss 1.8f
C6656 a_54992_17452# vss 1.66f
C6657 X2.X2.X2.X1.X2.X2.X3.vin2 vss 1.52f
C6658 X2.X2.X2.X1.X2.X2.X2.vin1 vss 1.8f
C6659 a_54606_17452# vss 0.884f
C6660 X2.X2.X1.X2.X1.X1.X1.vin2 vss 2.17f
C6661 X2.X2.X1.X2.X1.X1.X3.vin1 vss 0.912f
C6662 X2.X2.X1.X2.X1.X1.X1.vin1 vss 2.05f
C6663 a_46502_17540# vss 0.855f
C6664 a_46116_17540# vss 1.66f
C6665 a_40352_17452# vss 1.66f
C6666 X2.X1.X2.X1.X2.X2.X3.vin2 vss 1.52f
C6667 X2.X1.X2.X1.X2.X2.X2.vin1 vss 1.79f
C6668 a_39966_17452# vss 0.884f
C6669 X2.X1.X1.X2.X1.X1.X1.vin2 vss 2.17f
C6670 X2.X1.X1.X2.X1.X1.X3.vin1 vss 0.912f
C6671 X2.X1.X1.X2.X1.X1.X1.vin1 vss 2.05f
C6672 a_31862_17540# vss 0.855f
C6673 a_31476_17540# vss 1.66f
C6674 a_25712_17452# vss 1.66f
C6675 X1.X2.X2.X1.X2.X2.X3.vin2 vss 1.52f
C6676 X1.X2.X2.X1.X2.X2.X2.vin1 vss 1.79f
C6677 a_25326_17452# vss 0.884f
C6678 X1.X2.X1.X2.X1.X1.X1.vin2 vss 2.17f
C6679 X1.X2.X1.X2.X1.X1.X3.vin1 vss 0.912f
C6680 X1.X2.X1.X2.X1.X1.X1.vin1 vss 2.05f
C6681 a_17222_17540# vss 0.855f
C6682 a_16836_17540# vss 1.66f
C6683 a_11072_17452# vss 1.66f
C6684 X1.X1.X2.X1.X2.X2.X3.vin2 vss 1.52f
C6685 X1.X1.X2.X1.X2.X2.X2.vin1 vss 1.79f
C6686 a_10686_17452# vss 0.884f
C6687 X1.X1.X1.X2.X1.X1.X1.vin2 vss 2.18f
C6688 X1.X1.X1.X2.X1.X1.X3.vin1 vss 0.912f
C6689 X1.X1.X1.X2.X1.X1.X1.vin1 vss 2.05f
C6690 a_2582_17540# vss 0.855f
C6691 a_2196_17540# vss 1.66f
C6692 a_52492_18358# vss 1.67f
C6693 X2.X2.X3.vin2 vss 5.62f
C6694 X2.X2.X2.X3.vin1 vss 1.68f
C6695 a_52106_18358# vss 0.909f
C6696 X2.X2.X1.X3.vin2 vss 2.13f
C6697 X2.X2.X3.vin1 vss 4.8f
C6698 a_49002_18540# vss 0.91f
C6699 a_48616_18540# vss 1.67f
C6700 a_37852_18358# vss 1.67f
C6701 X2.X1.X3.vin2 vss 5.59f
C6702 X2.X1.X2.X3.vin1 vss 1.68f
C6703 a_37466_18358# vss 0.909f
C6704 X2.X1.X1.X3.vin2 vss 2.12f
C6705 X2.X1.X3.vin1 vss 4.78f
C6706 a_34362_18540# vss 0.91f
C6707 a_33976_18540# vss 1.67f
C6708 a_23212_18358# vss 1.67f
C6709 X1.X2.X3.vin2 vss 5.57f
C6710 X1.X2.X2.X3.vin1 vss 1.68f
C6711 a_22826_18358# vss 0.909f
C6712 X1.X2.X1.X3.vin2 vss 2.13f
C6713 X1.X2.X3.vin1 vss 4.78f
C6714 a_19722_18540# vss 0.91f
C6715 a_19336_18540# vss 1.67f
C6716 a_8572_18358# vss 1.67f
C6717 X1.X1.X3.vin2 vss 5.62f
C6718 X1.X1.X2.X3.vin1 vss 1.68f
C6719 a_8186_18358# vss 0.909f
C6720 X1.X1.X1.X3.vin2 vss 2.12f
C6721 X1.X1.X3.vin1 vss 4.8f
C6722 a_5082_18540# vss 0.91f
C6723 a_4696_18540# vss 1.67f
C6724 X2.X2.X2.X2.vrefh vss 4.21f
C6725 a_54992_19358# vss 1.66f
C6726 X2.X2.X2.X2.X1.X1.X1.vin1 vss 2.05f
C6727 a_54606_19358# vss 0.855f
C6728 X2.X2.X2.X2.X1.X1.X1.vin2 vss 2.18f
C6729 a_46502_19446# vss 0.884f
C6730 a_46116_19446# vss 1.66f
C6731 X2.X1.X2.X2.vrefh vss 4.05f
C6732 X2.X2.X1.X2.vrefh vss 4.05f
C6733 a_52792_20264# vss 1.67f
C6734 X2.X2.X2.X2.X1.X1.X3.vin1 vss 0.912f
C6735 a_52406_20264# vss 0.854f
C6736 X2.X2.X1.X1.X2.X2.X3.vin2 vss 1.52f
C6737 a_48702_20446# vss 0.945f
C6738 a_48316_20446# vss 1.67f
C6739 X2.X2.X1.X1.X2.X2.X2.vin1 vss 1.79f
C6740 a_40352_19358# vss 1.66f
C6741 X2.X1.X2.X2.X1.X1.X1.vin1 vss 2.05f
C6742 a_39966_19358# vss 0.855f
C6743 X2.X1.X2.X2.X1.X1.X1.vin2 vss 2.17f
C6744 a_31862_19446# vss 0.884f
C6745 a_31476_19446# vss 1.66f
C6746 X1.X2.X2.X2.vrefh vss 4.05f
C6747 X2.X1.X1.X2.vrefh vss 4.05f
C6748 a_38152_20264# vss 1.67f
C6749 X2.X1.X2.X2.X1.X1.X3.vin1 vss 0.912f
C6750 a_37766_20264# vss 0.854f
C6751 X2.X1.X1.X1.X2.X2.X3.vin2 vss 1.52f
C6752 a_34062_20446# vss 0.945f
C6753 a_33676_20446# vss 1.67f
C6754 X2.X1.X1.X1.X2.X2.X2.vin1 vss 1.79f
C6755 a_25712_19358# vss 1.66f
C6756 X1.X2.X2.X2.X1.X1.X1.vin1 vss 2.05f
C6757 a_25326_19358# vss 0.855f
C6758 X1.X2.X2.X2.X1.X1.X1.vin2 vss 2.17f
C6759 a_17222_19446# vss 0.884f
C6760 a_16836_19446# vss 1.66f
C6761 X1.X1.X2.X2.vrefh vss 4.05f
C6762 X1.X2.X1.X2.vrefh vss 4.05f
C6763 a_23512_20264# vss 1.67f
C6764 X1.X2.X2.X2.X1.X1.X3.vin1 vss 0.912f
C6765 a_23126_20264# vss 0.854f
C6766 X1.X2.X1.X1.X2.X2.X3.vin2 vss 1.52f
C6767 a_19422_20446# vss 0.945f
C6768 a_19036_20446# vss 1.67f
C6769 X1.X2.X1.X1.X2.X2.X2.vin1 vss 1.79f
C6770 a_11072_19358# vss 1.66f
C6771 X1.X1.X2.X2.X1.X1.X1.vin1 vss 2.05f
C6772 a_10686_19358# vss 0.855f
C6773 X1.X1.X2.X2.X1.X1.X1.vin2 vss 2.17f
C6774 a_2582_19446# vss 0.884f
C6775 a_2196_19446# vss 1.66f
C6776 X1.X1.X1.X2.vrefh vss 4.21f
C6777 a_8872_20264# vss 1.67f
C6778 X1.X1.X2.X2.X1.X1.X3.vin1 vss 0.912f
C6779 a_8486_20264# vss 0.854f
C6780 X1.X1.X1.X1.X2.X2.X3.vin2 vss 1.52f
C6781 a_4782_20446# vss 0.945f
C6782 a_4396_20446# vss 1.67f
C6783 X1.X1.X1.X1.X2.X2.X2.vin1 vss 1.8f
C6784 a_54992_21264# vss 1.66f
C6785 X2.X2.X2.X2.X1.X1.X3.vin2 vss 1.3f
C6786 X2.X2.X2.X2.X1.X1.X2.vin1 vss 1.8f
C6787 a_54606_21264# vss 0.883f
C6788 X2.X2.X1.X1.X2.X2.X1.vin2 vss 2.17f
C6789 X2.X2.X1.X1.X2.X2.X3.vin1 vss 0.888f
C6790 X2.X2.X1.X1.X2.X2.X1.vin1 vss 2.05f
C6791 a_46502_21352# vss 0.856f
C6792 a_46116_21352# vss 1.66f
C6793 a_40352_21264# vss 1.66f
C6794 X2.X1.X2.X2.X1.X1.X3.vin2 vss 1.3f
C6795 X2.X1.X2.X2.X1.X1.X2.vin1 vss 1.79f
C6796 a_39966_21264# vss 0.883f
C6797 X2.X1.X1.X1.X2.X2.X1.vin2 vss 2.17f
C6798 X2.X1.X1.X1.X2.X2.X3.vin1 vss 0.888f
C6799 X2.X1.X1.X1.X2.X2.X1.vin1 vss 2.05f
C6800 a_31862_21352# vss 0.856f
C6801 a_31476_21352# vss 1.66f
C6802 a_25712_21264# vss 1.66f
C6803 X1.X2.X2.X2.X1.X1.X3.vin2 vss 1.3f
C6804 X1.X2.X2.X2.X1.X1.X2.vin1 vss 1.79f
C6805 a_25326_21264# vss 0.883f
C6806 X1.X2.X1.X1.X2.X2.X1.vin2 vss 2.17f
C6807 X1.X2.X1.X1.X2.X2.X3.vin1 vss 0.888f
C6808 X1.X2.X1.X1.X2.X2.X1.vin1 vss 2.05f
C6809 a_17222_21352# vss 0.856f
C6810 a_16836_21352# vss 1.66f
C6811 a_11072_21264# vss 1.66f
C6812 X1.X1.X2.X2.X1.X1.X3.vin2 vss 1.3f
C6813 X1.X1.X2.X2.X1.X1.X2.vin1 vss 1.79f
C6814 a_10686_21264# vss 0.883f
C6815 X1.X1.X1.X1.X2.X2.X1.vin2 vss 2.18f
C6816 X1.X1.X1.X1.X2.X2.X3.vin1 vss 0.888f
C6817 X1.X1.X1.X1.X2.X2.X1.vin1 vss 2.05f
C6818 a_2582_21352# vss 0.856f
C6819 a_2196_21352# vss 1.66f
C6820 a_52492_22210# vss 1.66f
C6821 X2.X2.X2.X2.X1.X1.vout vss 0.841f
C6822 a_52106_22210# vss 0.909f
C6823 X2.X2.X1.X1.X2.X2.vout vss 1.04f
C6824 a_49002_22312# vss 0.876f
C6825 a_48616_22312# vss 1.66f
C6826 a_37852_22210# vss 1.66f
C6827 X2.X1.X2.X2.X1.X1.vout vss 0.842f
C6828 a_37466_22210# vss 0.909f
C6829 X2.X1.X1.X1.X2.X2.vout vss 1.04f
C6830 a_34362_22312# vss 0.876f
C6831 a_33976_22312# vss 1.66f
C6832 a_23212_22210# vss 1.66f
C6833 X1.X2.X2.X2.X1.X1.vout vss 0.841f
C6834 a_22826_22210# vss 0.909f
C6835 X1.X2.X1.X1.X2.X2.vout vss 1.04f
C6836 a_19722_22312# vss 0.876f
C6837 a_19336_22312# vss 1.66f
C6838 a_8572_22210# vss 1.66f
C6839 X1.X1.X2.X2.X1.X1.vout vss 0.842f
C6840 a_8186_22210# vss 0.909f
C6841 X1.X1.X1.X1.X2.X2.vout vss 1.04f
C6842 a_5082_22312# vss 0.876f
C6843 a_4696_22312# vss 1.66f
C6844 X2.X2.X2.X2.X1.X2.vrefh vss 4.21f
C6845 a_54992_23170# vss 1.66f
C6846 X2.X2.X2.X2.X1.X2.X1.vin1 vss 2.05f
C6847 a_54606_23170# vss 0.856f
C6848 X2.X2.X2.X2.X1.X2.X1.vin2 vss 2.19f
C6849 a_46502_23258# vss 0.883f
C6850 a_46116_23258# vss 1.66f
C6851 X2.X1.X2.X2.X1.X2.vrefh vss 4.05f
C6852 X2.X2.X1.X1.X2.X2.vrefh vss 4.05f
C6853 a_52792_24076# vss 1.67f
C6854 X2.X2.X2.X2.X1.X2.vout vss 1.04f
C6855 X2.X2.X2.X2.X1.X2.X3.vin1 vss 0.887f
C6856 a_52406_24076# vss 0.945f
C6857 X2.X2.X1.X1.X2.X1.X3.vin2 vss 1.28f
C6858 X2.X2.X1.X1.X2.X1.vout vss 0.789f
C6859 a_48702_24258# vss 0.854f
C6860 a_48316_24258# vss 1.67f
C6861 X2.X2.X1.X1.X2.X1.X2.vin1 vss 1.79f
C6862 a_40352_23170# vss 1.66f
C6863 X2.X1.X2.X2.X1.X2.X1.vin1 vss 2.05f
C6864 a_39966_23170# vss 0.856f
C6865 X2.X1.X2.X2.X1.X2.X1.vin2 vss 2.17f
C6866 a_31862_23258# vss 0.883f
C6867 a_31476_23258# vss 1.66f
C6868 X1.X2.X2.X2.X1.X2.vrefh vss 4.05f
C6869 X2.X1.X1.X1.X2.X2.vrefh vss 4.05f
C6870 a_38152_24076# vss 1.67f
C6871 X2.X1.X2.X2.X1.X2.vout vss 1.04f
C6872 X2.X1.X2.X2.X1.X2.X3.vin1 vss 0.887f
C6873 a_37766_24076# vss 0.945f
C6874 X2.X1.X1.X1.X2.X1.X3.vin2 vss 1.28f
C6875 X2.X1.X1.X1.X2.X1.vout vss 0.788f
C6876 a_34062_24258# vss 0.854f
C6877 a_33676_24258# vss 1.67f
C6878 X2.X1.X1.X1.X2.X1.X2.vin1 vss 1.79f
C6879 a_25712_23170# vss 1.66f
C6880 X1.X2.X2.X2.X1.X2.X1.vin1 vss 2.05f
C6881 a_25326_23170# vss 0.856f
C6882 X1.X2.X2.X2.X1.X2.X1.vin2 vss 2.17f
C6883 a_17222_23258# vss 0.883f
C6884 a_16836_23258# vss 1.66f
C6885 X1.X1.X2.X2.X1.X2.vrefh vss 4.05f
C6886 X1.X2.X1.X1.X2.X2.vrefh vss 4.05f
C6887 a_23512_24076# vss 1.67f
C6888 X1.X2.X2.X2.X1.X2.vout vss 1.04f
C6889 X1.X2.X2.X2.X1.X2.X3.vin1 vss 0.887f
C6890 a_23126_24076# vss 0.945f
C6891 X1.X2.X1.X1.X2.X1.X3.vin2 vss 1.28f
C6892 X1.X2.X1.X1.X2.X1.vout vss 0.789f
C6893 a_19422_24258# vss 0.854f
C6894 a_19036_24258# vss 1.67f
C6895 X1.X2.X1.X1.X2.X1.X2.vin1 vss 1.79f
C6896 a_11072_23170# vss 1.66f
C6897 X1.X1.X2.X2.X1.X2.X1.vin1 vss 2.05f
C6898 a_10686_23170# vss 0.856f
C6899 X1.X1.X2.X2.X1.X2.X1.vin2 vss 2.17f
C6900 a_2582_23258# vss 0.883f
C6901 a_2196_23258# vss 1.66f
C6902 X1.X1.X1.X1.X2.X2.vrefh vss 4.21f
C6903 a_8872_24076# vss 1.67f
C6904 X1.X1.X2.X2.X1.X2.vout vss 1.04f
C6905 X1.X1.X2.X2.X1.X2.X3.vin1 vss 0.887f
C6906 a_8486_24076# vss 0.945f
C6907 X1.X1.X1.X1.X2.X1.X3.vin2 vss 1.28f
C6908 X1.X1.X1.X1.X2.X1.vout vss 0.788f
C6909 a_4782_24258# vss 0.854f
C6910 a_4396_24258# vss 1.67f
C6911 X1.X1.X1.X1.X2.X1.X2.vin1 vss 1.8f
C6912 a_54992_25076# vss 1.66f
C6913 X2.X2.X2.X2.X1.X2.X3.vin2 vss 1.5f
C6914 X2.X2.X2.X2.X1.X2.X2.vin1 vss 1.8f
C6915 a_54606_25076# vss 0.884f
C6916 X2.X2.X1.X1.X2.X1.X1.vin2 vss 2.17f
C6917 X2.X2.X1.X1.X2.X1.X3.vin1 vss 0.905f
C6918 X2.X2.X1.X1.X2.X1.X1.vin1 vss 2.05f
C6919 a_46502_25164# vss 0.855f
C6920 a_46116_25164# vss 1.66f
C6921 a_40352_25076# vss 1.66f
C6922 X2.X1.X2.X2.X1.X2.X3.vin2 vss 1.5f
C6923 X2.X1.X2.X2.X1.X2.X2.vin1 vss 1.79f
C6924 a_39966_25076# vss 0.884f
C6925 X2.X1.X1.X1.X2.X1.X1.vin2 vss 2.17f
C6926 X2.X1.X1.X1.X2.X1.X3.vin1 vss 0.905f
C6927 X2.X1.X1.X1.X2.X1.X1.vin1 vss 2.05f
C6928 a_31862_25164# vss 0.855f
C6929 a_31476_25164# vss 1.66f
C6930 a_25712_25076# vss 1.66f
C6931 X1.X2.X2.X2.X1.X2.X3.vin2 vss 1.5f
C6932 X1.X2.X2.X2.X1.X2.X2.vin1 vss 1.79f
C6933 a_25326_25076# vss 0.884f
C6934 X1.X2.X1.X1.X2.X1.X1.vin2 vss 2.17f
C6935 X1.X2.X1.X1.X2.X1.X3.vin1 vss 0.905f
C6936 X1.X2.X1.X1.X2.X1.X1.vin1 vss 2.05f
C6937 a_17222_25164# vss 0.855f
C6938 a_16836_25164# vss 1.66f
C6939 a_11072_25076# vss 1.66f
C6940 X1.X1.X2.X2.X1.X2.X3.vin2 vss 1.5f
C6941 X1.X1.X2.X2.X1.X2.X2.vin1 vss 1.79f
C6942 a_10686_25076# vss 0.884f
C6943 X1.X1.X1.X1.X2.X1.X1.vin2 vss 2.18f
C6944 X1.X1.X1.X1.X2.X1.X3.vin1 vss 0.905f
C6945 X1.X1.X1.X1.X2.X1.X1.vin1 vss 2.05f
C6946 a_2582_25164# vss 0.855f
C6947 a_2196_25164# vss 1.66f
C6948 a_52492_25982# vss 1.67f
C6949 X2.X2.X2.X3.vin2 vss 2.05f
C6950 X2.X2.X2.X2.X3.vin1 vss 2.11f
C6951 a_52106_25982# vss 0.93f
C6952 X2.X2.X1.X1.X3.vin2 vss 1.73f
C6953 X2.X2.X1.X3.vin1 vss 1.91f
C6954 a_49002_26164# vss 0.926f
C6955 a_48616_26164# vss 1.67f
C6956 a_37852_25982# vss 1.67f
C6957 X2.X1.X2.X3.vin2 vss 2.29f
C6958 X2.X1.X2.X2.X3.vin1 vss 2.11f
C6959 a_37466_25982# vss 0.93f
C6960 X2.X1.X1.X1.X3.vin2 vss 1.74f
C6961 X2.X1.X1.X3.vin1 vss 1.67f
C6962 a_34362_26164# vss 0.926f
C6963 a_33976_26164# vss 1.67f
C6964 a_23212_25982# vss 1.67f
C6965 X1.X2.X2.X3.vin2 vss 2.05f
C6966 X1.X2.X2.X2.X3.vin1 vss 2.11f
C6967 a_22826_25982# vss 0.93f
C6968 X1.X2.X1.X1.X3.vin2 vss 1.73f
C6969 X1.X2.X1.X3.vin1 vss 1.91f
C6970 a_19722_26164# vss 0.926f
C6971 a_19336_26164# vss 1.67f
C6972 a_8572_25982# vss 1.67f
C6973 X1.X1.X2.X3.vin2 vss 2.29f
C6974 X1.X1.X2.X2.X3.vin1 vss 2.11f
C6975 a_8186_25982# vss 0.93f
C6976 X1.X1.X1.X1.X3.vin2 vss 1.74f
C6977 X1.X1.X1.X3.vin1 vss 1.67f
C6978 a_5082_26164# vss 0.926f
C6979 a_4696_26164# vss 1.67f
C6980 X2.X2.X2.X2.X2.vrefh vss 4.21f
C6981 a_54992_26982# vss 1.66f
C6982 X2.X2.X2.X2.X2.X1.X1.vin1 vss 2.05f
C6983 a_54606_26982# vss 0.855f
C6984 X2.X2.X2.X2.X2.X1.X1.vin2 vss 2.18f
C6985 a_46502_27070# vss 0.884f
C6986 a_46116_27070# vss 1.66f
C6987 X2.X1.X2.X2.X2.vrefh vss 4.06f
C6988 X2.X2.X1.X1.X2.vrefh vss 4.06f
C6989 a_52792_27888# vss 1.67f
C6990 X2.X2.X2.X2.X2.X1.X3.vin1 vss 0.91f
C6991 a_52406_27888# vss 0.854f
C6992 X2.X2.X1.X1.X1.X2.X3.vin2 vss 1.52f
C6993 a_48702_28070# vss 0.945f
C6994 a_48316_28070# vss 1.67f
C6995 X2.X2.X1.X1.X1.X2.X2.vin1 vss 1.79f
C6996 a_40352_26982# vss 1.66f
C6997 X2.X1.X2.X2.X2.X1.X1.vin1 vss 2.05f
C6998 a_39966_26982# vss 0.855f
C6999 X2.X1.X2.X2.X2.X1.X1.vin2 vss 2.17f
C7000 a_31862_27070# vss 0.884f
C7001 a_31476_27070# vss 1.66f
C7002 X1.X2.X2.X2.X2.vrefh vss 4.06f
C7003 X2.X1.X1.X1.X2.vrefh vss 4.06f
C7004 a_38152_27888# vss 1.67f
C7005 X2.X1.X2.X2.X2.X1.X3.vin1 vss 0.905f
C7006 a_37766_27888# vss 0.854f
C7007 X2.X1.X1.X1.X1.X2.X3.vin2 vss 1.54f
C7008 a_34062_28070# vss 0.945f
C7009 a_33676_28070# vss 1.67f
C7010 X2.X1.X1.X1.X1.X2.X2.vin1 vss 1.79f
C7011 a_25712_26982# vss 1.66f
C7012 X1.X2.X2.X2.X2.X1.X1.vin1 vss 2.05f
C7013 a_25326_26982# vss 0.855f
C7014 X1.X2.X2.X2.X2.X1.X1.vin2 vss 2.17f
C7015 a_17222_27070# vss 0.884f
C7016 a_16836_27070# vss 1.66f
C7017 X1.X1.X2.X2.X2.vrefh vss 4.06f
C7018 X1.X2.X1.X1.X2.vrefh vss 4.06f
C7019 a_23512_27888# vss 1.67f
C7020 X1.X2.X2.X2.X2.X1.X3.vin1 vss 0.91f
C7021 a_23126_27888# vss 0.854f
C7022 X1.X2.X1.X1.X1.X2.X3.vin2 vss 1.52f
C7023 a_19422_28070# vss 0.945f
C7024 a_19036_28070# vss 1.67f
C7025 X1.X2.X1.X1.X1.X2.X2.vin1 vss 1.79f
C7026 a_11072_26982# vss 1.66f
C7027 X1.X1.X2.X2.X2.X1.X1.vin1 vss 2.05f
C7028 a_10686_26982# vss 0.855f
C7029 X1.X1.X2.X2.X2.X1.X1.vin2 vss 2.17f
C7030 a_2582_27070# vss 0.884f
C7031 a_2196_27070# vss 1.66f
C7032 X1.X1.X1.X1.X2.vrefh vss 4.21f
C7033 a_8872_27888# vss 1.67f
C7034 X1.X1.X2.X2.X2.X1.X3.vin1 vss 0.905f
C7035 a_8486_27888# vss 0.854f
C7036 X1.X1.X1.X1.X1.X2.X3.vin2 vss 1.54f
C7037 a_4782_28070# vss 0.945f
C7038 a_4396_28070# vss 1.67f
C7039 X1.X1.X1.X1.X1.X2.X2.vin1 vss 1.8f
C7040 a_54992_28888# vss 1.66f
C7041 X2.X2.X2.X2.X2.X1.X3.vin2 vss 1.31f
C7042 X2.X2.X2.X2.X2.X1.X2.vin1 vss 1.8f
C7043 a_54606_28888# vss 0.883f
C7044 X2.X2.X1.X1.X1.X2.X1.vin2 vss 2.17f
C7045 X2.X2.X1.X1.X1.X2.X3.vin1 vss 0.89f
C7046 X2.X2.X1.X1.X1.X2.X1.vin1 vss 2.05f
C7047 a_46502_28976# vss 0.856f
C7048 a_46116_28976# vss 1.66f
C7049 a_40352_28888# vss 1.66f
C7050 X2.X1.X2.X2.X2.X1.X3.vin2 vss 1.28f
C7051 X2.X1.X2.X2.X2.X1.X2.vin1 vss 1.79f
C7052 a_39966_28888# vss 0.883f
C7053 X2.X1.X1.X1.X1.X2.X1.vin2 vss 2.17f
C7054 X2.X1.X1.X1.X1.X2.X3.vin1 vss 0.892f
C7055 X2.X1.X1.X1.X1.X2.X1.vin1 vss 2.05f
C7056 a_31862_28976# vss 0.856f
C7057 a_31476_28976# vss 1.66f
C7058 a_25712_28888# vss 1.66f
C7059 X1.X2.X2.X2.X2.X1.X3.vin2 vss 1.31f
C7060 X1.X2.X2.X2.X2.X1.X2.vin1 vss 1.79f
C7061 a_25326_28888# vss 0.883f
C7062 X1.X2.X1.X1.X1.X2.X1.vin2 vss 2.17f
C7063 X1.X2.X1.X1.X1.X2.X3.vin1 vss 0.89f
C7064 X1.X2.X1.X1.X1.X2.X1.vin1 vss 2.05f
C7065 a_17222_28976# vss 0.856f
C7066 a_16836_28976# vss 1.66f
C7067 a_11072_28888# vss 1.66f
C7068 X1.X1.X2.X2.X2.X1.X3.vin2 vss 1.28f
C7069 X1.X1.X2.X2.X2.X1.X2.vin1 vss 1.79f
C7070 a_10686_28888# vss 0.883f
C7071 X1.X1.X1.X1.X1.X2.X1.vin2 vss 2.19f
C7072 X1.X1.X1.X1.X1.X2.X3.vin1 vss 0.892f
C7073 X1.X1.X1.X1.X1.X2.X1.vin1 vss 2.05f
C7074 a_2582_28976# vss 0.856f
C7075 a_2196_28976# vss 1.66f
C7076 a_52492_29834# vss 1.66f
C7077 X2.X2.X2.X2.X3.vin2 vss 1.95f
C7078 X2.X2.X2.X2.X2.X1.vout vss 0.814f
C7079 a_52106_29834# vss 0.962f
C7080 X2.X2.X1.X1.X1.X2.vout vss 1.08f
C7081 X2.X2.X1.X1.X3.vin1 vss 2.31f
C7082 a_49002_29936# vss 0.96f
C7083 a_48616_29936# vss 1.66f
C7084 a_37852_29834# vss 1.66f
C7085 X2.X1.X2.X2.X3.vin2 vss 1.92f
C7086 X2.X1.X2.X2.X2.X1.vout vss 0.8f
C7087 a_37466_29834# vss 0.962f
C7088 X2.X1.X1.X1.X1.X2.vout vss 1.11f
C7089 X2.X1.X1.X1.X3.vin1 vss 2.32f
C7090 a_34362_29936# vss 0.96f
C7091 a_33976_29936# vss 1.66f
C7092 a_23212_29834# vss 1.66f
C7093 X1.X2.X2.X2.X3.vin2 vss 1.95f
C7094 X1.X2.X2.X2.X2.X1.vout vss 0.814f
C7095 a_22826_29834# vss 0.962f
C7096 X1.X2.X1.X1.X1.X2.vout vss 1.08f
C7097 X1.X2.X1.X1.X3.vin1 vss 2.31f
C7098 a_19722_29936# vss 0.96f
C7099 a_19336_29936# vss 1.66f
C7100 a_8572_29834# vss 1.66f
C7101 X1.X1.X2.X2.X3.vin2 vss 1.92f
C7102 X1.X1.X2.X2.X2.X1.vout vss 0.8f
C7103 a_8186_29834# vss 0.962f
C7104 X1.X1.X1.X1.X1.X2.vout vss 1.11f
C7105 X1.X1.X1.X1.X3.vin1 vss 2.32f
C7106 a_5082_29936# vss 0.96f
C7107 a_4696_29936# vss 1.66f
C7108 X2.X2.X2.X2.X2.X2.vrefh vss 4.21f
C7109 a_54992_30794# vss 1.66f
C7110 X2.X2.X2.X2.X2.X2.X1.vin1 vss 2.05f
C7111 a_54606_30794# vss 0.856f
C7112 X2.X2.X2.X2.X2.X2.X1.vin2 vss 2.24f
C7113 a_46502_30882# vss 0.883f
C7114 a_46116_30882# vss 1.66f
C7115 X2.X1.X2.X2.X2.X2.vrefh vss 4.05f
C7116 X2.X2.X1.X1.X1.X2.vrefh vss 4.07f
C7117 a_52792_31700# vss 1.67f
C7118 X2.X2.X2.X2.X2.X2.vout vss 1.17f
C7119 X2.X2.X2.X2.X2.X2.X3.vin1 vss 0.899f
C7120 a_52406_31700# vss 0.967f
C7121 X2.X2.X1.X1.X1.X1.X3.vin2 vss 1.32f
C7122 X2.X2.X1.X1.X1.X1.vout vss 0.853f
C7123 a_48702_31882# vss 0.879f
C7124 a_48316_31882# vss 1.67f
C7125 X2.X2.X1.X1.X1.X1.X2.vin1 vss 1.8f
C7126 a_40352_30794# vss 1.66f
C7127 X2.X1.X2.X2.X2.X2.X1.vin1 vss 2.05f
C7128 a_39966_30794# vss 0.856f
C7129 X2.X1.X2.X2.X2.X2.X1.vin2 vss 2.22f
C7130 a_31862_30882# vss 0.883f
C7131 a_31476_30882# vss 1.66f
C7132 X1.X2.X2.X2.X2.X2.vrefh vss 4.05f
C7133 X2.X1.X1.X1.X1.X2.vrefh vss 4.07f
C7134 a_38152_31700# vss 1.67f
C7135 X2.X1.X2.X2.X2.X2.vout vss 1.11f
C7136 X2.X1.X2.X2.X2.X2.X3.vin1 vss 0.894f
C7137 a_37766_31700# vss 0.967f
C7138 X2.X1.X1.X1.X1.X1.X3.vin2 vss 1.34f
C7139 X2.X1.X1.X1.X1.X1.vout vss 0.861f
C7140 a_34062_31882# vss 0.879f
C7141 a_33676_31882# vss 1.67f
C7142 X2.X1.X1.X1.X1.X1.X2.vin1 vss 1.8f
C7143 a_25712_30794# vss 1.66f
C7144 X1.X2.X2.X2.X2.X2.X1.vin1 vss 2.05f
C7145 a_25326_30794# vss 0.856f
C7146 X1.X2.X2.X2.X2.X2.X1.vin2 vss 2.22f
C7147 a_17222_30882# vss 0.883f
C7148 a_16836_30882# vss 1.66f
C7149 X1.X1.X2.X2.X2.X2.vrefh vss 4.05f
C7150 X1.X2.X1.X1.X1.X2.vrefh vss 4.07f
C7151 a_23512_31700# vss 1.67f
C7152 X1.X2.X2.X2.X2.X2.vout vss 1.17f
C7153 X1.X2.X2.X2.X2.X2.X3.vin1 vss 0.899f
C7154 a_23126_31700# vss 0.967f
C7155 X1.X2.X1.X1.X1.X1.X3.vin2 vss 1.32f
C7156 X1.X2.X1.X1.X1.X1.vout vss 0.853f
C7157 a_19422_31882# vss 0.879f
C7158 a_19036_31882# vss 1.67f
C7159 X1.X2.X1.X1.X1.X1.X2.vin1 vss 1.8f
C7160 a_11072_30794# vss 1.66f
C7161 X1.X1.X2.X2.X2.X2.X1.vin1 vss 2.05f
C7162 a_10686_30794# vss 0.856f
C7163 X1.X1.X2.X2.X2.X2.X1.vin2 vss 2.22f
C7164 a_2582_30882# vss 0.883f
C7165 a_2196_30882# vss 1.66f
C7166 X1.X1.X1.X1.X1.X2.vrefh vss 4.22f
C7167 a_8872_31700# vss 1.67f
C7168 X1.X1.X2.X2.X2.X2.vout vss 1.11f
C7169 X1.X1.X2.X2.X2.X2.X3.vin1 vss 0.894f
C7170 a_8486_31700# vss 0.967f
C7171 X1.X1.X1.X1.X1.X1.X3.vin2 vss 1.34f
C7172 X1.X1.X1.X1.X1.X1.vout vss 0.861f
C7173 a_4782_31882# vss 0.879f
C7174 a_4396_31882# vss 1.67f
C7175 X1.X1.X1.X1.X1.X1.X2.vin1 vss 1.8f
C7176 vrefh vss 1.34f
C7177 vrefl vss 3.21f
C7178 a_54992_32700# vss 1.66f
C7179 X2.X2.X2.X2.X2.X2.X3.vin2 vss 1.76f
C7180 X2.X2.X2.X2.X2.X2.X2.vin1 vss 1.83f
C7181 a_54606_32700# vss 0.887f
C7182 X2.X2.X1.X1.X1.X1.X1.vin2 vss 2.31f
C7183 X2.X2.X1.X1.X1.X1.X3.vin1 vss 0.999f
C7184 X2.X2.X1.X1.X1.X1.X1.vin1 vss 2.3f
C7185 a_46502_32788# vss 0.884f
C7186 a_46116_32788# vss 1.67f
C7187 X2.X2.vrefh vss 4.97f
C7188 a_40352_32700# vss 1.67f
C7189 X2.X1.X2.X2.X2.X2.X3.vin2 vss 1.69f
C7190 X2.X1.X2.X2.X2.X2.X2.vin1 vss 1.82f
C7191 a_39966_32700# vss 0.888f
C7192 X2.X1.X1.X1.X1.X1.X1.vin2 vss 2.31f
C7193 X2.X1.X1.X1.X1.X1.X3.vin1 vss 1f
C7194 X2.X1.X1.X1.X1.X1.X1.vin1 vss 2.3f
C7195 a_31862_32788# vss 0.884f
C7196 a_31476_32788# vss 1.67f
C7197 X2.vrefh vss 4.97f
C7198 a_25712_32700# vss 1.67f
C7199 X1.X2.X2.X2.X2.X2.X3.vin2 vss 1.74f
C7200 X1.X2.X2.X2.X2.X2.X2.vin1 vss 1.82f
C7201 a_25326_32700# vss 0.888f
C7202 X1.X2.X1.X1.X1.X1.X1.vin2 vss 2.31f
C7203 X1.X2.X1.X1.X1.X1.X3.vin1 vss 0.999f
C7204 X1.X2.X1.X1.X1.X1.X1.vin1 vss 2.3f
C7205 a_17222_32788# vss 0.884f
C7206 a_16836_32788# vss 1.67f
C7207 X1.X2.vrefh vss 4.97f
C7208 a_11072_32700# vss 1.67f
C7209 X1.X1.X2.X2.X2.X2.X3.vin2 vss 1.69f
C7210 X1.X1.X2.X2.X2.X2.X2.vin1 vss 1.82f
C7211 a_10686_32700# vss 0.888f
C7212 X1.X1.X1.X1.X1.X1.X1.vin2 vss 2.33f
C7213 X1.X1.X1.X1.X1.X1.X3.vin1 vss 1.01f
C7214 X1.X1.X1.X1.X1.X1.X1.vin1 vss 2.34f
C7215 a_2582_32788# vss 0.884f
C7216 a_2196_32788# vss 1.67f
C7217 X1.X1.X2.vrefh.t0 vss 0.0192f
C7218 X1.X1.X2.vrefh.t3 vss 7.12e-19
C7219 X1.X1.X2.vrefh.n0 vss 0.0125f
C7220 X1.X1.X2.vrefh.t1 vss 0.00866f
C7221 X1.X1.X2.vrefh.n1 vss 0.171f
C7222 X1.X1.X2.vrefh.n2 vss 0.425f
C7223 X1.X1.X2.vrefh.t2 vss 0.0179f
C7224 X1.X2.X2.vrefh.t0 vss 0.0183f
C7225 X1.X2.X2.vrefh.t2 vss 0.0196f
C7226 X1.X2.X2.vrefh.t3 vss 7.27e-19
C7227 X1.X2.X2.vrefh.n0 vss 0.0128f
C7228 X1.X2.X2.vrefh.t1 vss 0.00884f
C7229 X1.X2.X2.vrefh.n1 vss 0.174f
C7230 X1.X2.X2.vrefh.n2 vss 0.434f
C7231 X2.X1.X2.vrefh.t1 vss 0.0183f
C7232 X2.X1.X2.vrefh.t2 vss 0.0196f
C7233 X2.X1.X2.vrefh.t0 vss 7.27e-19
C7234 X2.X1.X2.vrefh.n0 vss 0.0128f
C7235 X2.X1.X2.vrefh.t3 vss 0.00884f
C7236 X2.X1.X2.vrefh.n1 vss 0.174f
C7237 X2.X1.X2.vrefh.n2 vss 0.434f
C7238 X2.X1.X3.vin1.t0 vss 0.00514f
C7239 X2.X1.X3.vin1.t1 vss 0.179f
C7240 X2.X1.X3.vin1.t2 vss 0.00574f
C7241 X2.X1.X3.vin1.t3 vss 0.00501f
C7242 X2.X1.X3.vin1.n0 vss 1.42f
C7243 X1.X1.X3.vin1.t3 vss 0.00514f
C7244 X1.X1.X3.vin1.t0 vss 0.179f
C7245 X1.X1.X3.vin1.t1 vss 0.00574f
C7246 X1.X1.X3.vin1.t2 vss 0.00501f
C7247 X1.X1.X3.vin1.n0 vss 1.42f
C7248 X3.vin2.t2 vss 0.0053f
C7249 X3.vin2.t1 vss 0.184f
C7250 X3.vin2.t3 vss 0.0148f
C7251 X3.vin2.t0 vss 0.00219f
C7252 X3.vin2.n0 vss 1.44f
C7253 X2.X1.X3.vin2.t1 vss 0.00205f
C7254 X2.X1.X3.vin2.t2 vss 0.0822f
C7255 X2.X1.X3.vin2.t3 vss 0.0133f
C7256 X2.X1.X3.vin2.t4 vss 0.00198f
C7257 X2.X1.X3.vin2.n0 vss 1.48f
C7258 X2.X1.X3.vin2.t0 vss 0.00478f
C7259 X1.X2.X3.vin2.t1 vss 0.00205f
C7260 X1.X2.X3.vin2.t0 vss 0.0822f
C7261 X1.X2.X3.vin2.t3 vss 0.0133f
C7262 X1.X2.X3.vin2.t2 vss 0.00198f
C7263 X1.X2.X3.vin2.n0 vss 1.48f
C7264 X2.X2.X3.vin2.t1 vss 0.00205f
C7265 X2.X2.X3.vin2.t0 vss 0.0822f
C7266 X2.X2.X3.vin2.t2 vss 0.0133f
C7267 X2.X2.X3.vin2.t3 vss 0.00198f
C7268 X2.X2.X3.vin2.n0 vss 1.48f
C7269 X3.vin1.t2 vss 0.00419f
C7270 X3.vin1.t0 vss 0.146f
C7271 X3.vin1.t1 vss 0.00408f
C7272 X3.vin1.t3 vss 0.00858f
C7273 d6.t3 vss 0.0335f
C7274 d6.t1 vss 0.0205f
C7275 d6.n0 vss 0.257f
C7276 d6.t0 vss 0.0335f
C7277 d6.t2 vss 0.0205f
C7278 d6.n1 vss 0.257f
C7279 X1.X1.X3.vin2.t3 vss 0.00205f
C7280 X1.X1.X3.vin2.t0 vss 0.0822f
C7281 X1.X1.X3.vin2.t1 vss 0.0133f
C7282 X1.X1.X3.vin2.t2 vss 0.00198f
C7283 X1.X1.X3.vin2.n0 vss 1.48f
C7284 d2.t30 vss 0.0587f
C7285 d2.t6 vss 0.036f
C7286 d2.t0 vss 0.036f
C7287 d2.t34 vss 0.0587f
C7288 d2.n0 vss 0.486f
C7289 d2.n1 vss 2.12f
C7290 d2.t3 vss 0.0587f
C7291 d2.t45 vss 0.036f
C7292 d2.n2 vss 0.497f
C7293 d2.n3 vss 2.13f
C7294 d2.t14 vss 0.0587f
C7295 d2.t54 vss 0.036f
C7296 d2.n4 vss 0.575f
C7297 d2.n5 vss 2.46f
C7298 d2.t16 vss 0.036f
C7299 d2.t52 vss 0.0587f
C7300 d2.n6 vss 0.564f
C7301 d2.t4 vss 0.036f
C7302 d2.t53 vss 0.0587f
C7303 d2.n7 vss 0.563f
C7304 d2.n8 vss 2.45f
C7305 d2.n9 vss 2.46f
C7306 d2.t51 vss 0.036f
C7307 d2.t48 vss 0.0587f
C7308 d2.n10 vss 0.486f
C7309 d2.n11 vss 1.75f
C7310 d2.t56 vss 0.036f
C7311 d2.t19 vss 0.0587f
C7312 d2.n12 vss 0.564f
C7313 d2.t40 vss 0.036f
C7314 d2.t20 vss 0.0587f
C7315 d2.n13 vss 0.563f
C7316 d2.t1 vss 0.036f
C7317 d2.t35 vss 0.0587f
C7318 d2.n14 vss 0.486f
C7319 d2.n15 vss 2.12f
C7320 d2.n16 vss 2.45f
C7321 d2.n17 vss 2.46f
C7322 d2.t17 vss 0.036f
C7323 d2.t12 vss 0.0587f
C7324 d2.n18 vss 0.486f
C7325 d2.n19 vss 1.79f
C7326 d2.t9 vss 0.0587f
C7327 d2.t10 vss 0.036f
C7328 d2.n20 vss 0.497f
C7329 d2.t61 vss 0.0587f
C7330 d2.t36 vss 0.036f
C7331 d2.n21 vss 0.497f
C7332 d2.n22 vss 2.13f
C7333 d2.t47 vss 0.0587f
C7334 d2.t11 vss 0.036f
C7335 d2.n23 vss 0.575f
C7336 d2.n24 vss 2.46f
C7337 d2.t63 vss 0.0587f
C7338 d2.t33 vss 0.036f
C7339 d2.n25 vss 0.574f
C7340 d2.n26 vss 2.46f
C7341 d2.n27 vss 1.68f
C7342 d2.n28 vss 3.67f
C7343 d2.t62 vss 0.036f
C7344 d2.t27 vss 0.0587f
C7345 d2.n29 vss 0.564f
C7346 d2.t44 vss 0.036f
C7347 d2.t28 vss 0.0587f
C7348 d2.n30 vss 0.563f
C7349 d2.t55 vss 0.036f
C7350 d2.t24 vss 0.0587f
C7351 d2.n31 vss 0.486f
C7352 d2.n32 vss 2.12f
C7353 d2.n33 vss 2.45f
C7354 d2.n34 vss 2.46f
C7355 d2.t25 vss 0.036f
C7356 d2.t22 vss 0.0587f
C7357 d2.n35 vss 0.486f
C7358 d2.n36 vss 1.75f
C7359 d2.t15 vss 0.0587f
C7360 d2.t23 vss 0.036f
C7361 d2.n37 vss 0.497f
C7362 d2.t58 vss 0.0587f
C7363 d2.t31 vss 0.036f
C7364 d2.n38 vss 0.497f
C7365 d2.n39 vss 2.13f
C7366 d2.t60 vss 0.0587f
C7367 d2.t29 vss 0.036f
C7368 d2.n40 vss 0.575f
C7369 d2.n41 vss 2.46f
C7370 d2.t8 vss 0.0587f
C7371 d2.t46 vss 0.036f
C7372 d2.n42 vss 0.574f
C7373 d2.n43 vss 2.46f
C7374 d2.n44 vss 1.73f
C7375 d2.n45 vss 1.43f
C7376 d2.n46 vss 5.83f
C7377 d2.t7 vss 0.036f
C7378 d2.t38 vss 0.0587f
C7379 d2.n47 vss 0.564f
C7380 d2.t59 vss 0.036f
C7381 d2.t39 vss 0.0587f
C7382 d2.n48 vss 0.563f
C7383 d2.t50 vss 0.036f
C7384 d2.t18 vss 0.0587f
C7385 d2.n49 vss 0.486f
C7386 d2.n50 vss 2.12f
C7387 d2.n51 vss 2.45f
C7388 d2.n52 vss 2.46f
C7389 d2.t37 vss 0.036f
C7390 d2.t32 vss 0.0587f
C7391 d2.n53 vss 0.486f
C7392 d2.n54 vss 1.79f
C7393 d2.t13 vss 0.0587f
C7394 d2.t21 vss 0.036f
C7395 d2.n55 vss 0.497f
C7396 d2.t2 vss 0.0587f
C7397 d2.t41 vss 0.036f
C7398 d2.n56 vss 0.497f
C7399 d2.n57 vss 2.13f
C7400 d2.t57 vss 0.0587f
C7401 d2.t26 vss 0.036f
C7402 d2.n58 vss 0.575f
C7403 d2.n59 vss 2.46f
C7404 d2.t5 vss 0.0587f
C7405 d2.t43 vss 0.036f
C7406 d2.n60 vss 0.574f
C7407 d2.n61 vss 2.46f
C7408 d2.n62 vss 1.68f
C7409 d2.n63 vss 1.43f
C7410 d2.n64 vss 5.83f
C7411 d2.n65 vss 3.67f
C7412 d2.t42 vss 0.0587f
C7413 d2.t49 vss 0.036f
C7414 d2.n66 vss 0.497f
C7415 d2.n67 vss 1.73f
C7416 d2.n68 vss 2.46f
C7417 d2.n69 vss 0.574f
C7418 d4.t5 vss 0.0229f
C7419 d4.t12 vss 0.0372f
C7420 d4.t14 vss 0.0229f
C7421 d4.n0 vss 0.135f
C7422 d4.t6 vss 0.0372f
C7423 d4.n1 vss 0.329f
C7424 d4.t4 vss 0.0373f
C7425 d4.t15 vss 0.0229f
C7426 d4.n2 vss 0.507f
C7427 d4.n3 vss 3.23f
C7428 d4.t0 vss 0.0229f
C7429 d4.n4 vss 0.135f
C7430 d4.t9 vss 0.0372f
C7431 d4.n5 vss 0.368f
C7432 d4.t10 vss 0.0373f
C7433 d4.t2 vss 0.0229f
C7434 d4.n6 vss 0.468f
C7435 d4.n7 vss 1.91f
C7436 d4.n8 vss 5.84f
C7437 d4.t3 vss 0.0229f
C7438 d4.n9 vss 0.135f
C7439 d4.t11 vss 0.0372f
C7440 d4.n10 vss 0.329f
C7441 d4.t7 vss 0.0373f
C7442 d4.t1 vss 0.0229f
C7443 d4.n11 vss 0.507f
C7444 d4.n12 vss 1.91f
C7445 d4.n13 vss 5.84f
C7446 d4.t13 vss 0.0373f
C7447 d4.t8 vss 0.0229f
C7448 d4.n14 vss 0.468f
C7449 d4.n15 vss 3.23f
C7450 d4.n16 vss 0.368f
C7451 d4.n17 vss 0.135f
C7452 X1.X2.X3.vin1.t3 vss 0.00514f
C7453 X1.X2.X3.vin1.t0 vss 0.179f
C7454 X1.X2.X3.vin1.t2 vss 0.00574f
C7455 X1.X2.X3.vin1.t1 vss 0.00501f
C7456 X1.X2.X3.vin1.n0 vss 1.42f
C7457 X2.X2.X2.vrefh.t0 vss 0.0192f
C7458 X2.X2.X2.vrefh.t1 vss 7.12e-19
C7459 X2.X2.X2.vrefh.n0 vss 0.0125f
C7460 X2.X2.X2.vrefh.t2 vss 0.00866f
C7461 X2.X2.X2.vrefh.n1 vss 0.171f
C7462 X2.X2.X2.vrefh.n2 vss 0.425f
C7463 X2.X2.X2.vrefh.t3 vss 0.0179f
C7464 d5.t5 vss 0.083f
C7465 d5.t7 vss 0.0509f
C7466 d5.n0 vss 0.638f
C7467 d5.t6 vss 0.083f
C7468 d5.t1 vss 0.0509f
C7469 d5.n1 vss 0.638f
C7470 d5.t3 vss 0.083f
C7471 d5.t2 vss 0.0509f
C7472 d5.n2 vss 0.638f
C7473 d5.n3 vss 6.2f
C7474 d5.t4 vss 0.083f
C7475 d5.t0 vss 0.0509f
C7476 d5.n4 vss 0.638f
C7477 d5.n5 vss 6.2f
C7478 d3.t7 vss 0.0303f
C7479 d3.t22 vss 0.0186f
C7480 d3.t17 vss 0.0304f
C7481 d3.t6 vss 0.0187f
C7482 d3.n0 vss 0.417f
C7483 d3.t13 vss 0.0304f
C7484 d3.t30 vss 0.0187f
C7485 d3.n1 vss 0.407f
C7486 d3.n2 vss 0.539f
C7487 d3.n3 vss 0.562f
C7488 d3.n4 vss 0.556f
C7489 d3.n5 vss 0.565f
C7490 d3.n6 vss 0.375f
C7491 d3.n7 vss 0.588f
C7492 d3.n8 vss 0.581f
C7493 d3.n9 vss 0.591f
C7494 d3.t8 vss 0.0187f
C7495 d3.t23 vss 0.0304f
C7496 d3.n10 vss 0.411f
C7497 d3.n11 vss 0.5f
C7498 d3.n12 vss 0.562f
C7499 d3.n13 vss 0.556f
C7500 d3.n14 vss 0.565f
C7501 d3.t27 vss 0.0187f
C7502 d3.t19 vss 0.0304f
C7503 d3.n15 vss 0.404f
C7504 d3.n16 vss 0.558f
C7505 d3.n17 vss 0.395f
C7506 d3.n18 vss 0.347f
C7507 d3.n19 vss 1.75f
C7508 d3.t31 vss 0.0187f
C7509 d3.t25 vss 0.0304f
C7510 d3.n20 vss 0.377f
C7511 d3.t10 vss 0.0187f
C7512 d3.t26 vss 0.0304f
C7513 d3.n21 vss 0.411f
C7514 d3.n22 vss 0.5f
C7515 d3.n23 vss 0.562f
C7516 d3.n24 vss 0.556f
C7517 d3.n25 vss 0.565f
C7518 d3.n26 vss 0.375f
C7519 d3.n27 vss 0.588f
C7520 d3.n28 vss 0.581f
C7521 d3.n29 vss 0.591f
C7522 d3.t18 vss 0.0304f
C7523 d3.t4 vss 0.0187f
C7524 d3.n30 vss 0.407f
C7525 d3.n31 vss 0.539f
C7526 d3.n32 vss 0.562f
C7527 d3.n33 vss 0.556f
C7528 d3.n34 vss 0.565f
C7529 d3.t21 vss 0.0304f
C7530 d3.t12 vss 0.0188f
C7531 d3.n35 vss 0.424f
C7532 d3.n36 vss 0.519f
C7533 d3.n37 vss 0.395f
C7534 d3.n38 vss 0.368f
C7535 d3.n39 vss 0.789f
C7536 d3.n40 vss 3.59f
C7537 d3.t20 vss 0.0304f
C7538 d3.t9 vss 0.0188f
C7539 d3.n41 vss 0.424f
C7540 d3.t15 vss 0.0306f
C7541 d3.t2 vss 0.0187f
C7542 d3.n42 vss 0.414f
C7543 d3.n43 vss 0.539f
C7544 d3.n44 vss 0.562f
C7545 d3.n45 vss 0.556f
C7546 d3.n46 vss 0.565f
C7547 d3.n47 vss 0.375f
C7548 d3.n48 vss 0.588f
C7549 d3.n49 vss 0.581f
C7550 d3.n50 vss 0.591f
C7551 d3.t14 vss 0.0187f
C7552 d3.t0 vss 0.0304f
C7553 d3.n51 vss 0.411f
C7554 d3.n52 vss 0.5f
C7555 d3.n53 vss 0.562f
C7556 d3.n54 vss 0.556f
C7557 d3.n55 vss 0.565f
C7558 d3.t5 vss 0.0187f
C7559 d3.t28 vss 0.0306f
C7560 d3.n56 vss 0.411f
C7561 d3.n57 vss 0.558f
C7562 d3.n58 vss 0.395f
C7563 d3.n59 vss 0.347f
C7564 d3.n60 vss 0.747f
C7565 d3.n61 vss 3.59f
C7566 d3.t11 vss 0.0187f
C7567 d3.t3 vss 0.0306f
C7568 d3.n62 vss 0.384f
C7569 d3.n63 vss 1.79f
C7570 d3.t1 vss 0.0304f
C7571 d3.t24 vss 0.0188f
C7572 d3.n64 vss 0.424f
C7573 d3.n65 vss 0.519f
C7574 d3.n66 vss 0.395f
C7575 d3.n67 vss 0.368f
C7576 d3.n68 vss 0.565f
C7577 d3.n69 vss 0.556f
C7578 d3.n70 vss 0.562f
C7579 d3.n71 vss 0.591f
C7580 d3.n72 vss 0.581f
C7581 d3.n73 vss 0.588f
C7582 d3.t16 vss 0.0186f
C7583 d3.t29 vss 0.0304f
C7584 d3.n74 vss 0.418f
C7585 d3.n75 vss 0.565f
C7586 d3.n76 vss 0.556f
C7587 d3.n77 vss 0.562f
C7588 d3.n78 vss 0.539f
C7589 d3.n79 vss 0.375f
C7590 d3.n80 vss 0.5f
C7591 d3.n81 vss 0.415f
C7592 d1.t127 vss 0.056f
C7593 d1.t78 vss 0.0343f
C7594 d1.n0 vss 0.425f
C7595 d1.t44 vss 0.056f
C7596 d1.t122 vss 0.0343f
C7597 d1.n1 vss 0.425f
C7598 d1.n2 vss 0.535f
C7599 d1.t15 vss 0.056f
C7600 d1.t63 vss 0.0343f
C7601 d1.n3 vss 0.425f
C7602 d1.n4 vss 0.0262f
C7603 d1.t2 vss 0.056f
C7604 d1.t81 vss 0.0343f
C7605 d1.n5 vss 0.425f
C7606 d1.n6 vss 0.0262f
C7607 d1.t85 vss 0.056f
C7608 d1.t29 vss 0.0343f
C7609 d1.n7 vss 0.425f
C7610 d1.n8 vss 0.0262f
C7611 d1.t104 vss 0.056f
C7612 d1.t49 vss 0.0343f
C7613 d1.n9 vss 0.425f
C7614 d1.n10 vss 0.0262f
C7615 d1.t120 vss 0.056f
C7616 d1.t72 vss 0.0343f
C7617 d1.n11 vss 0.425f
C7618 d1.n12 vss 0.0262f
C7619 d1.t11 vss 0.056f
C7620 d1.t87 vss 0.0343f
C7621 d1.n13 vss 0.425f
C7622 d1.n14 vss 0.0262f
C7623 d1.t6 vss 0.0343f
C7624 d1.t102 vss 0.056f
C7625 d1.n15 vss 0.425f
C7626 d1.t90 vss 0.0343f
C7627 d1.t53 vss 0.056f
C7628 d1.n16 vss 0.42f
C7629 d1.n17 vss 1.01f
C7630 d1.t113 vss 0.0343f
C7631 d1.t77 vss 0.056f
C7632 d1.n18 vss 0.425f
C7633 d1.n19 vss 1.07f
C7634 d1.t33 vss 0.0343f
C7635 d1.t101 vss 0.056f
C7636 d1.n20 vss 0.42f
C7637 d1.n21 vss 0.997f
C7638 d1.t75 vss 0.0343f
C7639 d1.t8 vss 0.056f
C7640 d1.n22 vss 0.425f
C7641 d1.n23 vss 0.997f
C7642 d1.t97 vss 0.0343f
C7643 d1.t26 vss 0.056f
C7644 d1.n24 vss 0.42f
C7645 d1.n25 vss 1.01f
C7646 d1.t16 vss 0.0343f
C7647 d1.t79 vss 0.056f
C7648 d1.n26 vss 0.425f
C7649 d1.n27 vss 1.07f
C7650 d1.t34 vss 0.0343f
C7651 d1.t107 vss 0.056f
C7652 d1.n28 vss 0.42f
C7653 d1.n29 vss 0.651f
C7654 d1.t74 vss 0.0343f
C7655 d1.t40 vss 0.056f
C7656 d1.n30 vss 0.425f
C7657 d1.t20 vss 0.0343f
C7658 d1.t119 vss 0.056f
C7659 d1.n31 vss 0.42f
C7660 d1.n32 vss 1.01f
C7661 d1.t55 vss 0.0343f
C7662 d1.t18 vss 0.056f
C7663 d1.n33 vss 0.425f
C7664 d1.n34 vss 1.07f
C7665 d1.t106 vss 0.0343f
C7666 d1.t36 vss 0.056f
C7667 d1.n35 vss 0.42f
C7668 d1.n36 vss 0.997f
C7669 d1.t14 vss 0.0343f
C7670 d1.t76 vss 0.056f
C7671 d1.n37 vss 0.425f
C7672 d1.n38 vss 0.997f
C7673 d1.t31 vss 0.0343f
C7674 d1.t99 vss 0.056f
C7675 d1.n39 vss 0.42f
C7676 d1.n40 vss 1.01f
C7677 d1.t17 vss 0.0343f
C7678 d1.t80 vss 0.056f
C7679 d1.n41 vss 0.425f
C7680 d1.n42 vss 1.07f
C7681 d1.t35 vss 0.0343f
C7682 d1.t108 vss 0.056f
C7683 d1.n43 vss 0.42f
C7684 d1.n44 vss 0.651f
C7685 d1.t103 vss 0.056f
C7686 d1.t48 vss 0.0343f
C7687 d1.n45 vss 0.425f
C7688 d1.n46 vss 0.535f
C7689 d1.t54 vss 0.056f
C7690 d1.t3 vss 0.0343f
C7691 d1.n47 vss 0.425f
C7692 d1.n48 vss 0.0262f
C7693 d1.n49 vss 1.07f
C7694 d1.t69 vss 0.056f
C7695 d1.t115 vss 0.0343f
C7696 d1.n50 vss 0.425f
C7697 d1.n51 vss 0.0262f
C7698 d1.n52 vss 1.01f
C7699 d1.t61 vss 0.056f
C7700 d1.t5 vss 0.0343f
C7701 d1.n53 vss 0.425f
C7702 d1.n54 vss 0.0262f
C7703 d1.n55 vss 0.997f
C7704 d1.t9 vss 0.056f
C7705 d1.t88 vss 0.0343f
C7706 d1.n56 vss 0.425f
C7707 d1.n57 vss 0.0262f
C7708 d1.n58 vss 0.997f
C7709 d1.t27 vss 0.056f
C7710 d1.t110 vss 0.0343f
C7711 d1.n59 vss 0.425f
C7712 d1.n60 vss 0.0262f
C7713 d1.n61 vss 1.07f
C7714 d1.t105 vss 0.056f
C7715 d1.t60 vss 0.0343f
C7716 d1.n62 vss 0.425f
C7717 d1.n63 vss 0.0262f
C7718 d1.n64 vss 1.01f
C7719 d1.t124 vss 0.056f
C7720 d1.t67 vss 0.0343f
C7721 d1.n65 vss 0.425f
C7722 d1.n66 vss 0.0262f
C7723 d1.n67 vss 1.42f
C7724 d1.n68 vss 3.26f
C7725 d1.t89 vss 0.0343f
C7726 d1.t52 vss 0.056f
C7727 d1.n69 vss 0.425f
C7728 d1.t38 vss 0.0343f
C7729 d1.t1 vss 0.056f
C7730 d1.n70 vss 0.42f
C7731 d1.n71 vss 1.01f
C7732 d1.t65 vss 0.0343f
C7733 d1.t23 vss 0.056f
C7734 d1.n72 vss 0.425f
C7735 d1.n73 vss 1.07f
C7736 d1.t114 vss 0.0343f
C7737 d1.t47 vss 0.056f
C7738 d1.n74 vss 0.42f
C7739 d1.n75 vss 0.997f
C7740 d1.t22 vss 0.0343f
C7741 d1.t91 vss 0.056f
C7742 d1.n76 vss 0.425f
C7743 d1.n77 vss 0.997f
C7744 d1.t46 vss 0.0343f
C7745 d1.t111 vss 0.056f
C7746 d1.n78 vss 0.42f
C7747 d1.n79 vss 1.01f
C7748 d1.t123 vss 0.0343f
C7749 d1.t58 vss 0.056f
C7750 d1.n80 vss 0.425f
C7751 d1.n81 vss 1.07f
C7752 d1.t13 vss 0.0343f
C7753 d1.t82 vss 0.056f
C7754 d1.n82 vss 0.42f
C7755 d1.n83 vss 0.651f
C7756 d1.t126 vss 0.056f
C7757 d1.t68 vss 0.0343f
C7758 d1.n84 vss 0.425f
C7759 d1.n85 vss 0.535f
C7760 d1.t73 vss 0.056f
C7761 d1.t24 vss 0.0343f
C7762 d1.n86 vss 0.425f
C7763 d1.n87 vss 0.0262f
C7764 d1.n88 vss 1.07f
C7765 d1.t95 vss 0.056f
C7766 d1.t7 vss 0.0343f
C7767 d1.n89 vss 0.425f
C7768 d1.n90 vss 0.0262f
C7769 d1.n91 vss 1.01f
C7770 d1.t83 vss 0.056f
C7771 d1.t25 vss 0.0343f
C7772 d1.n92 vss 0.425f
C7773 d1.n93 vss 0.0262f
C7774 d1.n94 vss 0.997f
C7775 d1.t30 vss 0.056f
C7776 d1.t112 vss 0.0343f
C7777 d1.n95 vss 0.425f
C7778 d1.n96 vss 0.0262f
C7779 d1.n97 vss 0.997f
C7780 d1.t56 vss 0.056f
C7781 d1.t0 vss 0.0343f
C7782 d1.n98 vss 0.425f
C7783 d1.n99 vss 0.0262f
C7784 d1.n100 vss 1.07f
C7785 d1.t98 vss 0.056f
C7786 d1.t51 vss 0.0343f
C7787 d1.n101 vss 0.425f
C7788 d1.n102 vss 0.0262f
C7789 d1.n103 vss 1.01f
C7790 d1.t116 vss 0.056f
C7791 d1.t64 vss 0.0343f
C7792 d1.n104 vss 0.425f
C7793 d1.n105 vss 0.0262f
C7794 d1.n106 vss 1.42f
C7795 d1.n107 vss 1.32f
C7796 d1.n108 vss 4.36f
C7797 d1.t96 vss 0.0343f
C7798 d1.t62 vss 0.056f
C7799 d1.n109 vss 0.425f
C7800 d1.t45 vss 0.0343f
C7801 d1.t10 vss 0.056f
C7802 d1.n110 vss 0.42f
C7803 d1.n111 vss 1.01f
C7804 d1.t70 vss 0.0343f
C7805 d1.t37 vss 0.056f
C7806 d1.n112 vss 0.425f
C7807 d1.n113 vss 1.07f
C7808 d1.t125 vss 0.0343f
C7809 d1.t59 vss 0.056f
C7810 d1.n114 vss 0.42f
C7811 d1.n115 vss 0.997f
C7812 d1.t32 vss 0.0343f
C7813 d1.t100 vss 0.056f
C7814 d1.n116 vss 0.425f
C7815 d1.n117 vss 0.997f
C7816 d1.t57 vss 0.0343f
C7817 d1.t117 vss 0.056f
C7818 d1.n118 vss 0.42f
C7819 d1.n119 vss 1.01f
C7820 d1.t28 vss 0.0343f
C7821 d1.t93 vss 0.056f
C7822 d1.n120 vss 0.425f
C7823 d1.n121 vss 1.07f
C7824 d1.t50 vss 0.0343f
C7825 d1.t118 vss 0.056f
C7826 d1.n122 vss 0.42f
C7827 d1.n123 vss 0.651f
C7828 d1.t4 vss 0.056f
C7829 d1.t84 vss 0.0343f
C7830 d1.n124 vss 0.425f
C7831 d1.n125 vss 0.535f
C7832 d1.t86 vss 0.056f
C7833 d1.t41 vss 0.0343f
C7834 d1.n126 vss 0.425f
C7835 d1.n127 vss 0.0262f
C7836 d1.n128 vss 1.07f
C7837 d1.t109 vss 0.056f
C7838 d1.t19 vss 0.0343f
C7839 d1.n129 vss 0.425f
C7840 d1.n130 vss 0.0262f
C7841 d1.n131 vss 1.01f
C7842 d1.t94 vss 0.056f
C7843 d1.t42 vss 0.0343f
C7844 d1.n132 vss 0.425f
C7845 d1.n133 vss 0.0262f
C7846 d1.n134 vss 0.997f
C7847 d1.t43 vss 0.056f
C7848 d1.t121 vss 0.0343f
C7849 d1.n135 vss 0.425f
C7850 d1.n136 vss 0.0262f
C7851 d1.n137 vss 0.997f
C7852 d1.t66 vss 0.056f
C7853 d1.t12 vss 0.0343f
C7854 d1.n138 vss 0.425f
C7855 d1.n139 vss 0.0262f
C7856 d1.n140 vss 1.07f
C7857 d1.t71 vss 0.056f
C7858 d1.t21 vss 0.0343f
C7859 d1.n141 vss 0.425f
C7860 d1.n142 vss 0.0262f
C7861 d1.n143 vss 1.01f
C7862 d1.t92 vss 0.056f
C7863 d1.t39 vss 0.0343f
C7864 d1.n144 vss 0.425f
C7865 d1.n145 vss 0.0262f
C7866 d1.n146 vss 1.42f
C7867 d1.n147 vss 1.32f
C7868 d1.n148 vss 4.36f
C7869 d1.n149 vss 3.26f
C7870 d1.n150 vss 1.42f
C7871 d1.n151 vss 1.01f
C7872 d1.n152 vss 1.07f
C7873 d1.n153 vss 0.997f
C7874 d1.n154 vss 0.997f
C7875 d1.n155 vss 1.01f
C7876 d1.n156 vss 1.07f
C7877 d1.n157 vss 0.0262f
C7878 d0.t245 vss 0.0286f
C7879 d0.t124 vss 0.0175f
C7880 d0.n0 vss 0.217f
C7881 d0.t135 vss 0.0286f
C7882 d0.t28 vss 0.0175f
C7883 d0.n1 vss 0.217f
C7884 d0.n2 vss 0.0134f
C7885 d0.t174 vss 0.0286f
C7886 d0.t81 vss 0.0175f
C7887 d0.n3 vss 0.217f
C7888 d0.n4 vss 0.0134f
C7889 d0.t216 vss 0.0286f
C7890 d0.t119 vss 0.0175f
C7891 d0.n5 vss 0.217f
C7892 d0.n6 vss 0.0134f
C7893 d0.t125 vss 0.0286f
C7894 d0.t21 vss 0.0175f
C7895 d0.n7 vss 0.217f
C7896 d0.n8 vss 0.0134f
C7897 d0.t165 vss 0.0286f
C7898 d0.t238 vss 0.0175f
C7899 d0.n9 vss 0.217f
C7900 d0.n10 vss 0.0134f
C7901 d0.t128 vss 0.0286f
C7902 d0.t136 vss 0.0175f
C7903 d0.n11 vss 0.217f
C7904 d0.n12 vss 0.0134f
C7905 d0.t15 vss 0.0286f
C7906 d0.t186 vss 0.0175f
C7907 d0.n13 vss 0.217f
C7908 d0.n14 vss 0.0134f
C7909 d0.t87 vss 0.0175f
C7910 d0.t9 vss 0.0286f
C7911 d0.n15 vss 0.217f
C7912 d0.t11 vss 0.0175f
C7913 d0.t200 vss 0.0286f
C7914 d0.n16 vss 0.217f
C7915 d0.n17 vss 0.46f
C7916 d0.t242 vss 0.0175f
C7917 d0.t176 vss 0.0286f
C7918 d0.n18 vss 0.214f
C7919 d0.n19 vss 0.459f
C7920 d0.t100 vss 0.0175f
C7921 d0.t38 vss 0.0286f
C7922 d0.n20 vss 0.217f
C7923 d0.n21 vss 0.457f
C7924 d0.t39 vss 0.0175f
C7925 d0.t218 vss 0.0286f
C7926 d0.n22 vss 0.217f
C7927 d0.n23 vss 0.459f
C7928 d0.t206 vss 0.0175f
C7929 d0.t77 vss 0.0286f
C7930 d0.n24 vss 0.217f
C7931 d0.n25 vss 0.457f
C7932 d0.t143 vss 0.0175f
C7933 d0.t6 vss 0.0286f
C7934 d0.n26 vss 0.214f
C7935 d0.n27 vss 0.459f
C7936 d0.t249 vss 0.0175f
C7937 d0.t233 vss 0.0286f
C7938 d0.n28 vss 0.217f
C7939 d0.n29 vss 0.457f
C7940 d0.t215 vss 0.0175f
C7941 d0.t92 vss 0.0286f
C7942 d0.n30 vss 0.217f
C7943 d0.n31 vss 0.459f
C7944 d0.t156 vss 0.0175f
C7945 d0.t17 vss 0.0286f
C7946 d0.n32 vss 0.217f
C7947 d0.n33 vss 0.457f
C7948 d0.t2 vss 0.0175f
C7949 d0.t129 vss 0.0286f
C7950 d0.n34 vss 0.214f
C7951 d0.n35 vss 0.459f
C7952 d0.t195 vss 0.0175f
C7953 d0.t63 vss 0.0286f
C7954 d0.n36 vss 0.217f
C7955 d0.n37 vss 0.457f
C7956 d0.t43 vss 0.0175f
C7957 d0.t229 vss 0.0286f
C7958 d0.n38 vss 0.217f
C7959 d0.n39 vss 0.459f
C7960 d0.t214 vss 0.0175f
C7961 d0.t107 vss 0.0286f
C7962 d0.n40 vss 0.217f
C7963 d0.n41 vss 0.457f
C7964 d0.t154 vss 0.0175f
C7965 d0.t33 vss 0.0286f
C7966 d0.n42 vss 0.214f
C7967 d0.n43 vss 0.459f
C7968 d0.t13 vss 0.0175f
C7969 d0.t146 vss 0.0286f
C7970 d0.n44 vss 0.214f
C7971 d0.n45 vss 1.26f
C7972 d0.t105 vss 0.0286f
C7973 d0.t232 vss 0.0175f
C7974 d0.n46 vss 0.217f
C7975 d0.n47 vss 0.143f
C7976 d0.t10 vss 0.0286f
C7977 d0.t168 vss 0.0175f
C7978 d0.n48 vss 0.217f
C7979 d0.n49 vss 0.0134f
C7980 d0.n50 vss 0.459f
C7981 d0.t243 vss 0.0286f
C7982 d0.t142 vss 0.0175f
C7983 d0.n51 vss 0.217f
C7984 d0.n52 vss 0.0134f
C7985 d0.n53 vss 0.457f
C7986 d0.t177 vss 0.0286f
C7987 d0.t82 vss 0.0175f
C7988 d0.n54 vss 0.217f
C7989 d0.n55 vss 0.0134f
C7990 d0.n56 vss 0.459f
C7991 d0.t26 vss 0.0286f
C7992 d0.t194 vss 0.0175f
C7993 d0.n57 vss 0.217f
C7994 d0.n58 vss 0.0134f
C7995 d0.n59 vss 0.457f
C7996 d0.t211 vss 0.0286f
C7997 d0.t44 vss 0.0175f
C7998 d0.n60 vss 0.217f
C7999 d0.n61 vss 0.0134f
C8000 d0.n62 vss 0.459f
C8001 d0.t79 vss 0.0286f
C8002 d0.t221 vss 0.0175f
C8003 d0.n63 vss 0.217f
C8004 d0.n64 vss 0.0134f
C8005 d0.n65 vss 0.457f
C8006 d0.t191 vss 0.0286f
C8007 d0.t203 vss 0.0175f
C8008 d0.n66 vss 0.217f
C8009 d0.n67 vss 0.0134f
C8010 d0.n68 vss 0.459f
C8011 d0.t234 vss 0.0286f
C8012 d0.t137 vss 0.0175f
C8013 d0.n69 vss 0.217f
C8014 d0.n70 vss 0.0134f
C8015 d0.n71 vss 0.457f
C8016 d0.t93 vss 0.0286f
C8017 d0.t241 vss 0.0175f
C8018 d0.n72 vss 0.217f
C8019 d0.n73 vss 0.0134f
C8020 d0.n74 vss 0.459f
C8021 d0.t18 vss 0.0286f
C8022 d0.t99 vss 0.0175f
C8023 d0.n75 vss 0.217f
C8024 d0.n76 vss 0.0134f
C8025 d0.n77 vss 0.457f
C8026 d0.t131 vss 0.0286f
C8027 d0.t23 vss 0.0175f
C8028 d0.n78 vss 0.217f
C8029 d0.n79 vss 0.0134f
C8030 d0.n80 vss 0.459f
C8031 d0.t236 vss 0.0286f
C8032 d0.t101 vss 0.0175f
C8033 d0.n81 vss 0.217f
C8034 d0.n82 vss 0.0134f
C8035 d0.n83 vss 0.457f
C8036 d0.t134 vss 0.0286f
C8037 d0.t40 vss 0.0175f
C8038 d0.n84 vss 0.217f
C8039 d0.n85 vss 0.0134f
C8040 d0.n86 vss 0.459f
C8041 d0.t239 vss 0.0286f
C8042 d0.t152 vss 0.0175f
C8043 d0.n87 vss 0.217f
C8044 d0.n88 vss 0.0134f
C8045 d0.n89 vss 0.457f
C8046 d0.t173 vss 0.0286f
C8047 d0.t67 vss 0.0175f
C8048 d0.n90 vss 0.217f
C8049 d0.n91 vss 0.0134f
C8050 d0.n92 vss 0.358f
C8051 d0.n93 vss 1.44f
C8052 d0.t192 vss 0.0175f
C8053 d0.t117 vss 0.0286f
C8054 d0.n94 vss 0.217f
C8055 d0.t118 vss 0.0175f
C8056 d0.t49 vss 0.0286f
C8057 d0.n95 vss 0.217f
C8058 d0.n96 vss 0.46f
C8059 d0.t94 vss 0.0175f
C8060 d0.t20 vss 0.0286f
C8061 d0.n97 vss 0.214f
C8062 d0.n98 vss 0.459f
C8063 d0.t201 vss 0.0175f
C8064 d0.t147 vss 0.0286f
C8065 d0.n99 vss 0.217f
C8066 d0.n100 vss 0.457f
C8067 d0.t148 vss 0.0175f
C8068 d0.t74 vss 0.0286f
C8069 d0.n101 vss 0.217f
C8070 d0.n102 vss 0.459f
C8071 d0.t61 vss 0.0175f
C8072 d0.t185 vss 0.0286f
C8073 d0.n103 vss 0.217f
C8074 d0.n104 vss 0.457f
C8075 d0.t244 vss 0.0175f
C8076 d0.t112 vss 0.0286f
C8077 d0.n105 vss 0.214f
C8078 d0.n106 vss 0.459f
C8079 d0.t102 vss 0.0175f
C8080 d0.t85 vss 0.0286f
C8081 d0.n107 vss 0.217f
C8082 d0.n108 vss 0.457f
C8083 d0.t70 vss 0.0175f
C8084 d0.t198 vss 0.0286f
C8085 d0.n109 vss 0.217f
C8086 d0.n110 vss 0.459f
C8087 d0.t252 vss 0.0175f
C8088 d0.t121 vss 0.0286f
C8089 d0.n111 vss 0.217f
C8090 d0.n112 vss 0.457f
C8091 d0.t110 vss 0.0175f
C8092 d0.t225 vss 0.0286f
C8093 d0.n113 vss 0.214f
C8094 d0.n114 vss 0.459f
C8095 d0.t37 vss 0.0175f
C8096 d0.t163 vss 0.0286f
C8097 d0.n115 vss 0.217f
C8098 d0.n116 vss 0.457f
C8099 d0.t151 vss 0.0175f
C8100 d0.t246 vss 0.0286f
C8101 d0.n117 vss 0.217f
C8102 d0.n118 vss 0.459f
C8103 d0.t224 vss 0.0175f
C8104 d0.t113 vss 0.0286f
C8105 d0.n119 vss 0.217f
C8106 d0.n120 vss 0.457f
C8107 d0.t162 vss 0.0175f
C8108 d0.t41 vss 0.0286f
C8109 d0.n121 vss 0.214f
C8110 d0.n122 vss 0.459f
C8111 d0.t30 vss 0.0175f
C8112 d0.t155 vss 0.0286f
C8113 d0.n123 vss 0.214f
C8114 d0.n124 vss 0.363f
C8115 d0.n125 vss 1.22f
C8116 d0.t149 vss 0.0286f
C8117 d0.t24 vss 0.0175f
C8118 d0.n126 vss 0.217f
C8119 d0.n127 vss 0.142f
C8120 d0.t65 vss 0.0286f
C8121 d0.t209 vss 0.0175f
C8122 d0.n128 vss 0.217f
C8123 d0.n129 vss 0.0134f
C8124 d0.n130 vss 0.459f
C8125 d0.t35 vss 0.0286f
C8126 d0.t187 vss 0.0175f
C8127 d0.n131 vss 0.217f
C8128 d0.n132 vss 0.0134f
C8129 d0.n133 vss 0.457f
C8130 d0.t213 vss 0.0286f
C8131 d0.t127 vss 0.0175f
C8132 d0.n134 vss 0.217f
C8133 d0.n135 vss 0.0134f
C8134 d0.n136 vss 0.459f
C8135 d0.t73 vss 0.0286f
C8136 d0.t231 vss 0.0175f
C8137 d0.n137 vss 0.217f
C8138 d0.n138 vss 0.0134f
C8139 d0.n139 vss 0.457f
C8140 d0.t255 vss 0.0286f
C8141 d0.t91 vss 0.0175f
C8142 d0.n140 vss 0.217f
C8143 d0.n141 vss 0.0134f
C8144 d0.n142 vss 0.459f
C8145 d0.t122 vss 0.0286f
C8146 d0.t16 vss 0.0175f
C8147 d0.n143 vss 0.217f
C8148 d0.n144 vss 0.0134f
C8149 d0.n145 vss 0.457f
C8150 d0.t226 vss 0.0286f
C8151 d0.t247 vss 0.0175f
C8152 d0.n146 vss 0.217f
C8153 d0.n147 vss 0.0134f
C8154 d0.n148 vss 0.459f
C8155 d0.t25 vss 0.0286f
C8156 d0.t180 vss 0.0175f
C8157 d0.n149 vss 0.217f
C8158 d0.n150 vss 0.0134f
C8159 d0.n151 vss 0.457f
C8160 d0.t138 vss 0.0286f
C8161 d0.t32 vss 0.0175f
C8162 d0.n152 vss 0.217f
C8163 d0.n153 vss 0.0134f
C8164 d0.n154 vss 0.459f
C8165 d0.t68 vss 0.0286f
C8166 d0.t145 vss 0.0175f
C8167 d0.n155 vss 0.217f
C8168 d0.n156 vss 0.0134f
C8169 d0.n157 vss 0.457f
C8170 d0.t178 vss 0.0286f
C8171 d0.t71 vss 0.0175f
C8172 d0.n158 vss 0.217f
C8173 d0.n159 vss 0.0134f
C8174 d0.n160 vss 0.459f
C8175 d0.t31 vss 0.0286f
C8176 d0.t86 vss 0.0175f
C8177 d0.n161 vss 0.217f
C8178 d0.n162 vss 0.0134f
C8179 d0.n163 vss 0.457f
C8180 d0.t120 vss 0.0286f
C8181 d0.t29 vss 0.0175f
C8182 d0.n164 vss 0.217f
C8183 d0.n165 vss 0.0134f
C8184 d0.n166 vss 0.459f
C8185 d0.t220 vss 0.0286f
C8186 d0.t140 vss 0.0175f
C8187 d0.n167 vss 0.217f
C8188 d0.n168 vss 0.0134f
C8189 d0.n169 vss 0.457f
C8190 d0.t158 vss 0.0286f
C8191 d0.t53 vss 0.0175f
C8192 d0.n170 vss 0.217f
C8193 d0.n171 vss 0.0134f
C8194 d0.n172 vss 0.358f
C8195 d0.n173 vss 1.21f
C8196 d0.t123 vss 0.0175f
C8197 d0.t55 vss 0.0286f
C8198 d0.n174 vss 0.217f
C8199 d0.t56 vss 0.0175f
C8200 d0.t237 vss 0.0286f
C8201 d0.n175 vss 0.217f
C8202 d0.n176 vss 0.46f
C8203 d0.t27 vss 0.0175f
C8204 d0.t210 vss 0.0286f
C8205 d0.n177 vss 0.214f
C8206 d0.n178 vss 0.459f
C8207 d0.t139 vss 0.0175f
C8208 d0.t78 vss 0.0286f
C8209 d0.n179 vss 0.217f
C8210 d0.n180 vss 0.457f
C8211 d0.t80 vss 0.0175f
C8212 d0.t7 vss 0.0286f
C8213 d0.n181 vss 0.217f
C8214 d0.n182 vss 0.459f
C8215 d0.t250 vss 0.0175f
C8216 d0.t116 vss 0.0286f
C8217 d0.n183 vss 0.217f
C8218 d0.n184 vss 0.457f
C8219 d0.t182 vss 0.0175f
C8220 d0.t48 vss 0.0286f
C8221 d0.n185 vss 0.214f
C8222 d0.n186 vss 0.459f
C8223 d0.t34 vss 0.0175f
C8224 d0.t19 vss 0.0286f
C8225 d0.n187 vss 0.217f
C8226 d0.n188 vss 0.457f
C8227 d0.t3 vss 0.0175f
C8228 d0.t132 vss 0.0286f
C8229 d0.n189 vss 0.217f
C8230 d0.n190 vss 0.459f
C8231 d0.t196 vss 0.0175f
C8232 d0.t64 vss 0.0286f
C8233 d0.n191 vss 0.217f
C8234 d0.n192 vss 0.457f
C8235 d0.t46 vss 0.0175f
C8236 d0.t171 vss 0.0286f
C8237 d0.n193 vss 0.214f
C8238 d0.n194 vss 0.459f
C8239 d0.t222 vss 0.0175f
C8240 d0.t103 vss 0.0286f
C8241 d0.n195 vss 0.217f
C8242 d0.n196 vss 0.457f
C8243 d0.t84 vss 0.0175f
C8244 d0.t5 vss 0.0286f
C8245 d0.n197 vss 0.217f
C8246 d0.n198 vss 0.459f
C8247 d0.t248 vss 0.0175f
C8248 d0.t130 vss 0.0286f
C8249 d0.n199 vss 0.217f
C8250 d0.n200 vss 0.457f
C8251 d0.t181 vss 0.0175f
C8252 d0.t62 vss 0.0286f
C8253 d0.n201 vss 0.214f
C8254 d0.n202 vss 0.459f
C8255 d0.t45 vss 0.0175f
C8256 d0.t170 vss 0.0286f
C8257 d0.n203 vss 0.214f
C8258 d0.n204 vss 0.363f
C8259 d0.n205 vss 1.22f
C8260 d0.t169 vss 0.0286f
C8261 d0.t50 vss 0.0175f
C8262 d0.n206 vss 0.217f
C8263 d0.n207 vss 0.143f
C8264 d0.t83 vss 0.0286f
C8265 d0.t227 vss 0.0175f
C8266 d0.n208 vss 0.217f
C8267 d0.n209 vss 0.0134f
C8268 d0.n210 vss 0.459f
C8269 d0.t59 vss 0.0286f
C8270 d0.t205 vss 0.0175f
C8271 d0.n211 vss 0.217f
C8272 d0.n212 vss 0.0134f
C8273 d0.n213 vss 0.457f
C8274 d0.t240 vss 0.0286f
C8275 d0.t153 vss 0.0175f
C8276 d0.n214 vss 0.217f
C8277 d0.n215 vss 0.0134f
C8278 d0.n216 vss 0.459f
C8279 d0.t98 vss 0.0286f
C8280 d0.t0 vss 0.0175f
C8281 d0.n217 vss 0.217f
C8282 d0.n218 vss 0.0134f
C8283 d0.n219 vss 0.457f
C8284 d0.t22 vss 0.0286f
C8285 d0.t114 vss 0.0175f
C8286 d0.n220 vss 0.217f
C8287 d0.n221 vss 0.0134f
C8288 d0.n222 vss 0.459f
C8289 d0.t150 vss 0.0286f
C8290 d0.t42 vss 0.0175f
C8291 d0.n223 vss 0.217f
C8292 d0.n224 vss 0.0134f
C8293 d0.n225 vss 0.457f
C8294 d0.t253 vss 0.0286f
C8295 d0.t12 vss 0.0175f
C8296 d0.n226 vss 0.217f
C8297 d0.n227 vss 0.0134f
C8298 d0.n228 vss 0.459f
C8299 d0.t51 vss 0.0286f
C8300 d0.t202 vss 0.0175f
C8301 d0.n229 vss 0.217f
C8302 d0.n230 vss 0.0134f
C8303 d0.n231 vss 0.457f
C8304 d0.t159 vss 0.0286f
C8305 d0.t57 vss 0.0175f
C8306 d0.n232 vss 0.217f
C8307 d0.n233 vss 0.0134f
C8308 d0.n234 vss 0.459f
C8309 d0.t88 vss 0.0286f
C8310 d0.t164 vss 0.0175f
C8311 d0.n235 vss 0.217f
C8312 d0.n236 vss 0.0134f
C8313 d0.n237 vss 0.457f
C8314 d0.t199 vss 0.0286f
C8315 d0.t97 vss 0.0175f
C8316 d0.n238 vss 0.217f
C8317 d0.n239 vss 0.0134f
C8318 d0.n240 vss 0.459f
C8319 d0.t52 vss 0.0286f
C8320 d0.t36 vss 0.0175f
C8321 d0.n241 vss 0.217f
C8322 d0.n242 vss 0.0134f
C8323 d0.n243 vss 0.457f
C8324 d0.t72 vss 0.0286f
C8325 d0.t230 vss 0.0175f
C8326 d0.n244 vss 0.217f
C8327 d0.n245 vss 0.0134f
C8328 d0.n246 vss 0.459f
C8329 d0.t184 vss 0.0286f
C8330 d0.t90 vss 0.0175f
C8331 d0.n247 vss 0.217f
C8332 d0.n248 vss 0.0134f
C8333 d0.n249 vss 0.457f
C8334 d0.t111 vss 0.0286f
C8335 d0.t1 vss 0.0175f
C8336 d0.n250 vss 0.217f
C8337 d0.n251 vss 0.0134f
C8338 d0.n252 vss 0.358f
C8339 d0.n253 vss 1.21f
C8340 d0.t254 vss 0.0175f
C8341 d0.t188 vss 0.0286f
C8342 d0.n254 vss 0.217f
C8343 d0.t189 vss 0.0175f
C8344 d0.t115 vss 0.0286f
C8345 d0.n255 vss 0.217f
C8346 d0.n256 vss 0.46f
C8347 d0.t161 vss 0.0175f
C8348 d0.t89 vss 0.0286f
C8349 d0.n257 vss 0.214f
C8350 d0.n258 vss 0.459f
C8351 d0.t8 vss 0.0175f
C8352 d0.t207 vss 0.0286f
C8353 d0.n259 vss 0.217f
C8354 d0.n260 vss 0.457f
C8355 d0.t208 vss 0.0175f
C8356 d0.t144 vss 0.0286f
C8357 d0.n261 vss 0.217f
C8358 d0.n262 vss 0.459f
C8359 d0.t126 vss 0.0175f
C8360 d0.t251 vss 0.0286f
C8361 d0.n263 vss 0.217f
C8362 d0.n264 vss 0.457f
C8363 d0.t60 vss 0.0175f
C8364 d0.t183 vss 0.0286f
C8365 d0.n265 vss 0.214f
C8366 d0.n266 vss 0.459f
C8367 d0.t166 vss 0.0175f
C8368 d0.t157 vss 0.0286f
C8369 d0.n267 vss 0.217f
C8370 d0.n268 vss 0.457f
C8371 d0.t141 vss 0.0175f
C8372 d0.t4 vss 0.0286f
C8373 d0.n269 vss 0.217f
C8374 d0.n270 vss 0.459f
C8375 d0.t69 vss 0.0175f
C8376 d0.t197 vss 0.0286f
C8377 d0.n271 vss 0.217f
C8378 d0.n272 vss 0.457f
C8379 d0.t179 vss 0.0175f
C8380 d0.t47 vss 0.0286f
C8381 d0.n273 vss 0.214f
C8382 d0.n274 vss 0.459f
C8383 d0.t109 vss 0.0175f
C8384 d0.t223 vss 0.0286f
C8385 d0.n275 vss 0.217f
C8386 d0.n276 vss 0.457f
C8387 d0.t212 vss 0.0175f
C8388 d0.t190 vss 0.0286f
C8389 d0.n277 vss 0.217f
C8390 d0.n278 vss 0.459f
C8391 d0.t175 vss 0.0175f
C8392 d0.t54 vss 0.0286f
C8393 d0.n279 vss 0.217f
C8394 d0.n280 vss 0.457f
C8395 d0.t108 vss 0.0175f
C8396 d0.t235 vss 0.0286f
C8397 d0.n281 vss 0.214f
C8398 d0.n282 vss 0.459f
C8399 d0.t217 vss 0.0175f
C8400 d0.t96 vss 0.0286f
C8401 d0.n283 vss 0.214f
C8402 d0.n284 vss 0.363f
C8403 d0.n285 vss 1.45f
C8404 d0.t204 vss 0.0286f
C8405 d0.t104 vss 0.0175f
C8406 d0.n286 vss 0.217f
C8407 d0.n287 vss 0.0134f
C8408 d0.n288 vss 1.25f
C8409 d0.n289 vss 0.457f
C8410 d0.t167 vss 0.0286f
C8411 d0.t75 vss 0.0175f
C8412 d0.n290 vss 0.217f
C8413 d0.n291 vss 0.0134f
C8414 d0.n292 vss 0.459f
C8415 d0.n293 vss 0.457f
C8416 d0.t14 vss 0.0286f
C8417 d0.t172 vss 0.0175f
C8418 d0.n294 vss 0.217f
C8419 d0.n295 vss 0.0134f
C8420 d0.n296 vss 0.459f
C8421 d0.n297 vss 0.457f
C8422 d0.t228 vss 0.0286f
C8423 d0.t133 vss 0.0175f
C8424 d0.n298 vss 0.217f
C8425 d0.n299 vss 0.0134f
C8426 d0.n300 vss 0.459f
C8427 d0.n301 vss 0.457f
C8428 d0.t76 vss 0.0286f
C8429 d0.t95 vss 0.0175f
C8430 d0.n302 vss 0.217f
C8431 d0.n303 vss 0.0134f
C8432 d0.n304 vss 0.459f
C8433 d0.n305 vss 0.457f
C8434 d0.t106 vss 0.0286f
C8435 d0.t193 vss 0.0175f
C8436 d0.n306 vss 0.217f
C8437 d0.n307 vss 0.0134f
C8438 d0.n308 vss 0.459f
C8439 d0.n309 vss 0.457f
C8440 d0.t66 vss 0.0286f
C8441 d0.t219 vss 0.0175f
C8442 d0.n310 vss 0.217f
C8443 d0.n311 vss 0.0134f
C8444 d0.n312 vss 0.459f
C8445 d0.n313 vss 0.457f
C8446 d0.t160 vss 0.0286f
C8447 d0.t58 vss 0.0175f
C8448 d0.n314 vss 0.217f
C8449 d0.n315 vss 0.0134f
C8450 d0.n316 vss 0.459f
C8451 d0.n317 vss 0.142f
C8452 X2.X2.X3.vin1.t0 vss 0.00514f
C8453 X2.X2.X3.vin1.t1 vss 0.179f
C8454 X2.X2.X3.vin1.t2 vss 0.00574f
C8455 X2.X2.X3.vin1.t3 vss 0.00501f
C8456 X2.X2.X3.vin1.n0 vss 1.42f
C8457 vdd.t1009 vss 0.0013f
C8458 vdd.t244 vss 0.00134f
C8459 vdd.n0 vss 0.00324f
C8460 vdd.n1 vss 0.0112f
C8461 vdd.n2 vss 0.0128f
C8462 vdd.n3 vss 0.00413f
C8463 vdd.n4 vss 0.00413f
C8464 vdd.n5 vss 0.0471f
C8465 vdd.n6 vss 0.00251f
C8466 vdd.t839 vss 0.0471f
C8467 vdd.n7 vss 0.00324f
C8468 vdd.n9 vss 0.00679f
C8469 vdd.n10 vss 0.00413f
C8470 vdd.n11 vss 0.00324f
C8471 vdd.n12 vss 0.00413f
C8472 vdd.n13 vss 0.0471f
C8473 vdd.n14 vss 0.00324f
C8474 vdd.n16 vss 0.00925f
C8475 vdd.t260 vss 0.0471f
C8476 vdd.n17 vss 0.00425f
C8477 vdd.n18 vss 0.0424f
C8478 vdd.n19 vss 0.0132f
C8479 vdd.n20 vss 0.00324f
C8480 vdd.n21 vss 0.0128f
C8481 vdd.n22 vss 0.02f
C8482 vdd.n23 vss 0.00425f
C8483 vdd.n24 vss 0.00413f
C8484 vdd.n25 vss 0.00251f
C8485 vdd.t653 vss 0.0471f
C8486 vdd.n26 vss 0.00251f
C8487 vdd.n27 vss 0.00517f
C8488 vdd.n28 vss 0.00679f
C8489 vdd.n29 vss 0.00517f
C8490 vdd.n30 vss 0.00679f
C8491 vdd.n31 vss 0.02f
C8492 vdd.n32 vss 0.00425f
C8493 vdd.n33 vss 0.0424f
C8494 vdd.n34 vss 0.0132f
C8495 vdd.n35 vss 0.00925f
C8496 vdd.n36 vss 0.00425f
C8497 vdd.n37 vss 0.00413f
C8498 vdd.n38 vss 0.00324f
C8499 vdd.n39 vss 0.0471f
C8500 vdd.t651 vss 0.0471f
C8501 vdd.n40 vss 0.00251f
C8502 vdd.n41 vss 0.0112f
C8503 vdd.n42 vss 0.0128f
C8504 vdd.t652 vss 0.00134f
C8505 vdd.t840 vss 0.0013f
C8506 vdd.n43 vss 0.0332f
C8507 vdd.n44 vss 0.0393f
C8508 vdd.n45 vss 0.119f
C8509 vdd.n46 vss 0.00324f
C8510 vdd.n47 vss 0.0112f
C8511 vdd.n48 vss 0.0128f
C8512 vdd.n49 vss 0.00413f
C8513 vdd.n50 vss 0.00413f
C8514 vdd.n51 vss 0.0471f
C8515 vdd.n52 vss 0.00251f
C8516 vdd.t1008 vss 0.0471f
C8517 vdd.n53 vss 0.00324f
C8518 vdd.n55 vss 0.00679f
C8519 vdd.n56 vss 0.00413f
C8520 vdd.n57 vss 0.00324f
C8521 vdd.n58 vss 0.00413f
C8522 vdd.n59 vss 0.0471f
C8523 vdd.n60 vss 0.00324f
C8524 vdd.n62 vss 0.00925f
C8525 vdd.t422 vss 0.0471f
C8526 vdd.n63 vss 0.00425f
C8527 vdd.n64 vss 0.0424f
C8528 vdd.n65 vss 0.0132f
C8529 vdd.n66 vss 0.00324f
C8530 vdd.n67 vss 0.0128f
C8531 vdd.n68 vss 0.02f
C8532 vdd.n69 vss 0.00425f
C8533 vdd.n70 vss 0.00413f
C8534 vdd.n71 vss 0.00251f
C8535 vdd.t242 vss 0.0471f
C8536 vdd.n72 vss 0.00251f
C8537 vdd.n73 vss 0.00517f
C8538 vdd.n74 vss 0.00679f
C8539 vdd.n75 vss 0.00517f
C8540 vdd.n76 vss 0.00679f
C8541 vdd.n77 vss 0.02f
C8542 vdd.n78 vss 0.00425f
C8543 vdd.n79 vss 0.0424f
C8544 vdd.n80 vss 0.0132f
C8545 vdd.n81 vss 0.00925f
C8546 vdd.n82 vss 0.00425f
C8547 vdd.n83 vss 0.00413f
C8548 vdd.n84 vss 0.00324f
C8549 vdd.n85 vss 0.0471f
C8550 vdd.t243 vss 0.0471f
C8551 vdd.n86 vss 0.00251f
C8552 vdd.n87 vss 0.0112f
C8553 vdd.n88 vss 0.0128f
C8554 vdd.n89 vss 0.118f
C8555 vdd.n90 vss 0.0393f
C8556 vdd.n91 vss 0.0332f
C8557 vdd.n92 vss 0.0596f
C8558 vdd.t508 vss 0.00134f
C8559 vdd.t1048 vss 0.0013f
C8560 vdd.n93 vss 0.032f
C8561 vdd.n94 vss 0.0393f
C8562 vdd.n95 vss 0.00324f
C8563 vdd.n96 vss 0.0112f
C8564 vdd.n97 vss 0.0128f
C8565 vdd.n98 vss 0.00413f
C8566 vdd.t509 vss 0.0471f
C8567 vdd.n99 vss 0.00324f
C8568 vdd.n101 vss 0.00925f
C8569 vdd.n102 vss 0.00413f
C8570 vdd.n103 vss 0.00679f
C8571 vdd.n104 vss 0.00413f
C8572 vdd.n105 vss 0.0471f
C8573 vdd.n106 vss 0.00324f
C8574 vdd.n107 vss 0.0471f
C8575 vdd.n108 vss 0.00324f
C8576 vdd.n109 vss 0.0424f
C8577 vdd.t1047 vss 0.0471f
C8578 vdd.n111 vss 0.00425f
C8579 vdd.n112 vss 0.00925f
C8580 vdd.n113 vss 0.0132f
C8581 vdd.n114 vss 0.00324f
C8582 vdd.n115 vss 0.0128f
C8583 vdd.n116 vss 0.02f
C8584 vdd.n117 vss 0.00425f
C8585 vdd.n118 vss 0.00413f
C8586 vdd.n119 vss 0.00251f
C8587 vdd.t507 vss 0.0471f
C8588 vdd.n120 vss 0.00251f
C8589 vdd.n121 vss 0.00517f
C8590 vdd.n122 vss 0.00679f
C8591 vdd.n123 vss 0.00324f
C8592 vdd.n124 vss 0.00679f
C8593 vdd.n125 vss 0.00517f
C8594 vdd.n126 vss 0.00251f
C8595 vdd.n127 vss 0.00413f
C8596 vdd.n128 vss 0.0471f
C8597 vdd.t1182 vss 0.0471f
C8598 vdd.n129 vss 0.00425f
C8599 vdd.n130 vss 0.0424f
C8600 vdd.n131 vss 0.0132f
C8601 vdd.n132 vss 0.02f
C8602 vdd.n133 vss 0.00425f
C8603 vdd.n134 vss 0.00413f
C8604 vdd.n135 vss 0.00251f
C8605 vdd.n136 vss 0.0112f
C8606 vdd.n137 vss 0.0128f
C8607 vdd.n138 vss 0.0418f
C8608 vdd.t914 vss 0.00134f
C8609 vdd.t8 vss 0.0013f
C8610 vdd.n139 vss 0.032f
C8611 vdd.n140 vss 0.0393f
C8612 vdd.n141 vss 0.00324f
C8613 vdd.n142 vss 0.0112f
C8614 vdd.n143 vss 0.0128f
C8615 vdd.n144 vss 0.00413f
C8616 vdd.t915 vss 0.0471f
C8617 vdd.n145 vss 0.00324f
C8618 vdd.n147 vss 0.00925f
C8619 vdd.n148 vss 0.00413f
C8620 vdd.n149 vss 0.00679f
C8621 vdd.n150 vss 0.00413f
C8622 vdd.n151 vss 0.0471f
C8623 vdd.n152 vss 0.00324f
C8624 vdd.n153 vss 0.0471f
C8625 vdd.n154 vss 0.00324f
C8626 vdd.n155 vss 0.0424f
C8627 vdd.t7 vss 0.0471f
C8628 vdd.n157 vss 0.00425f
C8629 vdd.n158 vss 0.00925f
C8630 vdd.n159 vss 0.0132f
C8631 vdd.n160 vss 0.00324f
C8632 vdd.n161 vss 0.0128f
C8633 vdd.n162 vss 0.02f
C8634 vdd.n163 vss 0.00425f
C8635 vdd.n164 vss 0.00413f
C8636 vdd.n165 vss 0.00251f
C8637 vdd.t913 vss 0.0471f
C8638 vdd.n166 vss 0.00251f
C8639 vdd.n167 vss 0.00517f
C8640 vdd.n168 vss 0.00679f
C8641 vdd.n169 vss 0.00324f
C8642 vdd.n170 vss 0.00679f
C8643 vdd.n171 vss 0.00517f
C8644 vdd.n172 vss 0.00251f
C8645 vdd.n173 vss 0.00413f
C8646 vdd.n174 vss 0.0471f
C8647 vdd.t977 vss 0.0471f
C8648 vdd.n175 vss 0.00425f
C8649 vdd.n176 vss 0.0424f
C8650 vdd.n177 vss 0.0132f
C8651 vdd.n178 vss 0.02f
C8652 vdd.n179 vss 0.00425f
C8653 vdd.n180 vss 0.00413f
C8654 vdd.n181 vss 0.00251f
C8655 vdd.n182 vss 0.0112f
C8656 vdd.n183 vss 0.0128f
C8657 vdd.n184 vss 0.0369f
C8658 vdd.n185 vss 0.00335f
C8659 vdd.t578 vss 0.0013f
C8660 vdd.n186 vss 0.0309f
C8661 vdd.n187 vss 0.0107f
C8662 vdd.n188 vss 0.0128f
C8663 vdd.n189 vss 0.0424f
C8664 vdd.t577 vss 0.0471f
C8665 vdd.n190 vss 0.00324f
C8666 vdd.n191 vss 0.0471f
C8667 vdd.t141 vss 0.0471f
C8668 vdd.n192 vss 0.00413f
C8669 vdd.n193 vss 0.00324f
C8670 vdd.t142 vss 0.00134f
C8671 vdd.n194 vss 0.0393f
C8672 vdd.n195 vss 0.0128f
C8673 vdd.t140 vss 0.0471f
C8674 vdd.n196 vss 0.00324f
C8675 vdd.n198 vss 0.00925f
C8676 vdd.n199 vss 0.0471f
C8677 vdd.n200 vss 0.00324f
C8678 vdd.n201 vss 0.00413f
C8679 vdd.n202 vss 0.00324f
C8680 vdd.n203 vss 0.00679f
C8681 vdd.n205 vss 0.00925f
C8682 vdd.n206 vss 0.00425f
C8683 vdd.n207 vss 0.00413f
C8684 vdd.n208 vss 0.00251f
C8685 vdd.n209 vss 0.00517f
C8686 vdd.n210 vss 0.00679f
C8687 vdd.n211 vss 0.00324f
C8688 vdd.n212 vss 0.00679f
C8689 vdd.n213 vss 0.00517f
C8690 vdd.n214 vss 0.00251f
C8691 vdd.n215 vss 0.00413f
C8692 vdd.n216 vss 0.0471f
C8693 vdd.t1381 vss 0.0471f
C8694 vdd.n217 vss 0.00425f
C8695 vdd.n218 vss 0.0424f
C8696 vdd.n219 vss 0.0132f
C8697 vdd.n220 vss 0.02f
C8698 vdd.n221 vss 0.00425f
C8699 vdd.n222 vss 0.00413f
C8700 vdd.n223 vss 0.00251f
C8701 vdd.n224 vss 0.0105f
C8702 vdd.n225 vss 0.0633f
C8703 vdd.n226 vss 0.00805f
C8704 vdd.n227 vss 0.0112f
C8705 vdd.n228 vss 0.00251f
C8706 vdd.n229 vss 0.00413f
C8707 vdd.n230 vss 0.00425f
C8708 vdd.n231 vss 0.00991f
C8709 vdd.n232 vss 0.0126f
C8710 vdd.n233 vss 9.89e-19
C8711 vdd.n234 vss 0.0011f
C8712 vdd.n235 vss 0.0271f
C8713 vdd.t737 vss 0.00134f
C8714 vdd.t1476 vss 0.0013f
C8715 vdd.n236 vss 0.032f
C8716 vdd.n237 vss 0.0393f
C8717 vdd.n238 vss 0.00324f
C8718 vdd.n239 vss 0.0112f
C8719 vdd.n240 vss 0.0128f
C8720 vdd.n241 vss 0.00413f
C8721 vdd.t738 vss 0.0471f
C8722 vdd.n242 vss 0.00324f
C8723 vdd.n244 vss 0.00925f
C8724 vdd.n245 vss 0.00413f
C8725 vdd.n246 vss 0.00679f
C8726 vdd.n247 vss 0.00413f
C8727 vdd.n248 vss 0.0471f
C8728 vdd.n249 vss 0.00324f
C8729 vdd.n250 vss 0.0471f
C8730 vdd.n251 vss 0.00324f
C8731 vdd.n252 vss 0.0424f
C8732 vdd.t1475 vss 0.0471f
C8733 vdd.n254 vss 0.00425f
C8734 vdd.n255 vss 0.00925f
C8735 vdd.n256 vss 0.0132f
C8736 vdd.n257 vss 0.00324f
C8737 vdd.n258 vss 0.0128f
C8738 vdd.n259 vss 0.02f
C8739 vdd.n260 vss 0.00425f
C8740 vdd.n261 vss 0.00413f
C8741 vdd.n262 vss 0.00251f
C8742 vdd.t736 vss 0.0471f
C8743 vdd.n263 vss 0.00251f
C8744 vdd.n264 vss 0.00517f
C8745 vdd.n265 vss 0.00679f
C8746 vdd.n266 vss 0.00324f
C8747 vdd.n267 vss 0.00679f
C8748 vdd.n268 vss 0.00517f
C8749 vdd.n269 vss 0.00251f
C8750 vdd.n270 vss 0.00413f
C8751 vdd.n271 vss 0.0471f
C8752 vdd.t527 vss 0.0471f
C8753 vdd.n272 vss 0.00425f
C8754 vdd.n273 vss 0.0424f
C8755 vdd.n274 vss 0.0132f
C8756 vdd.n275 vss 0.02f
C8757 vdd.n276 vss 0.00425f
C8758 vdd.n277 vss 0.00413f
C8759 vdd.n278 vss 0.00251f
C8760 vdd.n279 vss 0.0112f
C8761 vdd.n280 vss 0.0128f
C8762 vdd.n281 vss 0.0418f
C8763 vdd.t162 vss 0.00134f
C8764 vdd.t563 vss 0.0013f
C8765 vdd.n282 vss 0.032f
C8766 vdd.n283 vss 0.0393f
C8767 vdd.n284 vss 0.00324f
C8768 vdd.n285 vss 0.0112f
C8769 vdd.n286 vss 0.0128f
C8770 vdd.n287 vss 0.00413f
C8771 vdd.t163 vss 0.0471f
C8772 vdd.n288 vss 0.00324f
C8773 vdd.n290 vss 0.00925f
C8774 vdd.n291 vss 0.00413f
C8775 vdd.n292 vss 0.00679f
C8776 vdd.n293 vss 0.00413f
C8777 vdd.n294 vss 0.0471f
C8778 vdd.n295 vss 0.00324f
C8779 vdd.n296 vss 0.0471f
C8780 vdd.n297 vss 0.00324f
C8781 vdd.n298 vss 0.0424f
C8782 vdd.t562 vss 0.0471f
C8783 vdd.n300 vss 0.00425f
C8784 vdd.n301 vss 0.00925f
C8785 vdd.n302 vss 0.0132f
C8786 vdd.n303 vss 0.00324f
C8787 vdd.n304 vss 0.0128f
C8788 vdd.n305 vss 0.02f
C8789 vdd.n306 vss 0.00425f
C8790 vdd.n307 vss 0.00413f
C8791 vdd.n308 vss 0.00251f
C8792 vdd.t161 vss 0.0471f
C8793 vdd.n309 vss 0.00251f
C8794 vdd.n310 vss 0.00517f
C8795 vdd.n311 vss 0.00679f
C8796 vdd.n312 vss 0.00324f
C8797 vdd.n313 vss 0.00679f
C8798 vdd.n314 vss 0.00517f
C8799 vdd.n315 vss 0.00251f
C8800 vdd.n316 vss 0.00413f
C8801 vdd.n317 vss 0.0471f
C8802 vdd.t1238 vss 0.0471f
C8803 vdd.n318 vss 0.00425f
C8804 vdd.n319 vss 0.0424f
C8805 vdd.n320 vss 0.0132f
C8806 vdd.n321 vss 0.02f
C8807 vdd.n322 vss 0.00425f
C8808 vdd.n323 vss 0.00413f
C8809 vdd.n324 vss 0.00251f
C8810 vdd.n325 vss 0.0112f
C8811 vdd.n326 vss 0.0128f
C8812 vdd.n327 vss 0.0365f
C8813 vdd.t573 vss 0.00134f
C8814 vdd.t1299 vss 0.0013f
C8815 vdd.n328 vss 0.032f
C8816 vdd.n329 vss 0.0393f
C8817 vdd.n330 vss 0.00324f
C8818 vdd.n331 vss 0.0112f
C8819 vdd.n332 vss 0.0128f
C8820 vdd.n333 vss 0.00413f
C8821 vdd.t574 vss 0.0471f
C8822 vdd.n334 vss 0.00324f
C8823 vdd.n336 vss 0.00925f
C8824 vdd.n337 vss 0.00413f
C8825 vdd.n338 vss 0.00679f
C8826 vdd.n339 vss 0.00413f
C8827 vdd.n340 vss 0.0471f
C8828 vdd.n341 vss 0.00324f
C8829 vdd.n342 vss 0.0471f
C8830 vdd.n343 vss 0.00324f
C8831 vdd.n344 vss 0.0424f
C8832 vdd.t1298 vss 0.0471f
C8833 vdd.n346 vss 0.00425f
C8834 vdd.n347 vss 0.00925f
C8835 vdd.n348 vss 0.0132f
C8836 vdd.n349 vss 0.00324f
C8837 vdd.n350 vss 0.0128f
C8838 vdd.n351 vss 0.02f
C8839 vdd.n352 vss 0.00425f
C8840 vdd.n353 vss 0.00413f
C8841 vdd.n354 vss 0.00251f
C8842 vdd.t572 vss 0.0471f
C8843 vdd.n355 vss 0.00251f
C8844 vdd.n356 vss 0.00517f
C8845 vdd.n357 vss 0.00679f
C8846 vdd.n358 vss 0.00324f
C8847 vdd.n359 vss 0.00679f
C8848 vdd.n360 vss 0.00517f
C8849 vdd.n361 vss 0.00251f
C8850 vdd.n362 vss 0.00413f
C8851 vdd.n363 vss 0.0471f
C8852 vdd.t156 vss 0.0471f
C8853 vdd.n364 vss 0.00425f
C8854 vdd.n365 vss 0.0424f
C8855 vdd.n366 vss 0.0132f
C8856 vdd.n367 vss 0.02f
C8857 vdd.n368 vss 0.00425f
C8858 vdd.n369 vss 0.00413f
C8859 vdd.n370 vss 0.00251f
C8860 vdd.n371 vss 0.0112f
C8861 vdd.n372 vss 0.0128f
C8862 vdd.n373 vss 0.0418f
C8863 vdd.t1414 vss 0.00134f
C8864 vdd.t1486 vss 0.0013f
C8865 vdd.n374 vss 0.032f
C8866 vdd.n375 vss 0.0393f
C8867 vdd.n376 vss 0.00324f
C8868 vdd.n377 vss 0.0112f
C8869 vdd.n378 vss 0.0128f
C8870 vdd.n379 vss 0.00413f
C8871 vdd.t1415 vss 0.0471f
C8872 vdd.n380 vss 0.00324f
C8873 vdd.n382 vss 0.00925f
C8874 vdd.n383 vss 0.00413f
C8875 vdd.n384 vss 0.00679f
C8876 vdd.n385 vss 0.00413f
C8877 vdd.n386 vss 0.0471f
C8878 vdd.n387 vss 0.00324f
C8879 vdd.n388 vss 0.0471f
C8880 vdd.n389 vss 0.00324f
C8881 vdd.n390 vss 0.0424f
C8882 vdd.t1485 vss 0.0471f
C8883 vdd.n392 vss 0.00425f
C8884 vdd.n393 vss 0.00925f
C8885 vdd.n394 vss 0.0132f
C8886 vdd.n395 vss 0.00324f
C8887 vdd.n396 vss 0.0128f
C8888 vdd.n397 vss 0.02f
C8889 vdd.n398 vss 0.00425f
C8890 vdd.n399 vss 0.00413f
C8891 vdd.n400 vss 0.00251f
C8892 vdd.t1413 vss 0.0471f
C8893 vdd.n401 vss 0.00251f
C8894 vdd.n402 vss 0.00517f
C8895 vdd.n403 vss 0.00679f
C8896 vdd.n404 vss 0.00324f
C8897 vdd.n405 vss 0.00679f
C8898 vdd.n406 vss 0.00517f
C8899 vdd.n407 vss 0.00251f
C8900 vdd.n408 vss 0.00413f
C8901 vdd.n409 vss 0.0471f
C8902 vdd.t959 vss 0.0471f
C8903 vdd.n410 vss 0.00425f
C8904 vdd.n411 vss 0.0424f
C8905 vdd.n412 vss 0.0132f
C8906 vdd.n413 vss 0.02f
C8907 vdd.n414 vss 0.00425f
C8908 vdd.n415 vss 0.00413f
C8909 vdd.n416 vss 0.00251f
C8910 vdd.n417 vss 0.0112f
C8911 vdd.n418 vss 0.0128f
C8912 vdd.n419 vss 0.0369f
C8913 vdd.n420 vss 0.00335f
C8914 vdd.t580 vss 0.0013f
C8915 vdd.n421 vss 0.0309f
C8916 vdd.n422 vss 0.0107f
C8917 vdd.n423 vss 0.0128f
C8918 vdd.n424 vss 0.0424f
C8919 vdd.t579 vss 0.0471f
C8920 vdd.n425 vss 0.00324f
C8921 vdd.n426 vss 0.0471f
C8922 vdd.t740 vss 0.0471f
C8923 vdd.n427 vss 0.00413f
C8924 vdd.n428 vss 0.00324f
C8925 vdd.t741 vss 0.00134f
C8926 vdd.n429 vss 0.0393f
C8927 vdd.n430 vss 0.0128f
C8928 vdd.t739 vss 0.0471f
C8929 vdd.n431 vss 0.00324f
C8930 vdd.n433 vss 0.00925f
C8931 vdd.n434 vss 0.0471f
C8932 vdd.n435 vss 0.00324f
C8933 vdd.n436 vss 0.00413f
C8934 vdd.n437 vss 0.00324f
C8935 vdd.n438 vss 0.00679f
C8936 vdd.n440 vss 0.00925f
C8937 vdd.n441 vss 0.00425f
C8938 vdd.n442 vss 0.00413f
C8939 vdd.n443 vss 0.00251f
C8940 vdd.n444 vss 0.00517f
C8941 vdd.n445 vss 0.00679f
C8942 vdd.n446 vss 0.00324f
C8943 vdd.n447 vss 0.00679f
C8944 vdd.n448 vss 0.00517f
C8945 vdd.n449 vss 0.00251f
C8946 vdd.n450 vss 0.00413f
C8947 vdd.n451 vss 0.0471f
C8948 vdd.t1122 vss 0.0471f
C8949 vdd.n452 vss 0.00425f
C8950 vdd.n453 vss 0.0424f
C8951 vdd.n454 vss 0.0132f
C8952 vdd.n455 vss 0.02f
C8953 vdd.n456 vss 0.00425f
C8954 vdd.n457 vss 0.00413f
C8955 vdd.n458 vss 0.00251f
C8956 vdd.n459 vss 0.0105f
C8957 vdd.n460 vss 0.0633f
C8958 vdd.n461 vss 0.00805f
C8959 vdd.n462 vss 0.0112f
C8960 vdd.n463 vss 0.00251f
C8961 vdd.n464 vss 0.00413f
C8962 vdd.n465 vss 0.00425f
C8963 vdd.n466 vss 0.00991f
C8964 vdd.n467 vss 0.0126f
C8965 vdd.n468 vss 9.89e-19
C8966 vdd.n469 vss 0.0011f
C8967 vdd.n470 vss 0.0271f
C8968 vdd.t926 vss 0.00134f
C8969 vdd.t210 vss 0.0013f
C8970 vdd.n471 vss 0.032f
C8971 vdd.n472 vss 0.0393f
C8972 vdd.n473 vss 0.00324f
C8973 vdd.n474 vss 0.0112f
C8974 vdd.n475 vss 0.0128f
C8975 vdd.n476 vss 0.00413f
C8976 vdd.t927 vss 0.0471f
C8977 vdd.n477 vss 0.00324f
C8978 vdd.n479 vss 0.00925f
C8979 vdd.n480 vss 0.00413f
C8980 vdd.n481 vss 0.00679f
C8981 vdd.n482 vss 0.00413f
C8982 vdd.n483 vss 0.0471f
C8983 vdd.n484 vss 0.00324f
C8984 vdd.n485 vss 0.0471f
C8985 vdd.n486 vss 0.00324f
C8986 vdd.n487 vss 0.0424f
C8987 vdd.t209 vss 0.0471f
C8988 vdd.n489 vss 0.00425f
C8989 vdd.n490 vss 0.00925f
C8990 vdd.n491 vss 0.0132f
C8991 vdd.n492 vss 0.00324f
C8992 vdd.n493 vss 0.0128f
C8993 vdd.n494 vss 0.02f
C8994 vdd.n495 vss 0.00425f
C8995 vdd.n496 vss 0.00413f
C8996 vdd.n497 vss 0.00251f
C8997 vdd.t925 vss 0.0471f
C8998 vdd.n498 vss 0.00251f
C8999 vdd.n499 vss 0.00517f
C9000 vdd.n500 vss 0.00679f
C9001 vdd.n501 vss 0.00324f
C9002 vdd.n502 vss 0.00679f
C9003 vdd.n503 vss 0.00517f
C9004 vdd.n504 vss 0.00251f
C9005 vdd.n505 vss 0.00413f
C9006 vdd.n506 vss 0.0471f
C9007 vdd.t336 vss 0.0471f
C9008 vdd.n507 vss 0.00425f
C9009 vdd.n508 vss 0.0424f
C9010 vdd.n509 vss 0.0132f
C9011 vdd.n510 vss 0.02f
C9012 vdd.n511 vss 0.00425f
C9013 vdd.n512 vss 0.00413f
C9014 vdd.n513 vss 0.00251f
C9015 vdd.n514 vss 0.0112f
C9016 vdd.n515 vss 0.0128f
C9017 vdd.n516 vss 0.0418f
C9018 vdd.t128 vss 0.00134f
C9019 vdd.t376 vss 0.0013f
C9020 vdd.n517 vss 0.0315f
C9021 vdd.n518 vss 0.0393f
C9022 vdd.n519 vss 0.00324f
C9023 vdd.n520 vss 0.0112f
C9024 vdd.n521 vss 0.0128f
C9025 vdd.n522 vss 0.00413f
C9026 vdd.t126 vss 0.0471f
C9027 vdd.n523 vss 0.00324f
C9028 vdd.n525 vss 0.00925f
C9029 vdd.n526 vss 0.00413f
C9030 vdd.n527 vss 0.00679f
C9031 vdd.n528 vss 0.00413f
C9032 vdd.n529 vss 0.0471f
C9033 vdd.n530 vss 0.00324f
C9034 vdd.n531 vss 0.0471f
C9035 vdd.n532 vss 0.00324f
C9036 vdd.n533 vss 0.0424f
C9037 vdd.t375 vss 0.0471f
C9038 vdd.n535 vss 0.00425f
C9039 vdd.n536 vss 0.00925f
C9040 vdd.n537 vss 0.0132f
C9041 vdd.n538 vss 0.00324f
C9042 vdd.n539 vss 0.0128f
C9043 vdd.n540 vss 0.02f
C9044 vdd.n541 vss 0.00425f
C9045 vdd.n542 vss 0.00413f
C9046 vdd.n543 vss 0.00251f
C9047 vdd.t127 vss 0.0471f
C9048 vdd.n544 vss 0.00251f
C9049 vdd.n545 vss 0.00517f
C9050 vdd.n546 vss 0.00679f
C9051 vdd.n547 vss 0.00324f
C9052 vdd.n548 vss 0.00679f
C9053 vdd.n549 vss 0.00517f
C9054 vdd.n550 vss 0.00251f
C9055 vdd.n551 vss 0.00413f
C9056 vdd.n552 vss 0.0471f
C9057 vdd.t122 vss 0.0471f
C9058 vdd.n553 vss 0.00425f
C9059 vdd.n554 vss 0.0424f
C9060 vdd.n555 vss 0.0132f
C9061 vdd.n556 vss 0.02f
C9062 vdd.n557 vss 0.00425f
C9063 vdd.n558 vss 0.00413f
C9064 vdd.n559 vss 0.00251f
C9065 vdd.n560 vss 0.0112f
C9066 vdd.n561 vss 0.0128f
C9067 vdd.n562 vss 0.0365f
C9068 vdd.t27 vss 0.0013f
C9069 vdd.t911 vss 0.00134f
C9070 vdd.t985 vss 0.0013f
C9071 vdd.t1115 vss 0.00134f
C9072 vdd.t29 vss 0.0013f
C9073 vdd.t708 vss 0.00134f
C9074 vdd.t1187 vss 0.0013f
C9075 vdd.t551 vss 0.00134f
C9076 vdd.t25 vss 0.0013f
C9077 vdd.t1430 vss 0.00134f
C9078 vdd.t987 vss 0.0013f
C9079 vdd.t1174 vss 0.00134f
C9080 vdd.t31 vss 0.0013f
C9081 vdd.t1152 vss 0.00134f
C9082 vdd.n563 vss 0.00324f
C9083 vdd.n564 vss 0.0112f
C9084 vdd.n565 vss 0.0128f
C9085 vdd.n566 vss 0.00413f
C9086 vdd.n567 vss 0.00413f
C9087 vdd.n568 vss 0.0471f
C9088 vdd.n569 vss 0.00251f
C9089 vdd.t30 vss 0.0471f
C9090 vdd.n570 vss 0.00324f
C9091 vdd.n572 vss 0.00679f
C9092 vdd.n573 vss 0.00413f
C9093 vdd.n574 vss 0.00324f
C9094 vdd.n575 vss 0.00413f
C9095 vdd.n576 vss 0.0471f
C9096 vdd.n577 vss 0.00324f
C9097 vdd.n579 vss 0.00925f
C9098 vdd.t748 vss 0.0471f
C9099 vdd.n580 vss 0.00425f
C9100 vdd.n581 vss 0.0424f
C9101 vdd.n582 vss 0.0132f
C9102 vdd.n583 vss 0.00324f
C9103 vdd.n584 vss 0.0128f
C9104 vdd.n585 vss 0.02f
C9105 vdd.n586 vss 0.00425f
C9106 vdd.n587 vss 0.00413f
C9107 vdd.n588 vss 0.00251f
C9108 vdd.t1153 vss 0.0471f
C9109 vdd.n589 vss 0.00251f
C9110 vdd.n590 vss 0.00517f
C9111 vdd.n591 vss 0.00679f
C9112 vdd.n592 vss 0.00517f
C9113 vdd.n593 vss 0.00679f
C9114 vdd.n594 vss 0.02f
C9115 vdd.n595 vss 0.00425f
C9116 vdd.n596 vss 0.0424f
C9117 vdd.n597 vss 0.0132f
C9118 vdd.n598 vss 0.00925f
C9119 vdd.n599 vss 0.00425f
C9120 vdd.n600 vss 0.00413f
C9121 vdd.n601 vss 0.00324f
C9122 vdd.n602 vss 0.0471f
C9123 vdd.t1151 vss 0.0471f
C9124 vdd.n603 vss 0.00251f
C9125 vdd.n604 vss 0.0112f
C9126 vdd.n605 vss 0.0707f
C9127 vdd.n606 vss 0.0393f
C9128 vdd.n607 vss 0.0332f
C9129 vdd.t349 vss 0.00134f
C9130 vdd.t553 vss 0.0013f
C9131 vdd.n608 vss 0.0315f
C9132 vdd.n609 vss 0.0393f
C9133 vdd.n610 vss 0.00324f
C9134 vdd.n611 vss 0.0112f
C9135 vdd.n612 vss 0.0128f
C9136 vdd.n613 vss 0.00413f
C9137 vdd.t347 vss 0.0471f
C9138 vdd.n614 vss 0.00324f
C9139 vdd.n616 vss 0.00925f
C9140 vdd.n617 vss 0.00413f
C9141 vdd.n618 vss 0.00679f
C9142 vdd.n619 vss 0.00413f
C9143 vdd.n620 vss 0.0471f
C9144 vdd.n621 vss 0.00324f
C9145 vdd.n622 vss 0.0471f
C9146 vdd.n623 vss 0.00324f
C9147 vdd.n624 vss 0.0424f
C9148 vdd.t552 vss 0.0471f
C9149 vdd.n626 vss 0.00425f
C9150 vdd.n627 vss 0.00925f
C9151 vdd.n628 vss 0.0132f
C9152 vdd.n629 vss 0.00324f
C9153 vdd.n630 vss 0.0128f
C9154 vdd.n631 vss 0.02f
C9155 vdd.n632 vss 0.00425f
C9156 vdd.n633 vss 0.00413f
C9157 vdd.n634 vss 0.00251f
C9158 vdd.t348 vss 0.0471f
C9159 vdd.n635 vss 0.00251f
C9160 vdd.n636 vss 0.00517f
C9161 vdd.n637 vss 0.00679f
C9162 vdd.n638 vss 0.00324f
C9163 vdd.n639 vss 0.00679f
C9164 vdd.n640 vss 0.00517f
C9165 vdd.n641 vss 0.00251f
C9166 vdd.n642 vss 0.00413f
C9167 vdd.n643 vss 0.0471f
C9168 vdd.t893 vss 0.0471f
C9169 vdd.n644 vss 0.00425f
C9170 vdd.n645 vss 0.0424f
C9171 vdd.n646 vss 0.0132f
C9172 vdd.n647 vss 0.02f
C9173 vdd.n648 vss 0.00425f
C9174 vdd.n649 vss 0.00413f
C9175 vdd.n650 vss 0.00251f
C9176 vdd.n651 vss 0.0112f
C9177 vdd.n652 vss 0.0128f
C9178 vdd.n653 vss 0.0365f
C9179 vdd.n654 vss 0.202f
C9180 vdd.n655 vss 0.00324f
C9181 vdd.n656 vss 0.0112f
C9182 vdd.n657 vss 0.0128f
C9183 vdd.n658 vss 0.00413f
C9184 vdd.n659 vss 0.00413f
C9185 vdd.n660 vss 0.0471f
C9186 vdd.n661 vss 0.00251f
C9187 vdd.t1465 vss 0.0471f
C9188 vdd.n662 vss 0.00324f
C9189 vdd.n664 vss 0.00679f
C9190 vdd.n665 vss 0.00413f
C9191 vdd.n666 vss 0.00324f
C9192 vdd.n667 vss 0.00413f
C9193 vdd.n668 vss 0.0471f
C9194 vdd.n669 vss 0.00324f
C9195 vdd.n671 vss 0.00925f
C9196 vdd.t695 vss 0.0471f
C9197 vdd.n672 vss 0.00425f
C9198 vdd.n673 vss 0.0424f
C9199 vdd.n674 vss 0.0132f
C9200 vdd.n675 vss 0.00324f
C9201 vdd.n676 vss 0.0128f
C9202 vdd.n677 vss 0.02f
C9203 vdd.n678 vss 0.00425f
C9204 vdd.n679 vss 0.00413f
C9205 vdd.n680 vss 0.00251f
C9206 vdd.t46 vss 0.0471f
C9207 vdd.n681 vss 0.00251f
C9208 vdd.n682 vss 0.00517f
C9209 vdd.n683 vss 0.00679f
C9210 vdd.n684 vss 0.00517f
C9211 vdd.n685 vss 0.00679f
C9212 vdd.n686 vss 0.02f
C9213 vdd.n687 vss 0.00425f
C9214 vdd.n688 vss 0.0424f
C9215 vdd.n689 vss 0.0132f
C9216 vdd.n690 vss 0.00925f
C9217 vdd.n691 vss 0.00425f
C9218 vdd.n692 vss 0.00413f
C9219 vdd.n693 vss 0.00324f
C9220 vdd.n694 vss 0.0471f
C9221 vdd.t47 vss 0.0471f
C9222 vdd.n695 vss 0.00251f
C9223 vdd.n696 vss 0.0112f
C9224 vdd.n697 vss 0.0128f
C9225 vdd.t48 vss 0.00134f
C9226 vdd.t1466 vss 0.0013f
C9227 vdd.n698 vss 0.0332f
C9228 vdd.n699 vss 0.0393f
C9229 vdd.n700 vss 0.0418f
C9230 vdd.n701 vss 0.00324f
C9231 vdd.n702 vss 0.0112f
C9232 vdd.n703 vss 0.0128f
C9233 vdd.n704 vss 0.00413f
C9234 vdd.n705 vss 0.00413f
C9235 vdd.n706 vss 0.0471f
C9236 vdd.n707 vss 0.00251f
C9237 vdd.t1501 vss 0.0471f
C9238 vdd.n708 vss 0.00324f
C9239 vdd.n710 vss 0.00679f
C9240 vdd.n711 vss 0.00413f
C9241 vdd.n712 vss 0.00324f
C9242 vdd.n713 vss 0.00413f
C9243 vdd.n714 vss 0.0471f
C9244 vdd.n715 vss 0.00324f
C9245 vdd.n717 vss 0.00925f
C9246 vdd.t1406 vss 0.0471f
C9247 vdd.n718 vss 0.00425f
C9248 vdd.n719 vss 0.0424f
C9249 vdd.n720 vss 0.0132f
C9250 vdd.n721 vss 0.00324f
C9251 vdd.n722 vss 0.0128f
C9252 vdd.n723 vss 0.02f
C9253 vdd.n724 vss 0.00425f
C9254 vdd.n725 vss 0.00413f
C9255 vdd.n726 vss 0.00251f
C9256 vdd.t123 vss 0.0471f
C9257 vdd.n727 vss 0.00251f
C9258 vdd.n728 vss 0.00517f
C9259 vdd.n729 vss 0.00679f
C9260 vdd.n730 vss 0.00517f
C9261 vdd.n731 vss 0.00679f
C9262 vdd.n732 vss 0.02f
C9263 vdd.n733 vss 0.00425f
C9264 vdd.n734 vss 0.0424f
C9265 vdd.n735 vss 0.0132f
C9266 vdd.n736 vss 0.00925f
C9267 vdd.n737 vss 0.00425f
C9268 vdd.n738 vss 0.00413f
C9269 vdd.n739 vss 0.00324f
C9270 vdd.n740 vss 0.0471f
C9271 vdd.t124 vss 0.0471f
C9272 vdd.n741 vss 0.00251f
C9273 vdd.n742 vss 0.0112f
C9274 vdd.n743 vss 0.0128f
C9275 vdd.t125 vss 0.00134f
C9276 vdd.t1502 vss 0.0013f
C9277 vdd.n744 vss 0.0332f
C9278 vdd.n745 vss 0.0393f
C9279 vdd.n746 vss 0.0345f
C9280 vdd.n747 vss 0.00335f
C9281 vdd.t88 vss 0.0013f
C9282 vdd.n748 vss 0.0309f
C9283 vdd.n749 vss 0.00991f
C9284 vdd.n750 vss 0.0424f
C9285 vdd.n751 vss 0.00679f
C9286 vdd.n752 vss 0.00413f
C9287 vdd.n753 vss 0.0471f
C9288 vdd.n754 vss 0.00251f
C9289 vdd.n755 vss 0.00324f
C9290 vdd.n756 vss 0.0128f
C9291 vdd.n757 vss 0.00413f
C9292 vdd.n758 vss 0.00413f
C9293 vdd.n759 vss 0.0471f
C9294 vdd.n760 vss 0.00251f
C9295 vdd.n761 vss 0.00324f
C9296 vdd.n762 vss 0.00413f
C9297 vdd.n763 vss 0.00324f
C9298 vdd.n764 vss 0.0132f
C9299 vdd.n765 vss 0.0424f
C9300 vdd.n766 vss 0.00324f
C9301 vdd.n767 vss 0.00413f
C9302 vdd.n768 vss 0.02f
C9303 vdd.n769 vss 0.00425f
C9304 vdd.t1410 vss 0.0471f
C9305 vdd.n771 vss 0.00425f
C9306 vdd.n772 vss 0.00925f
C9307 vdd.n773 vss 0.00679f
C9308 vdd.n774 vss 0.00517f
C9309 vdd.n775 vss 0.00679f
C9310 vdd.n776 vss 0.00517f
C9311 vdd.n777 vss 0.00251f
C9312 vdd.t1431 vss 0.0471f
C9313 vdd.n778 vss 0.0471f
C9314 vdd.t1433 vss 0.0471f
C9315 vdd.n779 vss 0.00251f
C9316 vdd.n780 vss 0.0105f
C9317 vdd.t1432 vss 0.00134f
C9318 vdd.n781 vss 0.0393f
C9319 vdd.n782 vss 0.0633f
C9320 vdd.n783 vss 0.00805f
C9321 vdd.n784 vss 0.0112f
C9322 vdd.n785 vss 0.0128f
C9323 vdd.n786 vss 0.00324f
C9324 vdd.n787 vss 0.00324f
C9325 vdd.n788 vss 0.00413f
C9326 vdd.n789 vss 0.00425f
C9327 vdd.t87 vss 0.0471f
C9328 vdd.n791 vss 0.00425f
C9329 vdd.n792 vss 0.00925f
C9330 vdd.n793 vss 0.0107f
C9331 vdd.n794 vss 0.0126f
C9332 vdd.n795 vss 9.89e-19
C9333 vdd.n796 vss 0.00163f
C9334 vdd.n797 vss 0.00145f
C9335 vdd.n798 vss 0.0271f
C9336 vdd.n799 vss 0.00324f
C9337 vdd.n800 vss 0.0112f
C9338 vdd.n801 vss 0.0128f
C9339 vdd.n802 vss 0.00413f
C9340 vdd.n803 vss 0.00413f
C9341 vdd.n804 vss 0.0471f
C9342 vdd.n805 vss 0.00251f
C9343 vdd.t1358 vss 0.0471f
C9344 vdd.n806 vss 0.00324f
C9345 vdd.n808 vss 0.00679f
C9346 vdd.n809 vss 0.00413f
C9347 vdd.n810 vss 0.00324f
C9348 vdd.n811 vss 0.00413f
C9349 vdd.n812 vss 0.0471f
C9350 vdd.n813 vss 0.00324f
C9351 vdd.n815 vss 0.00925f
C9352 vdd.t1202 vss 0.0471f
C9353 vdd.n816 vss 0.00425f
C9354 vdd.n817 vss 0.0424f
C9355 vdd.n818 vss 0.0132f
C9356 vdd.n819 vss 0.00324f
C9357 vdd.n820 vss 0.0128f
C9358 vdd.n821 vss 0.02f
C9359 vdd.n822 vss 0.00425f
C9360 vdd.n823 vss 0.00413f
C9361 vdd.n824 vss 0.00251f
C9362 vdd.t291 vss 0.0471f
C9363 vdd.n825 vss 0.00251f
C9364 vdd.n826 vss 0.00517f
C9365 vdd.n827 vss 0.00679f
C9366 vdd.n828 vss 0.00517f
C9367 vdd.n829 vss 0.00679f
C9368 vdd.n830 vss 0.02f
C9369 vdd.n831 vss 0.00425f
C9370 vdd.n832 vss 0.0424f
C9371 vdd.n833 vss 0.0132f
C9372 vdd.n834 vss 0.00925f
C9373 vdd.n835 vss 0.00425f
C9374 vdd.n836 vss 0.00413f
C9375 vdd.n837 vss 0.00324f
C9376 vdd.n838 vss 0.0471f
C9377 vdd.t289 vss 0.0471f
C9378 vdd.n839 vss 0.00251f
C9379 vdd.n840 vss 0.0112f
C9380 vdd.n841 vss 0.0128f
C9381 vdd.t290 vss 0.00134f
C9382 vdd.t1359 vss 0.0013f
C9383 vdd.n842 vss 0.0332f
C9384 vdd.n843 vss 0.0393f
C9385 vdd.n844 vss 0.0418f
C9386 vdd.n845 vss 0.00324f
C9387 vdd.n846 vss 0.0112f
C9388 vdd.n847 vss 0.0128f
C9389 vdd.n848 vss 0.00413f
C9390 vdd.n849 vss 0.00413f
C9391 vdd.n850 vss 0.0471f
C9392 vdd.n851 vss 0.00251f
C9393 vdd.t1497 vss 0.0471f
C9394 vdd.n852 vss 0.00324f
C9395 vdd.n854 vss 0.00679f
C9396 vdd.n855 vss 0.00413f
C9397 vdd.n856 vss 0.00324f
C9398 vdd.n857 vss 0.00413f
C9399 vdd.n858 vss 0.0471f
C9400 vdd.n859 vss 0.00324f
C9401 vdd.n861 vss 0.00925f
C9402 vdd.t1383 vss 0.0471f
C9403 vdd.n862 vss 0.00425f
C9404 vdd.n863 vss 0.0424f
C9405 vdd.n864 vss 0.0132f
C9406 vdd.n865 vss 0.00324f
C9407 vdd.n866 vss 0.0128f
C9408 vdd.n867 vss 0.02f
C9409 vdd.n868 vss 0.00425f
C9410 vdd.n869 vss 0.00413f
C9411 vdd.n870 vss 0.00251f
C9412 vdd.t427 vss 0.0471f
C9413 vdd.n871 vss 0.00251f
C9414 vdd.n872 vss 0.00517f
C9415 vdd.n873 vss 0.00679f
C9416 vdd.n874 vss 0.00517f
C9417 vdd.n875 vss 0.00679f
C9418 vdd.n876 vss 0.02f
C9419 vdd.n877 vss 0.00425f
C9420 vdd.n878 vss 0.0424f
C9421 vdd.n879 vss 0.0132f
C9422 vdd.n880 vss 0.00925f
C9423 vdd.n881 vss 0.00425f
C9424 vdd.n882 vss 0.00413f
C9425 vdd.n883 vss 0.00324f
C9426 vdd.n884 vss 0.0471f
C9427 vdd.t425 vss 0.0471f
C9428 vdd.n885 vss 0.00251f
C9429 vdd.n886 vss 0.0112f
C9430 vdd.n887 vss 0.0128f
C9431 vdd.t426 vss 0.00134f
C9432 vdd.t1498 vss 0.0013f
C9433 vdd.n888 vss 0.0332f
C9434 vdd.n889 vss 0.0393f
C9435 vdd.n890 vss 0.0345f
C9436 vdd.n891 vss 0.00324f
C9437 vdd.n892 vss 0.0112f
C9438 vdd.n893 vss 0.0128f
C9439 vdd.n894 vss 0.00413f
C9440 vdd.n895 vss 0.00413f
C9441 vdd.n896 vss 0.0471f
C9442 vdd.n897 vss 0.00251f
C9443 vdd.t1312 vss 0.0471f
C9444 vdd.n898 vss 0.00324f
C9445 vdd.n900 vss 0.00679f
C9446 vdd.n901 vss 0.00413f
C9447 vdd.n902 vss 0.00324f
C9448 vdd.n903 vss 0.00413f
C9449 vdd.n904 vss 0.0471f
C9450 vdd.n905 vss 0.00324f
C9451 vdd.n907 vss 0.00925f
C9452 vdd.t361 vss 0.0471f
C9453 vdd.n908 vss 0.00425f
C9454 vdd.n909 vss 0.0424f
C9455 vdd.n910 vss 0.0132f
C9456 vdd.n911 vss 0.00324f
C9457 vdd.n912 vss 0.0128f
C9458 vdd.n913 vss 0.02f
C9459 vdd.n914 vss 0.00425f
C9460 vdd.n915 vss 0.00413f
C9461 vdd.n916 vss 0.00251f
C9462 vdd.t215 vss 0.0471f
C9463 vdd.n917 vss 0.00251f
C9464 vdd.n918 vss 0.00517f
C9465 vdd.n919 vss 0.00679f
C9466 vdd.n920 vss 0.00517f
C9467 vdd.n921 vss 0.00679f
C9468 vdd.n922 vss 0.02f
C9469 vdd.n923 vss 0.00425f
C9470 vdd.n924 vss 0.0424f
C9471 vdd.n925 vss 0.0132f
C9472 vdd.n926 vss 0.00925f
C9473 vdd.n927 vss 0.00425f
C9474 vdd.n928 vss 0.00413f
C9475 vdd.n929 vss 0.00324f
C9476 vdd.n930 vss 0.0471f
C9477 vdd.t213 vss 0.0471f
C9478 vdd.n931 vss 0.00251f
C9479 vdd.n932 vss 0.0112f
C9480 vdd.n933 vss 0.0128f
C9481 vdd.t214 vss 0.00134f
C9482 vdd.t1313 vss 0.0013f
C9483 vdd.n934 vss 0.0332f
C9484 vdd.n935 vss 0.0393f
C9485 vdd.n936 vss 0.0418f
C9486 vdd.n937 vss 0.00324f
C9487 vdd.n938 vss 0.0112f
C9488 vdd.n939 vss 0.0128f
C9489 vdd.n940 vss 0.00413f
C9490 vdd.n941 vss 0.00413f
C9491 vdd.n942 vss 0.0471f
C9492 vdd.n943 vss 0.00251f
C9493 vdd.t462 vss 0.0471f
C9494 vdd.n944 vss 0.00324f
C9495 vdd.n946 vss 0.00679f
C9496 vdd.n947 vss 0.00413f
C9497 vdd.n948 vss 0.00324f
C9498 vdd.n949 vss 0.00413f
C9499 vdd.n950 vss 0.0471f
C9500 vdd.n951 vss 0.00324f
C9501 vdd.n953 vss 0.00925f
C9502 vdd.t236 vss 0.0471f
C9503 vdd.n954 vss 0.00425f
C9504 vdd.n955 vss 0.0424f
C9505 vdd.n956 vss 0.0132f
C9506 vdd.n957 vss 0.00324f
C9507 vdd.n958 vss 0.0128f
C9508 vdd.n959 vss 0.02f
C9509 vdd.n960 vss 0.00425f
C9510 vdd.n961 vss 0.00413f
C9511 vdd.n962 vss 0.00251f
C9512 vdd.t923 vss 0.0471f
C9513 vdd.n963 vss 0.00251f
C9514 vdd.n964 vss 0.00517f
C9515 vdd.n965 vss 0.00679f
C9516 vdd.n966 vss 0.00517f
C9517 vdd.n967 vss 0.00679f
C9518 vdd.n968 vss 0.02f
C9519 vdd.n969 vss 0.00425f
C9520 vdd.n970 vss 0.0424f
C9521 vdd.n971 vss 0.0132f
C9522 vdd.n972 vss 0.00925f
C9523 vdd.n973 vss 0.00425f
C9524 vdd.n974 vss 0.00413f
C9525 vdd.n975 vss 0.00324f
C9526 vdd.n976 vss 0.0471f
C9527 vdd.t921 vss 0.0471f
C9528 vdd.n977 vss 0.00251f
C9529 vdd.n978 vss 0.0112f
C9530 vdd.n979 vss 0.0128f
C9531 vdd.t922 vss 0.00134f
C9532 vdd.t463 vss 0.0013f
C9533 vdd.n980 vss 0.0332f
C9534 vdd.n981 vss 0.0393f
C9535 vdd.n982 vss 0.0345f
C9536 vdd.n983 vss 0.00335f
C9537 vdd.t92 vss 0.0013f
C9538 vdd.n984 vss 0.0309f
C9539 vdd.n985 vss 0.00991f
C9540 vdd.n986 vss 0.0424f
C9541 vdd.n987 vss 0.00679f
C9542 vdd.n988 vss 0.00413f
C9543 vdd.n989 vss 0.0471f
C9544 vdd.n990 vss 0.00251f
C9545 vdd.n991 vss 0.00324f
C9546 vdd.n992 vss 0.0128f
C9547 vdd.n993 vss 0.00413f
C9548 vdd.n994 vss 0.00413f
C9549 vdd.n995 vss 0.0471f
C9550 vdd.n996 vss 0.00251f
C9551 vdd.n997 vss 0.00324f
C9552 vdd.n998 vss 0.00413f
C9553 vdd.n999 vss 0.00324f
C9554 vdd.n1000 vss 0.0132f
C9555 vdd.n1001 vss 0.0424f
C9556 vdd.n1002 vss 0.00324f
C9557 vdd.n1003 vss 0.00413f
C9558 vdd.n1004 vss 0.02f
C9559 vdd.n1005 vss 0.00425f
C9560 vdd.t1230 vss 0.0471f
C9561 vdd.n1007 vss 0.00425f
C9562 vdd.n1008 vss 0.00925f
C9563 vdd.n1009 vss 0.00679f
C9564 vdd.n1010 vss 0.00517f
C9565 vdd.n1011 vss 0.00679f
C9566 vdd.n1012 vss 0.00517f
C9567 vdd.n1013 vss 0.00251f
C9568 vdd.t402 vss 0.0471f
C9569 vdd.n1014 vss 0.0471f
C9570 vdd.t404 vss 0.0471f
C9571 vdd.n1015 vss 0.00251f
C9572 vdd.n1016 vss 0.0105f
C9573 vdd.t403 vss 0.00134f
C9574 vdd.n1017 vss 0.0393f
C9575 vdd.n1018 vss 0.0633f
C9576 vdd.n1019 vss 0.00805f
C9577 vdd.n1020 vss 0.0112f
C9578 vdd.n1021 vss 0.0128f
C9579 vdd.n1022 vss 0.00324f
C9580 vdd.n1023 vss 0.00324f
C9581 vdd.n1024 vss 0.00413f
C9582 vdd.n1025 vss 0.00425f
C9583 vdd.t91 vss 0.0471f
C9584 vdd.n1027 vss 0.00425f
C9585 vdd.n1028 vss 0.00925f
C9586 vdd.n1029 vss 0.0107f
C9587 vdd.n1030 vss 0.0126f
C9588 vdd.n1031 vss 9.89e-19
C9589 vdd.n1032 vss 0.00163f
C9590 vdd.n1033 vss 0.00145f
C9591 vdd.n1034 vss 0.0271f
C9592 vdd.n1035 vss 0.00324f
C9593 vdd.n1036 vss 0.0112f
C9594 vdd.n1037 vss 0.0128f
C9595 vdd.n1038 vss 0.00413f
C9596 vdd.n1039 vss 0.00413f
C9597 vdd.n1040 vss 0.0471f
C9598 vdd.n1041 vss 0.00251f
C9599 vdd.t1469 vss 0.0471f
C9600 vdd.n1042 vss 0.00324f
C9601 vdd.n1044 vss 0.00679f
C9602 vdd.n1045 vss 0.00413f
C9603 vdd.n1046 vss 0.00324f
C9604 vdd.n1047 vss 0.00413f
C9605 vdd.n1048 vss 0.0471f
C9606 vdd.n1049 vss 0.00324f
C9607 vdd.n1051 vss 0.00925f
C9608 vdd.t1259 vss 0.0471f
C9609 vdd.n1052 vss 0.00425f
C9610 vdd.n1053 vss 0.0424f
C9611 vdd.n1054 vss 0.0132f
C9612 vdd.n1055 vss 0.00324f
C9613 vdd.n1056 vss 0.0128f
C9614 vdd.n1057 vss 0.02f
C9615 vdd.n1058 vss 0.00425f
C9616 vdd.n1059 vss 0.00413f
C9617 vdd.n1060 vss 0.00251f
C9618 vdd.t957 vss 0.0471f
C9619 vdd.n1061 vss 0.00251f
C9620 vdd.n1062 vss 0.00517f
C9621 vdd.n1063 vss 0.00679f
C9622 vdd.n1064 vss 0.00517f
C9623 vdd.n1065 vss 0.00679f
C9624 vdd.n1066 vss 0.02f
C9625 vdd.n1067 vss 0.00425f
C9626 vdd.n1068 vss 0.0424f
C9627 vdd.n1069 vss 0.0132f
C9628 vdd.n1070 vss 0.00925f
C9629 vdd.n1071 vss 0.00425f
C9630 vdd.n1072 vss 0.00413f
C9631 vdd.n1073 vss 0.00324f
C9632 vdd.n1074 vss 0.0471f
C9633 vdd.t955 vss 0.0471f
C9634 vdd.n1075 vss 0.00251f
C9635 vdd.n1076 vss 0.0112f
C9636 vdd.n1077 vss 0.0128f
C9637 vdd.t956 vss 0.00134f
C9638 vdd.t1470 vss 0.0013f
C9639 vdd.n1078 vss 0.0332f
C9640 vdd.n1079 vss 0.0393f
C9641 vdd.n1080 vss 0.0418f
C9642 vdd.t112 vss 0.00134f
C9643 vdd.t4 vss 0.0013f
C9644 vdd.n1081 vss 0.032f
C9645 vdd.n1082 vss 0.0393f
C9646 vdd.n1083 vss 0.00324f
C9647 vdd.n1084 vss 0.0112f
C9648 vdd.n1085 vss 0.0128f
C9649 vdd.n1086 vss 0.00413f
C9650 vdd.t113 vss 0.0471f
C9651 vdd.n1087 vss 0.00324f
C9652 vdd.n1089 vss 0.00925f
C9653 vdd.n1090 vss 0.00413f
C9654 vdd.n1091 vss 0.00679f
C9655 vdd.n1092 vss 0.00413f
C9656 vdd.n1093 vss 0.0471f
C9657 vdd.n1094 vss 0.00324f
C9658 vdd.n1095 vss 0.0471f
C9659 vdd.n1096 vss 0.00324f
C9660 vdd.n1097 vss 0.0424f
C9661 vdd.t3 vss 0.0471f
C9662 vdd.n1099 vss 0.00425f
C9663 vdd.n1100 vss 0.00925f
C9664 vdd.n1101 vss 0.0132f
C9665 vdd.n1102 vss 0.00324f
C9666 vdd.n1103 vss 0.0128f
C9667 vdd.n1104 vss 0.02f
C9668 vdd.n1105 vss 0.00425f
C9669 vdd.n1106 vss 0.00413f
C9670 vdd.n1107 vss 0.00251f
C9671 vdd.t111 vss 0.0471f
C9672 vdd.n1108 vss 0.00251f
C9673 vdd.n1109 vss 0.00517f
C9674 vdd.n1110 vss 0.00679f
C9675 vdd.n1111 vss 0.00324f
C9676 vdd.n1112 vss 0.00679f
C9677 vdd.n1113 vss 0.00517f
C9678 vdd.n1114 vss 0.00251f
C9679 vdd.n1115 vss 0.00413f
C9680 vdd.n1116 vss 0.0471f
C9681 vdd.t947 vss 0.0471f
C9682 vdd.n1117 vss 0.00425f
C9683 vdd.n1118 vss 0.0424f
C9684 vdd.n1119 vss 0.0132f
C9685 vdd.n1120 vss 0.02f
C9686 vdd.n1121 vss 0.00425f
C9687 vdd.n1122 vss 0.00413f
C9688 vdd.n1123 vss 0.00251f
C9689 vdd.n1124 vss 0.0112f
C9690 vdd.n1125 vss 0.0128f
C9691 vdd.n1126 vss 0.0418f
C9692 vdd.t732 vss 0.00134f
C9693 vdd.t196 vss 0.0013f
C9694 vdd.n1127 vss 0.032f
C9695 vdd.n1128 vss 0.0393f
C9696 vdd.n1129 vss 0.00324f
C9697 vdd.n1130 vss 0.0112f
C9698 vdd.n1131 vss 0.0128f
C9699 vdd.n1132 vss 0.00413f
C9700 vdd.t730 vss 0.0471f
C9701 vdd.n1133 vss 0.00324f
C9702 vdd.n1135 vss 0.00925f
C9703 vdd.n1136 vss 0.00413f
C9704 vdd.n1137 vss 0.00679f
C9705 vdd.n1138 vss 0.00413f
C9706 vdd.n1139 vss 0.0471f
C9707 vdd.n1140 vss 0.00324f
C9708 vdd.n1141 vss 0.0471f
C9709 vdd.n1142 vss 0.00324f
C9710 vdd.n1143 vss 0.0424f
C9711 vdd.t195 vss 0.0471f
C9712 vdd.n1145 vss 0.00425f
C9713 vdd.n1146 vss 0.00925f
C9714 vdd.n1147 vss 0.0132f
C9715 vdd.n1148 vss 0.00324f
C9716 vdd.n1149 vss 0.0128f
C9717 vdd.n1150 vss 0.02f
C9718 vdd.n1151 vss 0.00425f
C9719 vdd.n1152 vss 0.00413f
C9720 vdd.n1153 vss 0.00251f
C9721 vdd.t731 vss 0.0471f
C9722 vdd.n1154 vss 0.00251f
C9723 vdd.n1155 vss 0.00517f
C9724 vdd.n1156 vss 0.00679f
C9725 vdd.n1157 vss 0.00324f
C9726 vdd.n1158 vss 0.00679f
C9727 vdd.n1159 vss 0.00517f
C9728 vdd.n1160 vss 0.00251f
C9729 vdd.n1161 vss 0.00413f
C9730 vdd.n1162 vss 0.0471f
C9731 vdd.t747 vss 0.0471f
C9732 vdd.n1163 vss 0.00425f
C9733 vdd.n1164 vss 0.0424f
C9734 vdd.n1165 vss 0.0132f
C9735 vdd.n1166 vss 0.02f
C9736 vdd.n1167 vss 0.00425f
C9737 vdd.n1168 vss 0.00413f
C9738 vdd.n1169 vss 0.00251f
C9739 vdd.n1170 vss 0.0112f
C9740 vdd.n1171 vss 0.0128f
C9741 vdd.n1172 vss 0.0369f
C9742 vdd.n1173 vss 0.00335f
C9743 vdd.t96 vss 0.0013f
C9744 vdd.n1174 vss 0.0309f
C9745 vdd.n1175 vss 0.0107f
C9746 vdd.n1176 vss 0.0128f
C9747 vdd.n1177 vss 0.0424f
C9748 vdd.t95 vss 0.0471f
C9749 vdd.n1178 vss 0.00324f
C9750 vdd.n1179 vss 0.0471f
C9751 vdd.t672 vss 0.0471f
C9752 vdd.n1180 vss 0.00413f
C9753 vdd.n1181 vss 0.00324f
C9754 vdd.t673 vss 0.00134f
C9755 vdd.n1182 vss 0.0393f
C9756 vdd.n1183 vss 0.0128f
C9757 vdd.t674 vss 0.0471f
C9758 vdd.n1184 vss 0.00324f
C9759 vdd.n1186 vss 0.00925f
C9760 vdd.n1187 vss 0.0471f
C9761 vdd.n1188 vss 0.00324f
C9762 vdd.n1189 vss 0.00413f
C9763 vdd.n1190 vss 0.00324f
C9764 vdd.n1191 vss 0.00679f
C9765 vdd.n1193 vss 0.00925f
C9766 vdd.n1194 vss 0.00425f
C9767 vdd.n1195 vss 0.00413f
C9768 vdd.n1196 vss 0.00251f
C9769 vdd.n1197 vss 0.00517f
C9770 vdd.n1198 vss 0.00679f
C9771 vdd.n1199 vss 0.00324f
C9772 vdd.n1200 vss 0.00679f
C9773 vdd.n1201 vss 0.00517f
C9774 vdd.n1202 vss 0.00251f
C9775 vdd.n1203 vss 0.00413f
C9776 vdd.n1204 vss 0.0471f
C9777 vdd.t1163 vss 0.0471f
C9778 vdd.n1205 vss 0.00425f
C9779 vdd.n1206 vss 0.0424f
C9780 vdd.n1207 vss 0.0132f
C9781 vdd.n1208 vss 0.02f
C9782 vdd.n1209 vss 0.00425f
C9783 vdd.n1210 vss 0.00413f
C9784 vdd.n1211 vss 0.00251f
C9785 vdd.n1212 vss 0.0105f
C9786 vdd.n1213 vss 0.0633f
C9787 vdd.n1214 vss 0.00805f
C9788 vdd.n1215 vss 0.0112f
C9789 vdd.n1216 vss 0.00251f
C9790 vdd.n1217 vss 0.00413f
C9791 vdd.n1218 vss 0.00425f
C9792 vdd.n1219 vss 0.00991f
C9793 vdd.n1220 vss 0.0126f
C9794 vdd.n1221 vss 9.89e-19
C9795 vdd.n1222 vss 0.0011f
C9796 vdd.n1223 vss 0.0271f
C9797 vdd.t1369 vss 0.00134f
C9798 vdd.t1309 vss 0.0013f
C9799 vdd.n1224 vss 0.032f
C9800 vdd.n1225 vss 0.0393f
C9801 vdd.n1226 vss 0.00324f
C9802 vdd.n1227 vss 0.0112f
C9803 vdd.n1228 vss 0.0128f
C9804 vdd.n1229 vss 0.00413f
C9805 vdd.t1370 vss 0.0471f
C9806 vdd.n1230 vss 0.00324f
C9807 vdd.n1232 vss 0.00925f
C9808 vdd.n1233 vss 0.00413f
C9809 vdd.n1234 vss 0.00679f
C9810 vdd.n1235 vss 0.00413f
C9811 vdd.n1236 vss 0.0471f
C9812 vdd.n1237 vss 0.00324f
C9813 vdd.n1238 vss 0.0471f
C9814 vdd.n1239 vss 0.00324f
C9815 vdd.n1240 vss 0.0424f
C9816 vdd.t1308 vss 0.0471f
C9817 vdd.n1242 vss 0.00425f
C9818 vdd.n1243 vss 0.00925f
C9819 vdd.n1244 vss 0.0132f
C9820 vdd.n1245 vss 0.00324f
C9821 vdd.n1246 vss 0.0128f
C9822 vdd.n1247 vss 0.02f
C9823 vdd.n1248 vss 0.00425f
C9824 vdd.n1249 vss 0.00413f
C9825 vdd.n1250 vss 0.00251f
C9826 vdd.t1368 vss 0.0471f
C9827 vdd.n1251 vss 0.00251f
C9828 vdd.n1252 vss 0.00517f
C9829 vdd.n1253 vss 0.00679f
C9830 vdd.n1254 vss 0.00324f
C9831 vdd.n1255 vss 0.00679f
C9832 vdd.n1256 vss 0.00517f
C9833 vdd.n1257 vss 0.00251f
C9834 vdd.n1258 vss 0.00413f
C9835 vdd.n1259 vss 0.0471f
C9836 vdd.t86 vss 0.0471f
C9837 vdd.n1260 vss 0.00425f
C9838 vdd.n1261 vss 0.0424f
C9839 vdd.n1262 vss 0.0132f
C9840 vdd.n1263 vss 0.02f
C9841 vdd.n1264 vss 0.00425f
C9842 vdd.n1265 vss 0.00413f
C9843 vdd.n1266 vss 0.00251f
C9844 vdd.n1267 vss 0.0112f
C9845 vdd.n1268 vss 0.0128f
C9846 vdd.n1269 vss 0.0418f
C9847 vdd.t1104 vss 0.00134f
C9848 vdd.t1496 vss 0.0013f
C9849 vdd.n1270 vss 0.032f
C9850 vdd.n1271 vss 0.0393f
C9851 vdd.n1272 vss 0.00324f
C9852 vdd.n1273 vss 0.0112f
C9853 vdd.n1274 vss 0.0128f
C9854 vdd.n1275 vss 0.00413f
C9855 vdd.t1105 vss 0.0471f
C9856 vdd.n1276 vss 0.00324f
C9857 vdd.n1278 vss 0.00925f
C9858 vdd.n1279 vss 0.00413f
C9859 vdd.n1280 vss 0.00679f
C9860 vdd.n1281 vss 0.00413f
C9861 vdd.n1282 vss 0.0471f
C9862 vdd.n1283 vss 0.00324f
C9863 vdd.n1284 vss 0.0471f
C9864 vdd.n1285 vss 0.00324f
C9865 vdd.n1286 vss 0.0424f
C9866 vdd.t1495 vss 0.0471f
C9867 vdd.n1288 vss 0.00425f
C9868 vdd.n1289 vss 0.00925f
C9869 vdd.n1290 vss 0.0132f
C9870 vdd.n1291 vss 0.00324f
C9871 vdd.n1292 vss 0.0128f
C9872 vdd.n1293 vss 0.02f
C9873 vdd.n1294 vss 0.00425f
C9874 vdd.n1295 vss 0.00413f
C9875 vdd.n1296 vss 0.00251f
C9876 vdd.t1103 vss 0.0471f
C9877 vdd.n1297 vss 0.00251f
C9878 vdd.n1298 vss 0.00517f
C9879 vdd.n1299 vss 0.00679f
C9880 vdd.n1300 vss 0.00324f
C9881 vdd.n1301 vss 0.00679f
C9882 vdd.n1302 vss 0.00517f
C9883 vdd.n1303 vss 0.00251f
C9884 vdd.n1304 vss 0.00413f
C9885 vdd.n1305 vss 0.0471f
C9886 vdd.t157 vss 0.0471f
C9887 vdd.n1306 vss 0.00425f
C9888 vdd.n1307 vss 0.0424f
C9889 vdd.n1308 vss 0.0132f
C9890 vdd.n1309 vss 0.02f
C9891 vdd.n1310 vss 0.00425f
C9892 vdd.n1311 vss 0.00413f
C9893 vdd.n1312 vss 0.00251f
C9894 vdd.n1313 vss 0.0112f
C9895 vdd.n1314 vss 0.0128f
C9896 vdd.n1315 vss 0.0365f
C9897 vdd.t312 vss 0.00134f
C9898 vdd.t1357 vss 0.0013f
C9899 vdd.n1316 vss 0.032f
C9900 vdd.n1317 vss 0.0393f
C9901 vdd.n1318 vss 0.00324f
C9902 vdd.n1319 vss 0.0112f
C9903 vdd.n1320 vss 0.0128f
C9904 vdd.n1321 vss 0.00413f
C9905 vdd.t313 vss 0.0471f
C9906 vdd.n1322 vss 0.00324f
C9907 vdd.n1324 vss 0.00925f
C9908 vdd.n1325 vss 0.00413f
C9909 vdd.n1326 vss 0.00679f
C9910 vdd.n1327 vss 0.00413f
C9911 vdd.n1328 vss 0.0471f
C9912 vdd.n1329 vss 0.00324f
C9913 vdd.n1330 vss 0.0471f
C9914 vdd.n1331 vss 0.00324f
C9915 vdd.n1332 vss 0.0424f
C9916 vdd.t1356 vss 0.0471f
C9917 vdd.n1334 vss 0.00425f
C9918 vdd.n1335 vss 0.00925f
C9919 vdd.n1336 vss 0.0132f
C9920 vdd.n1337 vss 0.00324f
C9921 vdd.n1338 vss 0.0128f
C9922 vdd.n1339 vss 0.02f
C9923 vdd.n1340 vss 0.00425f
C9924 vdd.n1341 vss 0.00413f
C9925 vdd.n1342 vss 0.00251f
C9926 vdd.t311 vss 0.0471f
C9927 vdd.n1343 vss 0.00251f
C9928 vdd.n1344 vss 0.00517f
C9929 vdd.n1345 vss 0.00679f
C9930 vdd.n1346 vss 0.00324f
C9931 vdd.n1347 vss 0.00679f
C9932 vdd.n1348 vss 0.00517f
C9933 vdd.n1349 vss 0.00251f
C9934 vdd.n1350 vss 0.00413f
C9935 vdd.n1351 vss 0.0471f
C9936 vdd.t65 vss 0.0471f
C9937 vdd.n1352 vss 0.00425f
C9938 vdd.n1353 vss 0.0424f
C9939 vdd.n1354 vss 0.0132f
C9940 vdd.n1355 vss 0.02f
C9941 vdd.n1356 vss 0.00425f
C9942 vdd.n1357 vss 0.00413f
C9943 vdd.n1358 vss 0.00251f
C9944 vdd.n1359 vss 0.0112f
C9945 vdd.n1360 vss 0.0128f
C9946 vdd.n1361 vss 0.0418f
C9947 vdd.t919 vss 0.00134f
C9948 vdd.t592 vss 0.0013f
C9949 vdd.n1362 vss 0.032f
C9950 vdd.n1363 vss 0.0393f
C9951 vdd.n1364 vss 0.00324f
C9952 vdd.n1365 vss 0.0112f
C9953 vdd.n1366 vss 0.0128f
C9954 vdd.n1367 vss 0.00413f
C9955 vdd.t917 vss 0.0471f
C9956 vdd.n1368 vss 0.00324f
C9957 vdd.n1370 vss 0.00925f
C9958 vdd.n1371 vss 0.00413f
C9959 vdd.n1372 vss 0.00679f
C9960 vdd.n1373 vss 0.00413f
C9961 vdd.n1374 vss 0.0471f
C9962 vdd.n1375 vss 0.00324f
C9963 vdd.n1376 vss 0.0471f
C9964 vdd.n1377 vss 0.00324f
C9965 vdd.n1378 vss 0.0424f
C9966 vdd.t591 vss 0.0471f
C9967 vdd.n1380 vss 0.00425f
C9968 vdd.n1381 vss 0.00925f
C9969 vdd.n1382 vss 0.0132f
C9970 vdd.n1383 vss 0.00324f
C9971 vdd.n1384 vss 0.0128f
C9972 vdd.n1385 vss 0.02f
C9973 vdd.n1386 vss 0.00425f
C9974 vdd.n1387 vss 0.00413f
C9975 vdd.n1388 vss 0.00251f
C9976 vdd.t918 vss 0.0471f
C9977 vdd.n1389 vss 0.00251f
C9978 vdd.n1390 vss 0.00517f
C9979 vdd.n1391 vss 0.00679f
C9980 vdd.n1392 vss 0.00324f
C9981 vdd.n1393 vss 0.00679f
C9982 vdd.n1394 vss 0.00517f
C9983 vdd.n1395 vss 0.00251f
C9984 vdd.n1396 vss 0.00413f
C9985 vdd.n1397 vss 0.0471f
C9986 vdd.t920 vss 0.0471f
C9987 vdd.n1398 vss 0.00425f
C9988 vdd.n1399 vss 0.0424f
C9989 vdd.n1400 vss 0.0132f
C9990 vdd.n1401 vss 0.02f
C9991 vdd.n1402 vss 0.00425f
C9992 vdd.n1403 vss 0.00413f
C9993 vdd.n1404 vss 0.00251f
C9994 vdd.n1405 vss 0.0112f
C9995 vdd.n1406 vss 0.0128f
C9996 vdd.n1407 vss 0.0369f
C9997 vdd.n1408 vss 0.00335f
C9998 vdd.t102 vss 0.0013f
C9999 vdd.n1409 vss 0.0309f
C10000 vdd.n1410 vss 0.0107f
C10001 vdd.n1411 vss 0.0128f
C10002 vdd.n1412 vss 0.0424f
C10003 vdd.t101 vss 0.0471f
C10004 vdd.n1413 vss 0.00324f
C10005 vdd.n1414 vss 0.0471f
C10006 vdd.t1072 vss 0.0471f
C10007 vdd.n1415 vss 0.00413f
C10008 vdd.n1416 vss 0.00324f
C10009 vdd.t1073 vss 0.00134f
C10010 vdd.n1417 vss 0.0393f
C10011 vdd.n1418 vss 0.0128f
C10012 vdd.t1074 vss 0.0471f
C10013 vdd.n1419 vss 0.00324f
C10014 vdd.n1421 vss 0.00925f
C10015 vdd.n1422 vss 0.0471f
C10016 vdd.n1423 vss 0.00324f
C10017 vdd.n1424 vss 0.00413f
C10018 vdd.n1425 vss 0.00324f
C10019 vdd.n1426 vss 0.00679f
C10020 vdd.n1428 vss 0.00925f
C10021 vdd.n1429 vss 0.00425f
C10022 vdd.n1430 vss 0.00413f
C10023 vdd.n1431 vss 0.00251f
C10024 vdd.n1432 vss 0.00517f
C10025 vdd.n1433 vss 0.00679f
C10026 vdd.n1434 vss 0.00324f
C10027 vdd.n1435 vss 0.00679f
C10028 vdd.n1436 vss 0.00517f
C10029 vdd.n1437 vss 0.00251f
C10030 vdd.n1438 vss 0.00413f
C10031 vdd.n1439 vss 0.0471f
C10032 vdd.t1443 vss 0.0471f
C10033 vdd.n1440 vss 0.00425f
C10034 vdd.n1441 vss 0.0424f
C10035 vdd.n1442 vss 0.0132f
C10036 vdd.n1443 vss 0.02f
C10037 vdd.n1444 vss 0.00425f
C10038 vdd.n1445 vss 0.00413f
C10039 vdd.n1446 vss 0.00251f
C10040 vdd.n1447 vss 0.0105f
C10041 vdd.n1448 vss 0.0633f
C10042 vdd.n1449 vss 0.00805f
C10043 vdd.n1450 vss 0.0112f
C10044 vdd.n1451 vss 0.00251f
C10045 vdd.n1452 vss 0.00413f
C10046 vdd.n1453 vss 0.00425f
C10047 vdd.n1454 vss 0.00991f
C10048 vdd.n1455 vss 0.0126f
C10049 vdd.n1456 vss 9.89e-19
C10050 vdd.n1457 vss 0.0011f
C10051 vdd.n1458 vss 0.0271f
C10052 vdd.t410 vss 0.00134f
C10053 vdd.t386 vss 0.0013f
C10054 vdd.n1459 vss 0.032f
C10055 vdd.n1460 vss 0.0393f
C10056 vdd.n1461 vss 0.00324f
C10057 vdd.n1462 vss 0.0112f
C10058 vdd.n1463 vss 0.0128f
C10059 vdd.n1464 vss 0.00413f
C10060 vdd.t408 vss 0.0471f
C10061 vdd.n1465 vss 0.00324f
C10062 vdd.n1467 vss 0.00925f
C10063 vdd.n1468 vss 0.00413f
C10064 vdd.n1469 vss 0.00679f
C10065 vdd.n1470 vss 0.00413f
C10066 vdd.n1471 vss 0.0471f
C10067 vdd.n1472 vss 0.00324f
C10068 vdd.n1473 vss 0.0471f
C10069 vdd.n1474 vss 0.00324f
C10070 vdd.n1475 vss 0.0424f
C10071 vdd.t385 vss 0.0471f
C10072 vdd.n1477 vss 0.00425f
C10073 vdd.n1478 vss 0.00925f
C10074 vdd.n1479 vss 0.0132f
C10075 vdd.n1480 vss 0.00324f
C10076 vdd.n1481 vss 0.0128f
C10077 vdd.n1482 vss 0.02f
C10078 vdd.n1483 vss 0.00425f
C10079 vdd.n1484 vss 0.00413f
C10080 vdd.n1485 vss 0.00251f
C10081 vdd.t409 vss 0.0471f
C10082 vdd.n1486 vss 0.00251f
C10083 vdd.n1487 vss 0.00517f
C10084 vdd.n1488 vss 0.00679f
C10085 vdd.n1489 vss 0.00324f
C10086 vdd.n1490 vss 0.00679f
C10087 vdd.n1491 vss 0.00517f
C10088 vdd.n1492 vss 0.00251f
C10089 vdd.n1493 vss 0.00413f
C10090 vdd.n1494 vss 0.0471f
C10091 vdd.t1447 vss 0.0471f
C10092 vdd.n1495 vss 0.00425f
C10093 vdd.n1496 vss 0.0424f
C10094 vdd.n1497 vss 0.0132f
C10095 vdd.n1498 vss 0.02f
C10096 vdd.n1499 vss 0.00425f
C10097 vdd.n1500 vss 0.00413f
C10098 vdd.n1501 vss 0.00251f
C10099 vdd.n1502 vss 0.0112f
C10100 vdd.n1503 vss 0.0128f
C10101 vdd.n1504 vss 0.0418f
C10102 vdd.t824 vss 0.0013f
C10103 vdd.t1223 vss 0.00134f
C10104 vdd.n1505 vss 0.00324f
C10105 vdd.n1506 vss 0.0112f
C10106 vdd.n1507 vss 0.0128f
C10107 vdd.n1508 vss 0.00413f
C10108 vdd.t1224 vss 0.0471f
C10109 vdd.n1509 vss 0.00324f
C10110 vdd.n1511 vss 0.00925f
C10111 vdd.n1512 vss 0.00413f
C10112 vdd.n1513 vss 0.00679f
C10113 vdd.n1514 vss 0.00413f
C10114 vdd.n1515 vss 0.0471f
C10115 vdd.n1516 vss 0.00324f
C10116 vdd.n1517 vss 0.0471f
C10117 vdd.n1518 vss 0.00324f
C10118 vdd.n1519 vss 0.0424f
C10119 vdd.t823 vss 0.0471f
C10120 vdd.n1521 vss 0.00425f
C10121 vdd.n1522 vss 0.00925f
C10122 vdd.n1523 vss 0.0132f
C10123 vdd.n1524 vss 0.00324f
C10124 vdd.n1525 vss 0.0128f
C10125 vdd.n1526 vss 0.02f
C10126 vdd.n1527 vss 0.00425f
C10127 vdd.n1528 vss 0.00413f
C10128 vdd.n1529 vss 0.00251f
C10129 vdd.t1222 vss 0.0471f
C10130 vdd.n1530 vss 0.00251f
C10131 vdd.n1531 vss 0.00517f
C10132 vdd.n1532 vss 0.00679f
C10133 vdd.n1533 vss 0.00324f
C10134 vdd.n1534 vss 0.00679f
C10135 vdd.n1535 vss 0.00517f
C10136 vdd.n1536 vss 0.00251f
C10137 vdd.n1537 vss 0.00413f
C10138 vdd.n1538 vss 0.0471f
C10139 vdd.t1142 vss 0.0471f
C10140 vdd.n1539 vss 0.00425f
C10141 vdd.n1540 vss 0.0424f
C10142 vdd.n1541 vss 0.0132f
C10143 vdd.n1542 vss 0.02f
C10144 vdd.n1543 vss 0.00425f
C10145 vdd.n1544 vss 0.00413f
C10146 vdd.n1545 vss 0.00251f
C10147 vdd.n1546 vss 0.0112f
C10148 vdd.n1547 vss 0.0128f
C10149 vdd.t1189 vss 0.00134f
C10150 vdd.t834 vss 0.0013f
C10151 vdd.n1548 vss 0.032f
C10152 vdd.n1549 vss 0.0393f
C10153 vdd.n1550 vss 0.00324f
C10154 vdd.n1551 vss 0.0112f
C10155 vdd.n1552 vss 0.0128f
C10156 vdd.n1553 vss 0.00413f
C10157 vdd.t1190 vss 0.0471f
C10158 vdd.n1554 vss 0.00324f
C10159 vdd.n1556 vss 0.00925f
C10160 vdd.n1557 vss 0.00413f
C10161 vdd.n1558 vss 0.00679f
C10162 vdd.n1559 vss 0.00413f
C10163 vdd.n1560 vss 0.0471f
C10164 vdd.n1561 vss 0.00324f
C10165 vdd.n1562 vss 0.0471f
C10166 vdd.n1563 vss 0.00324f
C10167 vdd.n1564 vss 0.0424f
C10168 vdd.t833 vss 0.0471f
C10169 vdd.n1566 vss 0.00425f
C10170 vdd.n1567 vss 0.00925f
C10171 vdd.n1568 vss 0.0132f
C10172 vdd.n1569 vss 0.00324f
C10173 vdd.n1570 vss 0.0128f
C10174 vdd.n1571 vss 0.02f
C10175 vdd.n1572 vss 0.00425f
C10176 vdd.n1573 vss 0.00413f
C10177 vdd.n1574 vss 0.00251f
C10178 vdd.t1188 vss 0.0471f
C10179 vdd.n1575 vss 0.00251f
C10180 vdd.n1576 vss 0.00517f
C10181 vdd.n1577 vss 0.00679f
C10182 vdd.n1578 vss 0.00324f
C10183 vdd.n1579 vss 0.00679f
C10184 vdd.n1580 vss 0.00517f
C10185 vdd.n1581 vss 0.00251f
C10186 vdd.n1582 vss 0.00413f
C10187 vdd.n1583 vss 0.0471f
C10188 vdd.t1121 vss 0.0471f
C10189 vdd.n1584 vss 0.00425f
C10190 vdd.n1585 vss 0.0424f
C10191 vdd.n1586 vss 0.0132f
C10192 vdd.n1587 vss 0.02f
C10193 vdd.n1588 vss 0.00425f
C10194 vdd.n1589 vss 0.00413f
C10195 vdd.n1590 vss 0.00251f
C10196 vdd.n1591 vss 0.0112f
C10197 vdd.n1592 vss 0.0128f
C10198 vdd.n1593 vss 0.119f
C10199 vdd.n1594 vss 0.118f
C10200 vdd.n1595 vss 0.0393f
C10201 vdd.n1596 vss 0.032f
C10202 vdd.n1597 vss 0.0608f
C10203 vdd.t1069 vss 0.00134f
C10204 vdd.t467 vss 0.0013f
C10205 vdd.n1598 vss 0.032f
C10206 vdd.n1599 vss 0.0393f
C10207 vdd.n1600 vss 0.00324f
C10208 vdd.n1601 vss 0.0112f
C10209 vdd.n1602 vss 0.0128f
C10210 vdd.n1603 vss 0.00413f
C10211 vdd.t1070 vss 0.0471f
C10212 vdd.n1604 vss 0.00324f
C10213 vdd.n1606 vss 0.00925f
C10214 vdd.n1607 vss 0.00413f
C10215 vdd.n1608 vss 0.00679f
C10216 vdd.n1609 vss 0.00413f
C10217 vdd.n1610 vss 0.0471f
C10218 vdd.n1611 vss 0.00324f
C10219 vdd.n1612 vss 0.0471f
C10220 vdd.n1613 vss 0.00324f
C10221 vdd.n1614 vss 0.0424f
C10222 vdd.t466 vss 0.0471f
C10223 vdd.n1616 vss 0.00425f
C10224 vdd.n1617 vss 0.00925f
C10225 vdd.n1618 vss 0.0132f
C10226 vdd.n1619 vss 0.00324f
C10227 vdd.n1620 vss 0.0128f
C10228 vdd.n1621 vss 0.02f
C10229 vdd.n1622 vss 0.00425f
C10230 vdd.n1623 vss 0.00413f
C10231 vdd.n1624 vss 0.00251f
C10232 vdd.t1068 vss 0.0471f
C10233 vdd.n1625 vss 0.00251f
C10234 vdd.n1626 vss 0.00517f
C10235 vdd.n1627 vss 0.00679f
C10236 vdd.n1628 vss 0.00324f
C10237 vdd.n1629 vss 0.00679f
C10238 vdd.n1630 vss 0.00517f
C10239 vdd.n1631 vss 0.00251f
C10240 vdd.n1632 vss 0.00413f
C10241 vdd.n1633 vss 0.0471f
C10242 vdd.t1033 vss 0.0471f
C10243 vdd.n1634 vss 0.00425f
C10244 vdd.n1635 vss 0.0424f
C10245 vdd.n1636 vss 0.0132f
C10246 vdd.n1637 vss 0.02f
C10247 vdd.n1638 vss 0.00425f
C10248 vdd.n1639 vss 0.00413f
C10249 vdd.n1640 vss 0.00251f
C10250 vdd.n1641 vss 0.0112f
C10251 vdd.n1642 vss 0.0128f
C10252 vdd.n1643 vss 0.0418f
C10253 vdd.n1644 vss 0.118f
C10254 vdd.n1645 vss 0.121f
C10255 vdd.t999 vss 0.0013f
C10256 vdd.t954 vss 0.00134f
C10257 vdd.n1646 vss 0.00324f
C10258 vdd.n1647 vss 0.0112f
C10259 vdd.n1648 vss 0.0128f
C10260 vdd.n1649 vss 0.00413f
C10261 vdd.t952 vss 0.0471f
C10262 vdd.n1650 vss 0.00324f
C10263 vdd.n1652 vss 0.00925f
C10264 vdd.n1653 vss 0.00413f
C10265 vdd.n1654 vss 0.00679f
C10266 vdd.n1655 vss 0.00413f
C10267 vdd.n1656 vss 0.0471f
C10268 vdd.n1657 vss 0.00324f
C10269 vdd.n1658 vss 0.0471f
C10270 vdd.n1659 vss 0.00324f
C10271 vdd.n1660 vss 0.0424f
C10272 vdd.t998 vss 0.0471f
C10273 vdd.n1662 vss 0.00425f
C10274 vdd.n1663 vss 0.00925f
C10275 vdd.n1664 vss 0.0132f
C10276 vdd.n1665 vss 0.00324f
C10277 vdd.n1666 vss 0.0128f
C10278 vdd.n1667 vss 0.02f
C10279 vdd.n1668 vss 0.00425f
C10280 vdd.n1669 vss 0.00413f
C10281 vdd.n1670 vss 0.00251f
C10282 vdd.t953 vss 0.0471f
C10283 vdd.n1671 vss 0.00251f
C10284 vdd.n1672 vss 0.00517f
C10285 vdd.n1673 vss 0.00679f
C10286 vdd.n1674 vss 0.00324f
C10287 vdd.n1675 vss 0.00679f
C10288 vdd.n1676 vss 0.00517f
C10289 vdd.n1677 vss 0.00251f
C10290 vdd.n1678 vss 0.00413f
C10291 vdd.n1679 vss 0.0471f
C10292 vdd.t309 vss 0.0471f
C10293 vdd.n1680 vss 0.00425f
C10294 vdd.n1681 vss 0.0424f
C10295 vdd.n1682 vss 0.0132f
C10296 vdd.n1683 vss 0.02f
C10297 vdd.n1684 vss 0.00425f
C10298 vdd.n1685 vss 0.00413f
C10299 vdd.n1686 vss 0.00251f
C10300 vdd.n1687 vss 0.0112f
C10301 vdd.n1688 vss 0.0707f
C10302 vdd.n1689 vss 0.0393f
C10303 vdd.n1690 vss 0.032f
C10304 vdd.n1691 vss 0.0608f
C10305 vdd.t84 vss 0.00134f
C10306 vdd.t1494 vss 0.0013f
C10307 vdd.n1692 vss 0.032f
C10308 vdd.n1693 vss 0.0393f
C10309 vdd.n1694 vss 0.00324f
C10310 vdd.n1695 vss 0.0112f
C10311 vdd.n1696 vss 0.0128f
C10312 vdd.n1697 vss 0.00413f
C10313 vdd.t85 vss 0.0471f
C10314 vdd.n1698 vss 0.00324f
C10315 vdd.n1700 vss 0.00925f
C10316 vdd.n1701 vss 0.00413f
C10317 vdd.n1702 vss 0.00679f
C10318 vdd.n1703 vss 0.00413f
C10319 vdd.n1704 vss 0.0471f
C10320 vdd.n1705 vss 0.00324f
C10321 vdd.n1706 vss 0.0471f
C10322 vdd.n1707 vss 0.00324f
C10323 vdd.n1708 vss 0.0424f
C10324 vdd.t1493 vss 0.0471f
C10325 vdd.n1710 vss 0.00425f
C10326 vdd.n1711 vss 0.00925f
C10327 vdd.n1712 vss 0.0132f
C10328 vdd.n1713 vss 0.00324f
C10329 vdd.n1714 vss 0.0128f
C10330 vdd.n1715 vss 0.02f
C10331 vdd.n1716 vss 0.00425f
C10332 vdd.n1717 vss 0.00413f
C10333 vdd.n1718 vss 0.00251f
C10334 vdd.t83 vss 0.0471f
C10335 vdd.n1719 vss 0.00251f
C10336 vdd.n1720 vss 0.00517f
C10337 vdd.n1721 vss 0.00679f
C10338 vdd.n1722 vss 0.00324f
C10339 vdd.n1723 vss 0.00679f
C10340 vdd.n1724 vss 0.00517f
C10341 vdd.n1725 vss 0.00251f
C10342 vdd.n1726 vss 0.00413f
C10343 vdd.n1727 vss 0.0471f
C10344 vdd.t1018 vss 0.0471f
C10345 vdd.n1728 vss 0.00425f
C10346 vdd.n1729 vss 0.0424f
C10347 vdd.n1730 vss 0.0132f
C10348 vdd.n1731 vss 0.02f
C10349 vdd.n1732 vss 0.00425f
C10350 vdd.n1733 vss 0.00413f
C10351 vdd.n1734 vss 0.00251f
C10352 vdd.n1735 vss 0.0112f
C10353 vdd.n1736 vss 0.0128f
C10354 vdd.n1737 vss 0.0418f
C10355 vdd.n1738 vss 0.0912f
C10356 vdd.n1739 vss 0.0824f
C10357 vdd.n1740 vss 0.0567f
C10358 vdd.t871 vss 0.0013f
C10359 vdd.t665 vss 0.00134f
C10360 vdd.n1741 vss 0.00324f
C10361 vdd.n1742 vss 0.0112f
C10362 vdd.n1743 vss 0.0128f
C10363 vdd.n1744 vss 0.00413f
C10364 vdd.t666 vss 0.0471f
C10365 vdd.n1745 vss 0.00324f
C10366 vdd.n1747 vss 0.00925f
C10367 vdd.n1748 vss 0.00413f
C10368 vdd.n1749 vss 0.00679f
C10369 vdd.n1750 vss 0.00413f
C10370 vdd.n1751 vss 0.0471f
C10371 vdd.n1752 vss 0.00324f
C10372 vdd.n1753 vss 0.0471f
C10373 vdd.n1754 vss 0.00324f
C10374 vdd.n1755 vss 0.0424f
C10375 vdd.t870 vss 0.0471f
C10376 vdd.n1757 vss 0.00425f
C10377 vdd.n1758 vss 0.00925f
C10378 vdd.n1759 vss 0.0132f
C10379 vdd.n1760 vss 0.00324f
C10380 vdd.n1761 vss 0.0128f
C10381 vdd.n1762 vss 0.02f
C10382 vdd.n1763 vss 0.00425f
C10383 vdd.n1764 vss 0.00413f
C10384 vdd.n1765 vss 0.00251f
C10385 vdd.t664 vss 0.0471f
C10386 vdd.n1766 vss 0.00251f
C10387 vdd.n1767 vss 0.00517f
C10388 vdd.n1768 vss 0.00679f
C10389 vdd.n1769 vss 0.00324f
C10390 vdd.n1770 vss 0.00679f
C10391 vdd.n1771 vss 0.00517f
C10392 vdd.n1772 vss 0.00251f
C10393 vdd.n1773 vss 0.00413f
C10394 vdd.n1774 vss 0.0471f
C10395 vdd.t683 vss 0.0471f
C10396 vdd.n1775 vss 0.00425f
C10397 vdd.n1776 vss 0.0424f
C10398 vdd.n1777 vss 0.0132f
C10399 vdd.n1778 vss 0.02f
C10400 vdd.n1779 vss 0.00425f
C10401 vdd.n1780 vss 0.00413f
C10402 vdd.n1781 vss 0.00251f
C10403 vdd.n1782 vss 0.0112f
C10404 vdd.n1783 vss 0.0128f
C10405 vdd.t369 vss 0.00134f
C10406 vdd.t171 vss 0.0013f
C10407 vdd.n1784 vss 0.032f
C10408 vdd.n1785 vss 0.0393f
C10409 vdd.n1786 vss 0.00324f
C10410 vdd.n1787 vss 0.0112f
C10411 vdd.n1788 vss 0.0128f
C10412 vdd.n1789 vss 0.00413f
C10413 vdd.t370 vss 0.0471f
C10414 vdd.n1790 vss 0.00324f
C10415 vdd.n1792 vss 0.00925f
C10416 vdd.n1793 vss 0.00413f
C10417 vdd.n1794 vss 0.00679f
C10418 vdd.n1795 vss 0.00413f
C10419 vdd.n1796 vss 0.0471f
C10420 vdd.n1797 vss 0.00324f
C10421 vdd.n1798 vss 0.0471f
C10422 vdd.n1799 vss 0.00324f
C10423 vdd.n1800 vss 0.0424f
C10424 vdd.t170 vss 0.0471f
C10425 vdd.n1802 vss 0.00425f
C10426 vdd.n1803 vss 0.00925f
C10427 vdd.n1804 vss 0.0132f
C10428 vdd.n1805 vss 0.00324f
C10429 vdd.n1806 vss 0.0128f
C10430 vdd.n1807 vss 0.02f
C10431 vdd.n1808 vss 0.00425f
C10432 vdd.n1809 vss 0.00413f
C10433 vdd.n1810 vss 0.00251f
C10434 vdd.t368 vss 0.0471f
C10435 vdd.n1811 vss 0.00251f
C10436 vdd.n1812 vss 0.00517f
C10437 vdd.n1813 vss 0.00679f
C10438 vdd.n1814 vss 0.00324f
C10439 vdd.n1815 vss 0.00679f
C10440 vdd.n1816 vss 0.00517f
C10441 vdd.n1817 vss 0.00251f
C10442 vdd.n1818 vss 0.00413f
C10443 vdd.n1819 vss 0.0471f
C10444 vdd.t132 vss 0.0471f
C10445 vdd.n1820 vss 0.00425f
C10446 vdd.n1821 vss 0.0424f
C10447 vdd.n1822 vss 0.0132f
C10448 vdd.n1823 vss 0.02f
C10449 vdd.n1824 vss 0.00425f
C10450 vdd.n1825 vss 0.00413f
C10451 vdd.n1826 vss 0.00251f
C10452 vdd.n1827 vss 0.0112f
C10453 vdd.n1828 vss 0.0128f
C10454 vdd.n1829 vss 0.0316f
C10455 vdd.t655 vss 0.00134f
C10456 vdd.t1128 vss 0.0013f
C10457 vdd.n1830 vss 0.032f
C10458 vdd.n1831 vss 0.0393f
C10459 vdd.n1832 vss 0.00324f
C10460 vdd.n1833 vss 0.0112f
C10461 vdd.n1834 vss 0.0128f
C10462 vdd.n1835 vss 0.00413f
C10463 vdd.t656 vss 0.0471f
C10464 vdd.n1836 vss 0.00324f
C10465 vdd.n1838 vss 0.00925f
C10466 vdd.n1839 vss 0.00413f
C10467 vdd.n1840 vss 0.00679f
C10468 vdd.n1841 vss 0.00413f
C10469 vdd.n1842 vss 0.0471f
C10470 vdd.n1843 vss 0.00324f
C10471 vdd.n1844 vss 0.0471f
C10472 vdd.n1845 vss 0.00324f
C10473 vdd.n1846 vss 0.0424f
C10474 vdd.t1127 vss 0.0471f
C10475 vdd.n1848 vss 0.00425f
C10476 vdd.n1849 vss 0.00925f
C10477 vdd.n1850 vss 0.0132f
C10478 vdd.n1851 vss 0.00324f
C10479 vdd.n1852 vss 0.0128f
C10480 vdd.n1853 vss 0.02f
C10481 vdd.n1854 vss 0.00425f
C10482 vdd.n1855 vss 0.00413f
C10483 vdd.n1856 vss 0.00251f
C10484 vdd.t654 vss 0.0471f
C10485 vdd.n1857 vss 0.00251f
C10486 vdd.n1858 vss 0.00517f
C10487 vdd.n1859 vss 0.00679f
C10488 vdd.n1860 vss 0.00324f
C10489 vdd.n1861 vss 0.00679f
C10490 vdd.n1862 vss 0.00517f
C10491 vdd.n1863 vss 0.00251f
C10492 vdd.n1864 vss 0.00413f
C10493 vdd.n1865 vss 0.0471f
C10494 vdd.t657 vss 0.0471f
C10495 vdd.n1866 vss 0.00425f
C10496 vdd.n1867 vss 0.0424f
C10497 vdd.n1868 vss 0.0132f
C10498 vdd.n1869 vss 0.02f
C10499 vdd.n1870 vss 0.00425f
C10500 vdd.n1871 vss 0.00413f
C10501 vdd.n1872 vss 0.00251f
C10502 vdd.n1873 vss 0.0112f
C10503 vdd.n1874 vss 0.0128f
C10504 vdd.n1875 vss 0.158f
C10505 vdd.n1876 vss 0.256f
C10506 vdd.n1877 vss 0.0953f
C10507 vdd.n1878 vss 0.0393f
C10508 vdd.n1879 vss 0.032f
C10509 vdd.n1880 vss 0.0608f
C10510 vdd.t788 vss 0.00134f
C10511 vdd.t1325 vss 0.0013f
C10512 vdd.n1881 vss 0.032f
C10513 vdd.n1882 vss 0.0393f
C10514 vdd.n1883 vss 0.00324f
C10515 vdd.n1884 vss 0.0112f
C10516 vdd.n1885 vss 0.0128f
C10517 vdd.n1886 vss 0.00413f
C10518 vdd.t789 vss 0.0471f
C10519 vdd.n1887 vss 0.00324f
C10520 vdd.n1889 vss 0.00925f
C10521 vdd.n1890 vss 0.00413f
C10522 vdd.n1891 vss 0.00679f
C10523 vdd.n1892 vss 0.00413f
C10524 vdd.n1893 vss 0.0471f
C10525 vdd.n1894 vss 0.00324f
C10526 vdd.n1895 vss 0.0471f
C10527 vdd.n1896 vss 0.00324f
C10528 vdd.n1897 vss 0.0424f
C10529 vdd.t1324 vss 0.0471f
C10530 vdd.n1899 vss 0.00425f
C10531 vdd.n1900 vss 0.00925f
C10532 vdd.n1901 vss 0.0132f
C10533 vdd.n1902 vss 0.00324f
C10534 vdd.n1903 vss 0.0128f
C10535 vdd.n1904 vss 0.02f
C10536 vdd.n1905 vss 0.00425f
C10537 vdd.n1906 vss 0.00413f
C10538 vdd.n1907 vss 0.00251f
C10539 vdd.t787 vss 0.0471f
C10540 vdd.n1908 vss 0.00251f
C10541 vdd.n1909 vss 0.00517f
C10542 vdd.n1910 vss 0.00679f
C10543 vdd.n1911 vss 0.00324f
C10544 vdd.n1912 vss 0.00679f
C10545 vdd.n1913 vss 0.00517f
C10546 vdd.n1914 vss 0.00251f
C10547 vdd.n1915 vss 0.00413f
C10548 vdd.n1916 vss 0.0471f
C10549 vdd.t1283 vss 0.0471f
C10550 vdd.n1917 vss 0.00425f
C10551 vdd.n1918 vss 0.0424f
C10552 vdd.n1919 vss 0.0132f
C10553 vdd.n1920 vss 0.02f
C10554 vdd.n1921 vss 0.00425f
C10555 vdd.n1922 vss 0.00413f
C10556 vdd.n1923 vss 0.00251f
C10557 vdd.n1924 vss 0.0112f
C10558 vdd.n1925 vss 0.0128f
C10559 vdd.n1926 vss 0.0418f
C10560 vdd.n1927 vss 0.118f
C10561 vdd.n1928 vss 0.121f
C10562 vdd.t993 vss 0.0013f
C10563 vdd.t389 vss 0.00134f
C10564 vdd.n1929 vss 0.00324f
C10565 vdd.n1930 vss 0.0112f
C10566 vdd.n1931 vss 0.0128f
C10567 vdd.n1932 vss 0.00413f
C10568 vdd.t390 vss 0.0471f
C10569 vdd.n1933 vss 0.00324f
C10570 vdd.n1935 vss 0.00925f
C10571 vdd.n1936 vss 0.00413f
C10572 vdd.n1937 vss 0.00679f
C10573 vdd.n1938 vss 0.00413f
C10574 vdd.n1939 vss 0.0471f
C10575 vdd.n1940 vss 0.00324f
C10576 vdd.n1941 vss 0.0471f
C10577 vdd.n1942 vss 0.00324f
C10578 vdd.n1943 vss 0.0424f
C10579 vdd.t992 vss 0.0471f
C10580 vdd.n1945 vss 0.00425f
C10581 vdd.n1946 vss 0.00925f
C10582 vdd.n1947 vss 0.0132f
C10583 vdd.n1948 vss 0.00324f
C10584 vdd.n1949 vss 0.0128f
C10585 vdd.n1950 vss 0.02f
C10586 vdd.n1951 vss 0.00425f
C10587 vdd.n1952 vss 0.00413f
C10588 vdd.n1953 vss 0.00251f
C10589 vdd.t388 vss 0.0471f
C10590 vdd.n1954 vss 0.00251f
C10591 vdd.n1955 vss 0.00517f
C10592 vdd.n1956 vss 0.00679f
C10593 vdd.n1957 vss 0.00324f
C10594 vdd.n1958 vss 0.00679f
C10595 vdd.n1959 vss 0.00517f
C10596 vdd.n1960 vss 0.00251f
C10597 vdd.n1961 vss 0.00413f
C10598 vdd.n1962 vss 0.0471f
C10599 vdd.t391 vss 0.0471f
C10600 vdd.n1963 vss 0.00425f
C10601 vdd.n1964 vss 0.0424f
C10602 vdd.n1965 vss 0.0132f
C10603 vdd.n1966 vss 0.02f
C10604 vdd.n1967 vss 0.00425f
C10605 vdd.n1968 vss 0.00413f
C10606 vdd.n1969 vss 0.00251f
C10607 vdd.n1970 vss 0.0112f
C10608 vdd.n1971 vss 0.0707f
C10609 vdd.n1972 vss 0.0393f
C10610 vdd.n1973 vss 0.032f
C10611 vdd.n1974 vss 0.0608f
C10612 vdd.t159 vss 0.00134f
C10613 vdd.t372 vss 0.0013f
C10614 vdd.n1975 vss 0.032f
C10615 vdd.n1976 vss 0.0393f
C10616 vdd.n1977 vss 0.00324f
C10617 vdd.n1978 vss 0.0112f
C10618 vdd.n1979 vss 0.0128f
C10619 vdd.n1980 vss 0.00413f
C10620 vdd.t160 vss 0.0471f
C10621 vdd.n1981 vss 0.00324f
C10622 vdd.n1983 vss 0.00925f
C10623 vdd.n1984 vss 0.00413f
C10624 vdd.n1985 vss 0.00679f
C10625 vdd.n1986 vss 0.00413f
C10626 vdd.n1987 vss 0.0471f
C10627 vdd.n1988 vss 0.00324f
C10628 vdd.n1989 vss 0.0471f
C10629 vdd.n1990 vss 0.00324f
C10630 vdd.n1991 vss 0.0424f
C10631 vdd.t371 vss 0.0471f
C10632 vdd.n1993 vss 0.00425f
C10633 vdd.n1994 vss 0.00925f
C10634 vdd.n1995 vss 0.0132f
C10635 vdd.n1996 vss 0.00324f
C10636 vdd.n1997 vss 0.0128f
C10637 vdd.n1998 vss 0.02f
C10638 vdd.n1999 vss 0.00425f
C10639 vdd.n2000 vss 0.00413f
C10640 vdd.n2001 vss 0.00251f
C10641 vdd.t158 vss 0.0471f
C10642 vdd.n2002 vss 0.00251f
C10643 vdd.n2003 vss 0.00517f
C10644 vdd.n2004 vss 0.00679f
C10645 vdd.n2005 vss 0.00324f
C10646 vdd.n2006 vss 0.00679f
C10647 vdd.n2007 vss 0.00517f
C10648 vdd.n2008 vss 0.00251f
C10649 vdd.n2009 vss 0.00413f
C10650 vdd.n2010 vss 0.0471f
C10651 vdd.t268 vss 0.0471f
C10652 vdd.n2011 vss 0.00425f
C10653 vdd.n2012 vss 0.0424f
C10654 vdd.n2013 vss 0.0132f
C10655 vdd.n2014 vss 0.02f
C10656 vdd.n2015 vss 0.00425f
C10657 vdd.n2016 vss 0.00413f
C10658 vdd.n2017 vss 0.00251f
C10659 vdd.n2018 vss 0.0112f
C10660 vdd.n2019 vss 0.0128f
C10661 vdd.n2020 vss 0.0418f
C10662 vdd.n2021 vss 0.118f
C10663 vdd.n2022 vss 0.0935f
C10664 vdd.t972 vss 0.0013f
C10665 vdd.t1219 vss 0.00134f
C10666 vdd.n2023 vss 0.00324f
C10667 vdd.n2024 vss 0.0112f
C10668 vdd.n2025 vss 0.0128f
C10669 vdd.n2026 vss 0.00413f
C10670 vdd.t1217 vss 0.0471f
C10671 vdd.n2027 vss 0.00324f
C10672 vdd.n2029 vss 0.00925f
C10673 vdd.n2030 vss 0.00413f
C10674 vdd.n2031 vss 0.00679f
C10675 vdd.n2032 vss 0.00413f
C10676 vdd.n2033 vss 0.0471f
C10677 vdd.n2034 vss 0.00324f
C10678 vdd.n2035 vss 0.0471f
C10679 vdd.n2036 vss 0.00324f
C10680 vdd.n2037 vss 0.0424f
C10681 vdd.t971 vss 0.0471f
C10682 vdd.n2039 vss 0.00425f
C10683 vdd.n2040 vss 0.00925f
C10684 vdd.n2041 vss 0.0132f
C10685 vdd.n2042 vss 0.00324f
C10686 vdd.n2043 vss 0.0128f
C10687 vdd.n2044 vss 0.02f
C10688 vdd.n2045 vss 0.00425f
C10689 vdd.n2046 vss 0.00413f
C10690 vdd.n2047 vss 0.00251f
C10691 vdd.t1218 vss 0.0471f
C10692 vdd.n2048 vss 0.00251f
C10693 vdd.n2049 vss 0.00517f
C10694 vdd.n2050 vss 0.00679f
C10695 vdd.n2051 vss 0.00324f
C10696 vdd.n2052 vss 0.00679f
C10697 vdd.n2053 vss 0.00517f
C10698 vdd.n2054 vss 0.00251f
C10699 vdd.n2055 vss 0.00413f
C10700 vdd.n2056 vss 0.0471f
C10701 vdd.t1220 vss 0.0471f
C10702 vdd.n2057 vss 0.00425f
C10703 vdd.n2058 vss 0.0424f
C10704 vdd.n2059 vss 0.0132f
C10705 vdd.n2060 vss 0.02f
C10706 vdd.n2061 vss 0.00425f
C10707 vdd.n2062 vss 0.00413f
C10708 vdd.n2063 vss 0.00251f
C10709 vdd.n2064 vss 0.0112f
C10710 vdd.n2065 vss 0.0128f
C10711 vdd.t842 vss 0.00134f
C10712 vdd.t169 vss 0.0013f
C10713 vdd.n2066 vss 0.032f
C10714 vdd.n2067 vss 0.0393f
C10715 vdd.n2068 vss 0.00324f
C10716 vdd.n2069 vss 0.0112f
C10717 vdd.n2070 vss 0.0128f
C10718 vdd.n2071 vss 0.00413f
C10719 vdd.t843 vss 0.0471f
C10720 vdd.n2072 vss 0.00324f
C10721 vdd.n2074 vss 0.00925f
C10722 vdd.n2075 vss 0.00413f
C10723 vdd.n2076 vss 0.00679f
C10724 vdd.n2077 vss 0.00413f
C10725 vdd.n2078 vss 0.0471f
C10726 vdd.n2079 vss 0.00324f
C10727 vdd.n2080 vss 0.0471f
C10728 vdd.n2081 vss 0.00324f
C10729 vdd.n2082 vss 0.0424f
C10730 vdd.t168 vss 0.0471f
C10731 vdd.n2084 vss 0.00425f
C10732 vdd.n2085 vss 0.00925f
C10733 vdd.n2086 vss 0.0132f
C10734 vdd.n2087 vss 0.00324f
C10735 vdd.n2088 vss 0.0128f
C10736 vdd.n2089 vss 0.02f
C10737 vdd.n2090 vss 0.00425f
C10738 vdd.n2091 vss 0.00413f
C10739 vdd.n2092 vss 0.00251f
C10740 vdd.t841 vss 0.0471f
C10741 vdd.n2093 vss 0.00251f
C10742 vdd.n2094 vss 0.00517f
C10743 vdd.n2095 vss 0.00679f
C10744 vdd.n2096 vss 0.00324f
C10745 vdd.n2097 vss 0.00679f
C10746 vdd.n2098 vss 0.00517f
C10747 vdd.n2099 vss 0.00251f
C10748 vdd.n2100 vss 0.00413f
C10749 vdd.n2101 vss 0.0471f
C10750 vdd.t226 vss 0.0471f
C10751 vdd.n2102 vss 0.00425f
C10752 vdd.n2103 vss 0.0424f
C10753 vdd.n2104 vss 0.0132f
C10754 vdd.n2105 vss 0.02f
C10755 vdd.n2106 vss 0.00425f
C10756 vdd.n2107 vss 0.00413f
C10757 vdd.n2108 vss 0.00251f
C10758 vdd.n2109 vss 0.0112f
C10759 vdd.n2110 vss 0.0128f
C10760 vdd.n2111 vss 0.119f
C10761 vdd.n2112 vss 0.118f
C10762 vdd.n2113 vss 0.0393f
C10763 vdd.n2114 vss 0.032f
C10764 vdd.n2115 vss 0.0608f
C10765 vdd.t636 vss 0.00134f
C10766 vdd.t1345 vss 0.0013f
C10767 vdd.n2116 vss 0.032f
C10768 vdd.n2117 vss 0.0393f
C10769 vdd.n2118 vss 0.00324f
C10770 vdd.n2119 vss 0.0112f
C10771 vdd.n2120 vss 0.0128f
C10772 vdd.n2121 vss 0.00413f
C10773 vdd.t637 vss 0.0471f
C10774 vdd.n2122 vss 0.00324f
C10775 vdd.n2124 vss 0.00925f
C10776 vdd.n2125 vss 0.00413f
C10777 vdd.n2126 vss 0.00679f
C10778 vdd.n2127 vss 0.00413f
C10779 vdd.n2128 vss 0.0471f
C10780 vdd.n2129 vss 0.00324f
C10781 vdd.n2130 vss 0.0471f
C10782 vdd.n2131 vss 0.00324f
C10783 vdd.n2132 vss 0.0424f
C10784 vdd.t1344 vss 0.0471f
C10785 vdd.n2134 vss 0.00425f
C10786 vdd.n2135 vss 0.00925f
C10787 vdd.n2136 vss 0.0132f
C10788 vdd.n2137 vss 0.00324f
C10789 vdd.n2138 vss 0.0128f
C10790 vdd.n2139 vss 0.02f
C10791 vdd.n2140 vss 0.00425f
C10792 vdd.n2141 vss 0.00413f
C10793 vdd.n2142 vss 0.00251f
C10794 vdd.t635 vss 0.0471f
C10795 vdd.n2143 vss 0.00251f
C10796 vdd.n2144 vss 0.00517f
C10797 vdd.n2145 vss 0.00679f
C10798 vdd.n2146 vss 0.00324f
C10799 vdd.n2147 vss 0.00679f
C10800 vdd.n2148 vss 0.00517f
C10801 vdd.n2149 vss 0.00251f
C10802 vdd.n2150 vss 0.00413f
C10803 vdd.n2151 vss 0.0471f
C10804 vdd.t110 vss 0.0471f
C10805 vdd.n2152 vss 0.00425f
C10806 vdd.n2153 vss 0.0424f
C10807 vdd.n2154 vss 0.0132f
C10808 vdd.n2155 vss 0.02f
C10809 vdd.n2156 vss 0.00425f
C10810 vdd.n2157 vss 0.00413f
C10811 vdd.n2158 vss 0.00251f
C10812 vdd.n2159 vss 0.0112f
C10813 vdd.n2160 vss 0.0128f
C10814 vdd.n2161 vss 0.0418f
C10815 vdd.n2162 vss 0.118f
C10816 vdd.n2163 vss 0.121f
C10817 vdd.t941 vss 0.0013f
C10818 vdd.t233 vss 0.00134f
C10819 vdd.n2164 vss 0.00324f
C10820 vdd.n2165 vss 0.0112f
C10821 vdd.n2166 vss 0.0128f
C10822 vdd.n2167 vss 0.00413f
C10823 vdd.t231 vss 0.0471f
C10824 vdd.n2168 vss 0.00324f
C10825 vdd.n2170 vss 0.00925f
C10826 vdd.n2171 vss 0.00413f
C10827 vdd.n2172 vss 0.00679f
C10828 vdd.n2173 vss 0.00413f
C10829 vdd.n2174 vss 0.0471f
C10830 vdd.n2175 vss 0.00324f
C10831 vdd.n2176 vss 0.0471f
C10832 vdd.n2177 vss 0.00324f
C10833 vdd.n2178 vss 0.0424f
C10834 vdd.t940 vss 0.0471f
C10835 vdd.n2180 vss 0.00425f
C10836 vdd.n2181 vss 0.00925f
C10837 vdd.n2182 vss 0.0132f
C10838 vdd.n2183 vss 0.00324f
C10839 vdd.n2184 vss 0.0128f
C10840 vdd.n2185 vss 0.02f
C10841 vdd.n2186 vss 0.00425f
C10842 vdd.n2187 vss 0.00413f
C10843 vdd.n2188 vss 0.00251f
C10844 vdd.t232 vss 0.0471f
C10845 vdd.n2189 vss 0.00251f
C10846 vdd.n2190 vss 0.00517f
C10847 vdd.n2191 vss 0.00679f
C10848 vdd.n2192 vss 0.00324f
C10849 vdd.n2193 vss 0.00679f
C10850 vdd.n2194 vss 0.00517f
C10851 vdd.n2195 vss 0.00251f
C10852 vdd.n2196 vss 0.00413f
C10853 vdd.n2197 vss 0.0471f
C10854 vdd.t1131 vss 0.0471f
C10855 vdd.n2198 vss 0.00425f
C10856 vdd.n2199 vss 0.0424f
C10857 vdd.n2200 vss 0.0132f
C10858 vdd.n2201 vss 0.02f
C10859 vdd.n2202 vss 0.00425f
C10860 vdd.n2203 vss 0.00413f
C10861 vdd.n2204 vss 0.00251f
C10862 vdd.n2205 vss 0.0112f
C10863 vdd.n2206 vss 0.0707f
C10864 vdd.n2207 vss 0.0393f
C10865 vdd.n2208 vss 0.032f
C10866 vdd.n2209 vss 0.0608f
C10867 vdd.t1117 vss 0.00134f
C10868 vdd.t1482 vss 0.0013f
C10869 vdd.n2210 vss 0.032f
C10870 vdd.n2211 vss 0.0393f
C10871 vdd.n2212 vss 0.00324f
C10872 vdd.n2213 vss 0.0112f
C10873 vdd.n2214 vss 0.0128f
C10874 vdd.n2215 vss 0.00413f
C10875 vdd.t1118 vss 0.0471f
C10876 vdd.n2216 vss 0.00324f
C10877 vdd.n2218 vss 0.00925f
C10878 vdd.n2219 vss 0.00413f
C10879 vdd.n2220 vss 0.00679f
C10880 vdd.n2221 vss 0.00413f
C10881 vdd.n2222 vss 0.0471f
C10882 vdd.n2223 vss 0.00324f
C10883 vdd.n2224 vss 0.0471f
C10884 vdd.n2225 vss 0.00324f
C10885 vdd.n2226 vss 0.0424f
C10886 vdd.t1481 vss 0.0471f
C10887 vdd.n2228 vss 0.00425f
C10888 vdd.n2229 vss 0.00925f
C10889 vdd.n2230 vss 0.0132f
C10890 vdd.n2231 vss 0.00324f
C10891 vdd.n2232 vss 0.0128f
C10892 vdd.n2233 vss 0.02f
C10893 vdd.n2234 vss 0.00425f
C10894 vdd.n2235 vss 0.00413f
C10895 vdd.n2236 vss 0.00251f
C10896 vdd.t1116 vss 0.0471f
C10897 vdd.n2237 vss 0.00251f
C10898 vdd.n2238 vss 0.00517f
C10899 vdd.n2239 vss 0.00679f
C10900 vdd.n2240 vss 0.00324f
C10901 vdd.n2241 vss 0.00679f
C10902 vdd.n2242 vss 0.00517f
C10903 vdd.n2243 vss 0.00251f
C10904 vdd.n2244 vss 0.00413f
C10905 vdd.n2245 vss 0.0471f
C10906 vdd.t1119 vss 0.0471f
C10907 vdd.n2246 vss 0.00425f
C10908 vdd.n2247 vss 0.0424f
C10909 vdd.n2248 vss 0.0132f
C10910 vdd.n2249 vss 0.02f
C10911 vdd.n2250 vss 0.00425f
C10912 vdd.n2251 vss 0.00413f
C10913 vdd.n2252 vss 0.00251f
C10914 vdd.n2253 vss 0.0112f
C10915 vdd.n2254 vss 0.0128f
C10916 vdd.n2255 vss 0.0418f
C10917 vdd.n2256 vss 0.0912f
C10918 vdd.n2257 vss 0.0824f
C10919 vdd.n2258 vss 0.0567f
C10920 vdd.t901 vss 0.0013f
C10921 vdd.t297 vss 0.00134f
C10922 vdd.n2259 vss 0.00324f
C10923 vdd.n2260 vss 0.0112f
C10924 vdd.n2261 vss 0.0128f
C10925 vdd.n2262 vss 0.00413f
C10926 vdd.t298 vss 0.0471f
C10927 vdd.n2263 vss 0.00324f
C10928 vdd.n2265 vss 0.00925f
C10929 vdd.n2266 vss 0.00413f
C10930 vdd.n2267 vss 0.00679f
C10931 vdd.n2268 vss 0.00413f
C10932 vdd.n2269 vss 0.0471f
C10933 vdd.n2270 vss 0.00324f
C10934 vdd.n2271 vss 0.0471f
C10935 vdd.n2272 vss 0.00324f
C10936 vdd.n2273 vss 0.0424f
C10937 vdd.t900 vss 0.0471f
C10938 vdd.n2275 vss 0.00425f
C10939 vdd.n2276 vss 0.00925f
C10940 vdd.n2277 vss 0.0132f
C10941 vdd.n2278 vss 0.00324f
C10942 vdd.n2279 vss 0.0128f
C10943 vdd.n2280 vss 0.02f
C10944 vdd.n2281 vss 0.00425f
C10945 vdd.n2282 vss 0.00413f
C10946 vdd.n2283 vss 0.00251f
C10947 vdd.t296 vss 0.0471f
C10948 vdd.n2284 vss 0.00251f
C10949 vdd.n2285 vss 0.00517f
C10950 vdd.n2286 vss 0.00679f
C10951 vdd.n2287 vss 0.00324f
C10952 vdd.n2288 vss 0.00679f
C10953 vdd.n2289 vss 0.00517f
C10954 vdd.n2290 vss 0.00251f
C10955 vdd.n2291 vss 0.00413f
C10956 vdd.n2292 vss 0.0471f
C10957 vdd.t929 vss 0.0471f
C10958 vdd.n2293 vss 0.00425f
C10959 vdd.n2294 vss 0.0424f
C10960 vdd.n2295 vss 0.0132f
C10961 vdd.n2296 vss 0.02f
C10962 vdd.n2297 vss 0.00425f
C10963 vdd.n2298 vss 0.00413f
C10964 vdd.n2299 vss 0.00251f
C10965 vdd.n2300 vss 0.0112f
C10966 vdd.n2301 vss 0.0128f
C10967 vdd.t117 vss 0.00134f
C10968 vdd.t772 vss 0.0013f
C10969 vdd.n2302 vss 0.032f
C10970 vdd.n2303 vss 0.0393f
C10971 vdd.n2304 vss 0.00324f
C10972 vdd.n2305 vss 0.0112f
C10973 vdd.n2306 vss 0.0128f
C10974 vdd.n2307 vss 0.00413f
C10975 vdd.t118 vss 0.0471f
C10976 vdd.n2308 vss 0.00324f
C10977 vdd.n2310 vss 0.00925f
C10978 vdd.n2311 vss 0.00413f
C10979 vdd.n2312 vss 0.00679f
C10980 vdd.n2313 vss 0.00413f
C10981 vdd.n2314 vss 0.0471f
C10982 vdd.n2315 vss 0.00324f
C10983 vdd.n2316 vss 0.0471f
C10984 vdd.n2317 vss 0.00324f
C10985 vdd.n2318 vss 0.0424f
C10986 vdd.t771 vss 0.0471f
C10987 vdd.n2320 vss 0.00425f
C10988 vdd.n2321 vss 0.00925f
C10989 vdd.n2322 vss 0.0132f
C10990 vdd.n2323 vss 0.00324f
C10991 vdd.n2324 vss 0.0128f
C10992 vdd.n2325 vss 0.02f
C10993 vdd.n2326 vss 0.00425f
C10994 vdd.n2327 vss 0.00413f
C10995 vdd.n2328 vss 0.00251f
C10996 vdd.t116 vss 0.0471f
C10997 vdd.n2329 vss 0.00251f
C10998 vdd.n2330 vss 0.00517f
C10999 vdd.n2331 vss 0.00679f
C11000 vdd.n2332 vss 0.00324f
C11001 vdd.n2333 vss 0.00679f
C11002 vdd.n2334 vss 0.00517f
C11003 vdd.n2335 vss 0.00251f
C11004 vdd.n2336 vss 0.00413f
C11005 vdd.n2337 vss 0.0471f
C11006 vdd.t516 vss 0.0471f
C11007 vdd.n2338 vss 0.00425f
C11008 vdd.n2339 vss 0.0424f
C11009 vdd.n2340 vss 0.0132f
C11010 vdd.n2341 vss 0.02f
C11011 vdd.n2342 vss 0.00425f
C11012 vdd.n2343 vss 0.00413f
C11013 vdd.n2344 vss 0.00251f
C11014 vdd.n2345 vss 0.0112f
C11015 vdd.n2346 vss 0.0128f
C11016 vdd.n2347 vss 0.119f
C11017 vdd.n2348 vss 0.118f
C11018 vdd.n2349 vss 0.0393f
C11019 vdd.n2350 vss 0.032f
C11020 vdd.n2351 vss 0.0608f
C11021 vdd.t1039 vss 0.00134f
C11022 vdd.t493 vss 0.0013f
C11023 vdd.n2352 vss 0.032f
C11024 vdd.n2353 vss 0.0393f
C11025 vdd.n2354 vss 0.00324f
C11026 vdd.n2355 vss 0.0112f
C11027 vdd.n2356 vss 0.0128f
C11028 vdd.n2357 vss 0.00413f
C11029 vdd.t1040 vss 0.0471f
C11030 vdd.n2358 vss 0.00324f
C11031 vdd.n2360 vss 0.00925f
C11032 vdd.n2361 vss 0.00413f
C11033 vdd.n2362 vss 0.00679f
C11034 vdd.n2363 vss 0.00413f
C11035 vdd.n2364 vss 0.0471f
C11036 vdd.n2365 vss 0.00324f
C11037 vdd.n2366 vss 0.0471f
C11038 vdd.n2367 vss 0.00324f
C11039 vdd.n2368 vss 0.0424f
C11040 vdd.t492 vss 0.0471f
C11041 vdd.n2370 vss 0.00425f
C11042 vdd.n2371 vss 0.00925f
C11043 vdd.n2372 vss 0.0132f
C11044 vdd.n2373 vss 0.00324f
C11045 vdd.n2374 vss 0.0128f
C11046 vdd.n2375 vss 0.02f
C11047 vdd.n2376 vss 0.00425f
C11048 vdd.n2377 vss 0.00413f
C11049 vdd.n2378 vss 0.00251f
C11050 vdd.t1038 vss 0.0471f
C11051 vdd.n2379 vss 0.00251f
C11052 vdd.n2380 vss 0.00517f
C11053 vdd.n2381 vss 0.00679f
C11054 vdd.n2382 vss 0.00324f
C11055 vdd.n2383 vss 0.00679f
C11056 vdd.n2384 vss 0.00517f
C11057 vdd.n2385 vss 0.00251f
C11058 vdd.n2386 vss 0.00413f
C11059 vdd.n2387 vss 0.0471f
C11060 vdd.t103 vss 0.0471f
C11061 vdd.n2388 vss 0.00425f
C11062 vdd.n2389 vss 0.0424f
C11063 vdd.n2390 vss 0.0132f
C11064 vdd.n2391 vss 0.02f
C11065 vdd.n2392 vss 0.00425f
C11066 vdd.n2393 vss 0.00413f
C11067 vdd.n2394 vss 0.00251f
C11068 vdd.n2395 vss 0.0112f
C11069 vdd.n2396 vss 0.0128f
C11070 vdd.n2397 vss 0.0418f
C11071 vdd.n2398 vss 0.118f
C11072 vdd.n2399 vss 0.121f
C11073 vdd.t976 vss 0.0013f
C11074 vdd.t876 vss 0.00134f
C11075 vdd.n2400 vss 0.00324f
C11076 vdd.n2401 vss 0.0112f
C11077 vdd.n2402 vss 0.0128f
C11078 vdd.n2403 vss 0.00413f
C11079 vdd.t877 vss 0.0471f
C11080 vdd.n2404 vss 0.00324f
C11081 vdd.n2406 vss 0.00925f
C11082 vdd.n2407 vss 0.00413f
C11083 vdd.n2408 vss 0.00679f
C11084 vdd.n2409 vss 0.00413f
C11085 vdd.n2410 vss 0.0471f
C11086 vdd.n2411 vss 0.00324f
C11087 vdd.n2412 vss 0.0471f
C11088 vdd.n2413 vss 0.00324f
C11089 vdd.n2414 vss 0.0424f
C11090 vdd.t975 vss 0.0471f
C11091 vdd.n2416 vss 0.00425f
C11092 vdd.n2417 vss 0.00925f
C11093 vdd.n2418 vss 0.0132f
C11094 vdd.n2419 vss 0.00324f
C11095 vdd.n2420 vss 0.0128f
C11096 vdd.n2421 vss 0.02f
C11097 vdd.n2422 vss 0.00425f
C11098 vdd.n2423 vss 0.00413f
C11099 vdd.n2424 vss 0.00251f
C11100 vdd.t875 vss 0.0471f
C11101 vdd.n2425 vss 0.00251f
C11102 vdd.n2426 vss 0.00517f
C11103 vdd.n2427 vss 0.00679f
C11104 vdd.n2428 vss 0.00324f
C11105 vdd.n2429 vss 0.00679f
C11106 vdd.n2430 vss 0.00517f
C11107 vdd.n2431 vss 0.00251f
C11108 vdd.n2432 vss 0.00413f
C11109 vdd.n2433 vss 0.0471f
C11110 vdd.t606 vss 0.0471f
C11111 vdd.n2434 vss 0.00425f
C11112 vdd.n2435 vss 0.0424f
C11113 vdd.n2436 vss 0.0132f
C11114 vdd.n2437 vss 0.02f
C11115 vdd.n2438 vss 0.00425f
C11116 vdd.n2439 vss 0.00413f
C11117 vdd.n2440 vss 0.00251f
C11118 vdd.n2441 vss 0.0112f
C11119 vdd.n2442 vss 0.0707f
C11120 vdd.n2443 vss 0.0393f
C11121 vdd.n2444 vss 0.032f
C11122 vdd.n2445 vss 0.0608f
C11123 vdd.t1445 vss 0.00134f
C11124 vdd.t1349 vss 0.0013f
C11125 vdd.n2446 vss 0.032f
C11126 vdd.n2447 vss 0.0393f
C11127 vdd.n2448 vss 0.00324f
C11128 vdd.n2449 vss 0.0112f
C11129 vdd.n2450 vss 0.0128f
C11130 vdd.n2451 vss 0.00413f
C11131 vdd.t1446 vss 0.0471f
C11132 vdd.n2452 vss 0.00324f
C11133 vdd.n2454 vss 0.00925f
C11134 vdd.n2455 vss 0.00413f
C11135 vdd.n2456 vss 0.00679f
C11136 vdd.n2457 vss 0.00413f
C11137 vdd.n2458 vss 0.0471f
C11138 vdd.n2459 vss 0.00324f
C11139 vdd.n2460 vss 0.0471f
C11140 vdd.n2461 vss 0.00324f
C11141 vdd.n2462 vss 0.0424f
C11142 vdd.t1348 vss 0.0471f
C11143 vdd.n2464 vss 0.00425f
C11144 vdd.n2465 vss 0.00925f
C11145 vdd.n2466 vss 0.0132f
C11146 vdd.n2467 vss 0.00324f
C11147 vdd.n2468 vss 0.0128f
C11148 vdd.n2469 vss 0.02f
C11149 vdd.n2470 vss 0.00425f
C11150 vdd.n2471 vss 0.00413f
C11151 vdd.n2472 vss 0.00251f
C11152 vdd.t1444 vss 0.0471f
C11153 vdd.n2473 vss 0.00251f
C11154 vdd.n2474 vss 0.00517f
C11155 vdd.n2475 vss 0.00679f
C11156 vdd.n2476 vss 0.00324f
C11157 vdd.n2477 vss 0.00679f
C11158 vdd.n2478 vss 0.00517f
C11159 vdd.n2479 vss 0.00251f
C11160 vdd.n2480 vss 0.00413f
C11161 vdd.n2481 vss 0.0471f
C11162 vdd.t1423 vss 0.0471f
C11163 vdd.n2482 vss 0.00425f
C11164 vdd.n2483 vss 0.0424f
C11165 vdd.n2484 vss 0.0132f
C11166 vdd.n2485 vss 0.02f
C11167 vdd.n2486 vss 0.00425f
C11168 vdd.n2487 vss 0.00413f
C11169 vdd.n2488 vss 0.00251f
C11170 vdd.n2489 vss 0.0112f
C11171 vdd.n2490 vss 0.0128f
C11172 vdd.n2491 vss 0.0418f
C11173 vdd.n2492 vss 0.299f
C11174 vdd.n2493 vss 0.00324f
C11175 vdd.n2494 vss 0.0112f
C11176 vdd.n2495 vss 0.0128f
C11177 vdd.n2496 vss 0.00413f
C11178 vdd.n2497 vss 0.00413f
C11179 vdd.n2498 vss 0.0471f
C11180 vdd.n2499 vss 0.00251f
C11181 vdd.t381 vss 0.0471f
C11182 vdd.n2500 vss 0.00324f
C11183 vdd.n2502 vss 0.00679f
C11184 vdd.n2503 vss 0.00413f
C11185 vdd.n2504 vss 0.00324f
C11186 vdd.n2505 vss 0.00413f
C11187 vdd.n2506 vss 0.0471f
C11188 vdd.n2507 vss 0.00324f
C11189 vdd.n2509 vss 0.00925f
C11190 vdd.t1213 vss 0.0471f
C11191 vdd.n2510 vss 0.00425f
C11192 vdd.n2511 vss 0.0424f
C11193 vdd.n2512 vss 0.0132f
C11194 vdd.n2513 vss 0.00324f
C11195 vdd.n2514 vss 0.0128f
C11196 vdd.n2515 vss 0.02f
C11197 vdd.n2516 vss 0.00425f
C11198 vdd.n2517 vss 0.00413f
C11199 vdd.n2518 vss 0.00251f
C11200 vdd.t181 vss 0.0471f
C11201 vdd.n2519 vss 0.00251f
C11202 vdd.n2520 vss 0.00517f
C11203 vdd.n2521 vss 0.00679f
C11204 vdd.n2522 vss 0.00517f
C11205 vdd.n2523 vss 0.00679f
C11206 vdd.n2524 vss 0.02f
C11207 vdd.n2525 vss 0.00425f
C11208 vdd.n2526 vss 0.0424f
C11209 vdd.n2527 vss 0.0132f
C11210 vdd.n2528 vss 0.00925f
C11211 vdd.n2529 vss 0.00425f
C11212 vdd.n2530 vss 0.00413f
C11213 vdd.n2531 vss 0.00324f
C11214 vdd.n2532 vss 0.0471f
C11215 vdd.t179 vss 0.0471f
C11216 vdd.n2533 vss 0.00251f
C11217 vdd.n2534 vss 0.0112f
C11218 vdd.n2535 vss 0.0128f
C11219 vdd.t180 vss 0.00134f
C11220 vdd.t382 vss 0.0013f
C11221 vdd.n2536 vss 0.0332f
C11222 vdd.n2537 vss 0.0393f
C11223 vdd.n2538 vss 0.0345f
C11224 vdd.n2539 vss 0.262f
C11225 vdd.t816 vss 0.0013f
C11226 vdd.t525 vss 0.00134f
C11227 vdd.n2540 vss 0.00324f
C11228 vdd.n2541 vss 0.0112f
C11229 vdd.n2542 vss 0.0128f
C11230 vdd.n2543 vss 0.00413f
C11231 vdd.n2544 vss 0.00413f
C11232 vdd.n2545 vss 0.0471f
C11233 vdd.n2546 vss 0.00251f
C11234 vdd.t769 vss 0.0471f
C11235 vdd.n2547 vss 0.00324f
C11236 vdd.n2549 vss 0.00679f
C11237 vdd.n2550 vss 0.00413f
C11238 vdd.n2551 vss 0.00324f
C11239 vdd.n2552 vss 0.00413f
C11240 vdd.n2553 vss 0.0471f
C11241 vdd.n2554 vss 0.00324f
C11242 vdd.n2556 vss 0.00925f
C11243 vdd.t1027 vss 0.0471f
C11244 vdd.n2557 vss 0.00425f
C11245 vdd.n2558 vss 0.0424f
C11246 vdd.n2559 vss 0.0132f
C11247 vdd.n2560 vss 0.00324f
C11248 vdd.n2561 vss 0.0128f
C11249 vdd.n2562 vss 0.02f
C11250 vdd.n2563 vss 0.00425f
C11251 vdd.n2564 vss 0.00413f
C11252 vdd.n2565 vss 0.00251f
C11253 vdd.t334 vss 0.0471f
C11254 vdd.n2566 vss 0.00251f
C11255 vdd.n2567 vss 0.00517f
C11256 vdd.n2568 vss 0.00679f
C11257 vdd.n2569 vss 0.00517f
C11258 vdd.n2570 vss 0.00679f
C11259 vdd.n2571 vss 0.02f
C11260 vdd.n2572 vss 0.00425f
C11261 vdd.n2573 vss 0.0424f
C11262 vdd.n2574 vss 0.0132f
C11263 vdd.n2575 vss 0.00925f
C11264 vdd.n2576 vss 0.00425f
C11265 vdd.n2577 vss 0.00413f
C11266 vdd.n2578 vss 0.00324f
C11267 vdd.n2579 vss 0.0471f
C11268 vdd.t332 vss 0.0471f
C11269 vdd.n2580 vss 0.00251f
C11270 vdd.n2581 vss 0.0112f
C11271 vdd.n2582 vss 0.0128f
C11272 vdd.t333 vss 0.00134f
C11273 vdd.t770 vss 0.0013f
C11274 vdd.n2583 vss 0.0332f
C11275 vdd.n2584 vss 0.0393f
C11276 vdd.n2585 vss 0.119f
C11277 vdd.n2586 vss 0.00324f
C11278 vdd.n2587 vss 0.0112f
C11279 vdd.n2588 vss 0.0128f
C11280 vdd.n2589 vss 0.00413f
C11281 vdd.n2590 vss 0.00413f
C11282 vdd.n2591 vss 0.0471f
C11283 vdd.n2592 vss 0.00251f
C11284 vdd.t815 vss 0.0471f
C11285 vdd.n2593 vss 0.00324f
C11286 vdd.n2595 vss 0.00679f
C11287 vdd.n2596 vss 0.00413f
C11288 vdd.n2597 vss 0.00324f
C11289 vdd.n2598 vss 0.00413f
C11290 vdd.n2599 vss 0.0471f
C11291 vdd.n2600 vss 0.00324f
C11292 vdd.n2602 vss 0.00925f
C11293 vdd.t423 vss 0.0471f
C11294 vdd.n2603 vss 0.00425f
C11295 vdd.n2604 vss 0.0424f
C11296 vdd.n2605 vss 0.0132f
C11297 vdd.n2606 vss 0.00324f
C11298 vdd.n2607 vss 0.0128f
C11299 vdd.n2608 vss 0.02f
C11300 vdd.n2609 vss 0.00425f
C11301 vdd.n2610 vss 0.00413f
C11302 vdd.n2611 vss 0.00251f
C11303 vdd.t526 vss 0.0471f
C11304 vdd.n2612 vss 0.00251f
C11305 vdd.n2613 vss 0.00517f
C11306 vdd.n2614 vss 0.00679f
C11307 vdd.n2615 vss 0.00517f
C11308 vdd.n2616 vss 0.00679f
C11309 vdd.n2617 vss 0.02f
C11310 vdd.n2618 vss 0.00425f
C11311 vdd.n2619 vss 0.0424f
C11312 vdd.n2620 vss 0.0132f
C11313 vdd.n2621 vss 0.00925f
C11314 vdd.n2622 vss 0.00425f
C11315 vdd.n2623 vss 0.00413f
C11316 vdd.n2624 vss 0.00324f
C11317 vdd.n2625 vss 0.0471f
C11318 vdd.t524 vss 0.0471f
C11319 vdd.n2626 vss 0.00251f
C11320 vdd.n2627 vss 0.0112f
C11321 vdd.n2628 vss 0.0128f
C11322 vdd.n2629 vss 0.118f
C11323 vdd.n2630 vss 0.0393f
C11324 vdd.n2631 vss 0.0332f
C11325 vdd.n2632 vss 0.0596f
C11326 vdd.n2633 vss 0.00324f
C11327 vdd.n2634 vss 0.0112f
C11328 vdd.n2635 vss 0.0128f
C11329 vdd.n2636 vss 0.00413f
C11330 vdd.n2637 vss 0.00413f
C11331 vdd.n2638 vss 0.0471f
C11332 vdd.n2639 vss 0.00251f
C11333 vdd.t1350 vss 0.0471f
C11334 vdd.n2640 vss 0.00324f
C11335 vdd.n2642 vss 0.00679f
C11336 vdd.n2643 vss 0.00413f
C11337 vdd.n2644 vss 0.00324f
C11338 vdd.n2645 vss 0.00413f
C11339 vdd.n2646 vss 0.0471f
C11340 vdd.n2647 vss 0.00324f
C11341 vdd.n2649 vss 0.00925f
C11342 vdd.t916 vss 0.0471f
C11343 vdd.n2650 vss 0.00425f
C11344 vdd.n2651 vss 0.0424f
C11345 vdd.n2652 vss 0.0132f
C11346 vdd.n2653 vss 0.00324f
C11347 vdd.n2654 vss 0.0128f
C11348 vdd.n2655 vss 0.02f
C11349 vdd.n2656 vss 0.00425f
C11350 vdd.n2657 vss 0.00413f
C11351 vdd.n2658 vss 0.00251f
C11352 vdd.t618 vss 0.0471f
C11353 vdd.n2659 vss 0.00251f
C11354 vdd.n2660 vss 0.00517f
C11355 vdd.n2661 vss 0.00679f
C11356 vdd.n2662 vss 0.00517f
C11357 vdd.n2663 vss 0.00679f
C11358 vdd.n2664 vss 0.02f
C11359 vdd.n2665 vss 0.00425f
C11360 vdd.n2666 vss 0.0424f
C11361 vdd.n2667 vss 0.0132f
C11362 vdd.n2668 vss 0.00925f
C11363 vdd.n2669 vss 0.00425f
C11364 vdd.n2670 vss 0.00413f
C11365 vdd.n2671 vss 0.00324f
C11366 vdd.n2672 vss 0.0471f
C11367 vdd.t616 vss 0.0471f
C11368 vdd.n2673 vss 0.00251f
C11369 vdd.n2674 vss 0.0112f
C11370 vdd.n2675 vss 0.0128f
C11371 vdd.t617 vss 0.00134f
C11372 vdd.t1351 vss 0.0013f
C11373 vdd.n2676 vss 0.0332f
C11374 vdd.n2677 vss 0.0393f
C11375 vdd.n2678 vss 0.0418f
C11376 vdd.n2679 vss 0.118f
C11377 vdd.n2680 vss 0.121f
C11378 vdd.t1017 vss 0.0013f
C11379 vdd.t1097 vss 0.00134f
C11380 vdd.n2681 vss 0.00324f
C11381 vdd.n2682 vss 0.0112f
C11382 vdd.n2683 vss 0.0128f
C11383 vdd.n2684 vss 0.00413f
C11384 vdd.n2685 vss 0.00413f
C11385 vdd.n2686 vss 0.0471f
C11386 vdd.n2687 vss 0.00251f
C11387 vdd.t1016 vss 0.0471f
C11388 vdd.n2688 vss 0.00324f
C11389 vdd.n2690 vss 0.00679f
C11390 vdd.n2691 vss 0.00413f
C11391 vdd.n2692 vss 0.00324f
C11392 vdd.n2693 vss 0.00413f
C11393 vdd.n2694 vss 0.0471f
C11394 vdd.n2695 vss 0.00324f
C11395 vdd.n2697 vss 0.00925f
C11396 vdd.t717 vss 0.0471f
C11397 vdd.n2698 vss 0.00425f
C11398 vdd.n2699 vss 0.0424f
C11399 vdd.n2700 vss 0.0132f
C11400 vdd.n2701 vss 0.00324f
C11401 vdd.n2702 vss 0.0128f
C11402 vdd.n2703 vss 0.02f
C11403 vdd.n2704 vss 0.00425f
C11404 vdd.n2705 vss 0.00413f
C11405 vdd.n2706 vss 0.00251f
C11406 vdd.t1098 vss 0.0471f
C11407 vdd.n2707 vss 0.00251f
C11408 vdd.n2708 vss 0.00517f
C11409 vdd.n2709 vss 0.00679f
C11410 vdd.n2710 vss 0.00517f
C11411 vdd.n2711 vss 0.00679f
C11412 vdd.n2712 vss 0.02f
C11413 vdd.n2713 vss 0.00425f
C11414 vdd.n2714 vss 0.0424f
C11415 vdd.n2715 vss 0.0132f
C11416 vdd.n2716 vss 0.00925f
C11417 vdd.n2717 vss 0.00425f
C11418 vdd.n2718 vss 0.00413f
C11419 vdd.n2719 vss 0.00324f
C11420 vdd.n2720 vss 0.0471f
C11421 vdd.t1096 vss 0.0471f
C11422 vdd.n2721 vss 0.00251f
C11423 vdd.n2722 vss 0.0112f
C11424 vdd.n2723 vss 0.0707f
C11425 vdd.n2724 vss 0.0393f
C11426 vdd.n2725 vss 0.0332f
C11427 vdd.n2726 vss 0.0596f
C11428 vdd.n2727 vss 0.00324f
C11429 vdd.n2728 vss 0.0112f
C11430 vdd.n2729 vss 0.0128f
C11431 vdd.n2730 vss 0.00413f
C11432 vdd.n2731 vss 0.00413f
C11433 vdd.n2732 vss 0.0471f
C11434 vdd.n2733 vss 0.00251f
C11435 vdd.t494 vss 0.0471f
C11436 vdd.n2734 vss 0.00324f
C11437 vdd.n2736 vss 0.00679f
C11438 vdd.n2737 vss 0.00413f
C11439 vdd.n2738 vss 0.00324f
C11440 vdd.n2739 vss 0.00413f
C11441 vdd.n2740 vss 0.0471f
C11442 vdd.n2741 vss 0.00324f
C11443 vdd.n2743 vss 0.00925f
C11444 vdd.t392 vss 0.0471f
C11445 vdd.n2744 vss 0.00425f
C11446 vdd.n2745 vss 0.0424f
C11447 vdd.n2746 vss 0.0132f
C11448 vdd.n2747 vss 0.00324f
C11449 vdd.n2748 vss 0.0128f
C11450 vdd.n2749 vss 0.02f
C11451 vdd.n2750 vss 0.00425f
C11452 vdd.n2751 vss 0.00413f
C11453 vdd.n2752 vss 0.00251f
C11454 vdd.t1141 vss 0.0471f
C11455 vdd.n2753 vss 0.00251f
C11456 vdd.n2754 vss 0.00517f
C11457 vdd.n2755 vss 0.00679f
C11458 vdd.n2756 vss 0.00517f
C11459 vdd.n2757 vss 0.00679f
C11460 vdd.n2758 vss 0.02f
C11461 vdd.n2759 vss 0.00425f
C11462 vdd.n2760 vss 0.0424f
C11463 vdd.n2761 vss 0.0132f
C11464 vdd.n2762 vss 0.00925f
C11465 vdd.n2763 vss 0.00425f
C11466 vdd.n2764 vss 0.00413f
C11467 vdd.n2765 vss 0.00324f
C11468 vdd.n2766 vss 0.0471f
C11469 vdd.t1139 vss 0.0471f
C11470 vdd.n2767 vss 0.00251f
C11471 vdd.n2768 vss 0.0112f
C11472 vdd.n2769 vss 0.0128f
C11473 vdd.t1140 vss 0.00134f
C11474 vdd.t495 vss 0.0013f
C11475 vdd.n2770 vss 0.0332f
C11476 vdd.n2771 vss 0.0393f
C11477 vdd.n2772 vss 0.0418f
C11478 vdd.n2773 vss 0.0912f
C11479 vdd.n2774 vss 0.0824f
C11480 vdd.n2775 vss 0.059f
C11481 vdd.t45 vss 0.0013f
C11482 vdd.t74 vss 0.00134f
C11483 vdd.n2776 vss 0.00324f
C11484 vdd.n2777 vss 0.0112f
C11485 vdd.n2778 vss 0.0128f
C11486 vdd.n2779 vss 0.00413f
C11487 vdd.n2780 vss 0.00413f
C11488 vdd.n2781 vss 0.0471f
C11489 vdd.n2782 vss 0.00251f
C11490 vdd.t1125 vss 0.0471f
C11491 vdd.n2783 vss 0.00324f
C11492 vdd.n2785 vss 0.00679f
C11493 vdd.n2786 vss 0.00413f
C11494 vdd.n2787 vss 0.00324f
C11495 vdd.n2788 vss 0.00413f
C11496 vdd.n2789 vss 0.0471f
C11497 vdd.n2790 vss 0.00324f
C11498 vdd.n2792 vss 0.00925f
C11499 vdd.t729 vss 0.0471f
C11500 vdd.n2793 vss 0.00425f
C11501 vdd.n2794 vss 0.0424f
C11502 vdd.n2795 vss 0.0132f
C11503 vdd.n2796 vss 0.00324f
C11504 vdd.n2797 vss 0.0128f
C11505 vdd.n2798 vss 0.02f
C11506 vdd.n2799 vss 0.00425f
C11507 vdd.n2800 vss 0.00413f
C11508 vdd.n2801 vss 0.00251f
C11509 vdd.t614 vss 0.0471f
C11510 vdd.n2802 vss 0.00251f
C11511 vdd.n2803 vss 0.00517f
C11512 vdd.n2804 vss 0.00679f
C11513 vdd.n2805 vss 0.00517f
C11514 vdd.n2806 vss 0.00679f
C11515 vdd.n2807 vss 0.02f
C11516 vdd.n2808 vss 0.00425f
C11517 vdd.n2809 vss 0.0424f
C11518 vdd.n2810 vss 0.0132f
C11519 vdd.n2811 vss 0.00925f
C11520 vdd.n2812 vss 0.00425f
C11521 vdd.n2813 vss 0.00413f
C11522 vdd.n2814 vss 0.00324f
C11523 vdd.n2815 vss 0.0471f
C11524 vdd.t612 vss 0.0471f
C11525 vdd.n2816 vss 0.00251f
C11526 vdd.n2817 vss 0.0112f
C11527 vdd.n2818 vss 0.0128f
C11528 vdd.t613 vss 0.00134f
C11529 vdd.t1126 vss 0.0013f
C11530 vdd.n2819 vss 0.0332f
C11531 vdd.n2820 vss 0.0393f
C11532 vdd.n2821 vss 0.158f
C11533 vdd.n2822 vss 0.00324f
C11534 vdd.n2823 vss 0.0112f
C11535 vdd.n2824 vss 0.0128f
C11536 vdd.n2825 vss 0.00413f
C11537 vdd.n2826 vss 0.00413f
C11538 vdd.n2827 vss 0.0471f
C11539 vdd.n2828 vss 0.00251f
C11540 vdd.t438 vss 0.0471f
C11541 vdd.n2829 vss 0.00324f
C11542 vdd.n2831 vss 0.00679f
C11543 vdd.n2832 vss 0.00413f
C11544 vdd.n2833 vss 0.00324f
C11545 vdd.n2834 vss 0.00413f
C11546 vdd.n2835 vss 0.0471f
C11547 vdd.n2836 vss 0.00324f
C11548 vdd.n2838 vss 0.00925f
C11549 vdd.t1106 vss 0.0471f
C11550 vdd.n2839 vss 0.00425f
C11551 vdd.n2840 vss 0.0424f
C11552 vdd.n2841 vss 0.0132f
C11553 vdd.n2842 vss 0.00324f
C11554 vdd.n2843 vss 0.0128f
C11555 vdd.n2844 vss 0.02f
C11556 vdd.n2845 vss 0.00425f
C11557 vdd.n2846 vss 0.00413f
C11558 vdd.n2847 vss 0.00251f
C11559 vdd.t133 vss 0.0471f
C11560 vdd.n2848 vss 0.00251f
C11561 vdd.n2849 vss 0.00517f
C11562 vdd.n2850 vss 0.00679f
C11563 vdd.n2851 vss 0.00517f
C11564 vdd.n2852 vss 0.00679f
C11565 vdd.n2853 vss 0.02f
C11566 vdd.n2854 vss 0.00425f
C11567 vdd.n2855 vss 0.0424f
C11568 vdd.n2856 vss 0.0132f
C11569 vdd.n2857 vss 0.00925f
C11570 vdd.n2858 vss 0.00425f
C11571 vdd.n2859 vss 0.00413f
C11572 vdd.n2860 vss 0.00324f
C11573 vdd.n2861 vss 0.0471f
C11574 vdd.t134 vss 0.0471f
C11575 vdd.n2862 vss 0.00251f
C11576 vdd.n2863 vss 0.0112f
C11577 vdd.n2864 vss 0.0128f
C11578 vdd.t135 vss 0.00134f
C11579 vdd.t439 vss 0.0013f
C11580 vdd.n2865 vss 0.0332f
C11581 vdd.n2866 vss 0.0393f
C11582 vdd.n2867 vss 0.0316f
C11583 vdd.n2868 vss 0.256f
C11584 vdd.n2869 vss 0.00324f
C11585 vdd.n2870 vss 0.0112f
C11586 vdd.n2871 vss 0.0128f
C11587 vdd.n2872 vss 0.00413f
C11588 vdd.n2873 vss 0.00413f
C11589 vdd.n2874 vss 0.0471f
C11590 vdd.n2875 vss 0.00251f
C11591 vdd.t44 vss 0.0471f
C11592 vdd.n2876 vss 0.00324f
C11593 vdd.n2878 vss 0.00679f
C11594 vdd.n2879 vss 0.00413f
C11595 vdd.n2880 vss 0.00324f
C11596 vdd.n2881 vss 0.00413f
C11597 vdd.n2882 vss 0.0471f
C11598 vdd.n2883 vss 0.00324f
C11599 vdd.n2885 vss 0.00925f
C11600 vdd.t445 vss 0.0471f
C11601 vdd.n2886 vss 0.00425f
C11602 vdd.n2887 vss 0.0424f
C11603 vdd.n2888 vss 0.0132f
C11604 vdd.n2889 vss 0.00324f
C11605 vdd.n2890 vss 0.0128f
C11606 vdd.n2891 vss 0.02f
C11607 vdd.n2892 vss 0.00425f
C11608 vdd.n2893 vss 0.00413f
C11609 vdd.n2894 vss 0.00251f
C11610 vdd.t75 vss 0.0471f
C11611 vdd.n2895 vss 0.00251f
C11612 vdd.n2896 vss 0.00517f
C11613 vdd.n2897 vss 0.00679f
C11614 vdd.n2898 vss 0.00517f
C11615 vdd.n2899 vss 0.00679f
C11616 vdd.n2900 vss 0.02f
C11617 vdd.n2901 vss 0.00425f
C11618 vdd.n2902 vss 0.0424f
C11619 vdd.n2903 vss 0.0132f
C11620 vdd.n2904 vss 0.00925f
C11621 vdd.n2905 vss 0.00425f
C11622 vdd.n2906 vss 0.00413f
C11623 vdd.n2907 vss 0.00324f
C11624 vdd.n2908 vss 0.0471f
C11625 vdd.t73 vss 0.0471f
C11626 vdd.n2909 vss 0.00251f
C11627 vdd.n2910 vss 0.0112f
C11628 vdd.n2911 vss 0.0128f
C11629 vdd.n2912 vss 0.0953f
C11630 vdd.n2913 vss 0.0393f
C11631 vdd.n2914 vss 0.0332f
C11632 vdd.n2915 vss 0.0596f
C11633 vdd.n2916 vss 0.00324f
C11634 vdd.n2917 vss 0.0112f
C11635 vdd.n2918 vss 0.0128f
C11636 vdd.n2919 vss 0.00413f
C11637 vdd.n2920 vss 0.00413f
C11638 vdd.n2921 vss 0.0471f
C11639 vdd.n2922 vss 0.00251f
C11640 vdd.t11 vss 0.0471f
C11641 vdd.n2923 vss 0.00324f
C11642 vdd.n2925 vss 0.00679f
C11643 vdd.n2926 vss 0.00413f
C11644 vdd.n2927 vss 0.00324f
C11645 vdd.n2928 vss 0.00413f
C11646 vdd.n2929 vss 0.0471f
C11647 vdd.n2930 vss 0.00324f
C11648 vdd.n2932 vss 0.00925f
C11649 vdd.t605 vss 0.0471f
C11650 vdd.n2933 vss 0.00425f
C11651 vdd.n2934 vss 0.0424f
C11652 vdd.n2935 vss 0.0132f
C11653 vdd.n2936 vss 0.00324f
C11654 vdd.n2937 vss 0.0128f
C11655 vdd.n2938 vss 0.02f
C11656 vdd.n2939 vss 0.00425f
C11657 vdd.n2940 vss 0.00413f
C11658 vdd.n2941 vss 0.00251f
C11659 vdd.t222 vss 0.0471f
C11660 vdd.n2942 vss 0.00251f
C11661 vdd.n2943 vss 0.00517f
C11662 vdd.n2944 vss 0.00679f
C11663 vdd.n2945 vss 0.00517f
C11664 vdd.n2946 vss 0.00679f
C11665 vdd.n2947 vss 0.02f
C11666 vdd.n2948 vss 0.00425f
C11667 vdd.n2949 vss 0.0424f
C11668 vdd.n2950 vss 0.0132f
C11669 vdd.n2951 vss 0.00925f
C11670 vdd.n2952 vss 0.00425f
C11671 vdd.n2953 vss 0.00413f
C11672 vdd.n2954 vss 0.00324f
C11673 vdd.n2955 vss 0.0471f
C11674 vdd.t220 vss 0.0471f
C11675 vdd.n2956 vss 0.00251f
C11676 vdd.n2957 vss 0.0112f
C11677 vdd.n2958 vss 0.0128f
C11678 vdd.t221 vss 0.00134f
C11679 vdd.t12 vss 0.0013f
C11680 vdd.n2959 vss 0.0332f
C11681 vdd.n2960 vss 0.0393f
C11682 vdd.n2961 vss 0.0418f
C11683 vdd.n2962 vss 0.118f
C11684 vdd.n2963 vss 0.121f
C11685 vdd.t39 vss 0.0013f
C11686 vdd.t1385 vss 0.00134f
C11687 vdd.n2964 vss 0.00324f
C11688 vdd.n2965 vss 0.0112f
C11689 vdd.n2966 vss 0.0128f
C11690 vdd.n2967 vss 0.00413f
C11691 vdd.n2968 vss 0.00413f
C11692 vdd.n2969 vss 0.0471f
C11693 vdd.n2970 vss 0.00251f
C11694 vdd.t38 vss 0.0471f
C11695 vdd.n2971 vss 0.00324f
C11696 vdd.n2973 vss 0.00679f
C11697 vdd.n2974 vss 0.00413f
C11698 vdd.n2975 vss 0.00324f
C11699 vdd.n2976 vss 0.00413f
C11700 vdd.n2977 vss 0.0471f
C11701 vdd.n2978 vss 0.00324f
C11702 vdd.n2980 vss 0.00925f
C11703 vdd.t1221 vss 0.0471f
C11704 vdd.n2981 vss 0.00425f
C11705 vdd.n2982 vss 0.0424f
C11706 vdd.n2983 vss 0.0132f
C11707 vdd.n2984 vss 0.00324f
C11708 vdd.n2985 vss 0.0128f
C11709 vdd.n2986 vss 0.02f
C11710 vdd.n2987 vss 0.00425f
C11711 vdd.n2988 vss 0.00413f
C11712 vdd.n2989 vss 0.00251f
C11713 vdd.t1386 vss 0.0471f
C11714 vdd.n2990 vss 0.00251f
C11715 vdd.n2991 vss 0.00517f
C11716 vdd.n2992 vss 0.00679f
C11717 vdd.n2993 vss 0.00517f
C11718 vdd.n2994 vss 0.00679f
C11719 vdd.n2995 vss 0.02f
C11720 vdd.n2996 vss 0.00425f
C11721 vdd.n2997 vss 0.0424f
C11722 vdd.n2998 vss 0.0132f
C11723 vdd.n2999 vss 0.00925f
C11724 vdd.n3000 vss 0.00425f
C11725 vdd.n3001 vss 0.00413f
C11726 vdd.n3002 vss 0.00324f
C11727 vdd.n3003 vss 0.0471f
C11728 vdd.t1384 vss 0.0471f
C11729 vdd.n3004 vss 0.00251f
C11730 vdd.n3005 vss 0.0112f
C11731 vdd.n3006 vss 0.0707f
C11732 vdd.n3007 vss 0.0393f
C11733 vdd.n3008 vss 0.0332f
C11734 vdd.n3009 vss 0.0596f
C11735 vdd.n3010 vss 0.00324f
C11736 vdd.n3011 vss 0.0112f
C11737 vdd.n3012 vss 0.0128f
C11738 vdd.n3013 vss 0.00413f
C11739 vdd.n3014 vss 0.00413f
C11740 vdd.n3015 vss 0.0471f
C11741 vdd.n3016 vss 0.00251f
C11742 vdd.t1296 vss 0.0471f
C11743 vdd.n3017 vss 0.00324f
C11744 vdd.n3019 vss 0.00679f
C11745 vdd.n3020 vss 0.00413f
C11746 vdd.n3021 vss 0.00324f
C11747 vdd.n3022 vss 0.00413f
C11748 vdd.n3023 vss 0.0471f
C11749 vdd.n3024 vss 0.00324f
C11750 vdd.n3026 vss 0.00925f
C11751 vdd.t1434 vss 0.0471f
C11752 vdd.n3027 vss 0.00425f
C11753 vdd.n3028 vss 0.0424f
C11754 vdd.n3029 vss 0.0132f
C11755 vdd.n3030 vss 0.00324f
C11756 vdd.n3031 vss 0.0128f
C11757 vdd.n3032 vss 0.02f
C11758 vdd.n3033 vss 0.00425f
C11759 vdd.n3034 vss 0.00413f
C11760 vdd.n3035 vss 0.00251f
C11761 vdd.t454 vss 0.0471f
C11762 vdd.n3036 vss 0.00251f
C11763 vdd.n3037 vss 0.00517f
C11764 vdd.n3038 vss 0.00679f
C11765 vdd.n3039 vss 0.00517f
C11766 vdd.n3040 vss 0.00679f
C11767 vdd.n3041 vss 0.02f
C11768 vdd.n3042 vss 0.00425f
C11769 vdd.n3043 vss 0.0424f
C11770 vdd.n3044 vss 0.0132f
C11771 vdd.n3045 vss 0.00925f
C11772 vdd.n3046 vss 0.00425f
C11773 vdd.n3047 vss 0.00413f
C11774 vdd.n3048 vss 0.00324f
C11775 vdd.n3049 vss 0.0471f
C11776 vdd.t452 vss 0.0471f
C11777 vdd.n3050 vss 0.00251f
C11778 vdd.n3051 vss 0.0112f
C11779 vdd.n3052 vss 0.0128f
C11780 vdd.t453 vss 0.00134f
C11781 vdd.t1297 vss 0.0013f
C11782 vdd.n3053 vss 0.0332f
C11783 vdd.n3054 vss 0.0393f
C11784 vdd.n3055 vss 0.0418f
C11785 vdd.n3056 vss 0.118f
C11786 vdd.n3057 vss 0.0951f
C11787 vdd.t853 vss 0.0013f
C11788 vdd.t800 vss 0.00134f
C11789 vdd.n3058 vss 0.00324f
C11790 vdd.n3059 vss 0.0112f
C11791 vdd.n3060 vss 0.0128f
C11792 vdd.n3061 vss 0.00413f
C11793 vdd.n3062 vss 0.00413f
C11794 vdd.n3063 vss 0.0471f
C11795 vdd.n3064 vss 0.00251f
C11796 vdd.t790 vss 0.0471f
C11797 vdd.n3065 vss 0.00324f
C11798 vdd.n3067 vss 0.00679f
C11799 vdd.n3068 vss 0.00413f
C11800 vdd.n3069 vss 0.00324f
C11801 vdd.n3070 vss 0.00413f
C11802 vdd.n3071 vss 0.0471f
C11803 vdd.n3072 vss 0.00324f
C11804 vdd.n3074 vss 0.00925f
C11805 vdd.t21 vss 0.0471f
C11806 vdd.n3075 vss 0.00425f
C11807 vdd.n3076 vss 0.0424f
C11808 vdd.n3077 vss 0.0132f
C11809 vdd.n3078 vss 0.00324f
C11810 vdd.n3079 vss 0.0128f
C11811 vdd.n3080 vss 0.02f
C11812 vdd.n3081 vss 0.00425f
C11813 vdd.n3082 vss 0.00413f
C11814 vdd.n3083 vss 0.00251f
C11815 vdd.t276 vss 0.0471f
C11816 vdd.n3084 vss 0.00251f
C11817 vdd.n3085 vss 0.00517f
C11818 vdd.n3086 vss 0.00679f
C11819 vdd.n3087 vss 0.00517f
C11820 vdd.n3088 vss 0.00679f
C11821 vdd.n3089 vss 0.02f
C11822 vdd.n3090 vss 0.00425f
C11823 vdd.n3091 vss 0.0424f
C11824 vdd.n3092 vss 0.0132f
C11825 vdd.n3093 vss 0.00925f
C11826 vdd.n3094 vss 0.00425f
C11827 vdd.n3095 vss 0.00413f
C11828 vdd.n3096 vss 0.00324f
C11829 vdd.n3097 vss 0.0471f
C11830 vdd.t274 vss 0.0471f
C11831 vdd.n3098 vss 0.00251f
C11832 vdd.n3099 vss 0.0112f
C11833 vdd.n3100 vss 0.0128f
C11834 vdd.t275 vss 0.00134f
C11835 vdd.t791 vss 0.0013f
C11836 vdd.n3101 vss 0.0332f
C11837 vdd.n3102 vss 0.0393f
C11838 vdd.n3103 vss 0.119f
C11839 vdd.n3104 vss 0.00324f
C11840 vdd.n3105 vss 0.0112f
C11841 vdd.n3106 vss 0.0128f
C11842 vdd.n3107 vss 0.00413f
C11843 vdd.n3108 vss 0.00413f
C11844 vdd.n3109 vss 0.0471f
C11845 vdd.n3110 vss 0.00251f
C11846 vdd.t852 vss 0.0471f
C11847 vdd.n3111 vss 0.00324f
C11848 vdd.n3113 vss 0.00679f
C11849 vdd.n3114 vss 0.00413f
C11850 vdd.n3115 vss 0.00324f
C11851 vdd.n3116 vss 0.00413f
C11852 vdd.n3117 vss 0.0471f
C11853 vdd.n3118 vss 0.00324f
C11854 vdd.n3120 vss 0.00925f
C11855 vdd.t1156 vss 0.0471f
C11856 vdd.n3121 vss 0.00425f
C11857 vdd.n3122 vss 0.0424f
C11858 vdd.n3123 vss 0.0132f
C11859 vdd.n3124 vss 0.00324f
C11860 vdd.n3125 vss 0.0128f
C11861 vdd.n3126 vss 0.02f
C11862 vdd.n3127 vss 0.00425f
C11863 vdd.n3128 vss 0.00413f
C11864 vdd.n3129 vss 0.00251f
C11865 vdd.t801 vss 0.0471f
C11866 vdd.n3130 vss 0.00251f
C11867 vdd.n3131 vss 0.00517f
C11868 vdd.n3132 vss 0.00679f
C11869 vdd.n3133 vss 0.00517f
C11870 vdd.n3134 vss 0.00679f
C11871 vdd.n3135 vss 0.02f
C11872 vdd.n3136 vss 0.00425f
C11873 vdd.n3137 vss 0.0424f
C11874 vdd.n3138 vss 0.0132f
C11875 vdd.n3139 vss 0.00925f
C11876 vdd.n3140 vss 0.00425f
C11877 vdd.n3141 vss 0.00413f
C11878 vdd.n3142 vss 0.00324f
C11879 vdd.n3143 vss 0.0471f
C11880 vdd.t799 vss 0.0471f
C11881 vdd.n3144 vss 0.00251f
C11882 vdd.n3145 vss 0.0112f
C11883 vdd.n3146 vss 0.0128f
C11884 vdd.n3147 vss 0.118f
C11885 vdd.n3148 vss 0.0393f
C11886 vdd.n3149 vss 0.0332f
C11887 vdd.n3150 vss 0.0596f
C11888 vdd.n3151 vss 0.00324f
C11889 vdd.n3152 vss 0.0112f
C11890 vdd.n3153 vss 0.0128f
C11891 vdd.n3154 vss 0.00413f
C11892 vdd.n3155 vss 0.00413f
C11893 vdd.n3156 vss 0.0471f
C11894 vdd.n3157 vss 0.00251f
C11895 vdd.t373 vss 0.0471f
C11896 vdd.n3158 vss 0.00324f
C11897 vdd.n3160 vss 0.00679f
C11898 vdd.n3161 vss 0.00413f
C11899 vdd.n3162 vss 0.00324f
C11900 vdd.n3163 vss 0.00413f
C11901 vdd.n3164 vss 0.0471f
C11902 vdd.n3165 vss 0.00324f
C11903 vdd.n3167 vss 0.00925f
C11904 vdd.t245 vss 0.0471f
C11905 vdd.n3168 vss 0.00425f
C11906 vdd.n3169 vss 0.0424f
C11907 vdd.n3170 vss 0.0132f
C11908 vdd.n3171 vss 0.00324f
C11909 vdd.n3172 vss 0.0128f
C11910 vdd.n3173 vss 0.02f
C11911 vdd.n3174 vss 0.00425f
C11912 vdd.n3175 vss 0.00413f
C11913 vdd.n3176 vss 0.00251f
C11914 vdd.t280 vss 0.0471f
C11915 vdd.n3177 vss 0.00251f
C11916 vdd.n3178 vss 0.00517f
C11917 vdd.n3179 vss 0.00679f
C11918 vdd.n3180 vss 0.00517f
C11919 vdd.n3181 vss 0.00679f
C11920 vdd.n3182 vss 0.02f
C11921 vdd.n3183 vss 0.00425f
C11922 vdd.n3184 vss 0.0424f
C11923 vdd.n3185 vss 0.0132f
C11924 vdd.n3186 vss 0.00925f
C11925 vdd.n3187 vss 0.00425f
C11926 vdd.n3188 vss 0.00413f
C11927 vdd.n3189 vss 0.00324f
C11928 vdd.n3190 vss 0.0471f
C11929 vdd.t278 vss 0.0471f
C11930 vdd.n3191 vss 0.00251f
C11931 vdd.n3192 vss 0.0112f
C11932 vdd.n3193 vss 0.0128f
C11933 vdd.t279 vss 0.00134f
C11934 vdd.t374 vss 0.0013f
C11935 vdd.n3194 vss 0.0332f
C11936 vdd.n3195 vss 0.0393f
C11937 vdd.n3196 vss 0.0418f
C11938 vdd.n3197 vss 0.118f
C11939 vdd.n3198 vss 0.121f
C11940 vdd.t968 vss 0.0013f
C11941 vdd.t1211 vss 0.00134f
C11942 vdd.n3199 vss 0.00324f
C11943 vdd.n3200 vss 0.0112f
C11944 vdd.n3201 vss 0.0128f
C11945 vdd.n3202 vss 0.00413f
C11946 vdd.n3203 vss 0.00413f
C11947 vdd.n3204 vss 0.0471f
C11948 vdd.n3205 vss 0.00251f
C11949 vdd.t967 vss 0.0471f
C11950 vdd.n3206 vss 0.00324f
C11951 vdd.n3208 vss 0.00679f
C11952 vdd.n3209 vss 0.00413f
C11953 vdd.n3210 vss 0.00324f
C11954 vdd.n3211 vss 0.00413f
C11955 vdd.n3212 vss 0.0471f
C11956 vdd.n3213 vss 0.00324f
C11957 vdd.n3215 vss 0.00925f
C11958 vdd.t1282 vss 0.0471f
C11959 vdd.n3216 vss 0.00425f
C11960 vdd.n3217 vss 0.0424f
C11961 vdd.n3218 vss 0.0132f
C11962 vdd.n3219 vss 0.00324f
C11963 vdd.n3220 vss 0.0128f
C11964 vdd.n3221 vss 0.02f
C11965 vdd.n3222 vss 0.00425f
C11966 vdd.n3223 vss 0.00413f
C11967 vdd.n3224 vss 0.00251f
C11968 vdd.t1212 vss 0.0471f
C11969 vdd.n3225 vss 0.00251f
C11970 vdd.n3226 vss 0.00517f
C11971 vdd.n3227 vss 0.00679f
C11972 vdd.n3228 vss 0.00517f
C11973 vdd.n3229 vss 0.00679f
C11974 vdd.n3230 vss 0.02f
C11975 vdd.n3231 vss 0.00425f
C11976 vdd.n3232 vss 0.0424f
C11977 vdd.n3233 vss 0.0132f
C11978 vdd.n3234 vss 0.00925f
C11979 vdd.n3235 vss 0.00425f
C11980 vdd.n3236 vss 0.00413f
C11981 vdd.n3237 vss 0.00324f
C11982 vdd.n3238 vss 0.0471f
C11983 vdd.t1210 vss 0.0471f
C11984 vdd.n3239 vss 0.00251f
C11985 vdd.n3240 vss 0.0112f
C11986 vdd.n3241 vss 0.0707f
C11987 vdd.n3242 vss 0.0393f
C11988 vdd.n3243 vss 0.0332f
C11989 vdd.n3244 vss 0.0596f
C11990 vdd.n3245 vss 0.00324f
C11991 vdd.n3246 vss 0.0112f
C11992 vdd.n3247 vss 0.0128f
C11993 vdd.n3248 vss 0.00413f
C11994 vdd.n3249 vss 0.00413f
C11995 vdd.n3250 vss 0.0471f
C11996 vdd.n3251 vss 0.00251f
C11997 vdd.t1328 vss 0.0471f
C11998 vdd.n3252 vss 0.00324f
C11999 vdd.n3254 vss 0.00679f
C12000 vdd.n3255 vss 0.00413f
C12001 vdd.n3256 vss 0.00324f
C12002 vdd.n3257 vss 0.00413f
C12003 vdd.n3258 vss 0.0471f
C12004 vdd.n3259 vss 0.00324f
C12005 vdd.n3261 vss 0.00925f
C12006 vdd.t798 vss 0.0471f
C12007 vdd.n3262 vss 0.00425f
C12008 vdd.n3263 vss 0.0424f
C12009 vdd.n3264 vss 0.0132f
C12010 vdd.n3265 vss 0.00324f
C12011 vdd.n3266 vss 0.0128f
C12012 vdd.n3267 vss 0.02f
C12013 vdd.n3268 vss 0.00425f
C12014 vdd.n3269 vss 0.00413f
C12015 vdd.n3270 vss 0.00251f
C12016 vdd.t1277 vss 0.0471f
C12017 vdd.n3271 vss 0.00251f
C12018 vdd.n3272 vss 0.00517f
C12019 vdd.n3273 vss 0.00679f
C12020 vdd.n3274 vss 0.00517f
C12021 vdd.n3275 vss 0.00679f
C12022 vdd.n3276 vss 0.02f
C12023 vdd.n3277 vss 0.00425f
C12024 vdd.n3278 vss 0.0424f
C12025 vdd.n3279 vss 0.0132f
C12026 vdd.n3280 vss 0.00925f
C12027 vdd.n3281 vss 0.00425f
C12028 vdd.n3282 vss 0.00413f
C12029 vdd.n3283 vss 0.00324f
C12030 vdd.n3284 vss 0.0471f
C12031 vdd.t1275 vss 0.0471f
C12032 vdd.n3285 vss 0.00251f
C12033 vdd.n3286 vss 0.0112f
C12034 vdd.n3287 vss 0.0128f
C12035 vdd.t1276 vss 0.00134f
C12036 vdd.t1329 vss 0.0013f
C12037 vdd.n3288 vss 0.0332f
C12038 vdd.n3289 vss 0.0393f
C12039 vdd.n3290 vss 0.0418f
C12040 vdd.n3291 vss 0.0912f
C12041 vdd.n3292 vss 0.0824f
C12042 vdd.n3293 vss 0.059f
C12043 vdd.t820 vss 0.0013f
C12044 vdd.t267 vss 0.00134f
C12045 vdd.n3294 vss 0.00324f
C12046 vdd.n3295 vss 0.0112f
C12047 vdd.n3296 vss 0.0128f
C12048 vdd.n3297 vss 0.00413f
C12049 vdd.n3298 vss 0.00413f
C12050 vdd.n3299 vss 0.0471f
C12051 vdd.n3300 vss 0.00251f
C12052 vdd.t436 vss 0.0471f
C12053 vdd.n3301 vss 0.00324f
C12054 vdd.n3303 vss 0.00679f
C12055 vdd.n3304 vss 0.00413f
C12056 vdd.n3305 vss 0.00324f
C12057 vdd.n3306 vss 0.00413f
C12058 vdd.n3307 vss 0.0471f
C12059 vdd.n3308 vss 0.00324f
C12060 vdd.n3310 vss 0.00925f
C12061 vdd.t310 vss 0.0471f
C12062 vdd.n3311 vss 0.00425f
C12063 vdd.n3312 vss 0.0424f
C12064 vdd.n3313 vss 0.0132f
C12065 vdd.n3314 vss 0.00324f
C12066 vdd.n3315 vss 0.0128f
C12067 vdd.n3316 vss 0.02f
C12068 vdd.n3317 vss 0.00425f
C12069 vdd.n3318 vss 0.00413f
C12070 vdd.n3319 vss 0.00251f
C12071 vdd.t1508 vss 0.0471f
C12072 vdd.n3320 vss 0.00251f
C12073 vdd.n3321 vss 0.00517f
C12074 vdd.n3322 vss 0.00679f
C12075 vdd.n3323 vss 0.00517f
C12076 vdd.n3324 vss 0.00679f
C12077 vdd.n3325 vss 0.02f
C12078 vdd.n3326 vss 0.00425f
C12079 vdd.n3327 vss 0.0424f
C12080 vdd.n3328 vss 0.0132f
C12081 vdd.n3329 vss 0.00925f
C12082 vdd.n3330 vss 0.00425f
C12083 vdd.n3331 vss 0.00413f
C12084 vdd.n3332 vss 0.00324f
C12085 vdd.n3333 vss 0.0471f
C12086 vdd.t1509 vss 0.0471f
C12087 vdd.n3334 vss 0.00251f
C12088 vdd.n3335 vss 0.0112f
C12089 vdd.n3336 vss 0.0128f
C12090 vdd.t1510 vss 0.00134f
C12091 vdd.t437 vss 0.0013f
C12092 vdd.n3337 vss 0.0332f
C12093 vdd.n3338 vss 0.0393f
C12094 vdd.n3339 vss 0.119f
C12095 vdd.n3340 vss 0.00324f
C12096 vdd.n3341 vss 0.0112f
C12097 vdd.n3342 vss 0.0128f
C12098 vdd.n3343 vss 0.00413f
C12099 vdd.n3344 vss 0.00413f
C12100 vdd.n3345 vss 0.0471f
C12101 vdd.n3346 vss 0.00251f
C12102 vdd.t819 vss 0.0471f
C12103 vdd.n3347 vss 0.00324f
C12104 vdd.n3349 vss 0.00679f
C12105 vdd.n3350 vss 0.00413f
C12106 vdd.n3351 vss 0.00324f
C12107 vdd.n3352 vss 0.00413f
C12108 vdd.n3353 vss 0.0471f
C12109 vdd.n3354 vss 0.00324f
C12110 vdd.n3356 vss 0.00925f
C12111 vdd.t1203 vss 0.0471f
C12112 vdd.n3357 vss 0.00425f
C12113 vdd.n3358 vss 0.0424f
C12114 vdd.n3359 vss 0.0132f
C12115 vdd.n3360 vss 0.00324f
C12116 vdd.n3361 vss 0.0128f
C12117 vdd.n3362 vss 0.02f
C12118 vdd.n3363 vss 0.00425f
C12119 vdd.n3364 vss 0.00413f
C12120 vdd.n3365 vss 0.00251f
C12121 vdd.t265 vss 0.0471f
C12122 vdd.n3366 vss 0.00251f
C12123 vdd.n3367 vss 0.00517f
C12124 vdd.n3368 vss 0.00679f
C12125 vdd.n3369 vss 0.00517f
C12126 vdd.n3370 vss 0.00679f
C12127 vdd.n3371 vss 0.02f
C12128 vdd.n3372 vss 0.00425f
C12129 vdd.n3373 vss 0.0424f
C12130 vdd.n3374 vss 0.0132f
C12131 vdd.n3375 vss 0.00925f
C12132 vdd.n3376 vss 0.00425f
C12133 vdd.n3377 vss 0.00413f
C12134 vdd.n3378 vss 0.00324f
C12135 vdd.n3379 vss 0.0471f
C12136 vdd.t266 vss 0.0471f
C12137 vdd.n3380 vss 0.00251f
C12138 vdd.n3381 vss 0.0112f
C12139 vdd.n3382 vss 0.0128f
C12140 vdd.n3383 vss 0.118f
C12141 vdd.n3384 vss 0.0393f
C12142 vdd.n3385 vss 0.0332f
C12143 vdd.n3386 vss 0.0596f
C12144 vdd.n3387 vss 0.00324f
C12145 vdd.n3388 vss 0.0112f
C12146 vdd.n3389 vss 0.0128f
C12147 vdd.n3390 vss 0.00413f
C12148 vdd.n3391 vss 0.00413f
C12149 vdd.n3392 vss 0.0471f
C12150 vdd.n3393 vss 0.00251f
C12151 vdd.t1332 vss 0.0471f
C12152 vdd.n3394 vss 0.00324f
C12153 vdd.n3396 vss 0.00679f
C12154 vdd.n3397 vss 0.00413f
C12155 vdd.n3398 vss 0.00324f
C12156 vdd.n3399 vss 0.00413f
C12157 vdd.n3400 vss 0.0471f
C12158 vdd.n3401 vss 0.00324f
C12159 vdd.n3403 vss 0.00925f
C12160 vdd.t1124 vss 0.0471f
C12161 vdd.n3404 vss 0.00425f
C12162 vdd.n3405 vss 0.0424f
C12163 vdd.n3406 vss 0.0132f
C12164 vdd.n3407 vss 0.00324f
C12165 vdd.n3408 vss 0.0128f
C12166 vdd.n3409 vss 0.02f
C12167 vdd.n3410 vss 0.00425f
C12168 vdd.n3411 vss 0.00413f
C12169 vdd.n3412 vss 0.00251f
C12170 vdd.t1137 vss 0.0471f
C12171 vdd.n3413 vss 0.00251f
C12172 vdd.n3414 vss 0.00517f
C12173 vdd.n3415 vss 0.00679f
C12174 vdd.n3416 vss 0.00517f
C12175 vdd.n3417 vss 0.00679f
C12176 vdd.n3418 vss 0.02f
C12177 vdd.n3419 vss 0.00425f
C12178 vdd.n3420 vss 0.0424f
C12179 vdd.n3421 vss 0.0132f
C12180 vdd.n3422 vss 0.00925f
C12181 vdd.n3423 vss 0.00425f
C12182 vdd.n3424 vss 0.00413f
C12183 vdd.n3425 vss 0.00324f
C12184 vdd.n3426 vss 0.0471f
C12185 vdd.t1135 vss 0.0471f
C12186 vdd.n3427 vss 0.00251f
C12187 vdd.n3428 vss 0.0112f
C12188 vdd.n3429 vss 0.0128f
C12189 vdd.t1136 vss 0.00134f
C12190 vdd.t1333 vss 0.0013f
C12191 vdd.n3430 vss 0.0332f
C12192 vdd.n3431 vss 0.0393f
C12193 vdd.n3432 vss 0.0418f
C12194 vdd.n3433 vss 0.118f
C12195 vdd.n3434 vss 0.121f
C12196 vdd.t905 vss 0.0013f
C12197 vdd.t650 vss 0.00134f
C12198 vdd.n3435 vss 0.00324f
C12199 vdd.n3436 vss 0.0112f
C12200 vdd.n3437 vss 0.0128f
C12201 vdd.n3438 vss 0.00413f
C12202 vdd.n3439 vss 0.00413f
C12203 vdd.n3440 vss 0.0471f
C12204 vdd.n3441 vss 0.00251f
C12205 vdd.t904 vss 0.0471f
C12206 vdd.n3442 vss 0.00324f
C12207 vdd.n3444 vss 0.00679f
C12208 vdd.n3445 vss 0.00413f
C12209 vdd.n3446 vss 0.00324f
C12210 vdd.n3447 vss 0.00413f
C12211 vdd.n3448 vss 0.0471f
C12212 vdd.n3449 vss 0.00324f
C12213 vdd.n3451 vss 0.00925f
C12214 vdd.t1061 vss 0.0471f
C12215 vdd.n3452 vss 0.00425f
C12216 vdd.n3453 vss 0.0424f
C12217 vdd.n3454 vss 0.0132f
C12218 vdd.n3455 vss 0.00324f
C12219 vdd.n3456 vss 0.0128f
C12220 vdd.n3457 vss 0.02f
C12221 vdd.n3458 vss 0.00425f
C12222 vdd.n3459 vss 0.00413f
C12223 vdd.n3460 vss 0.00251f
C12224 vdd.t648 vss 0.0471f
C12225 vdd.n3461 vss 0.00251f
C12226 vdd.n3462 vss 0.00517f
C12227 vdd.n3463 vss 0.00679f
C12228 vdd.n3464 vss 0.00517f
C12229 vdd.n3465 vss 0.00679f
C12230 vdd.n3466 vss 0.02f
C12231 vdd.n3467 vss 0.00425f
C12232 vdd.n3468 vss 0.0424f
C12233 vdd.n3469 vss 0.0132f
C12234 vdd.n3470 vss 0.00925f
C12235 vdd.n3471 vss 0.00425f
C12236 vdd.n3472 vss 0.00413f
C12237 vdd.n3473 vss 0.00324f
C12238 vdd.n3474 vss 0.0471f
C12239 vdd.t649 vss 0.0471f
C12240 vdd.n3475 vss 0.00251f
C12241 vdd.n3476 vss 0.0112f
C12242 vdd.n3477 vss 0.0707f
C12243 vdd.n3478 vss 0.0393f
C12244 vdd.n3479 vss 0.0332f
C12245 vdd.n3480 vss 0.0596f
C12246 vdd.n3481 vss 0.00324f
C12247 vdd.n3482 vss 0.0112f
C12248 vdd.n3483 vss 0.0128f
C12249 vdd.n3484 vss 0.00413f
C12250 vdd.n3485 vss 0.00413f
C12251 vdd.n3486 vss 0.0471f
C12252 vdd.n3487 vss 0.00251f
C12253 vdd.t488 vss 0.0471f
C12254 vdd.n3488 vss 0.00324f
C12255 vdd.n3490 vss 0.00679f
C12256 vdd.n3491 vss 0.00413f
C12257 vdd.n3492 vss 0.00324f
C12258 vdd.n3493 vss 0.00413f
C12259 vdd.n3494 vss 0.0471f
C12260 vdd.n3495 vss 0.00324f
C12261 vdd.n3497 vss 0.00925f
C12262 vdd.t1123 vss 0.0471f
C12263 vdd.n3498 vss 0.00425f
C12264 vdd.n3499 vss 0.0424f
C12265 vdd.n3500 vss 0.0132f
C12266 vdd.n3501 vss 0.00324f
C12267 vdd.n3502 vss 0.0128f
C12268 vdd.n3503 vss 0.02f
C12269 vdd.n3504 vss 0.00425f
C12270 vdd.n3505 vss 0.00413f
C12271 vdd.n3506 vss 0.00251f
C12272 vdd.t830 vss 0.0471f
C12273 vdd.n3507 vss 0.00251f
C12274 vdd.n3508 vss 0.00517f
C12275 vdd.n3509 vss 0.00679f
C12276 vdd.n3510 vss 0.00517f
C12277 vdd.n3511 vss 0.00679f
C12278 vdd.n3512 vss 0.02f
C12279 vdd.n3513 vss 0.00425f
C12280 vdd.n3514 vss 0.0424f
C12281 vdd.n3515 vss 0.0132f
C12282 vdd.n3516 vss 0.00925f
C12283 vdd.n3517 vss 0.00425f
C12284 vdd.n3518 vss 0.00413f
C12285 vdd.n3519 vss 0.00324f
C12286 vdd.n3520 vss 0.0471f
C12287 vdd.t831 vss 0.0471f
C12288 vdd.n3521 vss 0.00251f
C12289 vdd.n3522 vss 0.0112f
C12290 vdd.n3523 vss 0.0128f
C12291 vdd.t832 vss 0.00134f
C12292 vdd.t489 vss 0.0013f
C12293 vdd.n3524 vss 0.0332f
C12294 vdd.n3525 vss 0.0393f
C12295 vdd.n3526 vss 0.0418f
C12296 vdd.n3527 vss 0.121f
C12297 vdd.n3528 vss 0.291f
C12298 vdd.n3529 vss 0.227f
C12299 vdd.n3530 vss 0.00324f
C12300 vdd.n3531 vss 0.0112f
C12301 vdd.n3532 vss 0.0128f
C12302 vdd.n3533 vss 0.00413f
C12303 vdd.n3534 vss 0.00413f
C12304 vdd.n3535 vss 0.0471f
C12305 vdd.n3536 vss 0.00251f
C12306 vdd.t986 vss 0.0471f
C12307 vdd.n3537 vss 0.00324f
C12308 vdd.n3539 vss 0.00679f
C12309 vdd.n3540 vss 0.00413f
C12310 vdd.n3541 vss 0.00324f
C12311 vdd.n3542 vss 0.00413f
C12312 vdd.n3543 vss 0.0471f
C12313 vdd.n3544 vss 0.00324f
C12314 vdd.n3546 vss 0.00925f
C12315 vdd.t1150 vss 0.0471f
C12316 vdd.n3547 vss 0.00425f
C12317 vdd.n3548 vss 0.0424f
C12318 vdd.n3549 vss 0.0132f
C12319 vdd.n3550 vss 0.00324f
C12320 vdd.n3551 vss 0.0128f
C12321 vdd.n3552 vss 0.02f
C12322 vdd.n3553 vss 0.00425f
C12323 vdd.n3554 vss 0.00413f
C12324 vdd.n3555 vss 0.00251f
C12325 vdd.t1172 vss 0.0471f
C12326 vdd.n3556 vss 0.00251f
C12327 vdd.n3557 vss 0.00517f
C12328 vdd.n3558 vss 0.00679f
C12329 vdd.n3559 vss 0.00517f
C12330 vdd.n3560 vss 0.00679f
C12331 vdd.n3561 vss 0.02f
C12332 vdd.n3562 vss 0.00425f
C12333 vdd.n3563 vss 0.0424f
C12334 vdd.n3564 vss 0.0132f
C12335 vdd.n3565 vss 0.00925f
C12336 vdd.n3566 vss 0.00425f
C12337 vdd.n3567 vss 0.00413f
C12338 vdd.n3568 vss 0.00324f
C12339 vdd.n3569 vss 0.0471f
C12340 vdd.t1173 vss 0.0471f
C12341 vdd.n3570 vss 0.00251f
C12342 vdd.n3571 vss 0.0112f
C12343 vdd.n3572 vss 0.0128f
C12344 vdd.n3573 vss 0.152f
C12345 vdd.n3574 vss 0.0393f
C12346 vdd.n3575 vss 0.0332f
C12347 vdd.n3576 vss 0.00324f
C12348 vdd.n3577 vss 0.0112f
C12349 vdd.n3578 vss 0.0128f
C12350 vdd.n3579 vss 0.00413f
C12351 vdd.n3580 vss 0.00413f
C12352 vdd.n3581 vss 0.0471f
C12353 vdd.n3582 vss 0.00251f
C12354 vdd.t24 vss 0.0471f
C12355 vdd.n3583 vss 0.00324f
C12356 vdd.n3585 vss 0.00679f
C12357 vdd.n3586 vss 0.00413f
C12358 vdd.n3587 vss 0.00324f
C12359 vdd.n3588 vss 0.00413f
C12360 vdd.n3589 vss 0.0471f
C12361 vdd.n3590 vss 0.00324f
C12362 vdd.n3592 vss 0.00925f
C12363 vdd.t1382 vss 0.0471f
C12364 vdd.n3593 vss 0.00425f
C12365 vdd.n3594 vss 0.0424f
C12366 vdd.n3595 vss 0.0132f
C12367 vdd.n3596 vss 0.00324f
C12368 vdd.n3597 vss 0.0128f
C12369 vdd.n3598 vss 0.02f
C12370 vdd.n3599 vss 0.00425f
C12371 vdd.n3600 vss 0.00413f
C12372 vdd.n3601 vss 0.00251f
C12373 vdd.t1428 vss 0.0471f
C12374 vdd.n3602 vss 0.00251f
C12375 vdd.n3603 vss 0.00517f
C12376 vdd.n3604 vss 0.00679f
C12377 vdd.n3605 vss 0.00517f
C12378 vdd.n3606 vss 0.00679f
C12379 vdd.n3607 vss 0.02f
C12380 vdd.n3608 vss 0.00425f
C12381 vdd.n3609 vss 0.0424f
C12382 vdd.n3610 vss 0.0132f
C12383 vdd.n3611 vss 0.00925f
C12384 vdd.n3612 vss 0.00425f
C12385 vdd.n3613 vss 0.00413f
C12386 vdd.n3614 vss 0.00324f
C12387 vdd.n3615 vss 0.0471f
C12388 vdd.t1429 vss 0.0471f
C12389 vdd.n3616 vss 0.00251f
C12390 vdd.n3617 vss 0.0112f
C12391 vdd.n3618 vss 0.0128f
C12392 vdd.n3619 vss 0.221f
C12393 vdd.n3620 vss 0.0393f
C12394 vdd.n3621 vss 0.0332f
C12395 vdd.t1035 vss 0.00134f
C12396 vdd.t561 vss 0.0013f
C12397 vdd.n3622 vss 0.0315f
C12398 vdd.n3623 vss 0.0393f
C12399 vdd.n3624 vss 0.00324f
C12400 vdd.n3625 vss 0.0112f
C12401 vdd.n3626 vss 0.0128f
C12402 vdd.n3627 vss 0.00413f
C12403 vdd.t1036 vss 0.0471f
C12404 vdd.n3628 vss 0.00324f
C12405 vdd.n3630 vss 0.00925f
C12406 vdd.n3631 vss 0.00413f
C12407 vdd.n3632 vss 0.00679f
C12408 vdd.n3633 vss 0.00413f
C12409 vdd.n3634 vss 0.0471f
C12410 vdd.n3635 vss 0.00324f
C12411 vdd.n3636 vss 0.0471f
C12412 vdd.n3637 vss 0.00324f
C12413 vdd.n3638 vss 0.0424f
C12414 vdd.t560 vss 0.0471f
C12415 vdd.n3640 vss 0.00425f
C12416 vdd.n3641 vss 0.00925f
C12417 vdd.n3642 vss 0.0132f
C12418 vdd.n3643 vss 0.00324f
C12419 vdd.n3644 vss 0.0128f
C12420 vdd.n3645 vss 0.02f
C12421 vdd.n3646 vss 0.00425f
C12422 vdd.n3647 vss 0.00413f
C12423 vdd.n3648 vss 0.00251f
C12424 vdd.t1034 vss 0.0471f
C12425 vdd.n3649 vss 0.00251f
C12426 vdd.n3650 vss 0.00517f
C12427 vdd.n3651 vss 0.00679f
C12428 vdd.n3652 vss 0.00324f
C12429 vdd.n3653 vss 0.00679f
C12430 vdd.n3654 vss 0.00517f
C12431 vdd.n3655 vss 0.00251f
C12432 vdd.n3656 vss 0.00413f
C12433 vdd.n3657 vss 0.0471f
C12434 vdd.t230 vss 0.0471f
C12435 vdd.n3658 vss 0.00425f
C12436 vdd.n3659 vss 0.0424f
C12437 vdd.n3660 vss 0.0132f
C12438 vdd.n3661 vss 0.02f
C12439 vdd.n3662 vss 0.00425f
C12440 vdd.n3663 vss 0.00413f
C12441 vdd.n3664 vss 0.00251f
C12442 vdd.n3665 vss 0.0112f
C12443 vdd.n3666 vss 0.0128f
C12444 vdd.n3667 vss 0.0365f
C12445 vdd.n3668 vss 0.202f
C12446 vdd.n3669 vss 0.00324f
C12447 vdd.n3670 vss 0.0112f
C12448 vdd.n3671 vss 0.0128f
C12449 vdd.n3672 vss 0.00413f
C12450 vdd.n3673 vss 0.00413f
C12451 vdd.n3674 vss 0.0471f
C12452 vdd.n3675 vss 0.00251f
C12453 vdd.t1483 vss 0.0471f
C12454 vdd.n3676 vss 0.00324f
C12455 vdd.n3678 vss 0.00679f
C12456 vdd.n3679 vss 0.00413f
C12457 vdd.n3680 vss 0.00324f
C12458 vdd.n3681 vss 0.00413f
C12459 vdd.n3682 vss 0.0471f
C12460 vdd.n3683 vss 0.00324f
C12461 vdd.n3685 vss 0.00925f
C12462 vdd.t441 vss 0.0471f
C12463 vdd.n3686 vss 0.00425f
C12464 vdd.n3687 vss 0.0424f
C12465 vdd.n3688 vss 0.0132f
C12466 vdd.n3689 vss 0.00324f
C12467 vdd.n3690 vss 0.0128f
C12468 vdd.n3691 vss 0.02f
C12469 vdd.n3692 vss 0.00425f
C12470 vdd.n3693 vss 0.00413f
C12471 vdd.n3694 vss 0.00251f
C12472 vdd.t474 vss 0.0471f
C12473 vdd.n3695 vss 0.00251f
C12474 vdd.n3696 vss 0.00517f
C12475 vdd.n3697 vss 0.00679f
C12476 vdd.n3698 vss 0.00517f
C12477 vdd.n3699 vss 0.00679f
C12478 vdd.n3700 vss 0.02f
C12479 vdd.n3701 vss 0.00425f
C12480 vdd.n3702 vss 0.0424f
C12481 vdd.n3703 vss 0.0132f
C12482 vdd.n3704 vss 0.00925f
C12483 vdd.n3705 vss 0.00425f
C12484 vdd.n3706 vss 0.00413f
C12485 vdd.n3707 vss 0.00324f
C12486 vdd.n3708 vss 0.0471f
C12487 vdd.t475 vss 0.0471f
C12488 vdd.n3709 vss 0.00251f
C12489 vdd.n3710 vss 0.0112f
C12490 vdd.n3711 vss 0.0128f
C12491 vdd.t476 vss 0.00134f
C12492 vdd.t1484 vss 0.0013f
C12493 vdd.n3712 vss 0.0332f
C12494 vdd.n3713 vss 0.0393f
C12495 vdd.n3714 vss 0.0418f
C12496 vdd.n3715 vss 0.00324f
C12497 vdd.n3716 vss 0.0112f
C12498 vdd.n3717 vss 0.0128f
C12499 vdd.n3718 vss 0.00413f
C12500 vdd.n3719 vss 0.00413f
C12501 vdd.n3720 vss 0.0471f
C12502 vdd.n3721 vss 0.00251f
C12503 vdd.t464 vss 0.0471f
C12504 vdd.n3722 vss 0.00324f
C12505 vdd.n3724 vss 0.00679f
C12506 vdd.n3725 vss 0.00413f
C12507 vdd.n3726 vss 0.00324f
C12508 vdd.n3727 vss 0.00413f
C12509 vdd.n3728 vss 0.0471f
C12510 vdd.n3729 vss 0.00324f
C12511 vdd.n3731 vss 0.00925f
C12512 vdd.t234 vss 0.0471f
C12513 vdd.n3732 vss 0.00425f
C12514 vdd.n3733 vss 0.0424f
C12515 vdd.n3734 vss 0.0132f
C12516 vdd.n3735 vss 0.00324f
C12517 vdd.n3736 vss 0.0128f
C12518 vdd.n3737 vss 0.02f
C12519 vdd.n3738 vss 0.00425f
C12520 vdd.n3739 vss 0.00413f
C12521 vdd.n3740 vss 0.00251f
C12522 vdd.t680 vss 0.0471f
C12523 vdd.n3741 vss 0.00251f
C12524 vdd.n3742 vss 0.00517f
C12525 vdd.n3743 vss 0.00679f
C12526 vdd.n3744 vss 0.00517f
C12527 vdd.n3745 vss 0.00679f
C12528 vdd.n3746 vss 0.02f
C12529 vdd.n3747 vss 0.00425f
C12530 vdd.n3748 vss 0.0424f
C12531 vdd.n3749 vss 0.0132f
C12532 vdd.n3750 vss 0.00925f
C12533 vdd.n3751 vss 0.00425f
C12534 vdd.n3752 vss 0.00413f
C12535 vdd.n3753 vss 0.00324f
C12536 vdd.n3754 vss 0.0471f
C12537 vdd.t681 vss 0.0471f
C12538 vdd.n3755 vss 0.00251f
C12539 vdd.n3756 vss 0.0112f
C12540 vdd.n3757 vss 0.0128f
C12541 vdd.t682 vss 0.00134f
C12542 vdd.t465 vss 0.0013f
C12543 vdd.n3758 vss 0.0332f
C12544 vdd.n3759 vss 0.0393f
C12545 vdd.n3760 vss 0.0345f
C12546 vdd.n3761 vss 0.00335f
C12547 vdd.t94 vss 0.0013f
C12548 vdd.n3762 vss 0.0309f
C12549 vdd.n3763 vss 0.00991f
C12550 vdd.n3764 vss 0.0424f
C12551 vdd.n3765 vss 0.00679f
C12552 vdd.n3766 vss 0.00413f
C12553 vdd.n3767 vss 0.0471f
C12554 vdd.n3768 vss 0.00251f
C12555 vdd.n3769 vss 0.00324f
C12556 vdd.n3770 vss 0.0128f
C12557 vdd.n3771 vss 0.00413f
C12558 vdd.n3772 vss 0.00413f
C12559 vdd.n3773 vss 0.0471f
C12560 vdd.n3774 vss 0.00251f
C12561 vdd.n3775 vss 0.00324f
C12562 vdd.n3776 vss 0.00413f
C12563 vdd.n3777 vss 0.00324f
C12564 vdd.n3778 vss 0.0132f
C12565 vdd.n3779 vss 0.0424f
C12566 vdd.n3780 vss 0.00324f
C12567 vdd.n3781 vss 0.00413f
C12568 vdd.n3782 vss 0.02f
C12569 vdd.n3783 vss 0.00425f
C12570 vdd.t724 vss 0.0471f
C12571 vdd.n3785 vss 0.00425f
C12572 vdd.n3786 vss 0.00925f
C12573 vdd.n3787 vss 0.00679f
C12574 vdd.n3788 vss 0.00517f
C12575 vdd.n3789 vss 0.00679f
C12576 vdd.n3790 vss 0.00517f
C12577 vdd.n3791 vss 0.00251f
C12578 vdd.t722 vss 0.0471f
C12579 vdd.n3792 vss 0.0471f
C12580 vdd.t721 vss 0.0471f
C12581 vdd.n3793 vss 0.00251f
C12582 vdd.n3794 vss 0.0105f
C12583 vdd.t723 vss 0.00134f
C12584 vdd.n3795 vss 0.0393f
C12585 vdd.n3796 vss 0.0633f
C12586 vdd.n3797 vss 0.00805f
C12587 vdd.n3798 vss 0.0112f
C12588 vdd.n3799 vss 0.0128f
C12589 vdd.n3800 vss 0.00324f
C12590 vdd.n3801 vss 0.00324f
C12591 vdd.n3802 vss 0.00413f
C12592 vdd.n3803 vss 0.00425f
C12593 vdd.t93 vss 0.0471f
C12594 vdd.n3805 vss 0.00425f
C12595 vdd.n3806 vss 0.00925f
C12596 vdd.n3807 vss 0.0107f
C12597 vdd.n3808 vss 0.0126f
C12598 vdd.n3809 vss 9.89e-19
C12599 vdd.n3810 vss 0.00163f
C12600 vdd.n3811 vss 0.00145f
C12601 vdd.n3812 vss 0.0271f
C12602 vdd.n3813 vss 0.00324f
C12603 vdd.n3814 vss 0.0112f
C12604 vdd.n3815 vss 0.0128f
C12605 vdd.n3816 vss 0.00413f
C12606 vdd.n3817 vss 0.00413f
C12607 vdd.n3818 vss 0.0471f
C12608 vdd.n3819 vss 0.00251f
C12609 vdd.t599 vss 0.0471f
C12610 vdd.n3820 vss 0.00324f
C12611 vdd.n3822 vss 0.00679f
C12612 vdd.n3823 vss 0.00413f
C12613 vdd.n3824 vss 0.00324f
C12614 vdd.n3825 vss 0.00413f
C12615 vdd.n3826 vss 0.0471f
C12616 vdd.n3827 vss 0.00324f
C12617 vdd.n3829 vss 0.00925f
C12618 vdd.t503 vss 0.0471f
C12619 vdd.n3830 vss 0.00425f
C12620 vdd.n3831 vss 0.0424f
C12621 vdd.n3832 vss 0.0132f
C12622 vdd.n3833 vss 0.00324f
C12623 vdd.n3834 vss 0.0128f
C12624 vdd.n3835 vss 0.02f
C12625 vdd.n3836 vss 0.00425f
C12626 vdd.n3837 vss 0.00413f
C12627 vdd.n3838 vss 0.00251f
C12628 vdd.t192 vss 0.0471f
C12629 vdd.n3839 vss 0.00251f
C12630 vdd.n3840 vss 0.00517f
C12631 vdd.n3841 vss 0.00679f
C12632 vdd.n3842 vss 0.00517f
C12633 vdd.n3843 vss 0.00679f
C12634 vdd.n3844 vss 0.02f
C12635 vdd.n3845 vss 0.00425f
C12636 vdd.n3846 vss 0.0424f
C12637 vdd.n3847 vss 0.0132f
C12638 vdd.n3848 vss 0.00925f
C12639 vdd.n3849 vss 0.00425f
C12640 vdd.n3850 vss 0.00413f
C12641 vdd.n3851 vss 0.00324f
C12642 vdd.n3852 vss 0.0471f
C12643 vdd.t193 vss 0.0471f
C12644 vdd.n3853 vss 0.00251f
C12645 vdd.n3854 vss 0.0112f
C12646 vdd.n3855 vss 0.0128f
C12647 vdd.t194 vss 0.00134f
C12648 vdd.t600 vss 0.0013f
C12649 vdd.n3856 vss 0.0332f
C12650 vdd.n3857 vss 0.0393f
C12651 vdd.n3858 vss 0.0418f
C12652 vdd.n3859 vss 0.00324f
C12653 vdd.n3860 vss 0.0112f
C12654 vdd.n3861 vss 0.0128f
C12655 vdd.n3862 vss 0.00413f
C12656 vdd.n3863 vss 0.00413f
C12657 vdd.n3864 vss 0.0471f
C12658 vdd.n3865 vss 0.00251f
C12659 vdd.t460 vss 0.0471f
C12660 vdd.n3866 vss 0.00324f
C12661 vdd.n3868 vss 0.00679f
C12662 vdd.n3869 vss 0.00413f
C12663 vdd.n3870 vss 0.00324f
C12664 vdd.n3871 vss 0.00413f
C12665 vdd.n3872 vss 0.0471f
C12666 vdd.n3873 vss 0.00324f
C12667 vdd.n3875 vss 0.00925f
C12668 vdd.t136 vss 0.0471f
C12669 vdd.n3876 vss 0.00425f
C12670 vdd.n3877 vss 0.0424f
C12671 vdd.n3878 vss 0.0132f
C12672 vdd.n3879 vss 0.00324f
C12673 vdd.n3880 vss 0.0128f
C12674 vdd.n3881 vss 0.02f
C12675 vdd.n3882 vss 0.00425f
C12676 vdd.n3883 vss 0.00413f
C12677 vdd.n3884 vss 0.00251f
C12678 vdd.t1279 vss 0.0471f
C12679 vdd.n3885 vss 0.00251f
C12680 vdd.n3886 vss 0.00517f
C12681 vdd.n3887 vss 0.00679f
C12682 vdd.n3888 vss 0.00517f
C12683 vdd.n3889 vss 0.00679f
C12684 vdd.n3890 vss 0.02f
C12685 vdd.n3891 vss 0.00425f
C12686 vdd.n3892 vss 0.0424f
C12687 vdd.n3893 vss 0.0132f
C12688 vdd.n3894 vss 0.00925f
C12689 vdd.n3895 vss 0.00425f
C12690 vdd.n3896 vss 0.00413f
C12691 vdd.n3897 vss 0.00324f
C12692 vdd.n3898 vss 0.0471f
C12693 vdd.t1280 vss 0.0471f
C12694 vdd.n3899 vss 0.00251f
C12695 vdd.n3900 vss 0.0112f
C12696 vdd.n3901 vss 0.0128f
C12697 vdd.t1281 vss 0.00134f
C12698 vdd.t461 vss 0.0013f
C12699 vdd.n3902 vss 0.0332f
C12700 vdd.n3903 vss 0.0393f
C12701 vdd.n3904 vss 0.0345f
C12702 vdd.n3905 vss 0.00324f
C12703 vdd.n3906 vss 0.0112f
C12704 vdd.n3907 vss 0.0128f
C12705 vdd.n3908 vss 0.00413f
C12706 vdd.n3909 vss 0.00413f
C12707 vdd.n3910 vss 0.0471f
C12708 vdd.n3911 vss 0.00251f
C12709 vdd.t1057 vss 0.0471f
C12710 vdd.n3912 vss 0.00324f
C12711 vdd.n3914 vss 0.00679f
C12712 vdd.n3915 vss 0.00413f
C12713 vdd.n3916 vss 0.00324f
C12714 vdd.n3917 vss 0.00413f
C12715 vdd.n3918 vss 0.0471f
C12716 vdd.n3919 vss 0.00324f
C12717 vdd.n3921 vss 0.00925f
C12718 vdd.t611 vss 0.0471f
C12719 vdd.n3922 vss 0.00425f
C12720 vdd.n3923 vss 0.0424f
C12721 vdd.n3924 vss 0.0132f
C12722 vdd.n3925 vss 0.00324f
C12723 vdd.n3926 vss 0.0128f
C12724 vdd.n3927 vss 0.02f
C12725 vdd.n3928 vss 0.00425f
C12726 vdd.n3929 vss 0.00413f
C12727 vdd.n3930 vss 0.00251f
C12728 vdd.t1132 vss 0.0471f
C12729 vdd.n3931 vss 0.00251f
C12730 vdd.n3932 vss 0.00517f
C12731 vdd.n3933 vss 0.00679f
C12732 vdd.n3934 vss 0.00517f
C12733 vdd.n3935 vss 0.00679f
C12734 vdd.n3936 vss 0.02f
C12735 vdd.n3937 vss 0.00425f
C12736 vdd.n3938 vss 0.0424f
C12737 vdd.n3939 vss 0.0132f
C12738 vdd.n3940 vss 0.00925f
C12739 vdd.n3941 vss 0.00425f
C12740 vdd.n3942 vss 0.00413f
C12741 vdd.n3943 vss 0.00324f
C12742 vdd.n3944 vss 0.0471f
C12743 vdd.t1133 vss 0.0471f
C12744 vdd.n3945 vss 0.00251f
C12745 vdd.n3946 vss 0.0112f
C12746 vdd.n3947 vss 0.0128f
C12747 vdd.t1134 vss 0.00134f
C12748 vdd.t1058 vss 0.0013f
C12749 vdd.n3948 vss 0.0332f
C12750 vdd.n3949 vss 0.0393f
C12751 vdd.n3950 vss 0.0418f
C12752 vdd.n3951 vss 0.00324f
C12753 vdd.n3952 vss 0.0112f
C12754 vdd.n3953 vss 0.0128f
C12755 vdd.n3954 vss 0.00413f
C12756 vdd.n3955 vss 0.00413f
C12757 vdd.n3956 vss 0.0471f
C12758 vdd.n3957 vss 0.00251f
C12759 vdd.t603 vss 0.0471f
C12760 vdd.n3958 vss 0.00324f
C12761 vdd.n3960 vss 0.00679f
C12762 vdd.n3961 vss 0.00413f
C12763 vdd.n3962 vss 0.00324f
C12764 vdd.n3963 vss 0.00413f
C12765 vdd.n3964 vss 0.0471f
C12766 vdd.n3965 vss 0.00324f
C12767 vdd.n3967 vss 0.00925f
C12768 vdd.t802 vss 0.0471f
C12769 vdd.n3968 vss 0.00425f
C12770 vdd.n3969 vss 0.0424f
C12771 vdd.n3970 vss 0.0132f
C12772 vdd.n3971 vss 0.00324f
C12773 vdd.n3972 vss 0.0128f
C12774 vdd.n3973 vss 0.02f
C12775 vdd.n3974 vss 0.00425f
C12776 vdd.n3975 vss 0.00413f
C12777 vdd.n3976 vss 0.00251f
C12778 vdd.t1207 vss 0.0471f
C12779 vdd.n3977 vss 0.00251f
C12780 vdd.n3978 vss 0.00517f
C12781 vdd.n3979 vss 0.00679f
C12782 vdd.n3980 vss 0.00517f
C12783 vdd.n3981 vss 0.00679f
C12784 vdd.n3982 vss 0.02f
C12785 vdd.n3983 vss 0.00425f
C12786 vdd.n3984 vss 0.0424f
C12787 vdd.n3985 vss 0.0132f
C12788 vdd.n3986 vss 0.00925f
C12789 vdd.n3987 vss 0.00425f
C12790 vdd.n3988 vss 0.00413f
C12791 vdd.n3989 vss 0.00324f
C12792 vdd.n3990 vss 0.0471f
C12793 vdd.t1208 vss 0.0471f
C12794 vdd.n3991 vss 0.00251f
C12795 vdd.n3992 vss 0.0112f
C12796 vdd.n3993 vss 0.0128f
C12797 vdd.t1209 vss 0.00134f
C12798 vdd.t604 vss 0.0013f
C12799 vdd.n3994 vss 0.0332f
C12800 vdd.n3995 vss 0.0393f
C12801 vdd.n3996 vss 0.0345f
C12802 vdd.n3997 vss 0.00335f
C12803 vdd.t100 vss 0.0013f
C12804 vdd.n3998 vss 0.0309f
C12805 vdd.n3999 vss 0.00991f
C12806 vdd.n4000 vss 0.0424f
C12807 vdd.n4001 vss 0.00679f
C12808 vdd.n4002 vss 0.00413f
C12809 vdd.n4003 vss 0.0471f
C12810 vdd.n4004 vss 0.00251f
C12811 vdd.n4005 vss 0.00324f
C12812 vdd.n4006 vss 0.0128f
C12813 vdd.n4007 vss 0.00413f
C12814 vdd.n4008 vss 0.00413f
C12815 vdd.n4009 vss 0.0471f
C12816 vdd.n4010 vss 0.00251f
C12817 vdd.n4011 vss 0.00324f
C12818 vdd.n4012 vss 0.00413f
C12819 vdd.n4013 vss 0.00324f
C12820 vdd.n4014 vss 0.0132f
C12821 vdd.n4015 vss 0.0424f
C12822 vdd.n4016 vss 0.00324f
C12823 vdd.n4017 vss 0.00413f
C12824 vdd.n4018 vss 0.02f
C12825 vdd.n4019 vss 0.00425f
C12826 vdd.t1422 vss 0.0471f
C12827 vdd.n4021 vss 0.00425f
C12828 vdd.n4022 vss 0.00925f
C12829 vdd.n4023 vss 0.00679f
C12830 vdd.n4024 vss 0.00517f
C12831 vdd.n4025 vss 0.00679f
C12832 vdd.n4026 vss 0.00517f
C12833 vdd.n4027 vss 0.00251f
C12834 vdd.t1515 vss 0.0471f
C12835 vdd.n4028 vss 0.0471f
C12836 vdd.t1517 vss 0.0471f
C12837 vdd.n4029 vss 0.00251f
C12838 vdd.n4030 vss 0.0105f
C12839 vdd.t1516 vss 0.00134f
C12840 vdd.n4031 vss 0.0393f
C12841 vdd.n4032 vss 0.0633f
C12842 vdd.n4033 vss 0.00805f
C12843 vdd.n4034 vss 0.0112f
C12844 vdd.n4035 vss 0.0128f
C12845 vdd.n4036 vss 0.00324f
C12846 vdd.n4037 vss 0.00324f
C12847 vdd.n4038 vss 0.00413f
C12848 vdd.n4039 vss 0.00425f
C12849 vdd.t99 vss 0.0471f
C12850 vdd.n4041 vss 0.00425f
C12851 vdd.n4042 vss 0.00925f
C12852 vdd.n4043 vss 0.0107f
C12853 vdd.n4044 vss 0.0126f
C12854 vdd.n4045 vss 9.89e-19
C12855 vdd.n4046 vss 0.00163f
C12856 vdd.n4047 vss 0.00145f
C12857 vdd.n4048 vss 0.0271f
C12858 vdd.n4049 vss 0.00324f
C12859 vdd.n4050 vss 0.0112f
C12860 vdd.n4051 vss 0.0128f
C12861 vdd.n4052 vss 0.00413f
C12862 vdd.n4053 vss 0.00413f
C12863 vdd.n4054 vss 0.0471f
C12864 vdd.n4055 vss 0.00251f
C12865 vdd.t468 vss 0.0471f
C12866 vdd.n4056 vss 0.00324f
C12867 vdd.n4058 vss 0.00679f
C12868 vdd.n4059 vss 0.00413f
C12869 vdd.n4060 vss 0.00324f
C12870 vdd.n4061 vss 0.00413f
C12871 vdd.n4062 vss 0.0471f
C12872 vdd.n4063 vss 0.00324f
C12873 vdd.n4065 vss 0.00925f
C12874 vdd.t473 vss 0.0471f
C12875 vdd.n4066 vss 0.00425f
C12876 vdd.n4067 vss 0.0424f
C12877 vdd.n4068 vss 0.0132f
C12878 vdd.n4069 vss 0.00324f
C12879 vdd.n4070 vss 0.0128f
C12880 vdd.n4071 vss 0.02f
C12881 vdd.n4072 vss 0.00425f
C12882 vdd.n4073 vss 0.00413f
C12883 vdd.n4074 vss 0.00251f
C12884 vdd.t1407 vss 0.0471f
C12885 vdd.n4075 vss 0.00251f
C12886 vdd.n4076 vss 0.00517f
C12887 vdd.n4077 vss 0.00679f
C12888 vdd.n4078 vss 0.00517f
C12889 vdd.n4079 vss 0.00679f
C12890 vdd.n4080 vss 0.02f
C12891 vdd.n4081 vss 0.00425f
C12892 vdd.n4082 vss 0.0424f
C12893 vdd.n4083 vss 0.0132f
C12894 vdd.n4084 vss 0.00925f
C12895 vdd.n4085 vss 0.00425f
C12896 vdd.n4086 vss 0.00413f
C12897 vdd.n4087 vss 0.00324f
C12898 vdd.n4088 vss 0.0471f
C12899 vdd.t1408 vss 0.0471f
C12900 vdd.n4089 vss 0.00251f
C12901 vdd.n4090 vss 0.0112f
C12902 vdd.n4091 vss 0.0128f
C12903 vdd.t1409 vss 0.00134f
C12904 vdd.t469 vss 0.0013f
C12905 vdd.n4092 vss 0.0332f
C12906 vdd.n4093 vss 0.0393f
C12907 vdd.n4094 vss 0.0418f
C12908 vdd.t395 vss 0.00134f
C12909 vdd.t204 vss 0.0013f
C12910 vdd.n4095 vss 0.032f
C12911 vdd.n4096 vss 0.0393f
C12912 vdd.n4097 vss 0.00324f
C12913 vdd.n4098 vss 0.0112f
C12914 vdd.n4099 vss 0.0128f
C12915 vdd.n4100 vss 0.00413f
C12916 vdd.t393 vss 0.0471f
C12917 vdd.n4101 vss 0.00324f
C12918 vdd.n4103 vss 0.00925f
C12919 vdd.n4104 vss 0.00413f
C12920 vdd.n4105 vss 0.00679f
C12921 vdd.n4106 vss 0.00413f
C12922 vdd.n4107 vss 0.0471f
C12923 vdd.n4108 vss 0.00324f
C12924 vdd.n4109 vss 0.0471f
C12925 vdd.n4110 vss 0.00324f
C12926 vdd.n4111 vss 0.0424f
C12927 vdd.t203 vss 0.0471f
C12928 vdd.n4113 vss 0.00425f
C12929 vdd.n4114 vss 0.00925f
C12930 vdd.n4115 vss 0.0132f
C12931 vdd.n4116 vss 0.00324f
C12932 vdd.n4117 vss 0.0128f
C12933 vdd.n4118 vss 0.02f
C12934 vdd.n4119 vss 0.00425f
C12935 vdd.n4120 vss 0.00413f
C12936 vdd.n4121 vss 0.00251f
C12937 vdd.t394 vss 0.0471f
C12938 vdd.n4122 vss 0.00251f
C12939 vdd.n4123 vss 0.00517f
C12940 vdd.n4124 vss 0.00679f
C12941 vdd.n4125 vss 0.00324f
C12942 vdd.n4126 vss 0.00679f
C12943 vdd.n4127 vss 0.00517f
C12944 vdd.n4128 vss 0.00251f
C12945 vdd.n4129 vss 0.00413f
C12946 vdd.n4130 vss 0.0471f
C12947 vdd.t440 vss 0.0471f
C12948 vdd.n4131 vss 0.00425f
C12949 vdd.n4132 vss 0.0424f
C12950 vdd.n4133 vss 0.0132f
C12951 vdd.n4134 vss 0.02f
C12952 vdd.n4135 vss 0.00425f
C12953 vdd.n4136 vss 0.00413f
C12954 vdd.n4137 vss 0.00251f
C12955 vdd.n4138 vss 0.0112f
C12956 vdd.n4139 vss 0.0128f
C12957 vdd.n4140 vss 0.0418f
C12958 vdd.t622 vss 0.00134f
C12959 vdd.t555 vss 0.0013f
C12960 vdd.n4141 vss 0.032f
C12961 vdd.n4142 vss 0.0393f
C12962 vdd.n4143 vss 0.00324f
C12963 vdd.n4144 vss 0.0112f
C12964 vdd.n4145 vss 0.0128f
C12965 vdd.n4146 vss 0.00413f
C12966 vdd.t623 vss 0.0471f
C12967 vdd.n4147 vss 0.00324f
C12968 vdd.n4149 vss 0.00925f
C12969 vdd.n4150 vss 0.00413f
C12970 vdd.n4151 vss 0.00679f
C12971 vdd.n4152 vss 0.00413f
C12972 vdd.n4153 vss 0.0471f
C12973 vdd.n4154 vss 0.00324f
C12974 vdd.n4155 vss 0.0471f
C12975 vdd.n4156 vss 0.00324f
C12976 vdd.n4157 vss 0.0424f
C12977 vdd.t554 vss 0.0471f
C12978 vdd.n4159 vss 0.00425f
C12979 vdd.n4160 vss 0.00925f
C12980 vdd.n4161 vss 0.0132f
C12981 vdd.n4162 vss 0.00324f
C12982 vdd.n4163 vss 0.0128f
C12983 vdd.n4164 vss 0.02f
C12984 vdd.n4165 vss 0.00425f
C12985 vdd.n4166 vss 0.00413f
C12986 vdd.n4167 vss 0.00251f
C12987 vdd.t621 vss 0.0471f
C12988 vdd.n4168 vss 0.00251f
C12989 vdd.n4169 vss 0.00517f
C12990 vdd.n4170 vss 0.00679f
C12991 vdd.n4171 vss 0.00324f
C12992 vdd.n4172 vss 0.00679f
C12993 vdd.n4173 vss 0.00517f
C12994 vdd.n4174 vss 0.00251f
C12995 vdd.n4175 vss 0.00413f
C12996 vdd.n4176 vss 0.0471f
C12997 vdd.t477 vss 0.0471f
C12998 vdd.n4177 vss 0.00425f
C12999 vdd.n4178 vss 0.0424f
C13000 vdd.n4179 vss 0.0132f
C13001 vdd.n4180 vss 0.02f
C13002 vdd.n4181 vss 0.00425f
C13003 vdd.n4182 vss 0.00413f
C13004 vdd.n4183 vss 0.00251f
C13005 vdd.n4184 vss 0.0112f
C13006 vdd.n4185 vss 0.0128f
C13007 vdd.n4186 vss 0.0369f
C13008 vdd.n4187 vss 0.00335f
C13009 vdd.t1456 vss 0.0013f
C13010 vdd.n4188 vss 0.0309f
C13011 vdd.n4189 vss 0.0107f
C13012 vdd.n4190 vss 0.0128f
C13013 vdd.n4191 vss 0.0424f
C13014 vdd.t1455 vss 0.0471f
C13015 vdd.n4192 vss 0.00324f
C13016 vdd.n4193 vss 0.0471f
C13017 vdd.t710 vss 0.0471f
C13018 vdd.n4194 vss 0.00413f
C13019 vdd.n4195 vss 0.00324f
C13020 vdd.t711 vss 0.00134f
C13021 vdd.n4196 vss 0.0393f
C13022 vdd.n4197 vss 0.0128f
C13023 vdd.t712 vss 0.0471f
C13024 vdd.n4198 vss 0.00324f
C13025 vdd.n4200 vss 0.00925f
C13026 vdd.n4201 vss 0.0471f
C13027 vdd.n4202 vss 0.00324f
C13028 vdd.n4203 vss 0.00413f
C13029 vdd.n4204 vss 0.00324f
C13030 vdd.n4205 vss 0.00679f
C13031 vdd.n4207 vss 0.00925f
C13032 vdd.n4208 vss 0.00425f
C13033 vdd.n4209 vss 0.00413f
C13034 vdd.n4210 vss 0.00251f
C13035 vdd.n4211 vss 0.00517f
C13036 vdd.n4212 vss 0.00679f
C13037 vdd.n4213 vss 0.00324f
C13038 vdd.n4214 vss 0.00679f
C13039 vdd.n4215 vss 0.00517f
C13040 vdd.n4216 vss 0.00251f
C13041 vdd.n4217 vss 0.00413f
C13042 vdd.n4218 vss 0.0471f
C13043 vdd.t1067 vss 0.0471f
C13044 vdd.n4219 vss 0.00425f
C13045 vdd.n4220 vss 0.0424f
C13046 vdd.n4221 vss 0.0132f
C13047 vdd.n4222 vss 0.02f
C13048 vdd.n4223 vss 0.00425f
C13049 vdd.n4224 vss 0.00413f
C13050 vdd.n4225 vss 0.00251f
C13051 vdd.n4226 vss 0.0105f
C13052 vdd.n4227 vss 0.0633f
C13053 vdd.n4228 vss 0.00805f
C13054 vdd.n4229 vss 0.0112f
C13055 vdd.n4230 vss 0.00251f
C13056 vdd.n4231 vss 0.00413f
C13057 vdd.n4232 vss 0.00425f
C13058 vdd.n4233 vss 0.00991f
C13059 vdd.n4234 vss 0.0126f
C13060 vdd.n4235 vss 9.89e-19
C13061 vdd.n4236 vss 0.0011f
C13062 vdd.n4237 vss 0.0271f
C13063 vdd.t1184 vss 0.00134f
C13064 vdd.t1291 vss 0.0013f
C13065 vdd.n4238 vss 0.032f
C13066 vdd.n4239 vss 0.0393f
C13067 vdd.n4240 vss 0.00324f
C13068 vdd.n4241 vss 0.0112f
C13069 vdd.n4242 vss 0.0128f
C13070 vdd.n4243 vss 0.00413f
C13071 vdd.t1185 vss 0.0471f
C13072 vdd.n4244 vss 0.00324f
C13073 vdd.n4246 vss 0.00925f
C13074 vdd.n4247 vss 0.00413f
C13075 vdd.n4248 vss 0.00679f
C13076 vdd.n4249 vss 0.00413f
C13077 vdd.n4250 vss 0.0471f
C13078 vdd.n4251 vss 0.00324f
C13079 vdd.n4252 vss 0.0471f
C13080 vdd.n4253 vss 0.00324f
C13081 vdd.n4254 vss 0.0424f
C13082 vdd.t1290 vss 0.0471f
C13083 vdd.n4256 vss 0.00425f
C13084 vdd.n4257 vss 0.00925f
C13085 vdd.n4258 vss 0.0132f
C13086 vdd.n4259 vss 0.00324f
C13087 vdd.n4260 vss 0.0128f
C13088 vdd.n4261 vss 0.02f
C13089 vdd.n4262 vss 0.00425f
C13090 vdd.n4263 vss 0.00413f
C13091 vdd.n4264 vss 0.00251f
C13092 vdd.t1183 vss 0.0471f
C13093 vdd.n4265 vss 0.00251f
C13094 vdd.n4266 vss 0.00517f
C13095 vdd.n4267 vss 0.00679f
C13096 vdd.n4268 vss 0.00324f
C13097 vdd.n4269 vss 0.00679f
C13098 vdd.n4270 vss 0.00517f
C13099 vdd.n4271 vss 0.00251f
C13100 vdd.n4272 vss 0.00413f
C13101 vdd.n4273 vss 0.0471f
C13102 vdd.t114 vss 0.0471f
C13103 vdd.n4274 vss 0.00425f
C13104 vdd.n4275 vss 0.0424f
C13105 vdd.n4276 vss 0.0132f
C13106 vdd.n4277 vss 0.02f
C13107 vdd.n4278 vss 0.00425f
C13108 vdd.n4279 vss 0.00413f
C13109 vdd.n4280 vss 0.00251f
C13110 vdd.n4281 vss 0.0112f
C13111 vdd.n4282 vss 0.0128f
C13112 vdd.n4283 vss 0.0418f
C13113 vdd.t420 vss 0.00134f
C13114 vdd.t1317 vss 0.0013f
C13115 vdd.n4284 vss 0.032f
C13116 vdd.n4285 vss 0.0393f
C13117 vdd.n4286 vss 0.00324f
C13118 vdd.n4287 vss 0.0112f
C13119 vdd.n4288 vss 0.0128f
C13120 vdd.n4289 vss 0.00413f
C13121 vdd.t421 vss 0.0471f
C13122 vdd.n4290 vss 0.00324f
C13123 vdd.n4292 vss 0.00925f
C13124 vdd.n4293 vss 0.00413f
C13125 vdd.n4294 vss 0.00679f
C13126 vdd.n4295 vss 0.00413f
C13127 vdd.n4296 vss 0.0471f
C13128 vdd.n4297 vss 0.00324f
C13129 vdd.n4298 vss 0.0471f
C13130 vdd.n4299 vss 0.00324f
C13131 vdd.n4300 vss 0.0424f
C13132 vdd.t1316 vss 0.0471f
C13133 vdd.n4302 vss 0.00425f
C13134 vdd.n4303 vss 0.00925f
C13135 vdd.n4304 vss 0.0132f
C13136 vdd.n4305 vss 0.00324f
C13137 vdd.n4306 vss 0.0128f
C13138 vdd.n4307 vss 0.02f
C13139 vdd.n4308 vss 0.00425f
C13140 vdd.n4309 vss 0.00413f
C13141 vdd.n4310 vss 0.00251f
C13142 vdd.t419 vss 0.0471f
C13143 vdd.n4311 vss 0.00251f
C13144 vdd.n4312 vss 0.00517f
C13145 vdd.n4313 vss 0.00679f
C13146 vdd.n4314 vss 0.00324f
C13147 vdd.n4315 vss 0.00679f
C13148 vdd.n4316 vss 0.00517f
C13149 vdd.n4317 vss 0.00251f
C13150 vdd.n4318 vss 0.00413f
C13151 vdd.n4319 vss 0.0471f
C13152 vdd.t810 vss 0.0471f
C13153 vdd.n4320 vss 0.00425f
C13154 vdd.n4321 vss 0.0424f
C13155 vdd.n4322 vss 0.0132f
C13156 vdd.n4323 vss 0.02f
C13157 vdd.n4324 vss 0.00425f
C13158 vdd.n4325 vss 0.00413f
C13159 vdd.n4326 vss 0.00251f
C13160 vdd.n4327 vss 0.0112f
C13161 vdd.n4328 vss 0.0128f
C13162 vdd.n4329 vss 0.0365f
C13163 vdd.t1425 vss 0.00134f
C13164 vdd.t1056 vss 0.0013f
C13165 vdd.n4330 vss 0.032f
C13166 vdd.n4331 vss 0.0393f
C13167 vdd.n4332 vss 0.00324f
C13168 vdd.n4333 vss 0.0112f
C13169 vdd.n4334 vss 0.0128f
C13170 vdd.n4335 vss 0.00413f
C13171 vdd.t1426 vss 0.0471f
C13172 vdd.n4336 vss 0.00324f
C13173 vdd.n4338 vss 0.00925f
C13174 vdd.n4339 vss 0.00413f
C13175 vdd.n4340 vss 0.00679f
C13176 vdd.n4341 vss 0.00413f
C13177 vdd.n4342 vss 0.0471f
C13178 vdd.n4343 vss 0.00324f
C13179 vdd.n4344 vss 0.0471f
C13180 vdd.n4345 vss 0.00324f
C13181 vdd.n4346 vss 0.0424f
C13182 vdd.t1055 vss 0.0471f
C13183 vdd.n4348 vss 0.00425f
C13184 vdd.n4349 vss 0.00925f
C13185 vdd.n4350 vss 0.0132f
C13186 vdd.n4351 vss 0.00324f
C13187 vdd.n4352 vss 0.0128f
C13188 vdd.n4353 vss 0.02f
C13189 vdd.n4354 vss 0.00425f
C13190 vdd.n4355 vss 0.00413f
C13191 vdd.n4356 vss 0.00251f
C13192 vdd.t1424 vss 0.0471f
C13193 vdd.n4357 vss 0.00251f
C13194 vdd.n4358 vss 0.00517f
C13195 vdd.n4359 vss 0.00679f
C13196 vdd.n4360 vss 0.00324f
C13197 vdd.n4361 vss 0.00679f
C13198 vdd.n4362 vss 0.00517f
C13199 vdd.n4363 vss 0.00251f
C13200 vdd.n4364 vss 0.00413f
C13201 vdd.n4365 vss 0.0471f
C13202 vdd.t1427 vss 0.0471f
C13203 vdd.n4366 vss 0.00425f
C13204 vdd.n4367 vss 0.0424f
C13205 vdd.n4368 vss 0.0132f
C13206 vdd.n4369 vss 0.02f
C13207 vdd.n4370 vss 0.00425f
C13208 vdd.n4371 vss 0.00413f
C13209 vdd.n4372 vss 0.00251f
C13210 vdd.n4373 vss 0.0112f
C13211 vdd.n4374 vss 0.0128f
C13212 vdd.n4375 vss 0.0418f
C13213 vdd.t1436 vss 0.00134f
C13214 vdd.t571 vss 0.0013f
C13215 vdd.n4376 vss 0.032f
C13216 vdd.n4377 vss 0.0393f
C13217 vdd.n4378 vss 0.00324f
C13218 vdd.n4379 vss 0.0112f
C13219 vdd.n4380 vss 0.0128f
C13220 vdd.n4381 vss 0.00413f
C13221 vdd.t1437 vss 0.0471f
C13222 vdd.n4382 vss 0.00324f
C13223 vdd.n4384 vss 0.00925f
C13224 vdd.n4385 vss 0.00413f
C13225 vdd.n4386 vss 0.00679f
C13226 vdd.n4387 vss 0.00413f
C13227 vdd.n4388 vss 0.0471f
C13228 vdd.n4389 vss 0.00324f
C13229 vdd.n4390 vss 0.0471f
C13230 vdd.n4391 vss 0.00324f
C13231 vdd.n4392 vss 0.0424f
C13232 vdd.t570 vss 0.0471f
C13233 vdd.n4394 vss 0.00425f
C13234 vdd.n4395 vss 0.00925f
C13235 vdd.n4396 vss 0.0132f
C13236 vdd.n4397 vss 0.00324f
C13237 vdd.n4398 vss 0.0128f
C13238 vdd.n4399 vss 0.02f
C13239 vdd.n4400 vss 0.00425f
C13240 vdd.n4401 vss 0.00413f
C13241 vdd.n4402 vss 0.00251f
C13242 vdd.t1435 vss 0.0471f
C13243 vdd.n4403 vss 0.00251f
C13244 vdd.n4404 vss 0.00517f
C13245 vdd.n4405 vss 0.00679f
C13246 vdd.n4406 vss 0.00324f
C13247 vdd.n4407 vss 0.00679f
C13248 vdd.n4408 vss 0.00517f
C13249 vdd.n4409 vss 0.00251f
C13250 vdd.n4410 vss 0.00413f
C13251 vdd.n4411 vss 0.0471f
C13252 vdd.t1225 vss 0.0471f
C13253 vdd.n4412 vss 0.00425f
C13254 vdd.n4413 vss 0.0424f
C13255 vdd.n4414 vss 0.0132f
C13256 vdd.n4415 vss 0.02f
C13257 vdd.n4416 vss 0.00425f
C13258 vdd.n4417 vss 0.00413f
C13259 vdd.n4418 vss 0.00251f
C13260 vdd.n4419 vss 0.0112f
C13261 vdd.n4420 vss 0.0128f
C13262 vdd.n4421 vss 0.0369f
C13263 vdd.n4422 vss 0.00335f
C13264 vdd.t1458 vss 0.0013f
C13265 vdd.n4423 vss 0.0309f
C13266 vdd.n4424 vss 0.0107f
C13267 vdd.n4425 vss 0.0128f
C13268 vdd.n4426 vss 0.0424f
C13269 vdd.t1457 vss 0.0471f
C13270 vdd.n4427 vss 0.00324f
C13271 vdd.n4428 vss 0.0471f
C13272 vdd.t1239 vss 0.0471f
C13273 vdd.n4429 vss 0.00413f
C13274 vdd.n4430 vss 0.00324f
C13275 vdd.t1240 vss 0.00134f
C13276 vdd.n4431 vss 0.0393f
C13277 vdd.n4432 vss 0.0128f
C13278 vdd.t1241 vss 0.0471f
C13279 vdd.n4433 vss 0.00324f
C13280 vdd.n4435 vss 0.00925f
C13281 vdd.n4436 vss 0.0471f
C13282 vdd.n4437 vss 0.00324f
C13283 vdd.n4438 vss 0.00413f
C13284 vdd.n4439 vss 0.00324f
C13285 vdd.n4440 vss 0.00679f
C13286 vdd.n4442 vss 0.00925f
C13287 vdd.n4443 vss 0.00425f
C13288 vdd.n4444 vss 0.00413f
C13289 vdd.n4445 vss 0.00251f
C13290 vdd.n4446 vss 0.00517f
C13291 vdd.n4447 vss 0.00679f
C13292 vdd.n4448 vss 0.00324f
C13293 vdd.n4449 vss 0.00679f
C13294 vdd.n4450 vss 0.00517f
C13295 vdd.n4451 vss 0.00251f
C13296 vdd.n4452 vss 0.00413f
C13297 vdd.n4453 vss 0.0471f
C13298 vdd.t455 vss 0.0471f
C13299 vdd.n4454 vss 0.00425f
C13300 vdd.n4455 vss 0.0424f
C13301 vdd.n4456 vss 0.0132f
C13302 vdd.n4457 vss 0.02f
C13303 vdd.n4458 vss 0.00425f
C13304 vdd.n4459 vss 0.00413f
C13305 vdd.n4460 vss 0.00251f
C13306 vdd.n4461 vss 0.0105f
C13307 vdd.n4462 vss 0.0633f
C13308 vdd.n4463 vss 0.00805f
C13309 vdd.n4464 vss 0.0112f
C13310 vdd.n4465 vss 0.00251f
C13311 vdd.n4466 vss 0.00413f
C13312 vdd.n4467 vss 0.00425f
C13313 vdd.n4468 vss 0.00991f
C13314 vdd.n4469 vss 0.0126f
C13315 vdd.n4470 vss 9.89e-19
C13316 vdd.n4471 vss 0.0011f
C13317 vdd.n4472 vss 0.0271f
C13318 vdd.t1232 vss 0.00134f
C13319 vdd.t1046 vss 0.0013f
C13320 vdd.n4473 vss 0.032f
C13321 vdd.n4474 vss 0.0393f
C13322 vdd.n4475 vss 0.00324f
C13323 vdd.n4476 vss 0.0112f
C13324 vdd.n4477 vss 0.0128f
C13325 vdd.n4478 vss 0.00413f
C13326 vdd.t1233 vss 0.0471f
C13327 vdd.n4479 vss 0.00324f
C13328 vdd.n4481 vss 0.00925f
C13329 vdd.n4482 vss 0.00413f
C13330 vdd.n4483 vss 0.00679f
C13331 vdd.n4484 vss 0.00413f
C13332 vdd.n4485 vss 0.0471f
C13333 vdd.n4486 vss 0.00324f
C13334 vdd.n4487 vss 0.0471f
C13335 vdd.n4488 vss 0.00324f
C13336 vdd.n4489 vss 0.0424f
C13337 vdd.t1045 vss 0.0471f
C13338 vdd.n4491 vss 0.00425f
C13339 vdd.n4492 vss 0.00925f
C13340 vdd.n4493 vss 0.0132f
C13341 vdd.n4494 vss 0.00324f
C13342 vdd.n4495 vss 0.0128f
C13343 vdd.n4496 vss 0.02f
C13344 vdd.n4497 vss 0.00425f
C13345 vdd.n4498 vss 0.00413f
C13346 vdd.n4499 vss 0.00251f
C13347 vdd.t1231 vss 0.0471f
C13348 vdd.n4500 vss 0.00251f
C13349 vdd.n4501 vss 0.00517f
C13350 vdd.n4502 vss 0.00679f
C13351 vdd.n4503 vss 0.00324f
C13352 vdd.n4504 vss 0.00679f
C13353 vdd.n4505 vss 0.00517f
C13354 vdd.n4506 vss 0.00251f
C13355 vdd.n4507 vss 0.00413f
C13356 vdd.n4508 vss 0.0471f
C13357 vdd.t951 vss 0.0471f
C13358 vdd.n4509 vss 0.00425f
C13359 vdd.n4510 vss 0.0424f
C13360 vdd.n4511 vss 0.0132f
C13361 vdd.n4512 vss 0.02f
C13362 vdd.n4513 vss 0.00425f
C13363 vdd.n4514 vss 0.00413f
C13364 vdd.n4515 vss 0.00251f
C13365 vdd.n4516 vss 0.0112f
C13366 vdd.n4517 vss 0.0128f
C13367 vdd.n4518 vss 0.0418f
C13368 vdd.t1001 vss 0.0013f
C13369 vdd.t697 vss 0.00134f
C13370 vdd.n4519 vss 0.00324f
C13371 vdd.n4520 vss 0.0112f
C13372 vdd.n4521 vss 0.0128f
C13373 vdd.n4522 vss 0.00413f
C13374 vdd.t698 vss 0.0471f
C13375 vdd.n4523 vss 0.00324f
C13376 vdd.n4525 vss 0.00925f
C13377 vdd.n4526 vss 0.00413f
C13378 vdd.n4527 vss 0.00679f
C13379 vdd.n4528 vss 0.00413f
C13380 vdd.n4529 vss 0.0471f
C13381 vdd.n4530 vss 0.00324f
C13382 vdd.n4531 vss 0.0471f
C13383 vdd.n4532 vss 0.00324f
C13384 vdd.n4533 vss 0.0424f
C13385 vdd.t1000 vss 0.0471f
C13386 vdd.n4535 vss 0.00425f
C13387 vdd.n4536 vss 0.00925f
C13388 vdd.n4537 vss 0.0132f
C13389 vdd.n4538 vss 0.00324f
C13390 vdd.n4539 vss 0.0128f
C13391 vdd.n4540 vss 0.02f
C13392 vdd.n4541 vss 0.00425f
C13393 vdd.n4542 vss 0.00413f
C13394 vdd.n4543 vss 0.00251f
C13395 vdd.t696 vss 0.0471f
C13396 vdd.n4544 vss 0.00251f
C13397 vdd.n4545 vss 0.00517f
C13398 vdd.n4546 vss 0.00679f
C13399 vdd.n4547 vss 0.00324f
C13400 vdd.n4548 vss 0.00679f
C13401 vdd.n4549 vss 0.00517f
C13402 vdd.n4550 vss 0.00251f
C13403 vdd.n4551 vss 0.00413f
C13404 vdd.n4552 vss 0.0471f
C13405 vdd.t1148 vss 0.0471f
C13406 vdd.n4553 vss 0.00425f
C13407 vdd.n4554 vss 0.0424f
C13408 vdd.n4555 vss 0.0132f
C13409 vdd.n4556 vss 0.02f
C13410 vdd.n4557 vss 0.00425f
C13411 vdd.n4558 vss 0.00413f
C13412 vdd.n4559 vss 0.00251f
C13413 vdd.n4560 vss 0.0112f
C13414 vdd.n4561 vss 0.0128f
C13415 vdd.t448 vss 0.00134f
C13416 vdd.t175 vss 0.0013f
C13417 vdd.n4562 vss 0.032f
C13418 vdd.n4563 vss 0.0393f
C13419 vdd.n4564 vss 0.00324f
C13420 vdd.n4565 vss 0.0112f
C13421 vdd.n4566 vss 0.0128f
C13422 vdd.n4567 vss 0.00413f
C13423 vdd.t446 vss 0.0471f
C13424 vdd.n4568 vss 0.00324f
C13425 vdd.n4570 vss 0.00925f
C13426 vdd.n4571 vss 0.00413f
C13427 vdd.n4572 vss 0.00679f
C13428 vdd.n4573 vss 0.00413f
C13429 vdd.n4574 vss 0.0471f
C13430 vdd.n4575 vss 0.00324f
C13431 vdd.n4576 vss 0.0471f
C13432 vdd.n4577 vss 0.00324f
C13433 vdd.n4578 vss 0.0424f
C13434 vdd.t174 vss 0.0471f
C13435 vdd.n4580 vss 0.00425f
C13436 vdd.n4581 vss 0.00925f
C13437 vdd.n4582 vss 0.0132f
C13438 vdd.n4583 vss 0.00324f
C13439 vdd.n4584 vss 0.0128f
C13440 vdd.n4585 vss 0.02f
C13441 vdd.n4586 vss 0.00425f
C13442 vdd.n4587 vss 0.00413f
C13443 vdd.n4588 vss 0.00251f
C13444 vdd.t447 vss 0.0471f
C13445 vdd.n4589 vss 0.00251f
C13446 vdd.n4590 vss 0.00517f
C13447 vdd.n4591 vss 0.00679f
C13448 vdd.n4592 vss 0.00324f
C13449 vdd.n4593 vss 0.00679f
C13450 vdd.n4594 vss 0.00517f
C13451 vdd.n4595 vss 0.00251f
C13452 vdd.n4596 vss 0.00413f
C13453 vdd.n4597 vss 0.0471f
C13454 vdd.t145 vss 0.0471f
C13455 vdd.n4598 vss 0.00425f
C13456 vdd.n4599 vss 0.0424f
C13457 vdd.n4600 vss 0.0132f
C13458 vdd.n4601 vss 0.02f
C13459 vdd.n4602 vss 0.00425f
C13460 vdd.n4603 vss 0.00413f
C13461 vdd.n4604 vss 0.00251f
C13462 vdd.n4605 vss 0.0112f
C13463 vdd.n4606 vss 0.0128f
C13464 vdd.n4607 vss 0.119f
C13465 vdd.n4608 vss 0.118f
C13466 vdd.n4609 vss 0.0393f
C13467 vdd.n4610 vss 0.032f
C13468 vdd.n4611 vss 0.0608f
C13469 vdd.t150 vss 0.00134f
C13470 vdd.t198 vss 0.0013f
C13471 vdd.n4612 vss 0.032f
C13472 vdd.n4613 vss 0.0393f
C13473 vdd.n4614 vss 0.00324f
C13474 vdd.n4615 vss 0.0112f
C13475 vdd.n4616 vss 0.0128f
C13476 vdd.n4617 vss 0.00413f
C13477 vdd.t151 vss 0.0471f
C13478 vdd.n4618 vss 0.00324f
C13479 vdd.n4620 vss 0.00925f
C13480 vdd.n4621 vss 0.00413f
C13481 vdd.n4622 vss 0.00679f
C13482 vdd.n4623 vss 0.00413f
C13483 vdd.n4624 vss 0.0471f
C13484 vdd.n4625 vss 0.00324f
C13485 vdd.n4626 vss 0.0471f
C13486 vdd.n4627 vss 0.00324f
C13487 vdd.n4628 vss 0.0424f
C13488 vdd.t197 vss 0.0471f
C13489 vdd.n4630 vss 0.00425f
C13490 vdd.n4631 vss 0.00925f
C13491 vdd.n4632 vss 0.0132f
C13492 vdd.n4633 vss 0.00324f
C13493 vdd.n4634 vss 0.0128f
C13494 vdd.n4635 vss 0.02f
C13495 vdd.n4636 vss 0.00425f
C13496 vdd.n4637 vss 0.00413f
C13497 vdd.n4638 vss 0.00251f
C13498 vdd.t149 vss 0.0471f
C13499 vdd.n4639 vss 0.00251f
C13500 vdd.n4640 vss 0.00517f
C13501 vdd.n4641 vss 0.00679f
C13502 vdd.n4642 vss 0.00324f
C13503 vdd.n4643 vss 0.00679f
C13504 vdd.n4644 vss 0.00517f
C13505 vdd.n4645 vss 0.00251f
C13506 vdd.n4646 vss 0.00413f
C13507 vdd.n4647 vss 0.0471f
C13508 vdd.t1178 vss 0.0471f
C13509 vdd.n4648 vss 0.00425f
C13510 vdd.n4649 vss 0.0424f
C13511 vdd.n4650 vss 0.0132f
C13512 vdd.n4651 vss 0.02f
C13513 vdd.n4652 vss 0.00425f
C13514 vdd.n4653 vss 0.00413f
C13515 vdd.n4654 vss 0.00251f
C13516 vdd.n4655 vss 0.0112f
C13517 vdd.n4656 vss 0.0128f
C13518 vdd.n4657 vss 0.0418f
C13519 vdd.n4658 vss 0.118f
C13520 vdd.n4659 vss 0.121f
C13521 vdd.t35 vss 0.0013f
C13522 vdd.t669 vss 0.00134f
C13523 vdd.n4660 vss 0.00324f
C13524 vdd.n4661 vss 0.0112f
C13525 vdd.n4662 vss 0.0128f
C13526 vdd.n4663 vss 0.00413f
C13527 vdd.t667 vss 0.0471f
C13528 vdd.n4664 vss 0.00324f
C13529 vdd.n4666 vss 0.00925f
C13530 vdd.n4667 vss 0.00413f
C13531 vdd.n4668 vss 0.00679f
C13532 vdd.n4669 vss 0.00413f
C13533 vdd.n4670 vss 0.0471f
C13534 vdd.n4671 vss 0.00324f
C13535 vdd.n4672 vss 0.0471f
C13536 vdd.n4673 vss 0.00324f
C13537 vdd.n4674 vss 0.0424f
C13538 vdd.t34 vss 0.0471f
C13539 vdd.n4676 vss 0.00425f
C13540 vdd.n4677 vss 0.00925f
C13541 vdd.n4678 vss 0.0132f
C13542 vdd.n4679 vss 0.00324f
C13543 vdd.n4680 vss 0.0128f
C13544 vdd.n4681 vss 0.02f
C13545 vdd.n4682 vss 0.00425f
C13546 vdd.n4683 vss 0.00413f
C13547 vdd.n4684 vss 0.00251f
C13548 vdd.t668 vss 0.0471f
C13549 vdd.n4685 vss 0.00251f
C13550 vdd.n4686 vss 0.00517f
C13551 vdd.n4687 vss 0.00679f
C13552 vdd.n4688 vss 0.00324f
C13553 vdd.n4689 vss 0.00679f
C13554 vdd.n4690 vss 0.00517f
C13555 vdd.n4691 vss 0.00251f
C13556 vdd.n4692 vss 0.00413f
C13557 vdd.n4693 vss 0.0471f
C13558 vdd.t670 vss 0.0471f
C13559 vdd.n4694 vss 0.00425f
C13560 vdd.n4695 vss 0.0424f
C13561 vdd.n4696 vss 0.0132f
C13562 vdd.n4697 vss 0.02f
C13563 vdd.n4698 vss 0.00425f
C13564 vdd.n4699 vss 0.00413f
C13565 vdd.n4700 vss 0.00251f
C13566 vdd.n4701 vss 0.0112f
C13567 vdd.n4702 vss 0.0707f
C13568 vdd.n4703 vss 0.0393f
C13569 vdd.n4704 vss 0.032f
C13570 vdd.n4705 vss 0.0608f
C13571 vdd.t471 vss 0.00134f
C13572 vdd.t1474 vss 0.0013f
C13573 vdd.n4706 vss 0.032f
C13574 vdd.n4707 vss 0.0393f
C13575 vdd.n4708 vss 0.00324f
C13576 vdd.n4709 vss 0.0112f
C13577 vdd.n4710 vss 0.0128f
C13578 vdd.n4711 vss 0.00413f
C13579 vdd.t472 vss 0.0471f
C13580 vdd.n4712 vss 0.00324f
C13581 vdd.n4714 vss 0.00925f
C13582 vdd.n4715 vss 0.00413f
C13583 vdd.n4716 vss 0.00679f
C13584 vdd.n4717 vss 0.00413f
C13585 vdd.n4718 vss 0.0471f
C13586 vdd.n4719 vss 0.00324f
C13587 vdd.n4720 vss 0.0471f
C13588 vdd.n4721 vss 0.00324f
C13589 vdd.n4722 vss 0.0424f
C13590 vdd.t1473 vss 0.0471f
C13591 vdd.n4724 vss 0.00425f
C13592 vdd.n4725 vss 0.00925f
C13593 vdd.n4726 vss 0.0132f
C13594 vdd.n4727 vss 0.00324f
C13595 vdd.n4728 vss 0.0128f
C13596 vdd.n4729 vss 0.02f
C13597 vdd.n4730 vss 0.00425f
C13598 vdd.n4731 vss 0.00413f
C13599 vdd.n4732 vss 0.00251f
C13600 vdd.t470 vss 0.0471f
C13601 vdd.n4733 vss 0.00251f
C13602 vdd.n4734 vss 0.00517f
C13603 vdd.n4735 vss 0.00679f
C13604 vdd.n4736 vss 0.00324f
C13605 vdd.n4737 vss 0.00679f
C13606 vdd.n4738 vss 0.00517f
C13607 vdd.n4739 vss 0.00251f
C13608 vdd.n4740 vss 0.00413f
C13609 vdd.n4741 vss 0.0471f
C13610 vdd.t1032 vss 0.0471f
C13611 vdd.n4742 vss 0.00425f
C13612 vdd.n4743 vss 0.0424f
C13613 vdd.n4744 vss 0.0132f
C13614 vdd.n4745 vss 0.02f
C13615 vdd.n4746 vss 0.00425f
C13616 vdd.n4747 vss 0.00413f
C13617 vdd.n4748 vss 0.00251f
C13618 vdd.n4749 vss 0.0112f
C13619 vdd.n4750 vss 0.0128f
C13620 vdd.n4751 vss 0.0418f
C13621 vdd.n4752 vss 0.0912f
C13622 vdd.n4753 vss 0.0824f
C13623 vdd.n4754 vss 0.0567f
C13624 vdd.t828 vss 0.0013f
C13625 vdd.t228 vss 0.00134f
C13626 vdd.n4755 vss 0.00324f
C13627 vdd.n4756 vss 0.0112f
C13628 vdd.n4757 vss 0.0128f
C13629 vdd.n4758 vss 0.00413f
C13630 vdd.t229 vss 0.0471f
C13631 vdd.n4759 vss 0.00324f
C13632 vdd.n4761 vss 0.00925f
C13633 vdd.n4762 vss 0.00413f
C13634 vdd.n4763 vss 0.00679f
C13635 vdd.n4764 vss 0.00413f
C13636 vdd.n4765 vss 0.0471f
C13637 vdd.n4766 vss 0.00324f
C13638 vdd.n4767 vss 0.0471f
C13639 vdd.n4768 vss 0.00324f
C13640 vdd.n4769 vss 0.0424f
C13641 vdd.t827 vss 0.0471f
C13642 vdd.n4771 vss 0.00425f
C13643 vdd.n4772 vss 0.00925f
C13644 vdd.n4773 vss 0.0132f
C13645 vdd.n4774 vss 0.00324f
C13646 vdd.n4775 vss 0.0128f
C13647 vdd.n4776 vss 0.02f
C13648 vdd.n4777 vss 0.00425f
C13649 vdd.n4778 vss 0.00413f
C13650 vdd.n4779 vss 0.00251f
C13651 vdd.t227 vss 0.0471f
C13652 vdd.n4780 vss 0.00251f
C13653 vdd.n4781 vss 0.00517f
C13654 vdd.n4782 vss 0.00679f
C13655 vdd.n4783 vss 0.00324f
C13656 vdd.n4784 vss 0.00679f
C13657 vdd.n4785 vss 0.00517f
C13658 vdd.n4786 vss 0.00251f
C13659 vdd.n4787 vss 0.00413f
C13660 vdd.n4788 vss 0.0471f
C13661 vdd.t72 vss 0.0471f
C13662 vdd.n4789 vss 0.00425f
C13663 vdd.n4790 vss 0.0424f
C13664 vdd.n4791 vss 0.0132f
C13665 vdd.n4792 vss 0.02f
C13666 vdd.n4793 vss 0.00425f
C13667 vdd.n4794 vss 0.00413f
C13668 vdd.n4795 vss 0.00251f
C13669 vdd.n4796 vss 0.0112f
C13670 vdd.n4797 vss 0.0128f
C13671 vdd.t366 vss 0.00134f
C13672 vdd.t53 vss 0.0013f
C13673 vdd.n4798 vss 0.032f
C13674 vdd.n4799 vss 0.0393f
C13675 vdd.n4800 vss 0.00324f
C13676 vdd.n4801 vss 0.0112f
C13677 vdd.n4802 vss 0.0128f
C13678 vdd.n4803 vss 0.00413f
C13679 vdd.t367 vss 0.0471f
C13680 vdd.n4804 vss 0.00324f
C13681 vdd.n4806 vss 0.00925f
C13682 vdd.n4807 vss 0.00413f
C13683 vdd.n4808 vss 0.00679f
C13684 vdd.n4809 vss 0.00413f
C13685 vdd.n4810 vss 0.0471f
C13686 vdd.n4811 vss 0.00324f
C13687 vdd.n4812 vss 0.0471f
C13688 vdd.n4813 vss 0.00324f
C13689 vdd.n4814 vss 0.0424f
C13690 vdd.t52 vss 0.0471f
C13691 vdd.n4816 vss 0.00425f
C13692 vdd.n4817 vss 0.00925f
C13693 vdd.n4818 vss 0.0132f
C13694 vdd.n4819 vss 0.00324f
C13695 vdd.n4820 vss 0.0128f
C13696 vdd.n4821 vss 0.02f
C13697 vdd.n4822 vss 0.00425f
C13698 vdd.n4823 vss 0.00413f
C13699 vdd.n4824 vss 0.00251f
C13700 vdd.t365 vss 0.0471f
C13701 vdd.n4825 vss 0.00251f
C13702 vdd.n4826 vss 0.00517f
C13703 vdd.n4827 vss 0.00679f
C13704 vdd.n4828 vss 0.00324f
C13705 vdd.n4829 vss 0.00679f
C13706 vdd.n4830 vss 0.00517f
C13707 vdd.n4831 vss 0.00251f
C13708 vdd.n4832 vss 0.00413f
C13709 vdd.n4833 vss 0.0471f
C13710 vdd.t1256 vss 0.0471f
C13711 vdd.n4834 vss 0.00425f
C13712 vdd.n4835 vss 0.0424f
C13713 vdd.n4836 vss 0.0132f
C13714 vdd.n4837 vss 0.02f
C13715 vdd.n4838 vss 0.00425f
C13716 vdd.n4839 vss 0.00413f
C13717 vdd.n4840 vss 0.00251f
C13718 vdd.n4841 vss 0.0112f
C13719 vdd.n4842 vss 0.0128f
C13720 vdd.n4843 vss 0.0316f
C13721 vdd.t415 vss 0.00134f
C13722 vdd.t1372 vss 0.0013f
C13723 vdd.n4844 vss 0.032f
C13724 vdd.n4845 vss 0.0393f
C13725 vdd.n4846 vss 0.00324f
C13726 vdd.n4847 vss 0.0112f
C13727 vdd.n4848 vss 0.0128f
C13728 vdd.n4849 vss 0.00413f
C13729 vdd.t416 vss 0.0471f
C13730 vdd.n4850 vss 0.00324f
C13731 vdd.n4852 vss 0.00925f
C13732 vdd.n4853 vss 0.00413f
C13733 vdd.n4854 vss 0.00679f
C13734 vdd.n4855 vss 0.00413f
C13735 vdd.n4856 vss 0.0471f
C13736 vdd.n4857 vss 0.00324f
C13737 vdd.n4858 vss 0.0471f
C13738 vdd.n4859 vss 0.00324f
C13739 vdd.n4860 vss 0.0424f
C13740 vdd.t1371 vss 0.0471f
C13741 vdd.n4862 vss 0.00425f
C13742 vdd.n4863 vss 0.00925f
C13743 vdd.n4864 vss 0.0132f
C13744 vdd.n4865 vss 0.00324f
C13745 vdd.n4866 vss 0.0128f
C13746 vdd.n4867 vss 0.02f
C13747 vdd.n4868 vss 0.00425f
C13748 vdd.n4869 vss 0.00413f
C13749 vdd.n4870 vss 0.00251f
C13750 vdd.t414 vss 0.0471f
C13751 vdd.n4871 vss 0.00251f
C13752 vdd.n4872 vss 0.00517f
C13753 vdd.n4873 vss 0.00679f
C13754 vdd.n4874 vss 0.00324f
C13755 vdd.n4875 vss 0.00679f
C13756 vdd.n4876 vss 0.00517f
C13757 vdd.n4877 vss 0.00251f
C13758 vdd.n4878 vss 0.00413f
C13759 vdd.n4879 vss 0.0471f
C13760 vdd.t411 vss 0.0471f
C13761 vdd.n4880 vss 0.00425f
C13762 vdd.n4881 vss 0.0424f
C13763 vdd.n4882 vss 0.0132f
C13764 vdd.n4883 vss 0.02f
C13765 vdd.n4884 vss 0.00425f
C13766 vdd.n4885 vss 0.00413f
C13767 vdd.n4886 vss 0.00251f
C13768 vdd.n4887 vss 0.0112f
C13769 vdd.n4888 vss 0.0128f
C13770 vdd.n4889 vss 0.158f
C13771 vdd.n4890 vss 0.256f
C13772 vdd.n4891 vss 0.0953f
C13773 vdd.n4892 vss 0.0393f
C13774 vdd.n4893 vss 0.032f
C13775 vdd.n4894 vss 0.0608f
C13776 vdd.t1228 vss 0.00134f
C13777 vdd.t1488 vss 0.0013f
C13778 vdd.n4895 vss 0.032f
C13779 vdd.n4896 vss 0.0393f
C13780 vdd.n4897 vss 0.00324f
C13781 vdd.n4898 vss 0.0112f
C13782 vdd.n4899 vss 0.0128f
C13783 vdd.n4900 vss 0.00413f
C13784 vdd.t1229 vss 0.0471f
C13785 vdd.n4901 vss 0.00324f
C13786 vdd.n4903 vss 0.00925f
C13787 vdd.n4904 vss 0.00413f
C13788 vdd.n4905 vss 0.00679f
C13789 vdd.n4906 vss 0.00413f
C13790 vdd.n4907 vss 0.0471f
C13791 vdd.n4908 vss 0.00324f
C13792 vdd.n4909 vss 0.0471f
C13793 vdd.n4910 vss 0.00324f
C13794 vdd.n4911 vss 0.0424f
C13795 vdd.t1487 vss 0.0471f
C13796 vdd.n4913 vss 0.00425f
C13797 vdd.n4914 vss 0.00925f
C13798 vdd.n4915 vss 0.0132f
C13799 vdd.n4916 vss 0.00324f
C13800 vdd.n4917 vss 0.0128f
C13801 vdd.n4918 vss 0.02f
C13802 vdd.n4919 vss 0.00425f
C13803 vdd.n4920 vss 0.00413f
C13804 vdd.n4921 vss 0.00251f
C13805 vdd.t1227 vss 0.0471f
C13806 vdd.n4922 vss 0.00251f
C13807 vdd.n4923 vss 0.00517f
C13808 vdd.n4924 vss 0.00679f
C13809 vdd.n4925 vss 0.00324f
C13810 vdd.n4926 vss 0.00679f
C13811 vdd.n4927 vss 0.00517f
C13812 vdd.n4928 vss 0.00251f
C13813 vdd.n4929 vss 0.00413f
C13814 vdd.n4930 vss 0.0471f
C13815 vdd.t1090 vss 0.0471f
C13816 vdd.n4931 vss 0.00425f
C13817 vdd.n4932 vss 0.0424f
C13818 vdd.n4933 vss 0.0132f
C13819 vdd.n4934 vss 0.02f
C13820 vdd.n4935 vss 0.00425f
C13821 vdd.n4936 vss 0.00413f
C13822 vdd.n4937 vss 0.00251f
C13823 vdd.n4938 vss 0.0112f
C13824 vdd.n4939 vss 0.0128f
C13825 vdd.n4940 vss 0.0418f
C13826 vdd.n4941 vss 0.118f
C13827 vdd.n4942 vss 0.121f
C13828 vdd.t859 vss 0.0013f
C13829 vdd.t511 vss 0.00134f
C13830 vdd.n4943 vss 0.00324f
C13831 vdd.n4944 vss 0.0112f
C13832 vdd.n4945 vss 0.0128f
C13833 vdd.n4946 vss 0.00413f
C13834 vdd.t512 vss 0.0471f
C13835 vdd.n4947 vss 0.00324f
C13836 vdd.n4949 vss 0.00925f
C13837 vdd.n4950 vss 0.00413f
C13838 vdd.n4951 vss 0.00679f
C13839 vdd.n4952 vss 0.00413f
C13840 vdd.n4953 vss 0.0471f
C13841 vdd.n4954 vss 0.00324f
C13842 vdd.n4955 vss 0.0471f
C13843 vdd.n4956 vss 0.00324f
C13844 vdd.n4957 vss 0.0424f
C13845 vdd.t858 vss 0.0471f
C13846 vdd.n4959 vss 0.00425f
C13847 vdd.n4960 vss 0.00925f
C13848 vdd.n4961 vss 0.0132f
C13849 vdd.n4962 vss 0.00324f
C13850 vdd.n4963 vss 0.0128f
C13851 vdd.n4964 vss 0.02f
C13852 vdd.n4965 vss 0.00425f
C13853 vdd.n4966 vss 0.00413f
C13854 vdd.n4967 vss 0.00251f
C13855 vdd.t510 vss 0.0471f
C13856 vdd.n4968 vss 0.00251f
C13857 vdd.n4969 vss 0.00517f
C13858 vdd.n4970 vss 0.00679f
C13859 vdd.n4971 vss 0.00324f
C13860 vdd.n4972 vss 0.00679f
C13861 vdd.n4973 vss 0.00517f
C13862 vdd.n4974 vss 0.00251f
C13863 vdd.n4975 vss 0.00413f
C13864 vdd.n4976 vss 0.0471f
C13865 vdd.t1165 vss 0.0471f
C13866 vdd.n4977 vss 0.00425f
C13867 vdd.n4978 vss 0.0424f
C13868 vdd.n4979 vss 0.0132f
C13869 vdd.n4980 vss 0.02f
C13870 vdd.n4981 vss 0.00425f
C13871 vdd.n4982 vss 0.00413f
C13872 vdd.n4983 vss 0.00251f
C13873 vdd.n4984 vss 0.0112f
C13874 vdd.n4985 vss 0.0707f
C13875 vdd.n4986 vss 0.0393f
C13876 vdd.n4987 vss 0.032f
C13877 vdd.n4988 vss 0.0608f
C13878 vdd.t1100 vss 0.00134f
C13879 vdd.t1301 vss 0.0013f
C13880 vdd.n4989 vss 0.032f
C13881 vdd.n4990 vss 0.0393f
C13882 vdd.n4991 vss 0.00324f
C13883 vdd.n4992 vss 0.0112f
C13884 vdd.n4993 vss 0.0128f
C13885 vdd.n4994 vss 0.00413f
C13886 vdd.t1101 vss 0.0471f
C13887 vdd.n4995 vss 0.00324f
C13888 vdd.n4997 vss 0.00925f
C13889 vdd.n4998 vss 0.00413f
C13890 vdd.n4999 vss 0.00679f
C13891 vdd.n5000 vss 0.00413f
C13892 vdd.n5001 vss 0.0471f
C13893 vdd.n5002 vss 0.00324f
C13894 vdd.n5003 vss 0.0471f
C13895 vdd.n5004 vss 0.00324f
C13896 vdd.n5005 vss 0.0424f
C13897 vdd.t1300 vss 0.0471f
C13898 vdd.n5007 vss 0.00425f
C13899 vdd.n5008 vss 0.00925f
C13900 vdd.n5009 vss 0.0132f
C13901 vdd.n5010 vss 0.00324f
C13902 vdd.n5011 vss 0.0128f
C13903 vdd.n5012 vss 0.02f
C13904 vdd.n5013 vss 0.00425f
C13905 vdd.n5014 vss 0.00413f
C13906 vdd.n5015 vss 0.00251f
C13907 vdd.t1099 vss 0.0471f
C13908 vdd.n5016 vss 0.00251f
C13909 vdd.n5017 vss 0.00517f
C13910 vdd.n5018 vss 0.00679f
C13911 vdd.n5019 vss 0.00324f
C13912 vdd.n5020 vss 0.00679f
C13913 vdd.n5021 vss 0.00517f
C13914 vdd.n5022 vss 0.00251f
C13915 vdd.n5023 vss 0.00413f
C13916 vdd.n5024 vss 0.0471f
C13917 vdd.t308 vss 0.0471f
C13918 vdd.n5025 vss 0.00425f
C13919 vdd.n5026 vss 0.0424f
C13920 vdd.n5027 vss 0.0132f
C13921 vdd.n5028 vss 0.02f
C13922 vdd.n5029 vss 0.00425f
C13923 vdd.n5030 vss 0.00413f
C13924 vdd.n5031 vss 0.00251f
C13925 vdd.n5032 vss 0.0112f
C13926 vdd.n5033 vss 0.0128f
C13927 vdd.n5034 vss 0.0418f
C13928 vdd.n5035 vss 0.118f
C13929 vdd.n5036 vss 0.0935f
C13930 vdd.t1011 vss 0.0013f
C13931 vdd.t1168 vss 0.00134f
C13932 vdd.n5037 vss 0.00324f
C13933 vdd.n5038 vss 0.0112f
C13934 vdd.n5039 vss 0.0128f
C13935 vdd.n5040 vss 0.00413f
C13936 vdd.t1166 vss 0.0471f
C13937 vdd.n5041 vss 0.00324f
C13938 vdd.n5043 vss 0.00925f
C13939 vdd.n5044 vss 0.00413f
C13940 vdd.n5045 vss 0.00679f
C13941 vdd.n5046 vss 0.00413f
C13942 vdd.n5047 vss 0.0471f
C13943 vdd.n5048 vss 0.00324f
C13944 vdd.n5049 vss 0.0471f
C13945 vdd.n5050 vss 0.00324f
C13946 vdd.n5051 vss 0.0424f
C13947 vdd.t1010 vss 0.0471f
C13948 vdd.n5053 vss 0.00425f
C13949 vdd.n5054 vss 0.00925f
C13950 vdd.n5055 vss 0.0132f
C13951 vdd.n5056 vss 0.00324f
C13952 vdd.n5057 vss 0.0128f
C13953 vdd.n5058 vss 0.02f
C13954 vdd.n5059 vss 0.00425f
C13955 vdd.n5060 vss 0.00413f
C13956 vdd.n5061 vss 0.00251f
C13957 vdd.t1167 vss 0.0471f
C13958 vdd.n5062 vss 0.00251f
C13959 vdd.n5063 vss 0.00517f
C13960 vdd.n5064 vss 0.00679f
C13961 vdd.n5065 vss 0.00324f
C13962 vdd.n5066 vss 0.00679f
C13963 vdd.n5067 vss 0.00517f
C13964 vdd.n5068 vss 0.00251f
C13965 vdd.n5069 vss 0.00413f
C13966 vdd.n5070 vss 0.0471f
C13967 vdd.t1412 vss 0.0471f
C13968 vdd.n5071 vss 0.00425f
C13969 vdd.n5072 vss 0.0424f
C13970 vdd.n5073 vss 0.0132f
C13971 vdd.n5074 vss 0.02f
C13972 vdd.n5075 vss 0.00425f
C13973 vdd.n5076 vss 0.00413f
C13974 vdd.n5077 vss 0.00251f
C13975 vdd.n5078 vss 0.0112f
C13976 vdd.n5079 vss 0.0128f
C13977 vdd.t108 vss 0.00134f
C13978 vdd.t51 vss 0.0013f
C13979 vdd.n5080 vss 0.032f
C13980 vdd.n5081 vss 0.0393f
C13981 vdd.n5082 vss 0.00324f
C13982 vdd.n5083 vss 0.0112f
C13983 vdd.n5084 vss 0.0128f
C13984 vdd.n5085 vss 0.00413f
C13985 vdd.t109 vss 0.0471f
C13986 vdd.n5086 vss 0.00324f
C13987 vdd.n5088 vss 0.00925f
C13988 vdd.n5089 vss 0.00413f
C13989 vdd.n5090 vss 0.00679f
C13990 vdd.n5091 vss 0.00413f
C13991 vdd.n5092 vss 0.0471f
C13992 vdd.n5093 vss 0.00324f
C13993 vdd.n5094 vss 0.0471f
C13994 vdd.n5095 vss 0.00324f
C13995 vdd.n5096 vss 0.0424f
C13996 vdd.t50 vss 0.0471f
C13997 vdd.n5098 vss 0.00425f
C13998 vdd.n5099 vss 0.00925f
C13999 vdd.n5100 vss 0.0132f
C14000 vdd.n5101 vss 0.00324f
C14001 vdd.n5102 vss 0.0128f
C14002 vdd.n5103 vss 0.02f
C14003 vdd.n5104 vss 0.00425f
C14004 vdd.n5105 vss 0.00413f
C14005 vdd.n5106 vss 0.00251f
C14006 vdd.t107 vss 0.0471f
C14007 vdd.n5107 vss 0.00251f
C14008 vdd.n5108 vss 0.00517f
C14009 vdd.n5109 vss 0.00679f
C14010 vdd.n5110 vss 0.00324f
C14011 vdd.n5111 vss 0.00679f
C14012 vdd.n5112 vss 0.00517f
C14013 vdd.n5113 vss 0.00251f
C14014 vdd.n5114 vss 0.00413f
C14015 vdd.n5115 vss 0.0471f
C14016 vdd.t607 vss 0.0471f
C14017 vdd.n5116 vss 0.00425f
C14018 vdd.n5117 vss 0.0424f
C14019 vdd.n5118 vss 0.0132f
C14020 vdd.n5119 vss 0.02f
C14021 vdd.n5120 vss 0.00425f
C14022 vdd.n5121 vss 0.00413f
C14023 vdd.n5122 vss 0.00251f
C14024 vdd.n5123 vss 0.0112f
C14025 vdd.n5124 vss 0.0128f
C14026 vdd.n5125 vss 0.119f
C14027 vdd.n5126 vss 0.118f
C14028 vdd.n5127 vss 0.0393f
C14029 vdd.n5128 vss 0.032f
C14030 vdd.n5129 vss 0.0608f
C14031 vdd.t345 vss 0.00134f
C14032 vdd.t1044 vss 0.0013f
C14033 vdd.n5130 vss 0.032f
C14034 vdd.n5131 vss 0.0393f
C14035 vdd.n5132 vss 0.00324f
C14036 vdd.n5133 vss 0.0112f
C14037 vdd.n5134 vss 0.0128f
C14038 vdd.n5135 vss 0.00413f
C14039 vdd.t346 vss 0.0471f
C14040 vdd.n5136 vss 0.00324f
C14041 vdd.n5138 vss 0.00925f
C14042 vdd.n5139 vss 0.00413f
C14043 vdd.n5140 vss 0.00679f
C14044 vdd.n5141 vss 0.00413f
C14045 vdd.n5142 vss 0.0471f
C14046 vdd.n5143 vss 0.00324f
C14047 vdd.n5144 vss 0.0471f
C14048 vdd.n5145 vss 0.00324f
C14049 vdd.n5146 vss 0.0424f
C14050 vdd.t1043 vss 0.0471f
C14051 vdd.n5148 vss 0.00425f
C14052 vdd.n5149 vss 0.00925f
C14053 vdd.n5150 vss 0.0132f
C14054 vdd.n5151 vss 0.00324f
C14055 vdd.n5152 vss 0.0128f
C14056 vdd.n5153 vss 0.02f
C14057 vdd.n5154 vss 0.00425f
C14058 vdd.n5155 vss 0.00413f
C14059 vdd.n5156 vss 0.00251f
C14060 vdd.t344 vss 0.0471f
C14061 vdd.n5157 vss 0.00251f
C14062 vdd.n5158 vss 0.00517f
C14063 vdd.n5159 vss 0.00679f
C14064 vdd.n5160 vss 0.00324f
C14065 vdd.n5161 vss 0.00679f
C14066 vdd.n5162 vss 0.00517f
C14067 vdd.n5163 vss 0.00251f
C14068 vdd.n5164 vss 0.00413f
C14069 vdd.n5165 vss 0.0471f
C14070 vdd.t191 vss 0.0471f
C14071 vdd.n5166 vss 0.00425f
C14072 vdd.n5167 vss 0.0424f
C14073 vdd.n5168 vss 0.0132f
C14074 vdd.n5169 vss 0.02f
C14075 vdd.n5170 vss 0.00425f
C14076 vdd.n5171 vss 0.00413f
C14077 vdd.n5172 vss 0.00251f
C14078 vdd.n5173 vss 0.0112f
C14079 vdd.n5174 vss 0.0128f
C14080 vdd.n5175 vss 0.0418f
C14081 vdd.n5176 vss 0.118f
C14082 vdd.n5177 vss 0.121f
C14083 vdd.t943 vss 0.0013f
C14084 vdd.t323 vss 0.00134f
C14085 vdd.n5178 vss 0.00324f
C14086 vdd.n5179 vss 0.0112f
C14087 vdd.n5180 vss 0.0128f
C14088 vdd.n5181 vss 0.00413f
C14089 vdd.t321 vss 0.0471f
C14090 vdd.n5182 vss 0.00324f
C14091 vdd.n5184 vss 0.00925f
C14092 vdd.n5185 vss 0.00413f
C14093 vdd.n5186 vss 0.00679f
C14094 vdd.n5187 vss 0.00413f
C14095 vdd.n5188 vss 0.0471f
C14096 vdd.n5189 vss 0.00324f
C14097 vdd.n5190 vss 0.0471f
C14098 vdd.n5191 vss 0.00324f
C14099 vdd.n5192 vss 0.0424f
C14100 vdd.t942 vss 0.0471f
C14101 vdd.n5194 vss 0.00425f
C14102 vdd.n5195 vss 0.00925f
C14103 vdd.n5196 vss 0.0132f
C14104 vdd.n5197 vss 0.00324f
C14105 vdd.n5198 vss 0.0128f
C14106 vdd.n5199 vss 0.02f
C14107 vdd.n5200 vss 0.00425f
C14108 vdd.n5201 vss 0.00413f
C14109 vdd.n5202 vss 0.00251f
C14110 vdd.t322 vss 0.0471f
C14111 vdd.n5203 vss 0.00251f
C14112 vdd.n5204 vss 0.00517f
C14113 vdd.n5205 vss 0.00679f
C14114 vdd.n5206 vss 0.00324f
C14115 vdd.n5207 vss 0.00679f
C14116 vdd.n5208 vss 0.00517f
C14117 vdd.n5209 vss 0.00251f
C14118 vdd.n5210 vss 0.00413f
C14119 vdd.n5211 vss 0.0471f
C14120 vdd.t1278 vss 0.0471f
C14121 vdd.n5212 vss 0.00425f
C14122 vdd.n5213 vss 0.0424f
C14123 vdd.n5214 vss 0.0132f
C14124 vdd.n5215 vss 0.02f
C14125 vdd.n5216 vss 0.00425f
C14126 vdd.n5217 vss 0.00413f
C14127 vdd.n5218 vss 0.00251f
C14128 vdd.n5219 vss 0.0112f
C14129 vdd.n5220 vss 0.0707f
C14130 vdd.n5221 vss 0.0393f
C14131 vdd.n5222 vss 0.032f
C14132 vdd.n5223 vss 0.0608f
C14133 vdd.t701 vss 0.00134f
C14134 vdd.t1305 vss 0.0013f
C14135 vdd.n5224 vss 0.032f
C14136 vdd.n5225 vss 0.0393f
C14137 vdd.n5226 vss 0.00324f
C14138 vdd.n5227 vss 0.0112f
C14139 vdd.n5228 vss 0.0128f
C14140 vdd.n5229 vss 0.00413f
C14141 vdd.t699 vss 0.0471f
C14142 vdd.n5230 vss 0.00324f
C14143 vdd.n5232 vss 0.00925f
C14144 vdd.n5233 vss 0.00413f
C14145 vdd.n5234 vss 0.00679f
C14146 vdd.n5235 vss 0.00413f
C14147 vdd.n5236 vss 0.0471f
C14148 vdd.n5237 vss 0.00324f
C14149 vdd.n5238 vss 0.0471f
C14150 vdd.n5239 vss 0.00324f
C14151 vdd.n5240 vss 0.0424f
C14152 vdd.t1304 vss 0.0471f
C14153 vdd.n5242 vss 0.00425f
C14154 vdd.n5243 vss 0.00925f
C14155 vdd.n5244 vss 0.0132f
C14156 vdd.n5245 vss 0.00324f
C14157 vdd.n5246 vss 0.0128f
C14158 vdd.n5247 vss 0.02f
C14159 vdd.n5248 vss 0.00425f
C14160 vdd.n5249 vss 0.00413f
C14161 vdd.n5250 vss 0.00251f
C14162 vdd.t700 vss 0.0471f
C14163 vdd.n5251 vss 0.00251f
C14164 vdd.n5252 vss 0.00517f
C14165 vdd.n5253 vss 0.00679f
C14166 vdd.n5254 vss 0.00324f
C14167 vdd.n5255 vss 0.00679f
C14168 vdd.n5256 vss 0.00517f
C14169 vdd.n5257 vss 0.00251f
C14170 vdd.n5258 vss 0.00413f
C14171 vdd.n5259 vss 0.0471f
C14172 vdd.t537 vss 0.0471f
C14173 vdd.n5260 vss 0.00425f
C14174 vdd.n5261 vss 0.0424f
C14175 vdd.n5262 vss 0.0132f
C14176 vdd.n5263 vss 0.02f
C14177 vdd.n5264 vss 0.00425f
C14178 vdd.n5265 vss 0.00413f
C14179 vdd.n5266 vss 0.00251f
C14180 vdd.n5267 vss 0.0112f
C14181 vdd.n5268 vss 0.0128f
C14182 vdd.n5269 vss 0.0418f
C14183 vdd.n5270 vss 0.0912f
C14184 vdd.n5271 vss 0.0824f
C14185 vdd.n5272 vss 0.0567f
C14186 vdd.t845 vss 0.0013f
C14187 vdd.t1110 vss 0.00134f
C14188 vdd.n5273 vss 0.00324f
C14189 vdd.n5274 vss 0.0112f
C14190 vdd.n5275 vss 0.0128f
C14191 vdd.n5276 vss 0.00413f
C14192 vdd.t1111 vss 0.0471f
C14193 vdd.n5277 vss 0.00324f
C14194 vdd.n5279 vss 0.00925f
C14195 vdd.n5280 vss 0.00413f
C14196 vdd.n5281 vss 0.00679f
C14197 vdd.n5282 vss 0.00413f
C14198 vdd.n5283 vss 0.0471f
C14199 vdd.n5284 vss 0.00324f
C14200 vdd.n5285 vss 0.0471f
C14201 vdd.n5286 vss 0.00324f
C14202 vdd.n5287 vss 0.0424f
C14203 vdd.t844 vss 0.0471f
C14204 vdd.n5289 vss 0.00425f
C14205 vdd.n5290 vss 0.00925f
C14206 vdd.n5291 vss 0.0132f
C14207 vdd.n5292 vss 0.00324f
C14208 vdd.n5293 vss 0.0128f
C14209 vdd.n5294 vss 0.02f
C14210 vdd.n5295 vss 0.00425f
C14211 vdd.n5296 vss 0.00413f
C14212 vdd.n5297 vss 0.00251f
C14213 vdd.t1109 vss 0.0471f
C14214 vdd.n5298 vss 0.00251f
C14215 vdd.n5299 vss 0.00517f
C14216 vdd.n5300 vss 0.00679f
C14217 vdd.n5301 vss 0.00324f
C14218 vdd.n5302 vss 0.00679f
C14219 vdd.n5303 vss 0.00517f
C14220 vdd.n5304 vss 0.00251f
C14221 vdd.n5305 vss 0.00413f
C14222 vdd.n5306 vss 0.0471f
C14223 vdd.t888 vss 0.0471f
C14224 vdd.n5307 vss 0.00425f
C14225 vdd.n5308 vss 0.0424f
C14226 vdd.n5309 vss 0.0132f
C14227 vdd.n5310 vss 0.02f
C14228 vdd.n5311 vss 0.00425f
C14229 vdd.n5312 vss 0.00413f
C14230 vdd.n5313 vss 0.00251f
C14231 vdd.n5314 vss 0.0112f
C14232 vdd.n5315 vss 0.0128f
C14233 vdd.t1504 vss 0.00134f
C14234 vdd.t173 vss 0.0013f
C14235 vdd.n5316 vss 0.032f
C14236 vdd.n5317 vss 0.0393f
C14237 vdd.n5318 vss 0.00324f
C14238 vdd.n5319 vss 0.0112f
C14239 vdd.n5320 vss 0.0128f
C14240 vdd.n5321 vss 0.00413f
C14241 vdd.t1505 vss 0.0471f
C14242 vdd.n5322 vss 0.00324f
C14243 vdd.n5324 vss 0.00925f
C14244 vdd.n5325 vss 0.00413f
C14245 vdd.n5326 vss 0.00679f
C14246 vdd.n5327 vss 0.00413f
C14247 vdd.n5328 vss 0.0471f
C14248 vdd.n5329 vss 0.00324f
C14249 vdd.n5330 vss 0.0471f
C14250 vdd.n5331 vss 0.00324f
C14251 vdd.n5332 vss 0.0424f
C14252 vdd.t172 vss 0.0471f
C14253 vdd.n5334 vss 0.00425f
C14254 vdd.n5335 vss 0.00925f
C14255 vdd.n5336 vss 0.0132f
C14256 vdd.n5337 vss 0.00324f
C14257 vdd.n5338 vss 0.0128f
C14258 vdd.n5339 vss 0.02f
C14259 vdd.n5340 vss 0.00425f
C14260 vdd.n5341 vss 0.00413f
C14261 vdd.n5342 vss 0.00251f
C14262 vdd.t1503 vss 0.0471f
C14263 vdd.n5343 vss 0.00251f
C14264 vdd.n5344 vss 0.00517f
C14265 vdd.n5345 vss 0.00679f
C14266 vdd.n5346 vss 0.00324f
C14267 vdd.n5347 vss 0.00679f
C14268 vdd.n5348 vss 0.00517f
C14269 vdd.n5349 vss 0.00251f
C14270 vdd.n5350 vss 0.00413f
C14271 vdd.n5351 vss 0.0471f
C14272 vdd.t660 vss 0.0471f
C14273 vdd.n5352 vss 0.00425f
C14274 vdd.n5353 vss 0.0424f
C14275 vdd.n5354 vss 0.0132f
C14276 vdd.n5355 vss 0.02f
C14277 vdd.n5356 vss 0.00425f
C14278 vdd.n5357 vss 0.00413f
C14279 vdd.n5358 vss 0.00251f
C14280 vdd.n5359 vss 0.0112f
C14281 vdd.n5360 vss 0.0128f
C14282 vdd.n5361 vss 0.119f
C14283 vdd.n5362 vss 0.118f
C14284 vdd.n5363 vss 0.0393f
C14285 vdd.n5364 vss 0.032f
C14286 vdd.n5365 vss 0.0608f
C14287 vdd.t720 vss 0.00134f
C14288 vdd.t457 vss 0.0013f
C14289 vdd.n5366 vss 0.032f
C14290 vdd.n5367 vss 0.0393f
C14291 vdd.n5368 vss 0.00324f
C14292 vdd.n5369 vss 0.0112f
C14293 vdd.n5370 vss 0.0128f
C14294 vdd.n5371 vss 0.00413f
C14295 vdd.t718 vss 0.0471f
C14296 vdd.n5372 vss 0.00324f
C14297 vdd.n5374 vss 0.00925f
C14298 vdd.n5375 vss 0.00413f
C14299 vdd.n5376 vss 0.00679f
C14300 vdd.n5377 vss 0.00413f
C14301 vdd.n5378 vss 0.0471f
C14302 vdd.n5379 vss 0.00324f
C14303 vdd.n5380 vss 0.0471f
C14304 vdd.n5381 vss 0.00324f
C14305 vdd.n5382 vss 0.0424f
C14306 vdd.t456 vss 0.0471f
C14307 vdd.n5384 vss 0.00425f
C14308 vdd.n5385 vss 0.00925f
C14309 vdd.n5386 vss 0.0132f
C14310 vdd.n5387 vss 0.00324f
C14311 vdd.n5388 vss 0.0128f
C14312 vdd.n5389 vss 0.02f
C14313 vdd.n5390 vss 0.00425f
C14314 vdd.n5391 vss 0.00413f
C14315 vdd.n5392 vss 0.00251f
C14316 vdd.t719 vss 0.0471f
C14317 vdd.n5393 vss 0.00251f
C14318 vdd.n5394 vss 0.00517f
C14319 vdd.n5395 vss 0.00679f
C14320 vdd.n5396 vss 0.00324f
C14321 vdd.n5397 vss 0.00679f
C14322 vdd.n5398 vss 0.00517f
C14323 vdd.n5399 vss 0.00251f
C14324 vdd.n5400 vss 0.00413f
C14325 vdd.n5401 vss 0.0471f
C14326 vdd.t63 vss 0.0471f
C14327 vdd.n5402 vss 0.00425f
C14328 vdd.n5403 vss 0.0424f
C14329 vdd.n5404 vss 0.0132f
C14330 vdd.n5405 vss 0.02f
C14331 vdd.n5406 vss 0.00425f
C14332 vdd.n5407 vss 0.00413f
C14333 vdd.n5408 vss 0.00251f
C14334 vdd.n5409 vss 0.0112f
C14335 vdd.n5410 vss 0.0128f
C14336 vdd.n5411 vss 0.0418f
C14337 vdd.n5412 vss 0.118f
C14338 vdd.n5413 vss 0.121f
C14339 vdd.t1013 vss 0.0013f
C14340 vdd.t501 vss 0.00134f
C14341 vdd.n5414 vss 0.00324f
C14342 vdd.n5415 vss 0.0112f
C14343 vdd.n5416 vss 0.0128f
C14344 vdd.n5417 vss 0.00413f
C14345 vdd.t499 vss 0.0471f
C14346 vdd.n5418 vss 0.00324f
C14347 vdd.n5420 vss 0.00925f
C14348 vdd.n5421 vss 0.00413f
C14349 vdd.n5422 vss 0.00679f
C14350 vdd.n5423 vss 0.00413f
C14351 vdd.n5424 vss 0.0471f
C14352 vdd.n5425 vss 0.00324f
C14353 vdd.n5426 vss 0.0471f
C14354 vdd.n5427 vss 0.00324f
C14355 vdd.n5428 vss 0.0424f
C14356 vdd.t1012 vss 0.0471f
C14357 vdd.n5430 vss 0.00425f
C14358 vdd.n5431 vss 0.00925f
C14359 vdd.n5432 vss 0.0132f
C14360 vdd.n5433 vss 0.00324f
C14361 vdd.n5434 vss 0.0128f
C14362 vdd.n5435 vss 0.02f
C14363 vdd.n5436 vss 0.00425f
C14364 vdd.n5437 vss 0.00413f
C14365 vdd.n5438 vss 0.00251f
C14366 vdd.t500 vss 0.0471f
C14367 vdd.n5439 vss 0.00251f
C14368 vdd.n5440 vss 0.00517f
C14369 vdd.n5441 vss 0.00679f
C14370 vdd.n5442 vss 0.00324f
C14371 vdd.n5443 vss 0.00679f
C14372 vdd.n5444 vss 0.00517f
C14373 vdd.n5445 vss 0.00251f
C14374 vdd.n5446 vss 0.00413f
C14375 vdd.n5447 vss 0.0471f
C14376 vdd.t1411 vss 0.0471f
C14377 vdd.n5448 vss 0.00425f
C14378 vdd.n5449 vss 0.0424f
C14379 vdd.n5450 vss 0.0132f
C14380 vdd.n5451 vss 0.02f
C14381 vdd.n5452 vss 0.00425f
C14382 vdd.n5453 vss 0.00413f
C14383 vdd.n5454 vss 0.00251f
C14384 vdd.n5455 vss 0.0112f
C14385 vdd.n5456 vss 0.0707f
C14386 vdd.n5457 vss 0.0393f
C14387 vdd.n5458 vss 0.032f
C14388 vdd.n5459 vss 0.0608f
C14389 vdd.t505 vss 0.00134f
C14390 vdd.t1052 vss 0.0013f
C14391 vdd.n5460 vss 0.032f
C14392 vdd.n5461 vss 0.0393f
C14393 vdd.n5462 vss 0.00324f
C14394 vdd.n5463 vss 0.0112f
C14395 vdd.n5464 vss 0.0128f
C14396 vdd.n5465 vss 0.00413f
C14397 vdd.t506 vss 0.0471f
C14398 vdd.n5466 vss 0.00324f
C14399 vdd.n5468 vss 0.00925f
C14400 vdd.n5469 vss 0.00413f
C14401 vdd.n5470 vss 0.00679f
C14402 vdd.n5471 vss 0.00413f
C14403 vdd.n5472 vss 0.0471f
C14404 vdd.n5473 vss 0.00324f
C14405 vdd.n5474 vss 0.0471f
C14406 vdd.n5475 vss 0.00324f
C14407 vdd.n5476 vss 0.0424f
C14408 vdd.t1051 vss 0.0471f
C14409 vdd.n5478 vss 0.00425f
C14410 vdd.n5479 vss 0.00925f
C14411 vdd.n5480 vss 0.0132f
C14412 vdd.n5481 vss 0.00324f
C14413 vdd.n5482 vss 0.0128f
C14414 vdd.n5483 vss 0.02f
C14415 vdd.n5484 vss 0.00425f
C14416 vdd.n5485 vss 0.00413f
C14417 vdd.n5486 vss 0.00251f
C14418 vdd.t504 vss 0.0471f
C14419 vdd.n5487 vss 0.00251f
C14420 vdd.n5488 vss 0.00517f
C14421 vdd.n5489 vss 0.00679f
C14422 vdd.n5490 vss 0.00324f
C14423 vdd.n5491 vss 0.00679f
C14424 vdd.n5492 vss 0.00517f
C14425 vdd.n5493 vss 0.00251f
C14426 vdd.n5494 vss 0.00413f
C14427 vdd.n5495 vss 0.0471f
C14428 vdd.t269 vss 0.0471f
C14429 vdd.n5496 vss 0.00425f
C14430 vdd.n5497 vss 0.0424f
C14431 vdd.n5498 vss 0.0132f
C14432 vdd.n5499 vss 0.02f
C14433 vdd.n5500 vss 0.00425f
C14434 vdd.n5501 vss 0.00413f
C14435 vdd.n5502 vss 0.00251f
C14436 vdd.n5503 vss 0.0112f
C14437 vdd.n5504 vss 0.0128f
C14438 vdd.n5505 vss 0.0418f
C14439 vdd.n5506 vss 0.299f
C14440 vdd.n5507 vss 0.00324f
C14441 vdd.n5508 vss 0.0112f
C14442 vdd.n5509 vss 0.0128f
C14443 vdd.n5510 vss 0.00413f
C14444 vdd.n5511 vss 0.00413f
C14445 vdd.n5512 vss 0.0471f
C14446 vdd.n5513 vss 0.00251f
C14447 vdd.t556 vss 0.0471f
C14448 vdd.n5514 vss 0.00324f
C14449 vdd.n5516 vss 0.00679f
C14450 vdd.n5517 vss 0.00413f
C14451 vdd.n5518 vss 0.00324f
C14452 vdd.n5519 vss 0.00413f
C14453 vdd.n5520 vss 0.0471f
C14454 vdd.n5521 vss 0.00324f
C14455 vdd.n5523 vss 0.00925f
C14456 vdd.t327 vss 0.0471f
C14457 vdd.n5524 vss 0.00425f
C14458 vdd.n5525 vss 0.0424f
C14459 vdd.n5526 vss 0.0132f
C14460 vdd.n5527 vss 0.00324f
C14461 vdd.n5528 vss 0.0128f
C14462 vdd.n5529 vss 0.02f
C14463 vdd.n5530 vss 0.00425f
C14464 vdd.n5531 vss 0.00413f
C14465 vdd.n5532 vss 0.00251f
C14466 vdd.t759 vss 0.0471f
C14467 vdd.n5533 vss 0.00251f
C14468 vdd.n5534 vss 0.00517f
C14469 vdd.n5535 vss 0.00679f
C14470 vdd.n5536 vss 0.00517f
C14471 vdd.n5537 vss 0.00679f
C14472 vdd.n5538 vss 0.02f
C14473 vdd.n5539 vss 0.00425f
C14474 vdd.n5540 vss 0.0424f
C14475 vdd.n5541 vss 0.0132f
C14476 vdd.n5542 vss 0.00925f
C14477 vdd.n5543 vss 0.00425f
C14478 vdd.n5544 vss 0.00413f
C14479 vdd.n5545 vss 0.00324f
C14480 vdd.n5546 vss 0.0471f
C14481 vdd.t760 vss 0.0471f
C14482 vdd.n5547 vss 0.00251f
C14483 vdd.n5548 vss 0.0112f
C14484 vdd.n5549 vss 0.0128f
C14485 vdd.t761 vss 0.00134f
C14486 vdd.t557 vss 0.0013f
C14487 vdd.n5550 vss 0.0332f
C14488 vdd.n5551 vss 0.0393f
C14489 vdd.n5552 vss 0.0345f
C14490 vdd.n5553 vss 0.262f
C14491 vdd.t907 vss 0.0013f
C14492 vdd.t715 vss 0.00134f
C14493 vdd.n5554 vss 0.00324f
C14494 vdd.n5555 vss 0.0112f
C14495 vdd.n5556 vss 0.0128f
C14496 vdd.n5557 vss 0.00413f
C14497 vdd.n5558 vss 0.00413f
C14498 vdd.n5559 vss 0.0471f
C14499 vdd.n5560 vss 0.00251f
C14500 vdd.t164 vss 0.0471f
C14501 vdd.n5561 vss 0.00324f
C14502 vdd.n5563 vss 0.00679f
C14503 vdd.n5564 vss 0.00413f
C14504 vdd.n5565 vss 0.00324f
C14505 vdd.n5566 vss 0.00413f
C14506 vdd.n5567 vss 0.0471f
C14507 vdd.n5568 vss 0.00324f
C14508 vdd.n5570 vss 0.00925f
C14509 vdd.t1237 vss 0.0471f
C14510 vdd.n5571 vss 0.00425f
C14511 vdd.n5572 vss 0.0424f
C14512 vdd.n5573 vss 0.0132f
C14513 vdd.n5574 vss 0.00324f
C14514 vdd.n5575 vss 0.0128f
C14515 vdd.n5576 vss 0.02f
C14516 vdd.n5577 vss 0.00425f
C14517 vdd.n5578 vss 0.00413f
C14518 vdd.n5579 vss 0.00251f
C14519 vdd.t185 vss 0.0471f
C14520 vdd.n5580 vss 0.00251f
C14521 vdd.n5581 vss 0.00517f
C14522 vdd.n5582 vss 0.00679f
C14523 vdd.n5583 vss 0.00517f
C14524 vdd.n5584 vss 0.00679f
C14525 vdd.n5585 vss 0.02f
C14526 vdd.n5586 vss 0.00425f
C14527 vdd.n5587 vss 0.0424f
C14528 vdd.n5588 vss 0.0132f
C14529 vdd.n5589 vss 0.00925f
C14530 vdd.n5590 vss 0.00425f
C14531 vdd.n5591 vss 0.00413f
C14532 vdd.n5592 vss 0.00324f
C14533 vdd.n5593 vss 0.0471f
C14534 vdd.t186 vss 0.0471f
C14535 vdd.n5594 vss 0.00251f
C14536 vdd.n5595 vss 0.0112f
C14537 vdd.n5596 vss 0.0128f
C14538 vdd.t187 vss 0.00134f
C14539 vdd.t165 vss 0.0013f
C14540 vdd.n5597 vss 0.0332f
C14541 vdd.n5598 vss 0.0393f
C14542 vdd.n5599 vss 0.119f
C14543 vdd.n5600 vss 0.00324f
C14544 vdd.n5601 vss 0.0112f
C14545 vdd.n5602 vss 0.0128f
C14546 vdd.n5603 vss 0.00413f
C14547 vdd.n5604 vss 0.00413f
C14548 vdd.n5605 vss 0.0471f
C14549 vdd.n5606 vss 0.00251f
C14550 vdd.t906 vss 0.0471f
C14551 vdd.n5607 vss 0.00324f
C14552 vdd.n5609 vss 0.00679f
C14553 vdd.n5610 vss 0.00413f
C14554 vdd.n5611 vss 0.00324f
C14555 vdd.n5612 vss 0.00413f
C14556 vdd.n5613 vss 0.0471f
C14557 vdd.n5614 vss 0.00324f
C14558 vdd.n5616 vss 0.00925f
C14559 vdd.t716 vss 0.0471f
C14560 vdd.n5617 vss 0.00425f
C14561 vdd.n5618 vss 0.0424f
C14562 vdd.n5619 vss 0.0132f
C14563 vdd.n5620 vss 0.00324f
C14564 vdd.n5621 vss 0.0128f
C14565 vdd.n5622 vss 0.02f
C14566 vdd.n5623 vss 0.00425f
C14567 vdd.n5624 vss 0.00413f
C14568 vdd.n5625 vss 0.00251f
C14569 vdd.t713 vss 0.0471f
C14570 vdd.n5626 vss 0.00251f
C14571 vdd.n5627 vss 0.00517f
C14572 vdd.n5628 vss 0.00679f
C14573 vdd.n5629 vss 0.00517f
C14574 vdd.n5630 vss 0.00679f
C14575 vdd.n5631 vss 0.02f
C14576 vdd.n5632 vss 0.00425f
C14577 vdd.n5633 vss 0.0424f
C14578 vdd.n5634 vss 0.0132f
C14579 vdd.n5635 vss 0.00925f
C14580 vdd.n5636 vss 0.00425f
C14581 vdd.n5637 vss 0.00413f
C14582 vdd.n5638 vss 0.00324f
C14583 vdd.n5639 vss 0.0471f
C14584 vdd.t714 vss 0.0471f
C14585 vdd.n5640 vss 0.00251f
C14586 vdd.n5641 vss 0.0112f
C14587 vdd.n5642 vss 0.0128f
C14588 vdd.n5643 vss 0.118f
C14589 vdd.n5644 vss 0.0393f
C14590 vdd.n5645 vss 0.0332f
C14591 vdd.n5646 vss 0.0596f
C14592 vdd.n5647 vss 0.00324f
C14593 vdd.n5648 vss 0.0112f
C14594 vdd.n5649 vss 0.0128f
C14595 vdd.n5650 vss 0.00413f
C14596 vdd.n5651 vss 0.00413f
C14597 vdd.n5652 vss 0.0471f
C14598 vdd.n5653 vss 0.00251f
C14599 vdd.t595 vss 0.0471f
C14600 vdd.n5654 vss 0.00324f
C14601 vdd.n5656 vss 0.00679f
C14602 vdd.n5657 vss 0.00413f
C14603 vdd.n5658 vss 0.00324f
C14604 vdd.n5659 vss 0.00413f
C14605 vdd.n5660 vss 0.0471f
C14606 vdd.n5661 vss 0.00324f
C14607 vdd.n5663 vss 0.00925f
C14608 vdd.t144 vss 0.0471f
C14609 vdd.n5664 vss 0.00425f
C14610 vdd.n5665 vss 0.0424f
C14611 vdd.n5666 vss 0.0132f
C14612 vdd.n5667 vss 0.00324f
C14613 vdd.n5668 vss 0.0128f
C14614 vdd.n5669 vss 0.02f
C14615 vdd.n5670 vss 0.00425f
C14616 vdd.n5671 vss 0.00413f
C14617 vdd.n5672 vss 0.00251f
C14618 vdd.t396 vss 0.0471f
C14619 vdd.n5673 vss 0.00251f
C14620 vdd.n5674 vss 0.00517f
C14621 vdd.n5675 vss 0.00679f
C14622 vdd.n5676 vss 0.00517f
C14623 vdd.n5677 vss 0.00679f
C14624 vdd.n5678 vss 0.02f
C14625 vdd.n5679 vss 0.00425f
C14626 vdd.n5680 vss 0.0424f
C14627 vdd.n5681 vss 0.0132f
C14628 vdd.n5682 vss 0.00925f
C14629 vdd.n5683 vss 0.00425f
C14630 vdd.n5684 vss 0.00413f
C14631 vdd.n5685 vss 0.00324f
C14632 vdd.n5686 vss 0.0471f
C14633 vdd.t397 vss 0.0471f
C14634 vdd.n5687 vss 0.00251f
C14635 vdd.n5688 vss 0.0112f
C14636 vdd.n5689 vss 0.0128f
C14637 vdd.t398 vss 0.00134f
C14638 vdd.t596 vss 0.0013f
C14639 vdd.n5690 vss 0.0332f
C14640 vdd.n5691 vss 0.0393f
C14641 vdd.n5692 vss 0.0418f
C14642 vdd.n5693 vss 0.118f
C14643 vdd.n5694 vss 0.121f
C14644 vdd.t991 vss 0.0013f
C14645 vdd.t1216 vss 0.00134f
C14646 vdd.n5695 vss 0.00324f
C14647 vdd.n5696 vss 0.0112f
C14648 vdd.n5697 vss 0.0128f
C14649 vdd.n5698 vss 0.00413f
C14650 vdd.n5699 vss 0.00413f
C14651 vdd.n5700 vss 0.0471f
C14652 vdd.n5701 vss 0.00251f
C14653 vdd.t990 vss 0.0471f
C14654 vdd.n5702 vss 0.00324f
C14655 vdd.n5704 vss 0.00679f
C14656 vdd.n5705 vss 0.00413f
C14657 vdd.n5706 vss 0.00324f
C14658 vdd.n5707 vss 0.00413f
C14659 vdd.n5708 vss 0.0471f
C14660 vdd.n5709 vss 0.00324f
C14661 vdd.n5711 vss 0.00925f
C14662 vdd.t924 vss 0.0471f
C14663 vdd.n5712 vss 0.00425f
C14664 vdd.n5713 vss 0.0424f
C14665 vdd.n5714 vss 0.0132f
C14666 vdd.n5715 vss 0.00324f
C14667 vdd.n5716 vss 0.0128f
C14668 vdd.n5717 vss 0.02f
C14669 vdd.n5718 vss 0.00425f
C14670 vdd.n5719 vss 0.00413f
C14671 vdd.n5720 vss 0.00251f
C14672 vdd.t1214 vss 0.0471f
C14673 vdd.n5721 vss 0.00251f
C14674 vdd.n5722 vss 0.00517f
C14675 vdd.n5723 vss 0.00679f
C14676 vdd.n5724 vss 0.00517f
C14677 vdd.n5725 vss 0.00679f
C14678 vdd.n5726 vss 0.02f
C14679 vdd.n5727 vss 0.00425f
C14680 vdd.n5728 vss 0.0424f
C14681 vdd.n5729 vss 0.0132f
C14682 vdd.n5730 vss 0.00925f
C14683 vdd.n5731 vss 0.00425f
C14684 vdd.n5732 vss 0.00413f
C14685 vdd.n5733 vss 0.00324f
C14686 vdd.n5734 vss 0.0471f
C14687 vdd.t1215 vss 0.0471f
C14688 vdd.n5735 vss 0.00251f
C14689 vdd.n5736 vss 0.0112f
C14690 vdd.n5737 vss 0.0707f
C14691 vdd.n5738 vss 0.0393f
C14692 vdd.n5739 vss 0.0332f
C14693 vdd.n5740 vss 0.0596f
C14694 vdd.n5741 vss 0.00324f
C14695 vdd.n5742 vss 0.0112f
C14696 vdd.n5743 vss 0.0128f
C14697 vdd.n5744 vss 0.00413f
C14698 vdd.n5745 vss 0.00413f
C14699 vdd.n5746 vss 0.0471f
C14700 vdd.n5747 vss 0.00251f
C14701 vdd.t13 vss 0.0471f
C14702 vdd.n5748 vss 0.00324f
C14703 vdd.n5750 vss 0.00679f
C14704 vdd.n5751 vss 0.00413f
C14705 vdd.n5752 vss 0.00324f
C14706 vdd.n5753 vss 0.00413f
C14707 vdd.n5754 vss 0.0471f
C14708 vdd.n5755 vss 0.00324f
C14709 vdd.n5757 vss 0.00925f
C14710 vdd.t424 vss 0.0471f
C14711 vdd.n5758 vss 0.00425f
C14712 vdd.n5759 vss 0.0424f
C14713 vdd.n5760 vss 0.0132f
C14714 vdd.n5761 vss 0.00324f
C14715 vdd.n5762 vss 0.0128f
C14716 vdd.n5763 vss 0.02f
C14717 vdd.n5764 vss 0.00425f
C14718 vdd.n5765 vss 0.00413f
C14719 vdd.n5766 vss 0.00251f
C14720 vdd.t583 vss 0.0471f
C14721 vdd.n5767 vss 0.00251f
C14722 vdd.n5768 vss 0.00517f
C14723 vdd.n5769 vss 0.00679f
C14724 vdd.n5770 vss 0.00517f
C14725 vdd.n5771 vss 0.00679f
C14726 vdd.n5772 vss 0.02f
C14727 vdd.n5773 vss 0.00425f
C14728 vdd.n5774 vss 0.0424f
C14729 vdd.n5775 vss 0.0132f
C14730 vdd.n5776 vss 0.00925f
C14731 vdd.n5777 vss 0.00425f
C14732 vdd.n5778 vss 0.00413f
C14733 vdd.n5779 vss 0.00324f
C14734 vdd.n5780 vss 0.0471f
C14735 vdd.t581 vss 0.0471f
C14736 vdd.n5781 vss 0.00251f
C14737 vdd.n5782 vss 0.0112f
C14738 vdd.n5783 vss 0.0128f
C14739 vdd.t582 vss 0.00134f
C14740 vdd.t14 vss 0.0013f
C14741 vdd.n5784 vss 0.0332f
C14742 vdd.n5785 vss 0.0393f
C14743 vdd.n5786 vss 0.0418f
C14744 vdd.n5787 vss 0.0912f
C14745 vdd.n5788 vss 0.0824f
C14746 vdd.n5789 vss 0.059f
C14747 vdd.t867 vss 0.0013f
C14748 vdd.t329 vss 0.00134f
C14749 vdd.n5790 vss 0.00324f
C14750 vdd.n5791 vss 0.0112f
C14751 vdd.n5792 vss 0.0128f
C14752 vdd.n5793 vss 0.00413f
C14753 vdd.n5794 vss 0.00413f
C14754 vdd.n5795 vss 0.0471f
C14755 vdd.n5796 vss 0.00251f
C14756 vdd.t1373 vss 0.0471f
C14757 vdd.n5797 vss 0.00324f
C14758 vdd.n5799 vss 0.00679f
C14759 vdd.n5800 vss 0.00413f
C14760 vdd.n5801 vss 0.00324f
C14761 vdd.n5802 vss 0.00413f
C14762 vdd.n5803 vss 0.0471f
C14763 vdd.n5804 vss 0.00324f
C14764 vdd.n5806 vss 0.00925f
C14765 vdd.t928 vss 0.0471f
C14766 vdd.n5807 vss 0.00425f
C14767 vdd.n5808 vss 0.0424f
C14768 vdd.n5809 vss 0.0132f
C14769 vdd.n5810 vss 0.00324f
C14770 vdd.n5811 vss 0.0128f
C14771 vdd.n5812 vss 0.02f
C14772 vdd.n5813 vss 0.00425f
C14773 vdd.n5814 vss 0.00413f
C14774 vdd.n5815 vss 0.00251f
C14775 vdd.t777 vss 0.0471f
C14776 vdd.n5816 vss 0.00251f
C14777 vdd.n5817 vss 0.00517f
C14778 vdd.n5818 vss 0.00679f
C14779 vdd.n5819 vss 0.00517f
C14780 vdd.n5820 vss 0.00679f
C14781 vdd.n5821 vss 0.02f
C14782 vdd.n5822 vss 0.00425f
C14783 vdd.n5823 vss 0.0424f
C14784 vdd.n5824 vss 0.0132f
C14785 vdd.n5825 vss 0.00925f
C14786 vdd.n5826 vss 0.00425f
C14787 vdd.n5827 vss 0.00413f
C14788 vdd.n5828 vss 0.00324f
C14789 vdd.n5829 vss 0.0471f
C14790 vdd.t778 vss 0.0471f
C14791 vdd.n5830 vss 0.00251f
C14792 vdd.n5831 vss 0.0112f
C14793 vdd.n5832 vss 0.0128f
C14794 vdd.t779 vss 0.00134f
C14795 vdd.t1374 vss 0.0013f
C14796 vdd.n5833 vss 0.0332f
C14797 vdd.n5834 vss 0.0393f
C14798 vdd.n5835 vss 0.158f
C14799 vdd.n5836 vss 0.00324f
C14800 vdd.n5837 vss 0.0112f
C14801 vdd.n5838 vss 0.0128f
C14802 vdd.n5839 vss 0.00413f
C14803 vdd.n5840 vss 0.00413f
C14804 vdd.n5841 vss 0.0471f
C14805 vdd.n5842 vss 0.00251f
C14806 vdd.t767 vss 0.0471f
C14807 vdd.n5843 vss 0.00324f
C14808 vdd.n5845 vss 0.00679f
C14809 vdd.n5846 vss 0.00413f
C14810 vdd.n5847 vss 0.00324f
C14811 vdd.n5848 vss 0.00413f
C14812 vdd.n5849 vss 0.0471f
C14813 vdd.n5850 vss 0.00324f
C14814 vdd.n5852 vss 0.00925f
C14815 vdd.t786 vss 0.0471f
C14816 vdd.n5853 vss 0.00425f
C14817 vdd.n5854 vss 0.0424f
C14818 vdd.n5855 vss 0.0132f
C14819 vdd.n5856 vss 0.00324f
C14820 vdd.n5857 vss 0.0128f
C14821 vdd.n5858 vss 0.02f
C14822 vdd.n5859 vss 0.00425f
C14823 vdd.n5860 vss 0.00413f
C14824 vdd.n5861 vss 0.00251f
C14825 vdd.t1527 vss 0.0471f
C14826 vdd.n5862 vss 0.00251f
C14827 vdd.n5863 vss 0.00517f
C14828 vdd.n5864 vss 0.00679f
C14829 vdd.n5865 vss 0.00517f
C14830 vdd.n5866 vss 0.00679f
C14831 vdd.n5867 vss 0.02f
C14832 vdd.n5868 vss 0.00425f
C14833 vdd.n5869 vss 0.0424f
C14834 vdd.n5870 vss 0.0132f
C14835 vdd.n5871 vss 0.00925f
C14836 vdd.n5872 vss 0.00425f
C14837 vdd.n5873 vss 0.00413f
C14838 vdd.n5874 vss 0.00324f
C14839 vdd.n5875 vss 0.0471f
C14840 vdd.t1528 vss 0.0471f
C14841 vdd.n5876 vss 0.00251f
C14842 vdd.n5877 vss 0.0112f
C14843 vdd.n5878 vss 0.0128f
C14844 vdd.t1529 vss 0.00134f
C14845 vdd.t768 vss 0.0013f
C14846 vdd.n5879 vss 0.0332f
C14847 vdd.n5880 vss 0.0393f
C14848 vdd.n5881 vss 0.0316f
C14849 vdd.n5882 vss 0.256f
C14850 vdd.n5883 vss 0.00324f
C14851 vdd.n5884 vss 0.0112f
C14852 vdd.n5885 vss 0.0128f
C14853 vdd.n5886 vss 0.00413f
C14854 vdd.n5887 vss 0.00413f
C14855 vdd.n5888 vss 0.0471f
C14856 vdd.n5889 vss 0.00251f
C14857 vdd.t866 vss 0.0471f
C14858 vdd.n5890 vss 0.00324f
C14859 vdd.n5892 vss 0.00679f
C14860 vdd.n5893 vss 0.00413f
C14861 vdd.n5894 vss 0.00324f
C14862 vdd.n5895 vss 0.00413f
C14863 vdd.n5896 vss 0.0471f
C14864 vdd.n5897 vss 0.00324f
C14865 vdd.n5899 vss 0.00925f
C14866 vdd.t23 vss 0.0471f
C14867 vdd.n5900 vss 0.00425f
C14868 vdd.n5901 vss 0.0424f
C14869 vdd.n5902 vss 0.0132f
C14870 vdd.n5903 vss 0.00324f
C14871 vdd.n5904 vss 0.0128f
C14872 vdd.n5905 vss 0.02f
C14873 vdd.n5906 vss 0.00425f
C14874 vdd.n5907 vss 0.00413f
C14875 vdd.n5908 vss 0.00251f
C14876 vdd.t330 vss 0.0471f
C14877 vdd.n5909 vss 0.00251f
C14878 vdd.n5910 vss 0.00517f
C14879 vdd.n5911 vss 0.00679f
C14880 vdd.n5912 vss 0.00517f
C14881 vdd.n5913 vss 0.00679f
C14882 vdd.n5914 vss 0.02f
C14883 vdd.n5915 vss 0.00425f
C14884 vdd.n5916 vss 0.0424f
C14885 vdd.n5917 vss 0.0132f
C14886 vdd.n5918 vss 0.00925f
C14887 vdd.n5919 vss 0.00425f
C14888 vdd.n5920 vss 0.00413f
C14889 vdd.n5921 vss 0.00324f
C14890 vdd.n5922 vss 0.0471f
C14891 vdd.t328 vss 0.0471f
C14892 vdd.n5923 vss 0.00251f
C14893 vdd.n5924 vss 0.0112f
C14894 vdd.n5925 vss 0.0128f
C14895 vdd.n5926 vss 0.0953f
C14896 vdd.n5927 vss 0.0393f
C14897 vdd.n5928 vss 0.0332f
C14898 vdd.n5929 vss 0.0596f
C14899 vdd.n5930 vss 0.00324f
C14900 vdd.n5931 vss 0.0112f
C14901 vdd.n5932 vss 0.0128f
C14902 vdd.n5933 vss 0.00413f
C14903 vdd.n5934 vss 0.00413f
C14904 vdd.n5935 vss 0.0471f
C14905 vdd.n5936 vss 0.00251f
C14906 vdd.t1479 vss 0.0471f
C14907 vdd.n5937 vss 0.00324f
C14908 vdd.n5939 vss 0.00679f
C14909 vdd.n5940 vss 0.00413f
C14910 vdd.n5941 vss 0.00324f
C14911 vdd.n5942 vss 0.00413f
C14912 vdd.n5943 vss 0.0471f
C14913 vdd.n5944 vss 0.00324f
C14914 vdd.n5946 vss 0.00925f
C14915 vdd.t679 vss 0.0471f
C14916 vdd.n5947 vss 0.00425f
C14917 vdd.n5948 vss 0.0424f
C14918 vdd.n5949 vss 0.0132f
C14919 vdd.n5950 vss 0.00324f
C14920 vdd.n5951 vss 0.0128f
C14921 vdd.n5952 vss 0.02f
C14922 vdd.n5953 vss 0.00425f
C14923 vdd.n5954 vss 0.00413f
C14924 vdd.n5955 vss 0.00251f
C14925 vdd.t676 vss 0.0471f
C14926 vdd.n5956 vss 0.00251f
C14927 vdd.n5957 vss 0.00517f
C14928 vdd.n5958 vss 0.00679f
C14929 vdd.n5959 vss 0.00517f
C14930 vdd.n5960 vss 0.00679f
C14931 vdd.n5961 vss 0.02f
C14932 vdd.n5962 vss 0.00425f
C14933 vdd.n5963 vss 0.0424f
C14934 vdd.n5964 vss 0.0132f
C14935 vdd.n5965 vss 0.00925f
C14936 vdd.n5966 vss 0.00425f
C14937 vdd.n5967 vss 0.00413f
C14938 vdd.n5968 vss 0.00324f
C14939 vdd.n5969 vss 0.0471f
C14940 vdd.t677 vss 0.0471f
C14941 vdd.n5970 vss 0.00251f
C14942 vdd.n5971 vss 0.0112f
C14943 vdd.n5972 vss 0.0128f
C14944 vdd.t678 vss 0.00134f
C14945 vdd.t1480 vss 0.0013f
C14946 vdd.n5973 vss 0.0332f
C14947 vdd.n5974 vss 0.0393f
C14948 vdd.n5975 vss 0.0418f
C14949 vdd.n5976 vss 0.118f
C14950 vdd.n5977 vss 0.121f
C14951 vdd.t1003 vss 0.0013f
C14952 vdd.t1194 vss 0.00134f
C14953 vdd.n5978 vss 0.00324f
C14954 vdd.n5979 vss 0.0112f
C14955 vdd.n5980 vss 0.0128f
C14956 vdd.n5981 vss 0.00413f
C14957 vdd.n5982 vss 0.00413f
C14958 vdd.n5983 vss 0.0471f
C14959 vdd.n5984 vss 0.00251f
C14960 vdd.t1002 vss 0.0471f
C14961 vdd.n5985 vss 0.00324f
C14962 vdd.n5987 vss 0.00679f
C14963 vdd.n5988 vss 0.00413f
C14964 vdd.n5989 vss 0.00324f
C14965 vdd.n5990 vss 0.00413f
C14966 vdd.n5991 vss 0.0471f
C14967 vdd.n5992 vss 0.00324f
C14968 vdd.n5994 vss 0.00925f
C14969 vdd.t1258 vss 0.0471f
C14970 vdd.n5995 vss 0.00425f
C14971 vdd.n5996 vss 0.0424f
C14972 vdd.n5997 vss 0.0132f
C14973 vdd.n5998 vss 0.00324f
C14974 vdd.n5999 vss 0.0128f
C14975 vdd.n6000 vss 0.02f
C14976 vdd.n6001 vss 0.00425f
C14977 vdd.n6002 vss 0.00413f
C14978 vdd.n6003 vss 0.00251f
C14979 vdd.t1192 vss 0.0471f
C14980 vdd.n6004 vss 0.00251f
C14981 vdd.n6005 vss 0.00517f
C14982 vdd.n6006 vss 0.00679f
C14983 vdd.n6007 vss 0.00517f
C14984 vdd.n6008 vss 0.00679f
C14985 vdd.n6009 vss 0.02f
C14986 vdd.n6010 vss 0.00425f
C14987 vdd.n6011 vss 0.0424f
C14988 vdd.n6012 vss 0.0132f
C14989 vdd.n6013 vss 0.00925f
C14990 vdd.n6014 vss 0.00425f
C14991 vdd.n6015 vss 0.00413f
C14992 vdd.n6016 vss 0.00324f
C14993 vdd.n6017 vss 0.0471f
C14994 vdd.t1193 vss 0.0471f
C14995 vdd.n6018 vss 0.00251f
C14996 vdd.n6019 vss 0.0112f
C14997 vdd.n6020 vss 0.0707f
C14998 vdd.n6021 vss 0.0393f
C14999 vdd.n6022 vss 0.0332f
C15000 vdd.n6023 vss 0.0596f
C15001 vdd.n6024 vss 0.00324f
C15002 vdd.n6025 vss 0.0112f
C15003 vdd.n6026 vss 0.0128f
C15004 vdd.n6027 vss 0.00413f
C15005 vdd.n6028 vss 0.00413f
C15006 vdd.n6029 vss 0.0471f
C15007 vdd.n6030 vss 0.00251f
C15008 vdd.t1489 vss 0.0471f
C15009 vdd.n6031 vss 0.00324f
C15010 vdd.n6033 vss 0.00679f
C15011 vdd.n6034 vss 0.00413f
C15012 vdd.n6035 vss 0.00324f
C15013 vdd.n6036 vss 0.00413f
C15014 vdd.n6037 vss 0.0471f
C15015 vdd.n6038 vss 0.00324f
C15016 vdd.n6040 vss 0.00925f
C15017 vdd.t429 vss 0.0471f
C15018 vdd.n6041 vss 0.00425f
C15019 vdd.n6042 vss 0.0424f
C15020 vdd.n6043 vss 0.0132f
C15021 vdd.n6044 vss 0.00324f
C15022 vdd.n6045 vss 0.0128f
C15023 vdd.n6046 vss 0.02f
C15024 vdd.n6047 vss 0.00425f
C15025 vdd.n6048 vss 0.00413f
C15026 vdd.n6049 vss 0.00251f
C15027 vdd.t2 vss 0.0471f
C15028 vdd.n6050 vss 0.00251f
C15029 vdd.n6051 vss 0.00517f
C15030 vdd.n6052 vss 0.00679f
C15031 vdd.n6053 vss 0.00517f
C15032 vdd.n6054 vss 0.00679f
C15033 vdd.n6055 vss 0.02f
C15034 vdd.n6056 vss 0.00425f
C15035 vdd.n6057 vss 0.0424f
C15036 vdd.n6058 vss 0.0132f
C15037 vdd.n6059 vss 0.00925f
C15038 vdd.n6060 vss 0.00425f
C15039 vdd.n6061 vss 0.00413f
C15040 vdd.n6062 vss 0.00324f
C15041 vdd.n6063 vss 0.0471f
C15042 vdd.t0 vss 0.0471f
C15043 vdd.n6064 vss 0.00251f
C15044 vdd.n6065 vss 0.0112f
C15045 vdd.n6066 vss 0.0128f
C15046 vdd.t1 vss 0.00134f
C15047 vdd.t1490 vss 0.0013f
C15048 vdd.n6067 vss 0.0332f
C15049 vdd.n6068 vss 0.0393f
C15050 vdd.n6069 vss 0.0418f
C15051 vdd.n6070 vss 0.118f
C15052 vdd.n6071 vss 0.0951f
C15053 vdd.t970 vss 0.0013f
C15054 vdd.t633 vss 0.00134f
C15055 vdd.n6072 vss 0.00324f
C15056 vdd.n6073 vss 0.0112f
C15057 vdd.n6074 vss 0.0128f
C15058 vdd.n6075 vss 0.00413f
C15059 vdd.n6076 vss 0.00413f
C15060 vdd.n6077 vss 0.0471f
C15061 vdd.n6078 vss 0.00251f
C15062 vdd.t434 vss 0.0471f
C15063 vdd.n6079 vss 0.00324f
C15064 vdd.n6081 vss 0.00679f
C15065 vdd.n6082 vss 0.00413f
C15066 vdd.n6083 vss 0.00324f
C15067 vdd.n6084 vss 0.00413f
C15068 vdd.n6085 vss 0.0471f
C15069 vdd.n6086 vss 0.00324f
C15070 vdd.n6088 vss 0.00925f
C15071 vdd.t671 vss 0.0471f
C15072 vdd.n6089 vss 0.00425f
C15073 vdd.n6090 vss 0.0424f
C15074 vdd.n6091 vss 0.0132f
C15075 vdd.n6092 vss 0.00324f
C15076 vdd.n6093 vss 0.0128f
C15077 vdd.n6094 vss 0.02f
C15078 vdd.n6095 vss 0.00425f
C15079 vdd.n6096 vss 0.00413f
C15080 vdd.n6097 vss 0.00251f
C15081 vdd.t1206 vss 0.0471f
C15082 vdd.n6098 vss 0.00251f
C15083 vdd.n6099 vss 0.00517f
C15084 vdd.n6100 vss 0.00679f
C15085 vdd.n6101 vss 0.00517f
C15086 vdd.n6102 vss 0.00679f
C15087 vdd.n6103 vss 0.02f
C15088 vdd.n6104 vss 0.00425f
C15089 vdd.n6105 vss 0.0424f
C15090 vdd.n6106 vss 0.0132f
C15091 vdd.n6107 vss 0.00925f
C15092 vdd.n6108 vss 0.00425f
C15093 vdd.n6109 vss 0.00413f
C15094 vdd.n6110 vss 0.00324f
C15095 vdd.n6111 vss 0.0471f
C15096 vdd.t1204 vss 0.0471f
C15097 vdd.n6112 vss 0.00251f
C15098 vdd.n6113 vss 0.0112f
C15099 vdd.n6114 vss 0.0128f
C15100 vdd.t1205 vss 0.00134f
C15101 vdd.t435 vss 0.0013f
C15102 vdd.n6115 vss 0.0332f
C15103 vdd.n6116 vss 0.0393f
C15104 vdd.n6117 vss 0.119f
C15105 vdd.n6118 vss 0.00324f
C15106 vdd.n6119 vss 0.0112f
C15107 vdd.n6120 vss 0.0128f
C15108 vdd.n6121 vss 0.00413f
C15109 vdd.n6122 vss 0.00413f
C15110 vdd.n6123 vss 0.0471f
C15111 vdd.n6124 vss 0.00251f
C15112 vdd.t969 vss 0.0471f
C15113 vdd.n6125 vss 0.00324f
C15114 vdd.n6127 vss 0.00679f
C15115 vdd.n6128 vss 0.00413f
C15116 vdd.n6129 vss 0.00324f
C15117 vdd.n6130 vss 0.00413f
C15118 vdd.n6131 vss 0.0471f
C15119 vdd.n6132 vss 0.00324f
C15120 vdd.n6134 vss 0.00925f
C15121 vdd.t305 vss 0.0471f
C15122 vdd.n6135 vss 0.00425f
C15123 vdd.n6136 vss 0.0424f
C15124 vdd.n6137 vss 0.0132f
C15125 vdd.n6138 vss 0.00324f
C15126 vdd.n6139 vss 0.0128f
C15127 vdd.n6140 vss 0.02f
C15128 vdd.n6141 vss 0.00425f
C15129 vdd.n6142 vss 0.00413f
C15130 vdd.n6143 vss 0.00251f
C15131 vdd.t631 vss 0.0471f
C15132 vdd.n6144 vss 0.00251f
C15133 vdd.n6145 vss 0.00517f
C15134 vdd.n6146 vss 0.00679f
C15135 vdd.n6147 vss 0.00517f
C15136 vdd.n6148 vss 0.00679f
C15137 vdd.n6149 vss 0.02f
C15138 vdd.n6150 vss 0.00425f
C15139 vdd.n6151 vss 0.0424f
C15140 vdd.n6152 vss 0.0132f
C15141 vdd.n6153 vss 0.00925f
C15142 vdd.n6154 vss 0.00425f
C15143 vdd.n6155 vss 0.00413f
C15144 vdd.n6156 vss 0.00324f
C15145 vdd.n6157 vss 0.0471f
C15146 vdd.t632 vss 0.0471f
C15147 vdd.n6158 vss 0.00251f
C15148 vdd.n6159 vss 0.0112f
C15149 vdd.n6160 vss 0.0128f
C15150 vdd.n6161 vss 0.118f
C15151 vdd.n6162 vss 0.0393f
C15152 vdd.n6163 vss 0.0332f
C15153 vdd.n6164 vss 0.0596f
C15154 vdd.n6165 vss 0.00324f
C15155 vdd.n6166 vss 0.0112f
C15156 vdd.n6167 vss 0.0128f
C15157 vdd.n6168 vss 0.00413f
C15158 vdd.n6169 vss 0.00413f
C15159 vdd.n6170 vss 0.0471f
C15160 vdd.n6171 vss 0.00251f
C15161 vdd.t1336 vss 0.0471f
C15162 vdd.n6172 vss 0.00324f
C15163 vdd.n6174 vss 0.00679f
C15164 vdd.n6175 vss 0.00413f
C15165 vdd.n6176 vss 0.00324f
C15166 vdd.n6177 vss 0.00413f
C15167 vdd.n6178 vss 0.0471f
C15168 vdd.n6179 vss 0.00324f
C15169 vdd.n6181 vss 0.00925f
C15170 vdd.t387 vss 0.0471f
C15171 vdd.n6182 vss 0.00425f
C15172 vdd.n6183 vss 0.0424f
C15173 vdd.n6184 vss 0.0132f
C15174 vdd.n6185 vss 0.00324f
C15175 vdd.n6186 vss 0.0128f
C15176 vdd.n6187 vss 0.02f
C15177 vdd.n6188 vss 0.00425f
C15178 vdd.n6189 vss 0.00413f
C15179 vdd.n6190 vss 0.00251f
C15180 vdd.t1157 vss 0.0471f
C15181 vdd.n6191 vss 0.00251f
C15182 vdd.n6192 vss 0.00517f
C15183 vdd.n6193 vss 0.00679f
C15184 vdd.n6194 vss 0.00517f
C15185 vdd.n6195 vss 0.00679f
C15186 vdd.n6196 vss 0.02f
C15187 vdd.n6197 vss 0.00425f
C15188 vdd.n6198 vss 0.0424f
C15189 vdd.n6199 vss 0.0132f
C15190 vdd.n6200 vss 0.00925f
C15191 vdd.n6201 vss 0.00425f
C15192 vdd.n6202 vss 0.00413f
C15193 vdd.n6203 vss 0.00324f
C15194 vdd.n6204 vss 0.0471f
C15195 vdd.t1158 vss 0.0471f
C15196 vdd.n6205 vss 0.00251f
C15197 vdd.n6206 vss 0.0112f
C15198 vdd.n6207 vss 0.0128f
C15199 vdd.t1159 vss 0.00134f
C15200 vdd.t1337 vss 0.0013f
C15201 vdd.n6208 vss 0.0332f
C15202 vdd.n6209 vss 0.0393f
C15203 vdd.n6210 vss 0.0418f
C15204 vdd.n6211 vss 0.118f
C15205 vdd.n6212 vss 0.121f
C15206 vdd.t33 vss 0.0013f
C15207 vdd.t1405 vss 0.00134f
C15208 vdd.n6213 vss 0.00324f
C15209 vdd.n6214 vss 0.0112f
C15210 vdd.n6215 vss 0.0128f
C15211 vdd.n6216 vss 0.00413f
C15212 vdd.n6217 vss 0.00413f
C15213 vdd.n6218 vss 0.0471f
C15214 vdd.n6219 vss 0.00251f
C15215 vdd.t32 vss 0.0471f
C15216 vdd.n6220 vss 0.00324f
C15217 vdd.n6222 vss 0.00679f
C15218 vdd.n6223 vss 0.00413f
C15219 vdd.n6224 vss 0.00324f
C15220 vdd.n6225 vss 0.00413f
C15221 vdd.n6226 vss 0.0471f
C15222 vdd.n6227 vss 0.00324f
C15223 vdd.n6229 vss 0.00925f
C15224 vdd.t246 vss 0.0471f
C15225 vdd.n6230 vss 0.00425f
C15226 vdd.n6231 vss 0.0424f
C15227 vdd.n6232 vss 0.0132f
C15228 vdd.n6233 vss 0.00324f
C15229 vdd.n6234 vss 0.0128f
C15230 vdd.n6235 vss 0.02f
C15231 vdd.n6236 vss 0.00425f
C15232 vdd.n6237 vss 0.00413f
C15233 vdd.n6238 vss 0.00251f
C15234 vdd.t1403 vss 0.0471f
C15235 vdd.n6239 vss 0.00251f
C15236 vdd.n6240 vss 0.00517f
C15237 vdd.n6241 vss 0.00679f
C15238 vdd.n6242 vss 0.00517f
C15239 vdd.n6243 vss 0.00679f
C15240 vdd.n6244 vss 0.02f
C15241 vdd.n6245 vss 0.00425f
C15242 vdd.n6246 vss 0.0424f
C15243 vdd.n6247 vss 0.0132f
C15244 vdd.n6248 vss 0.00925f
C15245 vdd.n6249 vss 0.00425f
C15246 vdd.n6250 vss 0.00413f
C15247 vdd.n6251 vss 0.00324f
C15248 vdd.n6252 vss 0.0471f
C15249 vdd.t1404 vss 0.0471f
C15250 vdd.n6253 vss 0.00251f
C15251 vdd.n6254 vss 0.0112f
C15252 vdd.n6255 vss 0.0707f
C15253 vdd.n6256 vss 0.0393f
C15254 vdd.n6257 vss 0.0332f
C15255 vdd.n6258 vss 0.0596f
C15256 vdd.n6259 vss 0.00324f
C15257 vdd.n6260 vss 0.0112f
C15258 vdd.n6261 vss 0.0128f
C15259 vdd.n6262 vss 0.00413f
C15260 vdd.n6263 vss 0.00413f
C15261 vdd.n6264 vss 0.0471f
C15262 vdd.n6265 vss 0.00251f
C15263 vdd.t496 vss 0.0471f
C15264 vdd.n6266 vss 0.00324f
C15265 vdd.n6268 vss 0.00679f
C15266 vdd.n6269 vss 0.00413f
C15267 vdd.n6270 vss 0.00324f
C15268 vdd.n6271 vss 0.00413f
C15269 vdd.n6272 vss 0.0471f
C15270 vdd.n6273 vss 0.00324f
C15271 vdd.n6275 vss 0.00925f
C15272 vdd.t1026 vss 0.0471f
C15273 vdd.n6276 vss 0.00425f
C15274 vdd.n6277 vss 0.0424f
C15275 vdd.n6278 vss 0.0132f
C15276 vdd.n6279 vss 0.00324f
C15277 vdd.n6280 vss 0.0128f
C15278 vdd.n6281 vss 0.02f
C15279 vdd.n6282 vss 0.00425f
C15280 vdd.n6283 vss 0.00413f
C15281 vdd.n6284 vss 0.00251f
C15282 vdd.t944 vss 0.0471f
C15283 vdd.n6285 vss 0.00251f
C15284 vdd.n6286 vss 0.00517f
C15285 vdd.n6287 vss 0.00679f
C15286 vdd.n6288 vss 0.00517f
C15287 vdd.n6289 vss 0.00679f
C15288 vdd.n6290 vss 0.02f
C15289 vdd.n6291 vss 0.00425f
C15290 vdd.n6292 vss 0.0424f
C15291 vdd.n6293 vss 0.0132f
C15292 vdd.n6294 vss 0.00925f
C15293 vdd.n6295 vss 0.00425f
C15294 vdd.n6296 vss 0.00413f
C15295 vdd.n6297 vss 0.00324f
C15296 vdd.n6298 vss 0.0471f
C15297 vdd.t945 vss 0.0471f
C15298 vdd.n6299 vss 0.00251f
C15299 vdd.n6300 vss 0.0112f
C15300 vdd.n6301 vss 0.0128f
C15301 vdd.t946 vss 0.00134f
C15302 vdd.t497 vss 0.0013f
C15303 vdd.n6302 vss 0.0332f
C15304 vdd.n6303 vss 0.0393f
C15305 vdd.n6304 vss 0.0418f
C15306 vdd.n6305 vss 0.0912f
C15307 vdd.n6306 vss 0.0824f
C15308 vdd.n6307 vss 0.059f
C15309 vdd.t869 vss 0.0013f
C15310 vdd.t19 vss 0.00134f
C15311 vdd.n6308 vss 0.00324f
C15312 vdd.n6309 vss 0.0112f
C15313 vdd.n6310 vss 0.0128f
C15314 vdd.n6311 vss 0.00413f
C15315 vdd.n6312 vss 0.00413f
C15316 vdd.n6313 vss 0.0471f
C15317 vdd.n6314 vss 0.00251f
C15318 vdd.t432 vss 0.0471f
C15319 vdd.n6315 vss 0.00324f
C15320 vdd.n6317 vss 0.00679f
C15321 vdd.n6318 vss 0.00413f
C15322 vdd.n6319 vss 0.00324f
C15323 vdd.n6320 vss 0.00413f
C15324 vdd.n6321 vss 0.0471f
C15325 vdd.n6322 vss 0.00324f
C15326 vdd.n6324 vss 0.00925f
C15327 vdd.t331 vss 0.0471f
C15328 vdd.n6325 vss 0.00425f
C15329 vdd.n6326 vss 0.0424f
C15330 vdd.n6327 vss 0.0132f
C15331 vdd.n6328 vss 0.00324f
C15332 vdd.n6329 vss 0.0128f
C15333 vdd.n6330 vss 0.02f
C15334 vdd.n6331 vss 0.00425f
C15335 vdd.n6332 vss 0.00413f
C15336 vdd.n6333 vss 0.00251f
C15337 vdd.t749 vss 0.0471f
C15338 vdd.n6334 vss 0.00251f
C15339 vdd.n6335 vss 0.00517f
C15340 vdd.n6336 vss 0.00679f
C15341 vdd.n6337 vss 0.00517f
C15342 vdd.n6338 vss 0.00679f
C15343 vdd.n6339 vss 0.02f
C15344 vdd.n6340 vss 0.00425f
C15345 vdd.n6341 vss 0.0424f
C15346 vdd.n6342 vss 0.0132f
C15347 vdd.n6343 vss 0.00925f
C15348 vdd.n6344 vss 0.00425f
C15349 vdd.n6345 vss 0.00413f
C15350 vdd.n6346 vss 0.00324f
C15351 vdd.n6347 vss 0.0471f
C15352 vdd.t750 vss 0.0471f
C15353 vdd.n6348 vss 0.00251f
C15354 vdd.n6349 vss 0.0112f
C15355 vdd.n6350 vss 0.0128f
C15356 vdd.t751 vss 0.00134f
C15357 vdd.t433 vss 0.0013f
C15358 vdd.n6351 vss 0.0332f
C15359 vdd.n6352 vss 0.0393f
C15360 vdd.n6353 vss 0.119f
C15361 vdd.n6354 vss 0.00324f
C15362 vdd.n6355 vss 0.0112f
C15363 vdd.n6356 vss 0.0128f
C15364 vdd.n6357 vss 0.00413f
C15365 vdd.n6358 vss 0.00413f
C15366 vdd.n6359 vss 0.0471f
C15367 vdd.n6360 vss 0.00251f
C15368 vdd.t868 vss 0.0471f
C15369 vdd.n6361 vss 0.00324f
C15370 vdd.n6363 vss 0.00679f
C15371 vdd.n6364 vss 0.00413f
C15372 vdd.n6365 vss 0.00324f
C15373 vdd.n6366 vss 0.00413f
C15374 vdd.n6367 vss 0.0471f
C15375 vdd.n6368 vss 0.00324f
C15376 vdd.n6370 vss 0.00925f
C15377 vdd.t20 vss 0.0471f
C15378 vdd.n6371 vss 0.00425f
C15379 vdd.n6372 vss 0.0424f
C15380 vdd.n6373 vss 0.0132f
C15381 vdd.n6374 vss 0.00324f
C15382 vdd.n6375 vss 0.0128f
C15383 vdd.n6376 vss 0.02f
C15384 vdd.n6377 vss 0.00425f
C15385 vdd.n6378 vss 0.00413f
C15386 vdd.n6379 vss 0.00251f
C15387 vdd.t17 vss 0.0471f
C15388 vdd.n6380 vss 0.00251f
C15389 vdd.n6381 vss 0.00517f
C15390 vdd.n6382 vss 0.00679f
C15391 vdd.n6383 vss 0.00517f
C15392 vdd.n6384 vss 0.00679f
C15393 vdd.n6385 vss 0.02f
C15394 vdd.n6386 vss 0.00425f
C15395 vdd.n6387 vss 0.0424f
C15396 vdd.n6388 vss 0.0132f
C15397 vdd.n6389 vss 0.00925f
C15398 vdd.n6390 vss 0.00425f
C15399 vdd.n6391 vss 0.00413f
C15400 vdd.n6392 vss 0.00324f
C15401 vdd.n6393 vss 0.0471f
C15402 vdd.t18 vss 0.0471f
C15403 vdd.n6394 vss 0.00251f
C15404 vdd.n6395 vss 0.0112f
C15405 vdd.n6396 vss 0.0128f
C15406 vdd.n6397 vss 0.118f
C15407 vdd.n6398 vss 0.0393f
C15408 vdd.n6399 vss 0.0332f
C15409 vdd.n6400 vss 0.0596f
C15410 vdd.n6401 vss 0.00324f
C15411 vdd.n6402 vss 0.0112f
C15412 vdd.n6403 vss 0.0128f
C15413 vdd.n6404 vss 0.00413f
C15414 vdd.n6405 vss 0.00413f
C15415 vdd.n6406 vss 0.0471f
C15416 vdd.n6407 vss 0.00251f
C15417 vdd.t1053 vss 0.0471f
C15418 vdd.n6408 vss 0.00324f
C15419 vdd.n6410 vss 0.00679f
C15420 vdd.n6411 vss 0.00413f
C15421 vdd.n6412 vss 0.00324f
C15422 vdd.n6413 vss 0.00413f
C15423 vdd.n6414 vss 0.0471f
C15424 vdd.n6415 vss 0.00324f
C15425 vdd.n6417 vss 0.00925f
C15426 vdd.t615 vss 0.0471f
C15427 vdd.n6418 vss 0.00425f
C15428 vdd.n6419 vss 0.0424f
C15429 vdd.n6420 vss 0.0132f
C15430 vdd.n6421 vss 0.00324f
C15431 vdd.n6422 vss 0.0128f
C15432 vdd.n6423 vss 0.02f
C15433 vdd.n6424 vss 0.00425f
C15434 vdd.n6425 vss 0.00413f
C15435 vdd.n6426 vss 0.00251f
C15436 vdd.t686 vss 0.0471f
C15437 vdd.n6427 vss 0.00251f
C15438 vdd.n6428 vss 0.00517f
C15439 vdd.n6429 vss 0.00679f
C15440 vdd.n6430 vss 0.00517f
C15441 vdd.n6431 vss 0.00679f
C15442 vdd.n6432 vss 0.02f
C15443 vdd.n6433 vss 0.00425f
C15444 vdd.n6434 vss 0.0424f
C15445 vdd.n6435 vss 0.0132f
C15446 vdd.n6436 vss 0.00925f
C15447 vdd.n6437 vss 0.00425f
C15448 vdd.n6438 vss 0.00413f
C15449 vdd.n6439 vss 0.00324f
C15450 vdd.n6440 vss 0.0471f
C15451 vdd.t684 vss 0.0471f
C15452 vdd.n6441 vss 0.00251f
C15453 vdd.n6442 vss 0.0112f
C15454 vdd.n6443 vss 0.0128f
C15455 vdd.t685 vss 0.00134f
C15456 vdd.t1054 vss 0.0013f
C15457 vdd.n6444 vss 0.0332f
C15458 vdd.n6445 vss 0.0393f
C15459 vdd.n6446 vss 0.0418f
C15460 vdd.n6447 vss 0.118f
C15461 vdd.n6448 vss 0.121f
C15462 vdd.t895 vss 0.0013f
C15463 vdd.t1171 vss 0.00134f
C15464 vdd.n6449 vss 0.00324f
C15465 vdd.n6450 vss 0.0112f
C15466 vdd.n6451 vss 0.0128f
C15467 vdd.n6452 vss 0.00413f
C15468 vdd.n6453 vss 0.00413f
C15469 vdd.n6454 vss 0.0471f
C15470 vdd.n6455 vss 0.00251f
C15471 vdd.t894 vss 0.0471f
C15472 vdd.n6456 vss 0.00324f
C15473 vdd.n6458 vss 0.00679f
C15474 vdd.n6459 vss 0.00413f
C15475 vdd.n6460 vss 0.00324f
C15476 vdd.n6461 vss 0.00413f
C15477 vdd.n6462 vss 0.0471f
C15478 vdd.n6463 vss 0.00324f
C15479 vdd.n6465 vss 0.00925f
C15480 vdd.t1367 vss 0.0471f
C15481 vdd.n6466 vss 0.00425f
C15482 vdd.n6467 vss 0.0424f
C15483 vdd.n6468 vss 0.0132f
C15484 vdd.n6469 vss 0.00324f
C15485 vdd.n6470 vss 0.0128f
C15486 vdd.n6471 vss 0.02f
C15487 vdd.n6472 vss 0.00425f
C15488 vdd.n6473 vss 0.00413f
C15489 vdd.n6474 vss 0.00251f
C15490 vdd.t1169 vss 0.0471f
C15491 vdd.n6475 vss 0.00251f
C15492 vdd.n6476 vss 0.00517f
C15493 vdd.n6477 vss 0.00679f
C15494 vdd.n6478 vss 0.00517f
C15495 vdd.n6479 vss 0.00679f
C15496 vdd.n6480 vss 0.02f
C15497 vdd.n6481 vss 0.00425f
C15498 vdd.n6482 vss 0.0424f
C15499 vdd.n6483 vss 0.0132f
C15500 vdd.n6484 vss 0.00925f
C15501 vdd.n6485 vss 0.00425f
C15502 vdd.n6486 vss 0.00413f
C15503 vdd.n6487 vss 0.00324f
C15504 vdd.n6488 vss 0.0471f
C15505 vdd.t1170 vss 0.0471f
C15506 vdd.n6489 vss 0.00251f
C15507 vdd.n6490 vss 0.0112f
C15508 vdd.n6491 vss 0.0707f
C15509 vdd.n6492 vss 0.0393f
C15510 vdd.n6493 vss 0.0332f
C15511 vdd.n6494 vss 0.0596f
C15512 vdd.n6495 vss 0.00324f
C15513 vdd.n6496 vss 0.0112f
C15514 vdd.n6497 vss 0.0128f
C15515 vdd.n6498 vss 0.00413f
C15516 vdd.n6499 vss 0.00413f
C15517 vdd.n6500 vss 0.0471f
C15518 vdd.n6501 vss 0.00251f
C15519 vdd.t564 vss 0.0471f
C15520 vdd.n6502 vss 0.00324f
C15521 vdd.n6504 vss 0.00679f
C15522 vdd.n6505 vss 0.00413f
C15523 vdd.n6506 vss 0.00324f
C15524 vdd.n6507 vss 0.00413f
C15525 vdd.n6508 vss 0.0471f
C15526 vdd.n6509 vss 0.00324f
C15527 vdd.n6511 vss 0.00925f
C15528 vdd.t314 vss 0.0471f
C15529 vdd.n6512 vss 0.00425f
C15530 vdd.n6513 vss 0.0424f
C15531 vdd.n6514 vss 0.0132f
C15532 vdd.n6515 vss 0.00324f
C15533 vdd.n6516 vss 0.0128f
C15534 vdd.n6517 vss 0.02f
C15535 vdd.n6518 vss 0.00425f
C15536 vdd.n6519 vss 0.00413f
C15537 vdd.n6520 vss 0.00251f
C15538 vdd.t121 vss 0.0471f
C15539 vdd.n6521 vss 0.00251f
C15540 vdd.n6522 vss 0.00517f
C15541 vdd.n6523 vss 0.00679f
C15542 vdd.n6524 vss 0.00517f
C15543 vdd.n6525 vss 0.00679f
C15544 vdd.n6526 vss 0.02f
C15545 vdd.n6527 vss 0.00425f
C15546 vdd.n6528 vss 0.0424f
C15547 vdd.n6529 vss 0.0132f
C15548 vdd.n6530 vss 0.00925f
C15549 vdd.n6531 vss 0.00425f
C15550 vdd.n6532 vss 0.00413f
C15551 vdd.n6533 vss 0.00324f
C15552 vdd.n6534 vss 0.0471f
C15553 vdd.t119 vss 0.0471f
C15554 vdd.n6535 vss 0.00251f
C15555 vdd.n6536 vss 0.0112f
C15556 vdd.n6537 vss 0.0128f
C15557 vdd.t120 vss 0.00134f
C15558 vdd.t565 vss 0.0013f
C15559 vdd.n6538 vss 0.0332f
C15560 vdd.n6539 vss 0.0393f
C15561 vdd.n6540 vss 0.0418f
C15562 vdd.n6541 vss 0.121f
C15563 vdd.n6542 vss 0.291f
C15564 vdd.n6543 vss 0.234f
C15565 vdd.n6544 vss 0.00324f
C15566 vdd.n6545 vss 0.0112f
C15567 vdd.n6546 vss 0.0128f
C15568 vdd.n6547 vss 0.00413f
C15569 vdd.n6548 vss 0.00413f
C15570 vdd.n6549 vss 0.0471f
C15571 vdd.n6550 vss 0.00251f
C15572 vdd.t1186 vss 0.0471f
C15573 vdd.n6551 vss 0.00324f
C15574 vdd.n6553 vss 0.00679f
C15575 vdd.n6554 vss 0.00413f
C15576 vdd.n6555 vss 0.00324f
C15577 vdd.n6556 vss 0.00413f
C15578 vdd.n6557 vss 0.0471f
C15579 vdd.n6558 vss 0.00324f
C15580 vdd.n6560 vss 0.00925f
C15581 vdd.t1243 vss 0.0471f
C15582 vdd.n6561 vss 0.00425f
C15583 vdd.n6562 vss 0.0424f
C15584 vdd.n6563 vss 0.0132f
C15585 vdd.n6564 vss 0.00324f
C15586 vdd.n6565 vss 0.0128f
C15587 vdd.n6566 vss 0.02f
C15588 vdd.n6567 vss 0.00425f
C15589 vdd.n6568 vss 0.00413f
C15590 vdd.n6569 vss 0.00251f
C15591 vdd.t549 vss 0.0471f
C15592 vdd.n6570 vss 0.00251f
C15593 vdd.n6571 vss 0.00517f
C15594 vdd.n6572 vss 0.00679f
C15595 vdd.n6573 vss 0.00517f
C15596 vdd.n6574 vss 0.00679f
C15597 vdd.n6575 vss 0.02f
C15598 vdd.n6576 vss 0.00425f
C15599 vdd.n6577 vss 0.0424f
C15600 vdd.n6578 vss 0.0132f
C15601 vdd.n6579 vss 0.00925f
C15602 vdd.n6580 vss 0.00425f
C15603 vdd.n6581 vss 0.00413f
C15604 vdd.n6582 vss 0.00324f
C15605 vdd.n6583 vss 0.0471f
C15606 vdd.t550 vss 0.0471f
C15607 vdd.n6584 vss 0.00251f
C15608 vdd.n6585 vss 0.0112f
C15609 vdd.n6586 vss 0.0128f
C15610 vdd.n6587 vss 0.159f
C15611 vdd.n6588 vss 0.0393f
C15612 vdd.n6589 vss 0.0332f
C15613 vdd.n6590 vss 0.00324f
C15614 vdd.n6591 vss 0.0112f
C15615 vdd.n6592 vss 0.0128f
C15616 vdd.n6593 vss 0.00413f
C15617 vdd.n6594 vss 0.00413f
C15618 vdd.n6595 vss 0.0471f
C15619 vdd.n6596 vss 0.00251f
C15620 vdd.t28 vss 0.0471f
C15621 vdd.n6597 vss 0.00324f
C15622 vdd.n6599 vss 0.00679f
C15623 vdd.n6600 vss 0.00413f
C15624 vdd.n6601 vss 0.00324f
C15625 vdd.n6602 vss 0.00413f
C15626 vdd.n6603 vss 0.0471f
C15627 vdd.n6604 vss 0.00324f
C15628 vdd.n6606 vss 0.00925f
C15629 vdd.t1095 vss 0.0471f
C15630 vdd.n6607 vss 0.00425f
C15631 vdd.n6608 vss 0.0424f
C15632 vdd.n6609 vss 0.0132f
C15633 vdd.n6610 vss 0.00324f
C15634 vdd.n6611 vss 0.0128f
C15635 vdd.n6612 vss 0.02f
C15636 vdd.n6613 vss 0.00425f
C15637 vdd.n6614 vss 0.00413f
C15638 vdd.n6615 vss 0.00251f
C15639 vdd.t709 vss 0.0471f
C15640 vdd.n6616 vss 0.00251f
C15641 vdd.n6617 vss 0.00517f
C15642 vdd.n6618 vss 0.00679f
C15643 vdd.n6619 vss 0.00517f
C15644 vdd.n6620 vss 0.00679f
C15645 vdd.n6621 vss 0.02f
C15646 vdd.n6622 vss 0.00425f
C15647 vdd.n6623 vss 0.0424f
C15648 vdd.n6624 vss 0.0132f
C15649 vdd.n6625 vss 0.00925f
C15650 vdd.n6626 vss 0.00425f
C15651 vdd.n6627 vss 0.00413f
C15652 vdd.n6628 vss 0.00324f
C15653 vdd.n6629 vss 0.0471f
C15654 vdd.t707 vss 0.0471f
C15655 vdd.n6630 vss 0.00251f
C15656 vdd.n6631 vss 0.0112f
C15657 vdd.n6632 vss 0.0128f
C15658 vdd.n6633 vss 0.214f
C15659 vdd.n6634 vss 0.0393f
C15660 vdd.n6635 vss 0.0332f
C15661 vdd.t705 vss 0.00134f
C15662 vdd.t485 vss 0.0013f
C15663 vdd.n6636 vss 0.0315f
C15664 vdd.n6637 vss 0.0393f
C15665 vdd.n6638 vss 0.00324f
C15666 vdd.n6639 vss 0.0112f
C15667 vdd.n6640 vss 0.0128f
C15668 vdd.n6641 vss 0.00413f
C15669 vdd.t703 vss 0.0471f
C15670 vdd.n6642 vss 0.00324f
C15671 vdd.n6644 vss 0.00925f
C15672 vdd.n6645 vss 0.00413f
C15673 vdd.n6646 vss 0.00679f
C15674 vdd.n6647 vss 0.00413f
C15675 vdd.n6648 vss 0.0471f
C15676 vdd.n6649 vss 0.00324f
C15677 vdd.n6650 vss 0.0471f
C15678 vdd.n6651 vss 0.00324f
C15679 vdd.n6652 vss 0.0424f
C15680 vdd.t484 vss 0.0471f
C15681 vdd.n6654 vss 0.00425f
C15682 vdd.n6655 vss 0.00925f
C15683 vdd.n6656 vss 0.0132f
C15684 vdd.n6657 vss 0.00324f
C15685 vdd.n6658 vss 0.0128f
C15686 vdd.n6659 vss 0.02f
C15687 vdd.n6660 vss 0.00425f
C15688 vdd.n6661 vss 0.00413f
C15689 vdd.n6662 vss 0.00251f
C15690 vdd.t704 vss 0.0471f
C15691 vdd.n6663 vss 0.00251f
C15692 vdd.n6664 vss 0.00517f
C15693 vdd.n6665 vss 0.00679f
C15694 vdd.n6666 vss 0.00324f
C15695 vdd.n6667 vss 0.00679f
C15696 vdd.n6668 vss 0.00517f
C15697 vdd.n6669 vss 0.00251f
C15698 vdd.n6670 vss 0.00413f
C15699 vdd.n6671 vss 0.0471f
C15700 vdd.t1088 vss 0.0471f
C15701 vdd.n6672 vss 0.00425f
C15702 vdd.n6673 vss 0.0424f
C15703 vdd.n6674 vss 0.0132f
C15704 vdd.n6675 vss 0.02f
C15705 vdd.n6676 vss 0.00425f
C15706 vdd.n6677 vss 0.00413f
C15707 vdd.n6678 vss 0.00251f
C15708 vdd.n6679 vss 0.0112f
C15709 vdd.n6680 vss 0.0128f
C15710 vdd.n6681 vss 0.0365f
C15711 vdd.n6682 vss 0.202f
C15712 vdd.n6683 vss 0.00324f
C15713 vdd.n6684 vss 0.0112f
C15714 vdd.n6685 vss 0.0128f
C15715 vdd.n6686 vss 0.00413f
C15716 vdd.n6687 vss 0.00413f
C15717 vdd.n6688 vss 0.0471f
C15718 vdd.n6689 vss 0.00251f
C15719 vdd.t1288 vss 0.0471f
C15720 vdd.n6690 vss 0.00324f
C15721 vdd.n6692 vss 0.00679f
C15722 vdd.n6693 vss 0.00413f
C15723 vdd.n6694 vss 0.00324f
C15724 vdd.n6695 vss 0.00413f
C15725 vdd.n6696 vss 0.0471f
C15726 vdd.n6697 vss 0.00324f
C15727 vdd.n6699 vss 0.00925f
C15728 vdd.t728 vss 0.0471f
C15729 vdd.n6700 vss 0.00425f
C15730 vdd.n6701 vss 0.0424f
C15731 vdd.n6702 vss 0.0132f
C15732 vdd.n6703 vss 0.00324f
C15733 vdd.n6704 vss 0.0128f
C15734 vdd.n6705 vss 0.02f
C15735 vdd.n6706 vss 0.00425f
C15736 vdd.n6707 vss 0.00413f
C15737 vdd.n6708 vss 0.00251f
C15738 vdd.t362 vss 0.0471f
C15739 vdd.n6709 vss 0.00251f
C15740 vdd.n6710 vss 0.00517f
C15741 vdd.n6711 vss 0.00679f
C15742 vdd.n6712 vss 0.00517f
C15743 vdd.n6713 vss 0.00679f
C15744 vdd.n6714 vss 0.02f
C15745 vdd.n6715 vss 0.00425f
C15746 vdd.n6716 vss 0.0424f
C15747 vdd.n6717 vss 0.0132f
C15748 vdd.n6718 vss 0.00925f
C15749 vdd.n6719 vss 0.00425f
C15750 vdd.n6720 vss 0.00413f
C15751 vdd.n6721 vss 0.00324f
C15752 vdd.n6722 vss 0.0471f
C15753 vdd.t363 vss 0.0471f
C15754 vdd.n6723 vss 0.00251f
C15755 vdd.n6724 vss 0.0112f
C15756 vdd.n6725 vss 0.0128f
C15757 vdd.t364 vss 0.00134f
C15758 vdd.t1289 vss 0.0013f
C15759 vdd.n6726 vss 0.0332f
C15760 vdd.n6727 vss 0.0393f
C15761 vdd.n6728 vss 0.0418f
C15762 vdd.n6729 vss 0.00324f
C15763 vdd.n6730 vss 0.0112f
C15764 vdd.n6731 vss 0.0128f
C15765 vdd.n6732 vss 0.00413f
C15766 vdd.n6733 vss 0.00413f
C15767 vdd.n6734 vss 0.0471f
C15768 vdd.n6735 vss 0.00251f
C15769 vdd.t207 vss 0.0471f
C15770 vdd.n6736 vss 0.00324f
C15771 vdd.n6738 vss 0.00679f
C15772 vdd.n6739 vss 0.00413f
C15773 vdd.n6740 vss 0.00324f
C15774 vdd.n6741 vss 0.00413f
C15775 vdd.n6742 vss 0.0471f
C15776 vdd.n6743 vss 0.00324f
C15777 vdd.n6745 vss 0.00925f
C15778 vdd.t235 vss 0.0471f
C15779 vdd.n6746 vss 0.00425f
C15780 vdd.n6747 vss 0.0424f
C15781 vdd.n6748 vss 0.0132f
C15782 vdd.n6749 vss 0.00324f
C15783 vdd.n6750 vss 0.0128f
C15784 vdd.n6751 vss 0.02f
C15785 vdd.n6752 vss 0.00425f
C15786 vdd.n6753 vss 0.00413f
C15787 vdd.n6754 vss 0.00251f
C15788 vdd.t624 vss 0.0471f
C15789 vdd.n6755 vss 0.00251f
C15790 vdd.n6756 vss 0.00517f
C15791 vdd.n6757 vss 0.00679f
C15792 vdd.n6758 vss 0.00517f
C15793 vdd.n6759 vss 0.00679f
C15794 vdd.n6760 vss 0.02f
C15795 vdd.n6761 vss 0.00425f
C15796 vdd.n6762 vss 0.0424f
C15797 vdd.n6763 vss 0.0132f
C15798 vdd.n6764 vss 0.00925f
C15799 vdd.n6765 vss 0.00425f
C15800 vdd.n6766 vss 0.00413f
C15801 vdd.n6767 vss 0.00324f
C15802 vdd.n6768 vss 0.0471f
C15803 vdd.t625 vss 0.0471f
C15804 vdd.n6769 vss 0.00251f
C15805 vdd.n6770 vss 0.0112f
C15806 vdd.n6771 vss 0.0128f
C15807 vdd.t626 vss 0.00134f
C15808 vdd.t208 vss 0.0013f
C15809 vdd.n6772 vss 0.0332f
C15810 vdd.n6773 vss 0.0393f
C15811 vdd.n6774 vss 0.0345f
C15812 vdd.n6775 vss 0.00335f
C15813 vdd.t90 vss 0.0013f
C15814 vdd.n6776 vss 0.0309f
C15815 vdd.n6777 vss 0.00991f
C15816 vdd.n6778 vss 0.0424f
C15817 vdd.n6779 vss 0.00679f
C15818 vdd.n6780 vss 0.00413f
C15819 vdd.n6781 vss 0.0471f
C15820 vdd.n6782 vss 0.00251f
C15821 vdd.n6783 vss 0.00324f
C15822 vdd.n6784 vss 0.0128f
C15823 vdd.n6785 vss 0.00413f
C15824 vdd.n6786 vss 0.00413f
C15825 vdd.n6787 vss 0.0471f
C15826 vdd.n6788 vss 0.00251f
C15827 vdd.n6789 vss 0.00324f
C15828 vdd.n6790 vss 0.00413f
C15829 vdd.n6791 vss 0.00324f
C15830 vdd.n6792 vss 0.0132f
C15831 vdd.n6793 vss 0.0424f
C15832 vdd.n6794 vss 0.00324f
C15833 vdd.n6795 vss 0.00413f
C15834 vdd.n6796 vss 0.02f
C15835 vdd.n6797 vss 0.00425f
C15836 vdd.t1362 vss 0.0471f
C15837 vdd.n6799 vss 0.00425f
C15838 vdd.n6800 vss 0.00925f
C15839 vdd.n6801 vss 0.00679f
C15840 vdd.n6802 vss 0.00517f
C15841 vdd.n6803 vss 0.00679f
C15842 vdd.n6804 vss 0.00517f
C15843 vdd.n6805 vss 0.00251f
C15844 vdd.t691 vss 0.0471f
C15845 vdd.n6806 vss 0.0471f
C15846 vdd.t693 vss 0.0471f
C15847 vdd.n6807 vss 0.00251f
C15848 vdd.n6808 vss 0.0105f
C15849 vdd.t692 vss 0.00134f
C15850 vdd.n6809 vss 0.0393f
C15851 vdd.n6810 vss 0.0633f
C15852 vdd.n6811 vss 0.00805f
C15853 vdd.n6812 vss 0.0112f
C15854 vdd.n6813 vss 0.0128f
C15855 vdd.n6814 vss 0.00324f
C15856 vdd.n6815 vss 0.00324f
C15857 vdd.n6816 vss 0.00413f
C15858 vdd.n6817 vss 0.00425f
C15859 vdd.t89 vss 0.0471f
C15860 vdd.n6819 vss 0.00425f
C15861 vdd.n6820 vss 0.00925f
C15862 vdd.n6821 vss 0.0107f
C15863 vdd.n6822 vss 0.0126f
C15864 vdd.n6823 vss 9.89e-19
C15865 vdd.n6824 vss 0.00163f
C15866 vdd.n6825 vss 0.00145f
C15867 vdd.n6826 vss 0.0271f
C15868 vdd.n6827 vss 0.00324f
C15869 vdd.n6828 vss 0.0112f
C15870 vdd.n6829 vss 0.0128f
C15871 vdd.n6830 vss 0.00413f
C15872 vdd.n6831 vss 0.00413f
C15873 vdd.n6832 vss 0.0471f
C15874 vdd.n6833 vss 0.00251f
C15875 vdd.t1318 vss 0.0471f
C15876 vdd.n6834 vss 0.00324f
C15877 vdd.n6836 vss 0.00679f
C15878 vdd.n6837 vss 0.00413f
C15879 vdd.n6838 vss 0.00324f
C15880 vdd.n6839 vss 0.00413f
C15881 vdd.n6840 vss 0.0471f
C15882 vdd.n6841 vss 0.00324f
C15883 vdd.n6843 vss 0.00925f
C15884 vdd.t155 vss 0.0471f
C15885 vdd.n6844 vss 0.00425f
C15886 vdd.n6845 vss 0.0424f
C15887 vdd.n6846 vss 0.0132f
C15888 vdd.n6847 vss 0.00324f
C15889 vdd.n6848 vss 0.0128f
C15890 vdd.n6849 vss 0.02f
C15891 vdd.n6850 vss 0.00425f
C15892 vdd.n6851 vss 0.00413f
C15893 vdd.n6852 vss 0.00251f
C15894 vdd.t152 vss 0.0471f
C15895 vdd.n6853 vss 0.00251f
C15896 vdd.n6854 vss 0.00517f
C15897 vdd.n6855 vss 0.00679f
C15898 vdd.n6856 vss 0.00517f
C15899 vdd.n6857 vss 0.00679f
C15900 vdd.n6858 vss 0.02f
C15901 vdd.n6859 vss 0.00425f
C15902 vdd.n6860 vss 0.0424f
C15903 vdd.n6861 vss 0.0132f
C15904 vdd.n6862 vss 0.00925f
C15905 vdd.n6863 vss 0.00425f
C15906 vdd.n6864 vss 0.00413f
C15907 vdd.n6865 vss 0.00324f
C15908 vdd.n6866 vss 0.0471f
C15909 vdd.t153 vss 0.0471f
C15910 vdd.n6867 vss 0.00251f
C15911 vdd.n6868 vss 0.0112f
C15912 vdd.n6869 vss 0.0128f
C15913 vdd.t154 vss 0.00134f
C15914 vdd.t1319 vss 0.0013f
C15915 vdd.n6870 vss 0.0332f
C15916 vdd.n6871 vss 0.0393f
C15917 vdd.n6872 vss 0.0418f
C15918 vdd.n6873 vss 0.00324f
C15919 vdd.n6874 vss 0.0112f
C15920 vdd.n6875 vss 0.0128f
C15921 vdd.n6876 vss 0.00413f
C15922 vdd.n6877 vss 0.00413f
C15923 vdd.n6878 vss 0.0471f
C15924 vdd.n6879 vss 0.00251f
C15925 vdd.t205 vss 0.0471f
C15926 vdd.n6880 vss 0.00324f
C15927 vdd.n6882 vss 0.00679f
C15928 vdd.n6883 vss 0.00413f
C15929 vdd.n6884 vss 0.00324f
C15930 vdd.n6885 vss 0.00413f
C15931 vdd.n6886 vss 0.0471f
C15932 vdd.n6887 vss 0.00324f
C15933 vdd.n6889 vss 0.00925f
C15934 vdd.t413 vss 0.0471f
C15935 vdd.n6890 vss 0.00425f
C15936 vdd.n6891 vss 0.0424f
C15937 vdd.n6892 vss 0.0132f
C15938 vdd.n6893 vss 0.00324f
C15939 vdd.n6894 vss 0.0128f
C15940 vdd.n6895 vss 0.02f
C15941 vdd.n6896 vss 0.00425f
C15942 vdd.n6897 vss 0.00413f
C15943 vdd.n6898 vss 0.00251f
C15944 vdd.t217 vss 0.0471f
C15945 vdd.n6899 vss 0.00251f
C15946 vdd.n6900 vss 0.00517f
C15947 vdd.n6901 vss 0.00679f
C15948 vdd.n6902 vss 0.00517f
C15949 vdd.n6903 vss 0.00679f
C15950 vdd.n6904 vss 0.02f
C15951 vdd.n6905 vss 0.00425f
C15952 vdd.n6906 vss 0.0424f
C15953 vdd.n6907 vss 0.0132f
C15954 vdd.n6908 vss 0.00925f
C15955 vdd.n6909 vss 0.00425f
C15956 vdd.n6910 vss 0.00413f
C15957 vdd.n6911 vss 0.00324f
C15958 vdd.n6912 vss 0.0471f
C15959 vdd.t218 vss 0.0471f
C15960 vdd.n6913 vss 0.00251f
C15961 vdd.n6914 vss 0.0112f
C15962 vdd.n6915 vss 0.0128f
C15963 vdd.t219 vss 0.00134f
C15964 vdd.t206 vss 0.0013f
C15965 vdd.n6916 vss 0.0332f
C15966 vdd.n6917 vss 0.0393f
C15967 vdd.n6918 vss 0.0345f
C15968 vdd.n6919 vss 0.00324f
C15969 vdd.n6920 vss 0.0112f
C15970 vdd.n6921 vss 0.0128f
C15971 vdd.n6922 vss 0.00413f
C15972 vdd.n6923 vss 0.00413f
C15973 vdd.n6924 vss 0.0471f
C15974 vdd.n6925 vss 0.00251f
C15975 vdd.t558 vss 0.0471f
C15976 vdd.n6926 vss 0.00324f
C15977 vdd.n6928 vss 0.00679f
C15978 vdd.n6929 vss 0.00413f
C15979 vdd.n6930 vss 0.00324f
C15980 vdd.n6931 vss 0.00413f
C15981 vdd.n6932 vss 0.0471f
C15982 vdd.n6933 vss 0.00324f
C15983 vdd.n6935 vss 0.00925f
C15984 vdd.t983 vss 0.0471f
C15985 vdd.n6936 vss 0.00425f
C15986 vdd.n6937 vss 0.0424f
C15987 vdd.n6938 vss 0.0132f
C15988 vdd.n6939 vss 0.00324f
C15989 vdd.n6940 vss 0.0128f
C15990 vdd.n6941 vss 0.02f
C15991 vdd.n6942 vss 0.00425f
C15992 vdd.n6943 vss 0.00413f
C15993 vdd.n6944 vss 0.00251f
C15994 vdd.t980 vss 0.0471f
C15995 vdd.n6945 vss 0.00251f
C15996 vdd.n6946 vss 0.00517f
C15997 vdd.n6947 vss 0.00679f
C15998 vdd.n6948 vss 0.00517f
C15999 vdd.n6949 vss 0.00679f
C16000 vdd.n6950 vss 0.02f
C16001 vdd.n6951 vss 0.00425f
C16002 vdd.n6952 vss 0.0424f
C16003 vdd.n6953 vss 0.0132f
C16004 vdd.n6954 vss 0.00925f
C16005 vdd.n6955 vss 0.00425f
C16006 vdd.n6956 vss 0.00413f
C16007 vdd.n6957 vss 0.00324f
C16008 vdd.n6958 vss 0.0471f
C16009 vdd.t981 vss 0.0471f
C16010 vdd.n6959 vss 0.00251f
C16011 vdd.n6960 vss 0.0112f
C16012 vdd.n6961 vss 0.0128f
C16013 vdd.t982 vss 0.00134f
C16014 vdd.t559 vss 0.0013f
C16015 vdd.n6962 vss 0.0332f
C16016 vdd.n6963 vss 0.0393f
C16017 vdd.n6964 vss 0.0418f
C16018 vdd.n6965 vss 0.00324f
C16019 vdd.n6966 vss 0.0112f
C16020 vdd.n6967 vss 0.0128f
C16021 vdd.n6968 vss 0.00413f
C16022 vdd.n6969 vss 0.00413f
C16023 vdd.n6970 vss 0.0471f
C16024 vdd.n6971 vss 0.00251f
C16025 vdd.t377 vss 0.0471f
C16026 vdd.n6972 vss 0.00324f
C16027 vdd.n6974 vss 0.00679f
C16028 vdd.n6975 vss 0.00413f
C16029 vdd.n6976 vss 0.00324f
C16030 vdd.n6977 vss 0.00413f
C16031 vdd.n6978 vss 0.0471f
C16032 vdd.n6979 vss 0.00324f
C16033 vdd.n6981 vss 0.00925f
C16034 vdd.t1107 vss 0.0471f
C16035 vdd.n6982 vss 0.00425f
C16036 vdd.n6983 vss 0.0424f
C16037 vdd.n6984 vss 0.0132f
C16038 vdd.n6985 vss 0.00324f
C16039 vdd.n6986 vss 0.0128f
C16040 vdd.n6987 vss 0.02f
C16041 vdd.n6988 vss 0.00425f
C16042 vdd.n6989 vss 0.00413f
C16043 vdd.n6990 vss 0.00251f
C16044 vdd.t806 vss 0.0471f
C16045 vdd.n6991 vss 0.00251f
C16046 vdd.n6992 vss 0.00517f
C16047 vdd.n6993 vss 0.00679f
C16048 vdd.n6994 vss 0.00517f
C16049 vdd.n6995 vss 0.00679f
C16050 vdd.n6996 vss 0.02f
C16051 vdd.n6997 vss 0.00425f
C16052 vdd.n6998 vss 0.0424f
C16053 vdd.n6999 vss 0.0132f
C16054 vdd.n7000 vss 0.00925f
C16055 vdd.n7001 vss 0.00425f
C16056 vdd.n7002 vss 0.00413f
C16057 vdd.n7003 vss 0.00324f
C16058 vdd.n7004 vss 0.0471f
C16059 vdd.t807 vss 0.0471f
C16060 vdd.n7005 vss 0.00251f
C16061 vdd.n7006 vss 0.0112f
C16062 vdd.n7007 vss 0.0128f
C16063 vdd.t808 vss 0.00134f
C16064 vdd.t378 vss 0.0013f
C16065 vdd.n7008 vss 0.0332f
C16066 vdd.n7009 vss 0.0393f
C16067 vdd.n7010 vss 0.0345f
C16068 vdd.n7011 vss 0.00335f
C16069 vdd.t98 vss 0.0013f
C16070 vdd.n7012 vss 0.0309f
C16071 vdd.n7013 vss 0.00991f
C16072 vdd.n7014 vss 0.0424f
C16073 vdd.n7015 vss 0.00679f
C16074 vdd.n7016 vss 0.00413f
C16075 vdd.n7017 vss 0.0471f
C16076 vdd.n7018 vss 0.00251f
C16077 vdd.n7019 vss 0.00324f
C16078 vdd.n7020 vss 0.0128f
C16079 vdd.n7021 vss 0.00413f
C16080 vdd.n7022 vss 0.00413f
C16081 vdd.n7023 vss 0.0471f
C16082 vdd.n7024 vss 0.00251f
C16083 vdd.n7025 vss 0.00324f
C16084 vdd.n7026 vss 0.00413f
C16085 vdd.n7027 vss 0.00324f
C16086 vdd.n7028 vss 0.0132f
C16087 vdd.n7029 vss 0.0424f
C16088 vdd.n7030 vss 0.00324f
C16089 vdd.n7031 vss 0.00413f
C16090 vdd.n7032 vss 0.02f
C16091 vdd.n7033 vss 0.00425f
C16092 vdd.t1089 vss 0.0471f
C16093 vdd.n7035 vss 0.00425f
C16094 vdd.n7036 vss 0.00925f
C16095 vdd.n7037 vss 0.00679f
C16096 vdd.n7038 vss 0.00517f
C16097 vdd.n7039 vss 0.00679f
C16098 vdd.n7040 vss 0.00517f
C16099 vdd.n7041 vss 0.00251f
C16100 vdd.t80 vss 0.0471f
C16101 vdd.n7042 vss 0.0471f
C16102 vdd.t82 vss 0.0471f
C16103 vdd.n7043 vss 0.00251f
C16104 vdd.n7044 vss 0.0105f
C16105 vdd.t81 vss 0.00134f
C16106 vdd.n7045 vss 0.0393f
C16107 vdd.n7046 vss 0.0633f
C16108 vdd.n7047 vss 0.00805f
C16109 vdd.n7048 vss 0.0112f
C16110 vdd.n7049 vss 0.0128f
C16111 vdd.n7050 vss 0.00324f
C16112 vdd.n7051 vss 0.00324f
C16113 vdd.n7052 vss 0.00413f
C16114 vdd.n7053 vss 0.00425f
C16115 vdd.t97 vss 0.0471f
C16116 vdd.n7055 vss 0.00425f
C16117 vdd.n7056 vss 0.00925f
C16118 vdd.n7057 vss 0.0107f
C16119 vdd.n7058 vss 0.0126f
C16120 vdd.n7059 vss 9.89e-19
C16121 vdd.n7060 vss 0.00163f
C16122 vdd.n7061 vss 0.00145f
C16123 vdd.n7062 vss 0.0271f
C16124 vdd.n7063 vss 0.00324f
C16125 vdd.n7064 vss 0.0112f
C16126 vdd.n7065 vss 0.0128f
C16127 vdd.n7066 vss 0.00413f
C16128 vdd.n7067 vss 0.00413f
C16129 vdd.n7068 vss 0.0471f
C16130 vdd.n7069 vss 0.00251f
C16131 vdd.t587 vss 0.0471f
C16132 vdd.n7070 vss 0.00324f
C16133 vdd.n7072 vss 0.00679f
C16134 vdd.n7073 vss 0.00413f
C16135 vdd.n7074 vss 0.00324f
C16136 vdd.n7075 vss 0.00413f
C16137 vdd.n7076 vss 0.0471f
C16138 vdd.n7077 vss 0.00324f
C16139 vdd.n7079 vss 0.00925f
C16140 vdd.t353 vss 0.0471f
C16141 vdd.n7080 vss 0.00425f
C16142 vdd.n7081 vss 0.0424f
C16143 vdd.n7082 vss 0.0132f
C16144 vdd.n7083 vss 0.00324f
C16145 vdd.n7084 vss 0.0128f
C16146 vdd.n7085 vss 0.02f
C16147 vdd.n7086 vss 0.00425f
C16148 vdd.n7087 vss 0.00413f
C16149 vdd.n7088 vss 0.00251f
C16150 vdd.t302 vss 0.0471f
C16151 vdd.n7089 vss 0.00251f
C16152 vdd.n7090 vss 0.00517f
C16153 vdd.n7091 vss 0.00679f
C16154 vdd.n7092 vss 0.00517f
C16155 vdd.n7093 vss 0.00679f
C16156 vdd.n7094 vss 0.02f
C16157 vdd.n7095 vss 0.00425f
C16158 vdd.n7096 vss 0.0424f
C16159 vdd.n7097 vss 0.0132f
C16160 vdd.n7098 vss 0.00925f
C16161 vdd.n7099 vss 0.00425f
C16162 vdd.n7100 vss 0.00413f
C16163 vdd.n7101 vss 0.00324f
C16164 vdd.n7102 vss 0.0471f
C16165 vdd.t303 vss 0.0471f
C16166 vdd.n7103 vss 0.00251f
C16167 vdd.n7104 vss 0.0112f
C16168 vdd.n7105 vss 0.0128f
C16169 vdd.t304 vss 0.00134f
C16170 vdd.t588 vss 0.0013f
C16171 vdd.n7106 vss 0.0332f
C16172 vdd.n7107 vss 0.0393f
C16173 vdd.n7108 vss 0.0418f
C16174 vdd.t522 vss 0.00134f
C16175 vdd.t1464 vss 0.0013f
C16176 vdd.n7109 vss 0.032f
C16177 vdd.n7110 vss 0.0393f
C16178 vdd.n7111 vss 0.00324f
C16179 vdd.n7112 vss 0.0112f
C16180 vdd.n7113 vss 0.0128f
C16181 vdd.n7114 vss 0.00413f
C16182 vdd.t520 vss 0.0471f
C16183 vdd.n7115 vss 0.00324f
C16184 vdd.n7117 vss 0.00925f
C16185 vdd.n7118 vss 0.00413f
C16186 vdd.n7119 vss 0.00679f
C16187 vdd.n7120 vss 0.00413f
C16188 vdd.n7121 vss 0.0471f
C16189 vdd.n7122 vss 0.00324f
C16190 vdd.n7123 vss 0.0471f
C16191 vdd.n7124 vss 0.00324f
C16192 vdd.n7125 vss 0.0424f
C16193 vdd.t1463 vss 0.0471f
C16194 vdd.n7127 vss 0.00425f
C16195 vdd.n7128 vss 0.00925f
C16196 vdd.n7129 vss 0.0132f
C16197 vdd.n7130 vss 0.00324f
C16198 vdd.n7131 vss 0.0128f
C16199 vdd.n7132 vss 0.02f
C16200 vdd.n7133 vss 0.00425f
C16201 vdd.n7134 vss 0.00413f
C16202 vdd.n7135 vss 0.00251f
C16203 vdd.t521 vss 0.0471f
C16204 vdd.n7136 vss 0.00251f
C16205 vdd.n7137 vss 0.00517f
C16206 vdd.n7138 vss 0.00679f
C16207 vdd.n7139 vss 0.00324f
C16208 vdd.n7140 vss 0.00679f
C16209 vdd.n7141 vss 0.00517f
C16210 vdd.n7142 vss 0.00251f
C16211 vdd.n7143 vss 0.00413f
C16212 vdd.n7144 vss 0.0471f
C16213 vdd.t1025 vss 0.0471f
C16214 vdd.n7145 vss 0.00425f
C16215 vdd.n7146 vss 0.0424f
C16216 vdd.n7147 vss 0.0132f
C16217 vdd.n7148 vss 0.02f
C16218 vdd.n7149 vss 0.00425f
C16219 vdd.n7150 vss 0.00413f
C16220 vdd.n7151 vss 0.00251f
C16221 vdd.n7152 vss 0.0112f
C16222 vdd.n7153 vss 0.0128f
C16223 vdd.n7154 vss 0.0418f
C16224 vdd.t184 vss 0.00134f
C16225 vdd.t1311 vss 0.0013f
C16226 vdd.n7155 vss 0.032f
C16227 vdd.n7156 vss 0.0393f
C16228 vdd.n7157 vss 0.00324f
C16229 vdd.n7158 vss 0.0112f
C16230 vdd.n7159 vss 0.0128f
C16231 vdd.n7160 vss 0.00413f
C16232 vdd.t182 vss 0.0471f
C16233 vdd.n7161 vss 0.00324f
C16234 vdd.n7163 vss 0.00925f
C16235 vdd.n7164 vss 0.00413f
C16236 vdd.n7165 vss 0.00679f
C16237 vdd.n7166 vss 0.00413f
C16238 vdd.n7167 vss 0.0471f
C16239 vdd.n7168 vss 0.00324f
C16240 vdd.n7169 vss 0.0471f
C16241 vdd.n7170 vss 0.00324f
C16242 vdd.n7171 vss 0.0424f
C16243 vdd.t1310 vss 0.0471f
C16244 vdd.n7173 vss 0.00425f
C16245 vdd.n7174 vss 0.00925f
C16246 vdd.n7175 vss 0.0132f
C16247 vdd.n7176 vss 0.00324f
C16248 vdd.n7177 vss 0.0128f
C16249 vdd.n7178 vss 0.02f
C16250 vdd.n7179 vss 0.00425f
C16251 vdd.n7180 vss 0.00413f
C16252 vdd.n7181 vss 0.00251f
C16253 vdd.t183 vss 0.0471f
C16254 vdd.n7182 vss 0.00251f
C16255 vdd.n7183 vss 0.00517f
C16256 vdd.n7184 vss 0.00679f
C16257 vdd.n7185 vss 0.00324f
C16258 vdd.n7186 vss 0.00679f
C16259 vdd.n7187 vss 0.00517f
C16260 vdd.n7188 vss 0.00251f
C16261 vdd.n7189 vss 0.00413f
C16262 vdd.n7190 vss 0.0471f
C16263 vdd.t979 vss 0.0471f
C16264 vdd.n7191 vss 0.00425f
C16265 vdd.n7192 vss 0.0424f
C16266 vdd.n7193 vss 0.0132f
C16267 vdd.n7194 vss 0.02f
C16268 vdd.n7195 vss 0.00425f
C16269 vdd.n7196 vss 0.00413f
C16270 vdd.n7197 vss 0.00251f
C16271 vdd.n7198 vss 0.0112f
C16272 vdd.n7199 vss 0.0128f
C16273 vdd.n7200 vss 0.0369f
C16274 vdd.n7201 vss 0.00335f
C16275 vdd.t1460 vss 0.0013f
C16276 vdd.n7202 vss 0.0309f
C16277 vdd.n7203 vss 0.0107f
C16278 vdd.n7204 vss 0.0128f
C16279 vdd.n7205 vss 0.0424f
C16280 vdd.t1459 vss 0.0471f
C16281 vdd.n7206 vss 0.00324f
C16282 vdd.n7207 vss 0.0471f
C16283 vdd.t1394 vss 0.0471f
C16284 vdd.n7208 vss 0.00413f
C16285 vdd.n7209 vss 0.00324f
C16286 vdd.t1395 vss 0.00134f
C16287 vdd.n7210 vss 0.0393f
C16288 vdd.n7211 vss 0.0128f
C16289 vdd.t1393 vss 0.0471f
C16290 vdd.n7212 vss 0.00324f
C16291 vdd.n7214 vss 0.00925f
C16292 vdd.n7215 vss 0.0471f
C16293 vdd.n7216 vss 0.00324f
C16294 vdd.n7217 vss 0.00413f
C16295 vdd.n7218 vss 0.00324f
C16296 vdd.n7219 vss 0.00679f
C16297 vdd.n7221 vss 0.00925f
C16298 vdd.n7222 vss 0.00425f
C16299 vdd.n7223 vss 0.00413f
C16300 vdd.n7224 vss 0.00251f
C16301 vdd.n7225 vss 0.00517f
C16302 vdd.n7226 vss 0.00679f
C16303 vdd.n7227 vss 0.00324f
C16304 vdd.n7228 vss 0.00679f
C16305 vdd.n7229 vss 0.00517f
C16306 vdd.n7230 vss 0.00251f
C16307 vdd.n7231 vss 0.00413f
C16308 vdd.n7232 vss 0.0471f
C16309 vdd.t277 vss 0.0471f
C16310 vdd.n7233 vss 0.00425f
C16311 vdd.n7234 vss 0.0424f
C16312 vdd.n7235 vss 0.0132f
C16313 vdd.n7236 vss 0.02f
C16314 vdd.n7237 vss 0.00425f
C16315 vdd.n7238 vss 0.00413f
C16316 vdd.n7239 vss 0.00251f
C16317 vdd.n7240 vss 0.0105f
C16318 vdd.n7241 vss 0.0633f
C16319 vdd.n7242 vss 0.00805f
C16320 vdd.n7243 vss 0.0112f
C16321 vdd.n7244 vss 0.00251f
C16322 vdd.n7245 vss 0.00413f
C16323 vdd.n7246 vss 0.00425f
C16324 vdd.n7247 vss 0.00991f
C16325 vdd.n7248 vss 0.0126f
C16326 vdd.n7249 vss 9.89e-19
C16327 vdd.n7250 vss 0.0011f
C16328 vdd.n7251 vss 0.0271f
C16329 vdd.t884 vss 0.00134f
C16330 vdd.t1050 vss 0.0013f
C16331 vdd.n7252 vss 0.032f
C16332 vdd.n7253 vss 0.0393f
C16333 vdd.n7254 vss 0.00324f
C16334 vdd.n7255 vss 0.0112f
C16335 vdd.n7256 vss 0.0128f
C16336 vdd.n7257 vss 0.00413f
C16337 vdd.t882 vss 0.0471f
C16338 vdd.n7258 vss 0.00324f
C16339 vdd.n7260 vss 0.00925f
C16340 vdd.n7261 vss 0.00413f
C16341 vdd.n7262 vss 0.00679f
C16342 vdd.n7263 vss 0.00413f
C16343 vdd.n7264 vss 0.0471f
C16344 vdd.n7265 vss 0.00324f
C16345 vdd.n7266 vss 0.0471f
C16346 vdd.n7267 vss 0.00324f
C16347 vdd.n7268 vss 0.0424f
C16348 vdd.t1049 vss 0.0471f
C16349 vdd.n7270 vss 0.00425f
C16350 vdd.n7271 vss 0.00925f
C16351 vdd.n7272 vss 0.0132f
C16352 vdd.n7273 vss 0.00324f
C16353 vdd.n7274 vss 0.0128f
C16354 vdd.n7275 vss 0.02f
C16355 vdd.n7276 vss 0.00425f
C16356 vdd.n7277 vss 0.00413f
C16357 vdd.n7278 vss 0.00251f
C16358 vdd.t883 vss 0.0471f
C16359 vdd.n7279 vss 0.00251f
C16360 vdd.n7280 vss 0.00517f
C16361 vdd.n7281 vss 0.00679f
C16362 vdd.n7282 vss 0.00324f
C16363 vdd.n7283 vss 0.00679f
C16364 vdd.n7284 vss 0.00517f
C16365 vdd.n7285 vss 0.00251f
C16366 vdd.n7286 vss 0.00413f
C16367 vdd.n7287 vss 0.0471f
C16368 vdd.t1285 vss 0.0471f
C16369 vdd.n7288 vss 0.00425f
C16370 vdd.n7289 vss 0.0424f
C16371 vdd.n7290 vss 0.0132f
C16372 vdd.n7291 vss 0.02f
C16373 vdd.n7292 vss 0.00425f
C16374 vdd.n7293 vss 0.00413f
C16375 vdd.n7294 vss 0.00251f
C16376 vdd.n7295 vss 0.0112f
C16377 vdd.n7296 vss 0.0128f
C16378 vdd.n7297 vss 0.0418f
C16379 vdd.t533 vss 0.00134f
C16380 vdd.t1361 vss 0.0013f
C16381 vdd.n7298 vss 0.032f
C16382 vdd.n7299 vss 0.0393f
C16383 vdd.n7300 vss 0.00324f
C16384 vdd.n7301 vss 0.0112f
C16385 vdd.n7302 vss 0.0128f
C16386 vdd.n7303 vss 0.00413f
C16387 vdd.t534 vss 0.0471f
C16388 vdd.n7304 vss 0.00324f
C16389 vdd.n7306 vss 0.00925f
C16390 vdd.n7307 vss 0.00413f
C16391 vdd.n7308 vss 0.00679f
C16392 vdd.n7309 vss 0.00413f
C16393 vdd.n7310 vss 0.0471f
C16394 vdd.n7311 vss 0.00324f
C16395 vdd.n7312 vss 0.0471f
C16396 vdd.n7313 vss 0.00324f
C16397 vdd.n7314 vss 0.0424f
C16398 vdd.t1360 vss 0.0471f
C16399 vdd.n7316 vss 0.00425f
C16400 vdd.n7317 vss 0.00925f
C16401 vdd.n7318 vss 0.0132f
C16402 vdd.n7319 vss 0.00324f
C16403 vdd.n7320 vss 0.0128f
C16404 vdd.n7321 vss 0.02f
C16405 vdd.n7322 vss 0.00425f
C16406 vdd.n7323 vss 0.00413f
C16407 vdd.n7324 vss 0.00251f
C16408 vdd.t532 vss 0.0471f
C16409 vdd.n7325 vss 0.00251f
C16410 vdd.n7326 vss 0.00517f
C16411 vdd.n7327 vss 0.00679f
C16412 vdd.n7328 vss 0.00324f
C16413 vdd.n7329 vss 0.00679f
C16414 vdd.n7330 vss 0.00517f
C16415 vdd.n7331 vss 0.00251f
C16416 vdd.n7332 vss 0.00413f
C16417 vdd.n7333 vss 0.0471f
C16418 vdd.t536 vss 0.0471f
C16419 vdd.n7334 vss 0.00425f
C16420 vdd.n7335 vss 0.0424f
C16421 vdd.n7336 vss 0.0132f
C16422 vdd.n7337 vss 0.02f
C16423 vdd.n7338 vss 0.00425f
C16424 vdd.n7339 vss 0.00413f
C16425 vdd.n7340 vss 0.00251f
C16426 vdd.n7341 vss 0.0112f
C16427 vdd.n7342 vss 0.0128f
C16428 vdd.n7343 vss 0.0365f
C16429 vdd.t1093 vss 0.00134f
C16430 vdd.t594 vss 0.0013f
C16431 vdd.n7344 vss 0.032f
C16432 vdd.n7345 vss 0.0393f
C16433 vdd.n7346 vss 0.00324f
C16434 vdd.n7347 vss 0.0112f
C16435 vdd.n7348 vss 0.0128f
C16436 vdd.n7349 vss 0.00413f
C16437 vdd.t1091 vss 0.0471f
C16438 vdd.n7350 vss 0.00324f
C16439 vdd.n7352 vss 0.00925f
C16440 vdd.n7353 vss 0.00413f
C16441 vdd.n7354 vss 0.00679f
C16442 vdd.n7355 vss 0.00413f
C16443 vdd.n7356 vss 0.0471f
C16444 vdd.n7357 vss 0.00324f
C16445 vdd.n7358 vss 0.0471f
C16446 vdd.n7359 vss 0.00324f
C16447 vdd.n7360 vss 0.0424f
C16448 vdd.t593 vss 0.0471f
C16449 vdd.n7362 vss 0.00425f
C16450 vdd.n7363 vss 0.00925f
C16451 vdd.n7364 vss 0.0132f
C16452 vdd.n7365 vss 0.00324f
C16453 vdd.n7366 vss 0.0128f
C16454 vdd.n7367 vss 0.02f
C16455 vdd.n7368 vss 0.00425f
C16456 vdd.n7369 vss 0.00413f
C16457 vdd.n7370 vss 0.00251f
C16458 vdd.t1092 vss 0.0471f
C16459 vdd.n7371 vss 0.00251f
C16460 vdd.n7372 vss 0.00517f
C16461 vdd.n7373 vss 0.00679f
C16462 vdd.n7374 vss 0.00324f
C16463 vdd.n7375 vss 0.00679f
C16464 vdd.n7376 vss 0.00517f
C16465 vdd.n7377 vss 0.00251f
C16466 vdd.n7378 vss 0.00413f
C16467 vdd.n7379 vss 0.0471f
C16468 vdd.t1094 vss 0.0471f
C16469 vdd.n7380 vss 0.00425f
C16470 vdd.n7381 vss 0.0424f
C16471 vdd.n7382 vss 0.0132f
C16472 vdd.n7383 vss 0.02f
C16473 vdd.n7384 vss 0.00425f
C16474 vdd.n7385 vss 0.00413f
C16475 vdd.n7386 vss 0.00251f
C16476 vdd.n7387 vss 0.0112f
C16477 vdd.n7388 vss 0.0128f
C16478 vdd.n7389 vss 0.0418f
C16479 vdd.t1254 vss 0.00134f
C16480 vdd.t380 vss 0.0013f
C16481 vdd.n7390 vss 0.032f
C16482 vdd.n7391 vss 0.0393f
C16483 vdd.n7392 vss 0.00324f
C16484 vdd.n7393 vss 0.0112f
C16485 vdd.n7394 vss 0.0128f
C16486 vdd.n7395 vss 0.00413f
C16487 vdd.t1252 vss 0.0471f
C16488 vdd.n7396 vss 0.00324f
C16489 vdd.n7398 vss 0.00925f
C16490 vdd.n7399 vss 0.00413f
C16491 vdd.n7400 vss 0.00679f
C16492 vdd.n7401 vss 0.00413f
C16493 vdd.n7402 vss 0.0471f
C16494 vdd.n7403 vss 0.00324f
C16495 vdd.n7404 vss 0.0471f
C16496 vdd.n7405 vss 0.00324f
C16497 vdd.n7406 vss 0.0424f
C16498 vdd.t379 vss 0.0471f
C16499 vdd.n7408 vss 0.00425f
C16500 vdd.n7409 vss 0.00925f
C16501 vdd.n7410 vss 0.0132f
C16502 vdd.n7411 vss 0.00324f
C16503 vdd.n7412 vss 0.0128f
C16504 vdd.n7413 vss 0.02f
C16505 vdd.n7414 vss 0.00425f
C16506 vdd.n7415 vss 0.00413f
C16507 vdd.n7416 vss 0.00251f
C16508 vdd.t1253 vss 0.0471f
C16509 vdd.n7417 vss 0.00251f
C16510 vdd.n7418 vss 0.00517f
C16511 vdd.n7419 vss 0.00679f
C16512 vdd.n7420 vss 0.00324f
C16513 vdd.n7421 vss 0.00679f
C16514 vdd.n7422 vss 0.00517f
C16515 vdd.n7423 vss 0.00251f
C16516 vdd.n7424 vss 0.00413f
C16517 vdd.n7425 vss 0.0471f
C16518 vdd.t1255 vss 0.0471f
C16519 vdd.n7426 vss 0.00425f
C16520 vdd.n7427 vss 0.0424f
C16521 vdd.n7428 vss 0.0132f
C16522 vdd.n7429 vss 0.02f
C16523 vdd.n7430 vss 0.00425f
C16524 vdd.n7431 vss 0.00413f
C16525 vdd.n7432 vss 0.00251f
C16526 vdd.n7433 vss 0.0112f
C16527 vdd.n7434 vss 0.0128f
C16528 vdd.n7435 vss 0.0369f
C16529 vdd.n7436 vss 0.00335f
C16530 vdd.t1155 vss 0.0013f
C16531 vdd.n7437 vss 0.0309f
C16532 vdd.n7438 vss 0.0107f
C16533 vdd.n7439 vss 0.0128f
C16534 vdd.n7440 vss 0.0424f
C16535 vdd.t1154 vss 0.0471f
C16536 vdd.n7441 vss 0.00324f
C16537 vdd.n7442 vss 0.0471f
C16538 vdd.t443 vss 0.0471f
C16539 vdd.n7443 vss 0.00413f
C16540 vdd.n7444 vss 0.00324f
C16541 vdd.t444 vss 0.00134f
C16542 vdd.n7445 vss 0.0393f
C16543 vdd.n7446 vss 0.0128f
C16544 vdd.t442 vss 0.0471f
C16545 vdd.n7447 vss 0.00324f
C16546 vdd.n7449 vss 0.00925f
C16547 vdd.n7450 vss 0.0471f
C16548 vdd.n7451 vss 0.00324f
C16549 vdd.n7452 vss 0.00413f
C16550 vdd.n7453 vss 0.00324f
C16551 vdd.n7454 vss 0.00679f
C16552 vdd.n7456 vss 0.00925f
C16553 vdd.n7457 vss 0.00425f
C16554 vdd.n7458 vss 0.00413f
C16555 vdd.n7459 vss 0.00251f
C16556 vdd.n7460 vss 0.00517f
C16557 vdd.n7461 vss 0.00679f
C16558 vdd.n7462 vss 0.00324f
C16559 vdd.n7463 vss 0.00679f
C16560 vdd.n7464 vss 0.00517f
C16561 vdd.n7465 vss 0.00251f
C16562 vdd.n7466 vss 0.00413f
C16563 vdd.n7467 vss 0.0471f
C16564 vdd.t892 vss 0.0471f
C16565 vdd.n7468 vss 0.00425f
C16566 vdd.n7469 vss 0.0424f
C16567 vdd.n7470 vss 0.0132f
C16568 vdd.n7471 vss 0.02f
C16569 vdd.n7472 vss 0.00425f
C16570 vdd.n7473 vss 0.00413f
C16571 vdd.n7474 vss 0.00251f
C16572 vdd.n7475 vss 0.0105f
C16573 vdd.n7476 vss 0.0633f
C16574 vdd.n7477 vss 0.00805f
C16575 vdd.n7478 vss 0.0112f
C16576 vdd.n7479 vss 0.00251f
C16577 vdd.n7480 vss 0.00413f
C16578 vdd.n7481 vss 0.00425f
C16579 vdd.n7482 vss 0.00991f
C16580 vdd.n7483 vss 0.0126f
C16581 vdd.n7484 vss 9.89e-19
C16582 vdd.n7485 vss 0.0011f
C16583 vdd.n7486 vss 0.0271f
C16584 vdd.t932 vss 0.00134f
C16585 vdd.t1327 vss 0.0013f
C16586 vdd.n7487 vss 0.032f
C16587 vdd.n7488 vss 0.0393f
C16588 vdd.n7489 vss 0.00324f
C16589 vdd.n7490 vss 0.0112f
C16590 vdd.n7491 vss 0.0128f
C16591 vdd.n7492 vss 0.00413f
C16592 vdd.t930 vss 0.0471f
C16593 vdd.n7493 vss 0.00324f
C16594 vdd.n7495 vss 0.00925f
C16595 vdd.n7496 vss 0.00413f
C16596 vdd.n7497 vss 0.00679f
C16597 vdd.n7498 vss 0.00413f
C16598 vdd.n7499 vss 0.0471f
C16599 vdd.n7500 vss 0.00324f
C16600 vdd.n7501 vss 0.0471f
C16601 vdd.n7502 vss 0.00324f
C16602 vdd.n7503 vss 0.0424f
C16603 vdd.t1326 vss 0.0471f
C16604 vdd.n7505 vss 0.00425f
C16605 vdd.n7506 vss 0.00925f
C16606 vdd.n7507 vss 0.0132f
C16607 vdd.n7508 vss 0.00324f
C16608 vdd.n7509 vss 0.0128f
C16609 vdd.n7510 vss 0.02f
C16610 vdd.n7511 vss 0.00425f
C16611 vdd.n7512 vss 0.00413f
C16612 vdd.n7513 vss 0.00251f
C16613 vdd.t931 vss 0.0471f
C16614 vdd.n7514 vss 0.00251f
C16615 vdd.n7515 vss 0.00517f
C16616 vdd.n7516 vss 0.00679f
C16617 vdd.n7517 vss 0.00324f
C16618 vdd.n7518 vss 0.00679f
C16619 vdd.n7519 vss 0.00517f
C16620 vdd.n7520 vss 0.00251f
C16621 vdd.n7521 vss 0.00413f
C16622 vdd.n7522 vss 0.0471f
C16623 vdd.t143 vss 0.0471f
C16624 vdd.n7523 vss 0.00425f
C16625 vdd.n7524 vss 0.0424f
C16626 vdd.n7525 vss 0.0132f
C16627 vdd.n7526 vss 0.02f
C16628 vdd.n7527 vss 0.00425f
C16629 vdd.n7528 vss 0.00413f
C16630 vdd.n7529 vss 0.00251f
C16631 vdd.n7530 vss 0.0112f
C16632 vdd.n7531 vss 0.0128f
C16633 vdd.n7532 vss 0.0418f
C16634 vdd.t899 vss 0.0013f
C16635 vdd.t1274 vss 0.00134f
C16636 vdd.n7533 vss 0.00324f
C16637 vdd.n7534 vss 0.0112f
C16638 vdd.n7535 vss 0.0128f
C16639 vdd.n7536 vss 0.00413f
C16640 vdd.t1272 vss 0.0471f
C16641 vdd.n7537 vss 0.00324f
C16642 vdd.n7539 vss 0.00925f
C16643 vdd.n7540 vss 0.00413f
C16644 vdd.n7541 vss 0.00679f
C16645 vdd.n7542 vss 0.00413f
C16646 vdd.n7543 vss 0.0471f
C16647 vdd.n7544 vss 0.00324f
C16648 vdd.n7545 vss 0.0471f
C16649 vdd.n7546 vss 0.00324f
C16650 vdd.n7547 vss 0.0424f
C16651 vdd.t898 vss 0.0471f
C16652 vdd.n7549 vss 0.00425f
C16653 vdd.n7550 vss 0.00925f
C16654 vdd.n7551 vss 0.0132f
C16655 vdd.n7552 vss 0.00324f
C16656 vdd.n7553 vss 0.0128f
C16657 vdd.n7554 vss 0.02f
C16658 vdd.n7555 vss 0.00425f
C16659 vdd.n7556 vss 0.00413f
C16660 vdd.n7557 vss 0.00251f
C16661 vdd.t1273 vss 0.0471f
C16662 vdd.n7558 vss 0.00251f
C16663 vdd.n7559 vss 0.00517f
C16664 vdd.n7560 vss 0.00679f
C16665 vdd.n7561 vss 0.00324f
C16666 vdd.n7562 vss 0.00679f
C16667 vdd.n7563 vss 0.00517f
C16668 vdd.n7564 vss 0.00251f
C16669 vdd.n7565 vss 0.00413f
C16670 vdd.n7566 vss 0.0471f
C16671 vdd.t1263 vss 0.0471f
C16672 vdd.n7567 vss 0.00425f
C16673 vdd.n7568 vss 0.0424f
C16674 vdd.n7569 vss 0.0132f
C16675 vdd.n7570 vss 0.02f
C16676 vdd.n7571 vss 0.00425f
C16677 vdd.n7572 vss 0.00413f
C16678 vdd.n7573 vss 0.00251f
C16679 vdd.n7574 vss 0.0112f
C16680 vdd.n7575 vss 0.0128f
C16681 vdd.t887 vss 0.00134f
C16682 vdd.t167 vss 0.0013f
C16683 vdd.n7576 vss 0.032f
C16684 vdd.n7577 vss 0.0393f
C16685 vdd.n7578 vss 0.00324f
C16686 vdd.n7579 vss 0.0112f
C16687 vdd.n7580 vss 0.0128f
C16688 vdd.n7581 vss 0.00413f
C16689 vdd.t885 vss 0.0471f
C16690 vdd.n7582 vss 0.00324f
C16691 vdd.n7584 vss 0.00925f
C16692 vdd.n7585 vss 0.00413f
C16693 vdd.n7586 vss 0.00679f
C16694 vdd.n7587 vss 0.00413f
C16695 vdd.n7588 vss 0.0471f
C16696 vdd.n7589 vss 0.00324f
C16697 vdd.n7590 vss 0.0471f
C16698 vdd.n7591 vss 0.00324f
C16699 vdd.n7592 vss 0.0424f
C16700 vdd.t166 vss 0.0471f
C16701 vdd.n7594 vss 0.00425f
C16702 vdd.n7595 vss 0.00925f
C16703 vdd.n7596 vss 0.0132f
C16704 vdd.n7597 vss 0.00324f
C16705 vdd.n7598 vss 0.0128f
C16706 vdd.n7599 vss 0.02f
C16707 vdd.n7600 vss 0.00425f
C16708 vdd.n7601 vss 0.00413f
C16709 vdd.n7602 vss 0.00251f
C16710 vdd.t886 vss 0.0471f
C16711 vdd.n7603 vss 0.00251f
C16712 vdd.n7604 vss 0.00517f
C16713 vdd.n7605 vss 0.00679f
C16714 vdd.n7606 vss 0.00324f
C16715 vdd.n7607 vss 0.00679f
C16716 vdd.n7608 vss 0.00517f
C16717 vdd.n7609 vss 0.00251f
C16718 vdd.n7610 vss 0.00413f
C16719 vdd.n7611 vss 0.0471f
C16720 vdd.t809 vss 0.0471f
C16721 vdd.n7612 vss 0.00425f
C16722 vdd.n7613 vss 0.0424f
C16723 vdd.n7614 vss 0.0132f
C16724 vdd.n7615 vss 0.02f
C16725 vdd.n7616 vss 0.00425f
C16726 vdd.n7617 vss 0.00413f
C16727 vdd.n7618 vss 0.00251f
C16728 vdd.n7619 vss 0.0112f
C16729 vdd.n7620 vss 0.0128f
C16730 vdd.n7621 vss 0.119f
C16731 vdd.n7622 vss 0.118f
C16732 vdd.n7623 vss 0.0393f
C16733 vdd.n7624 vss 0.032f
C16734 vdd.n7625 vss 0.0608f
C16735 vdd.t224 vss 0.00134f
C16736 vdd.t590 vss 0.0013f
C16737 vdd.n7626 vss 0.032f
C16738 vdd.n7627 vss 0.0393f
C16739 vdd.n7628 vss 0.00324f
C16740 vdd.n7629 vss 0.0112f
C16741 vdd.n7630 vss 0.0128f
C16742 vdd.n7631 vss 0.00413f
C16743 vdd.t225 vss 0.0471f
C16744 vdd.n7632 vss 0.00324f
C16745 vdd.n7634 vss 0.00925f
C16746 vdd.n7635 vss 0.00413f
C16747 vdd.n7636 vss 0.00679f
C16748 vdd.n7637 vss 0.00413f
C16749 vdd.n7638 vss 0.0471f
C16750 vdd.n7639 vss 0.00324f
C16751 vdd.n7640 vss 0.0471f
C16752 vdd.n7641 vss 0.00324f
C16753 vdd.n7642 vss 0.0424f
C16754 vdd.t589 vss 0.0471f
C16755 vdd.n7644 vss 0.00425f
C16756 vdd.n7645 vss 0.00925f
C16757 vdd.n7646 vss 0.0132f
C16758 vdd.n7647 vss 0.00324f
C16759 vdd.n7648 vss 0.0128f
C16760 vdd.n7649 vss 0.02f
C16761 vdd.n7650 vss 0.00425f
C16762 vdd.n7651 vss 0.00413f
C16763 vdd.n7652 vss 0.00251f
C16764 vdd.t223 vss 0.0471f
C16765 vdd.n7653 vss 0.00251f
C16766 vdd.n7654 vss 0.00517f
C16767 vdd.n7655 vss 0.00679f
C16768 vdd.n7656 vss 0.00324f
C16769 vdd.n7657 vss 0.00679f
C16770 vdd.n7658 vss 0.00517f
C16771 vdd.n7659 vss 0.00251f
C16772 vdd.n7660 vss 0.00413f
C16773 vdd.n7661 vss 0.0471f
C16774 vdd.t1226 vss 0.0471f
C16775 vdd.n7662 vss 0.00425f
C16776 vdd.n7663 vss 0.0424f
C16777 vdd.n7664 vss 0.0132f
C16778 vdd.n7665 vss 0.02f
C16779 vdd.n7666 vss 0.00425f
C16780 vdd.n7667 vss 0.00413f
C16781 vdd.n7668 vss 0.00251f
C16782 vdd.n7669 vss 0.0112f
C16783 vdd.n7670 vss 0.0128f
C16784 vdd.n7671 vss 0.0418f
C16785 vdd.n7672 vss 0.118f
C16786 vdd.n7673 vss 0.121f
C16787 vdd.t863 vss 0.0013f
C16788 vdd.t252 vss 0.00134f
C16789 vdd.n7674 vss 0.00324f
C16790 vdd.n7675 vss 0.0112f
C16791 vdd.n7676 vss 0.0128f
C16792 vdd.n7677 vss 0.00413f
C16793 vdd.t250 vss 0.0471f
C16794 vdd.n7678 vss 0.00324f
C16795 vdd.n7680 vss 0.00925f
C16796 vdd.n7681 vss 0.00413f
C16797 vdd.n7682 vss 0.00679f
C16798 vdd.n7683 vss 0.00413f
C16799 vdd.n7684 vss 0.0471f
C16800 vdd.n7685 vss 0.00324f
C16801 vdd.n7686 vss 0.0471f
C16802 vdd.n7687 vss 0.00324f
C16803 vdd.n7688 vss 0.0424f
C16804 vdd.t862 vss 0.0471f
C16805 vdd.n7690 vss 0.00425f
C16806 vdd.n7691 vss 0.00925f
C16807 vdd.n7692 vss 0.0132f
C16808 vdd.n7693 vss 0.00324f
C16809 vdd.n7694 vss 0.0128f
C16810 vdd.n7695 vss 0.02f
C16811 vdd.n7696 vss 0.00425f
C16812 vdd.n7697 vss 0.00413f
C16813 vdd.n7698 vss 0.00251f
C16814 vdd.t251 vss 0.0471f
C16815 vdd.n7699 vss 0.00251f
C16816 vdd.n7700 vss 0.00517f
C16817 vdd.n7701 vss 0.00679f
C16818 vdd.n7702 vss 0.00324f
C16819 vdd.n7703 vss 0.00679f
C16820 vdd.n7704 vss 0.00517f
C16821 vdd.n7705 vss 0.00251f
C16822 vdd.n7706 vss 0.00413f
C16823 vdd.n7707 vss 0.0471f
C16824 vdd.t874 vss 0.0471f
C16825 vdd.n7708 vss 0.00425f
C16826 vdd.n7709 vss 0.0424f
C16827 vdd.n7710 vss 0.0132f
C16828 vdd.n7711 vss 0.02f
C16829 vdd.n7712 vss 0.00425f
C16830 vdd.n7713 vss 0.00413f
C16831 vdd.n7714 vss 0.00251f
C16832 vdd.n7715 vss 0.0112f
C16833 vdd.n7716 vss 0.0707f
C16834 vdd.n7717 vss 0.0393f
C16835 vdd.n7718 vss 0.032f
C16836 vdd.n7719 vss 0.0608f
C16837 vdd.t1266 vss 0.00134f
C16838 vdd.t1343 vss 0.0013f
C16839 vdd.n7720 vss 0.032f
C16840 vdd.n7721 vss 0.0393f
C16841 vdd.n7722 vss 0.00324f
C16842 vdd.n7723 vss 0.0112f
C16843 vdd.n7724 vss 0.0128f
C16844 vdd.n7725 vss 0.00413f
C16845 vdd.t1264 vss 0.0471f
C16846 vdd.n7726 vss 0.00324f
C16847 vdd.n7728 vss 0.00925f
C16848 vdd.n7729 vss 0.00413f
C16849 vdd.n7730 vss 0.00679f
C16850 vdd.n7731 vss 0.00413f
C16851 vdd.n7732 vss 0.0471f
C16852 vdd.n7733 vss 0.00324f
C16853 vdd.n7734 vss 0.0471f
C16854 vdd.n7735 vss 0.00324f
C16855 vdd.n7736 vss 0.0424f
C16856 vdd.t1342 vss 0.0471f
C16857 vdd.n7738 vss 0.00425f
C16858 vdd.n7739 vss 0.00925f
C16859 vdd.n7740 vss 0.0132f
C16860 vdd.n7741 vss 0.00324f
C16861 vdd.n7742 vss 0.0128f
C16862 vdd.n7743 vss 0.02f
C16863 vdd.n7744 vss 0.00425f
C16864 vdd.n7745 vss 0.00413f
C16865 vdd.n7746 vss 0.00251f
C16866 vdd.t1265 vss 0.0471f
C16867 vdd.n7747 vss 0.00251f
C16868 vdd.n7748 vss 0.00517f
C16869 vdd.n7749 vss 0.00679f
C16870 vdd.n7750 vss 0.00324f
C16871 vdd.n7751 vss 0.00679f
C16872 vdd.n7752 vss 0.00517f
C16873 vdd.n7753 vss 0.00251f
C16874 vdd.n7754 vss 0.00413f
C16875 vdd.n7755 vss 0.0471f
C16876 vdd.t1078 vss 0.0471f
C16877 vdd.n7756 vss 0.00425f
C16878 vdd.n7757 vss 0.0424f
C16879 vdd.n7758 vss 0.0132f
C16880 vdd.n7759 vss 0.02f
C16881 vdd.n7760 vss 0.00425f
C16882 vdd.n7761 vss 0.00413f
C16883 vdd.n7762 vss 0.00251f
C16884 vdd.n7763 vss 0.0112f
C16885 vdd.n7764 vss 0.0128f
C16886 vdd.n7765 vss 0.0418f
C16887 vdd.n7766 vss 0.0912f
C16888 vdd.n7767 vss 0.0824f
C16889 vdd.n7768 vss 0.0567f
C16890 vdd.t897 vss 0.0013f
C16891 vdd.t519 vss 0.00134f
C16892 vdd.n7769 vss 0.00324f
C16893 vdd.n7770 vss 0.0112f
C16894 vdd.n7771 vss 0.0128f
C16895 vdd.n7772 vss 0.00413f
C16896 vdd.t517 vss 0.0471f
C16897 vdd.n7773 vss 0.00324f
C16898 vdd.n7775 vss 0.00925f
C16899 vdd.n7776 vss 0.00413f
C16900 vdd.n7777 vss 0.00679f
C16901 vdd.n7778 vss 0.00413f
C16902 vdd.n7779 vss 0.0471f
C16903 vdd.n7780 vss 0.00324f
C16904 vdd.n7781 vss 0.0471f
C16905 vdd.n7782 vss 0.00324f
C16906 vdd.n7783 vss 0.0424f
C16907 vdd.t896 vss 0.0471f
C16908 vdd.n7785 vss 0.00425f
C16909 vdd.n7786 vss 0.00925f
C16910 vdd.n7787 vss 0.0132f
C16911 vdd.n7788 vss 0.00324f
C16912 vdd.n7789 vss 0.0128f
C16913 vdd.n7790 vss 0.02f
C16914 vdd.n7791 vss 0.00425f
C16915 vdd.n7792 vss 0.00413f
C16916 vdd.n7793 vss 0.00251f
C16917 vdd.t518 vss 0.0471f
C16918 vdd.n7794 vss 0.00251f
C16919 vdd.n7795 vss 0.00517f
C16920 vdd.n7796 vss 0.00679f
C16921 vdd.n7797 vss 0.00324f
C16922 vdd.n7798 vss 0.00679f
C16923 vdd.n7799 vss 0.00517f
C16924 vdd.n7800 vss 0.00251f
C16925 vdd.n7801 vss 0.00413f
C16926 vdd.n7802 vss 0.0471f
C16927 vdd.t1506 vss 0.0471f
C16928 vdd.n7803 vss 0.00425f
C16929 vdd.n7804 vss 0.0424f
C16930 vdd.n7805 vss 0.0132f
C16931 vdd.n7806 vss 0.02f
C16932 vdd.n7807 vss 0.00425f
C16933 vdd.n7808 vss 0.00413f
C16934 vdd.n7809 vss 0.00251f
C16935 vdd.n7810 vss 0.0112f
C16936 vdd.n7811 vss 0.0128f
C16937 vdd.t240 vss 0.00134f
C16938 vdd.t838 vss 0.0013f
C16939 vdd.n7812 vss 0.032f
C16940 vdd.n7813 vss 0.0393f
C16941 vdd.n7814 vss 0.00324f
C16942 vdd.n7815 vss 0.0112f
C16943 vdd.n7816 vss 0.0128f
C16944 vdd.n7817 vss 0.00413f
C16945 vdd.t238 vss 0.0471f
C16946 vdd.n7818 vss 0.00324f
C16947 vdd.n7820 vss 0.00925f
C16948 vdd.n7821 vss 0.00413f
C16949 vdd.n7822 vss 0.00679f
C16950 vdd.n7823 vss 0.00413f
C16951 vdd.n7824 vss 0.0471f
C16952 vdd.n7825 vss 0.00324f
C16953 vdd.n7826 vss 0.0471f
C16954 vdd.n7827 vss 0.00324f
C16955 vdd.n7828 vss 0.0424f
C16956 vdd.t837 vss 0.0471f
C16957 vdd.n7830 vss 0.00425f
C16958 vdd.n7831 vss 0.00925f
C16959 vdd.n7832 vss 0.0132f
C16960 vdd.n7833 vss 0.00324f
C16961 vdd.n7834 vss 0.0128f
C16962 vdd.n7835 vss 0.02f
C16963 vdd.n7836 vss 0.00425f
C16964 vdd.n7837 vss 0.00413f
C16965 vdd.n7838 vss 0.00251f
C16966 vdd.t239 vss 0.0471f
C16967 vdd.n7839 vss 0.00251f
C16968 vdd.n7840 vss 0.00517f
C16969 vdd.n7841 vss 0.00679f
C16970 vdd.n7842 vss 0.00324f
C16971 vdd.n7843 vss 0.00679f
C16972 vdd.n7844 vss 0.00517f
C16973 vdd.n7845 vss 0.00251f
C16974 vdd.n7846 vss 0.00413f
C16975 vdd.n7847 vss 0.0471f
C16976 vdd.t241 vss 0.0471f
C16977 vdd.n7848 vss 0.00425f
C16978 vdd.n7849 vss 0.0424f
C16979 vdd.n7850 vss 0.0132f
C16980 vdd.n7851 vss 0.02f
C16981 vdd.n7852 vss 0.00425f
C16982 vdd.n7853 vss 0.00413f
C16983 vdd.n7854 vss 0.00251f
C16984 vdd.n7855 vss 0.0112f
C16985 vdd.n7856 vss 0.0128f
C16986 vdd.n7857 vss 0.0316f
C16987 vdd.t542 vss 0.00134f
C16988 vdd.t1376 vss 0.0013f
C16989 vdd.n7858 vss 0.032f
C16990 vdd.n7859 vss 0.0393f
C16991 vdd.n7860 vss 0.00324f
C16992 vdd.n7861 vss 0.0112f
C16993 vdd.n7862 vss 0.0128f
C16994 vdd.n7863 vss 0.00413f
C16995 vdd.t540 vss 0.0471f
C16996 vdd.n7864 vss 0.00324f
C16997 vdd.n7866 vss 0.00925f
C16998 vdd.n7867 vss 0.00413f
C16999 vdd.n7868 vss 0.00679f
C17000 vdd.n7869 vss 0.00413f
C17001 vdd.n7870 vss 0.0471f
C17002 vdd.n7871 vss 0.00324f
C17003 vdd.n7872 vss 0.0471f
C17004 vdd.n7873 vss 0.00324f
C17005 vdd.n7874 vss 0.0424f
C17006 vdd.t1375 vss 0.0471f
C17007 vdd.n7876 vss 0.00425f
C17008 vdd.n7877 vss 0.00925f
C17009 vdd.n7878 vss 0.0132f
C17010 vdd.n7879 vss 0.00324f
C17011 vdd.n7880 vss 0.0128f
C17012 vdd.n7881 vss 0.02f
C17013 vdd.n7882 vss 0.00425f
C17014 vdd.n7883 vss 0.00413f
C17015 vdd.n7884 vss 0.00251f
C17016 vdd.t541 vss 0.0471f
C17017 vdd.n7885 vss 0.00251f
C17018 vdd.n7886 vss 0.00517f
C17019 vdd.n7887 vss 0.00679f
C17020 vdd.n7888 vss 0.00324f
C17021 vdd.n7889 vss 0.00679f
C17022 vdd.n7890 vss 0.00517f
C17023 vdd.n7891 vss 0.00251f
C17024 vdd.n7892 vss 0.00413f
C17025 vdd.n7893 vss 0.0471f
C17026 vdd.t543 vss 0.0471f
C17027 vdd.n7894 vss 0.00425f
C17028 vdd.n7895 vss 0.0424f
C17029 vdd.n7896 vss 0.0132f
C17030 vdd.n7897 vss 0.02f
C17031 vdd.n7898 vss 0.00425f
C17032 vdd.n7899 vss 0.00413f
C17033 vdd.n7900 vss 0.00251f
C17034 vdd.n7901 vss 0.0112f
C17035 vdd.n7902 vss 0.0128f
C17036 vdd.n7903 vss 0.158f
C17037 vdd.n7904 vss 0.256f
C17038 vdd.n7905 vss 0.0953f
C17039 vdd.n7906 vss 0.0393f
C17040 vdd.n7907 vss 0.032f
C17041 vdd.n7908 vss 0.0608f
C17042 vdd.t69 vss 0.00134f
C17043 vdd.t487 vss 0.0013f
C17044 vdd.n7909 vss 0.032f
C17045 vdd.n7910 vss 0.0393f
C17046 vdd.n7911 vss 0.00324f
C17047 vdd.n7912 vss 0.0112f
C17048 vdd.n7913 vss 0.0128f
C17049 vdd.n7914 vss 0.00413f
C17050 vdd.t67 vss 0.0471f
C17051 vdd.n7915 vss 0.00324f
C17052 vdd.n7917 vss 0.00925f
C17053 vdd.n7918 vss 0.00413f
C17054 vdd.n7919 vss 0.00679f
C17055 vdd.n7920 vss 0.00413f
C17056 vdd.n7921 vss 0.0471f
C17057 vdd.n7922 vss 0.00324f
C17058 vdd.n7923 vss 0.0471f
C17059 vdd.n7924 vss 0.00324f
C17060 vdd.n7925 vss 0.0424f
C17061 vdd.t486 vss 0.0471f
C17062 vdd.n7927 vss 0.00425f
C17063 vdd.n7928 vss 0.00925f
C17064 vdd.n7929 vss 0.0132f
C17065 vdd.n7930 vss 0.00324f
C17066 vdd.n7931 vss 0.0128f
C17067 vdd.n7932 vss 0.02f
C17068 vdd.n7933 vss 0.00425f
C17069 vdd.n7934 vss 0.00413f
C17070 vdd.n7935 vss 0.00251f
C17071 vdd.t68 vss 0.0471f
C17072 vdd.n7936 vss 0.00251f
C17073 vdd.n7937 vss 0.00517f
C17074 vdd.n7938 vss 0.00679f
C17075 vdd.n7939 vss 0.00324f
C17076 vdd.n7940 vss 0.00679f
C17077 vdd.n7941 vss 0.00517f
C17078 vdd.n7942 vss 0.00251f
C17079 vdd.n7943 vss 0.00413f
C17080 vdd.n7944 vss 0.0471f
C17081 vdd.t306 vss 0.0471f
C17082 vdd.n7945 vss 0.00425f
C17083 vdd.n7946 vss 0.0424f
C17084 vdd.n7947 vss 0.0132f
C17085 vdd.n7948 vss 0.02f
C17086 vdd.n7949 vss 0.00425f
C17087 vdd.n7950 vss 0.00413f
C17088 vdd.n7951 vss 0.00251f
C17089 vdd.n7952 vss 0.0112f
C17090 vdd.n7953 vss 0.0128f
C17091 vdd.n7954 vss 0.0418f
C17092 vdd.n7955 vss 0.118f
C17093 vdd.n7956 vss 0.121f
C17094 vdd.t873 vss 0.0013f
C17095 vdd.t320 vss 0.00134f
C17096 vdd.n7957 vss 0.00324f
C17097 vdd.n7958 vss 0.0112f
C17098 vdd.n7959 vss 0.0128f
C17099 vdd.n7960 vss 0.00413f
C17100 vdd.t318 vss 0.0471f
C17101 vdd.n7961 vss 0.00324f
C17102 vdd.n7963 vss 0.00925f
C17103 vdd.n7964 vss 0.00413f
C17104 vdd.n7965 vss 0.00679f
C17105 vdd.n7966 vss 0.00413f
C17106 vdd.n7967 vss 0.0471f
C17107 vdd.n7968 vss 0.00324f
C17108 vdd.n7969 vss 0.0471f
C17109 vdd.n7970 vss 0.00324f
C17110 vdd.n7971 vss 0.0424f
C17111 vdd.t872 vss 0.0471f
C17112 vdd.n7973 vss 0.00425f
C17113 vdd.n7974 vss 0.00925f
C17114 vdd.n7975 vss 0.0132f
C17115 vdd.n7976 vss 0.00324f
C17116 vdd.n7977 vss 0.0128f
C17117 vdd.n7978 vss 0.02f
C17118 vdd.n7979 vss 0.00425f
C17119 vdd.n7980 vss 0.00413f
C17120 vdd.n7981 vss 0.00251f
C17121 vdd.t319 vss 0.0471f
C17122 vdd.n7982 vss 0.00251f
C17123 vdd.n7983 vss 0.00517f
C17124 vdd.n7984 vss 0.00679f
C17125 vdd.n7985 vss 0.00324f
C17126 vdd.n7986 vss 0.00679f
C17127 vdd.n7987 vss 0.00517f
C17128 vdd.n7988 vss 0.00251f
C17129 vdd.n7989 vss 0.00413f
C17130 vdd.n7990 vss 0.0471f
C17131 vdd.t620 vss 0.0471f
C17132 vdd.n7991 vss 0.00425f
C17133 vdd.n7992 vss 0.0424f
C17134 vdd.n7993 vss 0.0132f
C17135 vdd.n7994 vss 0.02f
C17136 vdd.n7995 vss 0.00425f
C17137 vdd.n7996 vss 0.00413f
C17138 vdd.n7997 vss 0.00251f
C17139 vdd.n7998 vss 0.0112f
C17140 vdd.n7999 vss 0.0707f
C17141 vdd.n8000 vss 0.0393f
C17142 vdd.n8001 vss 0.032f
C17143 vdd.n8002 vss 0.0608f
C17144 vdd.t963 vss 0.00134f
C17145 vdd.t1331 vss 0.0013f
C17146 vdd.n8003 vss 0.032f
C17147 vdd.n8004 vss 0.0393f
C17148 vdd.n8005 vss 0.00324f
C17149 vdd.n8006 vss 0.0112f
C17150 vdd.n8007 vss 0.0128f
C17151 vdd.n8008 vss 0.00413f
C17152 vdd.t961 vss 0.0471f
C17153 vdd.n8009 vss 0.00324f
C17154 vdd.n8011 vss 0.00925f
C17155 vdd.n8012 vss 0.00413f
C17156 vdd.n8013 vss 0.00679f
C17157 vdd.n8014 vss 0.00413f
C17158 vdd.n8015 vss 0.0471f
C17159 vdd.n8016 vss 0.00324f
C17160 vdd.n8017 vss 0.0471f
C17161 vdd.n8018 vss 0.00324f
C17162 vdd.n8019 vss 0.0424f
C17163 vdd.t1330 vss 0.0471f
C17164 vdd.n8021 vss 0.00425f
C17165 vdd.n8022 vss 0.00925f
C17166 vdd.n8023 vss 0.0132f
C17167 vdd.n8024 vss 0.00324f
C17168 vdd.n8025 vss 0.0128f
C17169 vdd.n8026 vss 0.02f
C17170 vdd.n8027 vss 0.00425f
C17171 vdd.n8028 vss 0.00413f
C17172 vdd.n8029 vss 0.00251f
C17173 vdd.t962 vss 0.0471f
C17174 vdd.n8030 vss 0.00251f
C17175 vdd.n8031 vss 0.00517f
C17176 vdd.n8032 vss 0.00679f
C17177 vdd.n8033 vss 0.00324f
C17178 vdd.n8034 vss 0.00679f
C17179 vdd.n8035 vss 0.00517f
C17180 vdd.n8036 vss 0.00251f
C17181 vdd.n8037 vss 0.00413f
C17182 vdd.n8038 vss 0.0471f
C17183 vdd.t978 vss 0.0471f
C17184 vdd.n8039 vss 0.00425f
C17185 vdd.n8040 vss 0.0424f
C17186 vdd.n8041 vss 0.0132f
C17187 vdd.n8042 vss 0.02f
C17188 vdd.n8043 vss 0.00425f
C17189 vdd.n8044 vss 0.00413f
C17190 vdd.n8045 vss 0.00251f
C17191 vdd.n8046 vss 0.0112f
C17192 vdd.n8047 vss 0.0128f
C17193 vdd.n8048 vss 0.0418f
C17194 vdd.n8049 vss 0.118f
C17195 vdd.n8050 vss 0.0935f
C17196 vdd.t37 vss 0.0013f
C17197 vdd.t644 vss 0.00134f
C17198 vdd.n8051 vss 0.00324f
C17199 vdd.n8052 vss 0.0112f
C17200 vdd.n8053 vss 0.0128f
C17201 vdd.n8054 vss 0.00413f
C17202 vdd.t642 vss 0.0471f
C17203 vdd.n8055 vss 0.00324f
C17204 vdd.n8057 vss 0.00925f
C17205 vdd.n8058 vss 0.00413f
C17206 vdd.n8059 vss 0.00679f
C17207 vdd.n8060 vss 0.00413f
C17208 vdd.n8061 vss 0.0471f
C17209 vdd.n8062 vss 0.00324f
C17210 vdd.n8063 vss 0.0471f
C17211 vdd.n8064 vss 0.00324f
C17212 vdd.n8065 vss 0.0424f
C17213 vdd.t36 vss 0.0471f
C17214 vdd.n8067 vss 0.00425f
C17215 vdd.n8068 vss 0.00925f
C17216 vdd.n8069 vss 0.0132f
C17217 vdd.n8070 vss 0.00324f
C17218 vdd.n8071 vss 0.0128f
C17219 vdd.n8072 vss 0.02f
C17220 vdd.n8073 vss 0.00425f
C17221 vdd.n8074 vss 0.00413f
C17222 vdd.n8075 vss 0.00251f
C17223 vdd.t643 vss 0.0471f
C17224 vdd.n8076 vss 0.00251f
C17225 vdd.n8077 vss 0.00517f
C17226 vdd.n8078 vss 0.00679f
C17227 vdd.n8079 vss 0.00324f
C17228 vdd.n8080 vss 0.00679f
C17229 vdd.n8081 vss 0.00517f
C17230 vdd.n8082 vss 0.00251f
C17231 vdd.n8083 vss 0.00413f
C17232 vdd.n8084 vss 0.0471f
C17233 vdd.t22 vss 0.0471f
C17234 vdd.n8085 vss 0.00425f
C17235 vdd.n8086 vss 0.0424f
C17236 vdd.n8087 vss 0.0132f
C17237 vdd.n8088 vss 0.02f
C17238 vdd.n8089 vss 0.00425f
C17239 vdd.n8090 vss 0.00413f
C17240 vdd.n8091 vss 0.00251f
C17241 vdd.n8092 vss 0.0112f
C17242 vdd.n8093 vss 0.0128f
C17243 vdd.t131 vss 0.00134f
C17244 vdd.t836 vss 0.0013f
C17245 vdd.n8094 vss 0.032f
C17246 vdd.n8095 vss 0.0393f
C17247 vdd.n8096 vss 0.00324f
C17248 vdd.n8097 vss 0.0112f
C17249 vdd.n8098 vss 0.0128f
C17250 vdd.n8099 vss 0.00413f
C17251 vdd.t129 vss 0.0471f
C17252 vdd.n8100 vss 0.00324f
C17253 vdd.n8102 vss 0.00925f
C17254 vdd.n8103 vss 0.00413f
C17255 vdd.n8104 vss 0.00679f
C17256 vdd.n8105 vss 0.00413f
C17257 vdd.n8106 vss 0.0471f
C17258 vdd.n8107 vss 0.00324f
C17259 vdd.n8108 vss 0.0471f
C17260 vdd.n8109 vss 0.00324f
C17261 vdd.n8110 vss 0.0424f
C17262 vdd.t835 vss 0.0471f
C17263 vdd.n8112 vss 0.00425f
C17264 vdd.n8113 vss 0.00925f
C17265 vdd.n8114 vss 0.0132f
C17266 vdd.n8115 vss 0.00324f
C17267 vdd.n8116 vss 0.0128f
C17268 vdd.n8117 vss 0.02f
C17269 vdd.n8118 vss 0.00425f
C17270 vdd.n8119 vss 0.00413f
C17271 vdd.n8120 vss 0.00251f
C17272 vdd.t130 vss 0.0471f
C17273 vdd.n8121 vss 0.00251f
C17274 vdd.n8122 vss 0.00517f
C17275 vdd.n8123 vss 0.00679f
C17276 vdd.n8124 vss 0.00324f
C17277 vdd.n8125 vss 0.00679f
C17278 vdd.n8126 vss 0.00517f
C17279 vdd.n8127 vss 0.00251f
C17280 vdd.n8128 vss 0.00413f
C17281 vdd.n8129 vss 0.0471f
C17282 vdd.t335 vss 0.0471f
C17283 vdd.n8130 vss 0.00425f
C17284 vdd.n8131 vss 0.0424f
C17285 vdd.n8132 vss 0.0132f
C17286 vdd.n8133 vss 0.02f
C17287 vdd.n8134 vss 0.00425f
C17288 vdd.n8135 vss 0.00413f
C17289 vdd.n8136 vss 0.00251f
C17290 vdd.n8137 vss 0.0112f
C17291 vdd.n8138 vss 0.0128f
C17292 vdd.n8139 vss 0.119f
C17293 vdd.n8140 vss 0.118f
C17294 vdd.n8141 vss 0.0393f
C17295 vdd.n8142 vss 0.032f
C17296 vdd.n8143 vss 0.0608f
C17297 vdd.t326 vss 0.00134f
C17298 vdd.t202 vss 0.0013f
C17299 vdd.n8144 vss 0.032f
C17300 vdd.n8145 vss 0.0393f
C17301 vdd.n8146 vss 0.00324f
C17302 vdd.n8147 vss 0.0112f
C17303 vdd.n8148 vss 0.0128f
C17304 vdd.n8149 vss 0.00413f
C17305 vdd.t324 vss 0.0471f
C17306 vdd.n8150 vss 0.00324f
C17307 vdd.n8152 vss 0.00925f
C17308 vdd.n8153 vss 0.00413f
C17309 vdd.n8154 vss 0.00679f
C17310 vdd.n8155 vss 0.00413f
C17311 vdd.n8156 vss 0.0471f
C17312 vdd.n8157 vss 0.00324f
C17313 vdd.n8158 vss 0.0471f
C17314 vdd.n8159 vss 0.00324f
C17315 vdd.n8160 vss 0.0424f
C17316 vdd.t201 vss 0.0471f
C17317 vdd.n8162 vss 0.00425f
C17318 vdd.n8163 vss 0.00925f
C17319 vdd.n8164 vss 0.0132f
C17320 vdd.n8165 vss 0.00324f
C17321 vdd.n8166 vss 0.0128f
C17322 vdd.n8167 vss 0.02f
C17323 vdd.n8168 vss 0.00425f
C17324 vdd.n8169 vss 0.00413f
C17325 vdd.n8170 vss 0.00251f
C17326 vdd.t325 vss 0.0471f
C17327 vdd.n8171 vss 0.00251f
C17328 vdd.n8172 vss 0.00517f
C17329 vdd.n8173 vss 0.00679f
C17330 vdd.n8174 vss 0.00324f
C17331 vdd.n8175 vss 0.00679f
C17332 vdd.n8176 vss 0.00517f
C17333 vdd.n8177 vss 0.00251f
C17334 vdd.n8178 vss 0.00413f
C17335 vdd.n8179 vss 0.0471f
C17336 vdd.t70 vss 0.0471f
C17337 vdd.n8180 vss 0.00425f
C17338 vdd.n8181 vss 0.0424f
C17339 vdd.n8182 vss 0.0132f
C17340 vdd.n8183 vss 0.02f
C17341 vdd.n8184 vss 0.00425f
C17342 vdd.n8185 vss 0.00413f
C17343 vdd.n8186 vss 0.00251f
C17344 vdd.n8187 vss 0.0112f
C17345 vdd.n8188 vss 0.0128f
C17346 vdd.n8189 vss 0.0418f
C17347 vdd.n8190 vss 0.118f
C17348 vdd.n8191 vss 0.121f
C17349 vdd.t974 vss 0.0013f
C17350 vdd.t249 vss 0.00134f
C17351 vdd.n8192 vss 0.00324f
C17352 vdd.n8193 vss 0.0112f
C17353 vdd.n8194 vss 0.0128f
C17354 vdd.n8195 vss 0.00413f
C17355 vdd.t247 vss 0.0471f
C17356 vdd.n8196 vss 0.00324f
C17357 vdd.n8198 vss 0.00925f
C17358 vdd.n8199 vss 0.00413f
C17359 vdd.n8200 vss 0.00679f
C17360 vdd.n8201 vss 0.00413f
C17361 vdd.n8202 vss 0.0471f
C17362 vdd.n8203 vss 0.00324f
C17363 vdd.n8204 vss 0.0471f
C17364 vdd.n8205 vss 0.00324f
C17365 vdd.n8206 vss 0.0424f
C17366 vdd.t973 vss 0.0471f
C17367 vdd.n8208 vss 0.00425f
C17368 vdd.n8209 vss 0.00925f
C17369 vdd.n8210 vss 0.0132f
C17370 vdd.n8211 vss 0.00324f
C17371 vdd.n8212 vss 0.0128f
C17372 vdd.n8213 vss 0.02f
C17373 vdd.n8214 vss 0.00425f
C17374 vdd.n8215 vss 0.00413f
C17375 vdd.n8216 vss 0.00251f
C17376 vdd.t248 vss 0.0471f
C17377 vdd.n8217 vss 0.00251f
C17378 vdd.n8218 vss 0.00517f
C17379 vdd.n8219 vss 0.00679f
C17380 vdd.n8220 vss 0.00324f
C17381 vdd.n8221 vss 0.00679f
C17382 vdd.n8222 vss 0.00517f
C17383 vdd.n8223 vss 0.00251f
C17384 vdd.n8224 vss 0.00413f
C17385 vdd.n8225 vss 0.0471f
C17386 vdd.t1442 vss 0.0471f
C17387 vdd.n8226 vss 0.00425f
C17388 vdd.n8227 vss 0.0424f
C17389 vdd.n8228 vss 0.0132f
C17390 vdd.n8229 vss 0.02f
C17391 vdd.n8230 vss 0.00425f
C17392 vdd.n8231 vss 0.00413f
C17393 vdd.n8232 vss 0.00251f
C17394 vdd.n8233 vss 0.0112f
C17395 vdd.n8234 vss 0.0707f
C17396 vdd.n8235 vss 0.0393f
C17397 vdd.n8236 vss 0.032f
C17398 vdd.n8237 vss 0.0608f
C17399 vdd.t1449 vss 0.00134f
C17400 vdd.t1347 vss 0.0013f
C17401 vdd.n8238 vss 0.032f
C17402 vdd.n8239 vss 0.0393f
C17403 vdd.n8240 vss 0.00324f
C17404 vdd.n8241 vss 0.0112f
C17405 vdd.n8242 vss 0.0128f
C17406 vdd.n8243 vss 0.00413f
C17407 vdd.t1450 vss 0.0471f
C17408 vdd.n8244 vss 0.00324f
C17409 vdd.n8246 vss 0.00925f
C17410 vdd.n8247 vss 0.00413f
C17411 vdd.n8248 vss 0.00679f
C17412 vdd.n8249 vss 0.00413f
C17413 vdd.n8250 vss 0.0471f
C17414 vdd.n8251 vss 0.00324f
C17415 vdd.n8252 vss 0.0471f
C17416 vdd.n8253 vss 0.00324f
C17417 vdd.n8254 vss 0.0424f
C17418 vdd.t1346 vss 0.0471f
C17419 vdd.n8256 vss 0.00425f
C17420 vdd.n8257 vss 0.00925f
C17421 vdd.n8258 vss 0.0132f
C17422 vdd.n8259 vss 0.00324f
C17423 vdd.n8260 vss 0.0128f
C17424 vdd.n8261 vss 0.02f
C17425 vdd.n8262 vss 0.00425f
C17426 vdd.n8263 vss 0.00413f
C17427 vdd.n8264 vss 0.00251f
C17428 vdd.t1448 vss 0.0471f
C17429 vdd.n8265 vss 0.00251f
C17430 vdd.n8266 vss 0.00517f
C17431 vdd.n8267 vss 0.00679f
C17432 vdd.n8268 vss 0.00324f
C17433 vdd.n8269 vss 0.00679f
C17434 vdd.n8270 vss 0.00517f
C17435 vdd.n8271 vss 0.00251f
C17436 vdd.n8272 vss 0.00413f
C17437 vdd.n8273 vss 0.0471f
C17438 vdd.t743 vss 0.0471f
C17439 vdd.n8274 vss 0.00425f
C17440 vdd.n8275 vss 0.0424f
C17441 vdd.n8276 vss 0.0132f
C17442 vdd.n8277 vss 0.02f
C17443 vdd.n8278 vss 0.00425f
C17444 vdd.n8279 vss 0.00413f
C17445 vdd.n8280 vss 0.00251f
C17446 vdd.n8281 vss 0.0112f
C17447 vdd.n8282 vss 0.0128f
C17448 vdd.n8283 vss 0.0418f
C17449 vdd.n8284 vss 0.0912f
C17450 vdd.n8285 vss 0.0824f
C17451 vdd.n8286 vss 0.0567f
C17452 vdd.t855 vss 0.0013f
C17453 vdd.t1177 vss 0.00134f
C17454 vdd.n8287 vss 0.00324f
C17455 vdd.n8288 vss 0.0112f
C17456 vdd.n8289 vss 0.0128f
C17457 vdd.n8290 vss 0.00413f
C17458 vdd.t1175 vss 0.0471f
C17459 vdd.n8291 vss 0.00324f
C17460 vdd.n8293 vss 0.00925f
C17461 vdd.n8294 vss 0.00413f
C17462 vdd.n8295 vss 0.00679f
C17463 vdd.n8296 vss 0.00413f
C17464 vdd.n8297 vss 0.0471f
C17465 vdd.n8298 vss 0.00324f
C17466 vdd.n8299 vss 0.0471f
C17467 vdd.n8300 vss 0.00324f
C17468 vdd.n8301 vss 0.0424f
C17469 vdd.t854 vss 0.0471f
C17470 vdd.n8303 vss 0.00425f
C17471 vdd.n8304 vss 0.00925f
C17472 vdd.n8305 vss 0.0132f
C17473 vdd.n8306 vss 0.00324f
C17474 vdd.n8307 vss 0.0128f
C17475 vdd.n8308 vss 0.02f
C17476 vdd.n8309 vss 0.00425f
C17477 vdd.n8310 vss 0.00413f
C17478 vdd.n8311 vss 0.00251f
C17479 vdd.t1176 vss 0.0471f
C17480 vdd.n8312 vss 0.00251f
C17481 vdd.n8313 vss 0.00517f
C17482 vdd.n8314 vss 0.00679f
C17483 vdd.n8315 vss 0.00324f
C17484 vdd.n8316 vss 0.00679f
C17485 vdd.n8317 vss 0.00517f
C17486 vdd.n8318 vss 0.00251f
C17487 vdd.n8319 vss 0.00413f
C17488 vdd.n8320 vss 0.0471f
C17489 vdd.t1112 vss 0.0471f
C17490 vdd.n8321 vss 0.00425f
C17491 vdd.n8322 vss 0.0424f
C17492 vdd.n8323 vss 0.0132f
C17493 vdd.n8324 vss 0.02f
C17494 vdd.n8325 vss 0.00425f
C17495 vdd.n8326 vss 0.00413f
C17496 vdd.n8327 vss 0.00251f
C17497 vdd.n8328 vss 0.0112f
C17498 vdd.n8329 vss 0.0128f
C17499 vdd.t451 vss 0.00134f
C17500 vdd.t57 vss 0.0013f
C17501 vdd.n8330 vss 0.032f
C17502 vdd.n8331 vss 0.0393f
C17503 vdd.n8332 vss 0.00324f
C17504 vdd.n8333 vss 0.0112f
C17505 vdd.n8334 vss 0.0128f
C17506 vdd.n8335 vss 0.00413f
C17507 vdd.t449 vss 0.0471f
C17508 vdd.n8336 vss 0.00324f
C17509 vdd.n8338 vss 0.00925f
C17510 vdd.n8339 vss 0.00413f
C17511 vdd.n8340 vss 0.00679f
C17512 vdd.n8341 vss 0.00413f
C17513 vdd.n8342 vss 0.0471f
C17514 vdd.n8343 vss 0.00324f
C17515 vdd.n8344 vss 0.0471f
C17516 vdd.n8345 vss 0.00324f
C17517 vdd.n8346 vss 0.0424f
C17518 vdd.t56 vss 0.0471f
C17519 vdd.n8348 vss 0.00425f
C17520 vdd.n8349 vss 0.00925f
C17521 vdd.n8350 vss 0.0132f
C17522 vdd.n8351 vss 0.00324f
C17523 vdd.n8352 vss 0.0128f
C17524 vdd.n8353 vss 0.02f
C17525 vdd.n8354 vss 0.00425f
C17526 vdd.n8355 vss 0.00413f
C17527 vdd.n8356 vss 0.00251f
C17528 vdd.t450 vss 0.0471f
C17529 vdd.n8357 vss 0.00251f
C17530 vdd.n8358 vss 0.00517f
C17531 vdd.n8359 vss 0.00679f
C17532 vdd.n8360 vss 0.00324f
C17533 vdd.n8361 vss 0.00679f
C17534 vdd.n8362 vss 0.00517f
C17535 vdd.n8363 vss 0.00251f
C17536 vdd.n8364 vss 0.00413f
C17537 vdd.n8365 vss 0.0471f
C17538 vdd.t343 vss 0.0471f
C17539 vdd.n8366 vss 0.00425f
C17540 vdd.n8367 vss 0.0424f
C17541 vdd.n8368 vss 0.0132f
C17542 vdd.n8369 vss 0.02f
C17543 vdd.n8370 vss 0.00425f
C17544 vdd.n8371 vss 0.00413f
C17545 vdd.n8372 vss 0.00251f
C17546 vdd.n8373 vss 0.0112f
C17547 vdd.n8374 vss 0.0128f
C17548 vdd.n8375 vss 0.119f
C17549 vdd.n8376 vss 0.118f
C17550 vdd.n8377 vss 0.0393f
C17551 vdd.n8378 vss 0.032f
C17552 vdd.n8379 vss 0.0608f
C17553 vdd.t880 vss 0.00134f
C17554 vdd.t10 vss 0.0013f
C17555 vdd.n8380 vss 0.032f
C17556 vdd.n8381 vss 0.0393f
C17557 vdd.n8382 vss 0.00324f
C17558 vdd.n8383 vss 0.0112f
C17559 vdd.n8384 vss 0.0128f
C17560 vdd.n8385 vss 0.00413f
C17561 vdd.t878 vss 0.0471f
C17562 vdd.n8386 vss 0.00324f
C17563 vdd.n8388 vss 0.00925f
C17564 vdd.n8389 vss 0.00413f
C17565 vdd.n8390 vss 0.00679f
C17566 vdd.n8391 vss 0.00413f
C17567 vdd.n8392 vss 0.0471f
C17568 vdd.n8393 vss 0.00324f
C17569 vdd.n8394 vss 0.0471f
C17570 vdd.n8395 vss 0.00324f
C17571 vdd.n8396 vss 0.0424f
C17572 vdd.t9 vss 0.0471f
C17573 vdd.n8398 vss 0.00425f
C17574 vdd.n8399 vss 0.00925f
C17575 vdd.n8400 vss 0.0132f
C17576 vdd.n8401 vss 0.00324f
C17577 vdd.n8402 vss 0.0128f
C17578 vdd.n8403 vss 0.02f
C17579 vdd.n8404 vss 0.00425f
C17580 vdd.n8405 vss 0.00413f
C17581 vdd.n8406 vss 0.00251f
C17582 vdd.t879 vss 0.0471f
C17583 vdd.n8407 vss 0.00251f
C17584 vdd.n8408 vss 0.00517f
C17585 vdd.n8409 vss 0.00679f
C17586 vdd.n8410 vss 0.00324f
C17587 vdd.n8411 vss 0.00679f
C17588 vdd.n8412 vss 0.00517f
C17589 vdd.n8413 vss 0.00251f
C17590 vdd.n8414 vss 0.00413f
C17591 vdd.n8415 vss 0.0471f
C17592 vdd.t881 vss 0.0471f
C17593 vdd.n8416 vss 0.00425f
C17594 vdd.n8417 vss 0.0424f
C17595 vdd.n8418 vss 0.0132f
C17596 vdd.n8419 vss 0.02f
C17597 vdd.n8420 vss 0.00425f
C17598 vdd.n8421 vss 0.00413f
C17599 vdd.n8422 vss 0.00251f
C17600 vdd.n8423 vss 0.0112f
C17601 vdd.n8424 vss 0.0128f
C17602 vdd.n8425 vss 0.0418f
C17603 vdd.n8426 vss 0.118f
C17604 vdd.n8427 vss 0.121f
C17605 vdd.t41 vss 0.0013f
C17606 vdd.t1421 vss 0.00134f
C17607 vdd.n8428 vss 0.00324f
C17608 vdd.n8429 vss 0.0112f
C17609 vdd.n8430 vss 0.0128f
C17610 vdd.n8431 vss 0.00413f
C17611 vdd.t1419 vss 0.0471f
C17612 vdd.n8432 vss 0.00324f
C17613 vdd.n8434 vss 0.00925f
C17614 vdd.n8435 vss 0.00413f
C17615 vdd.n8436 vss 0.00679f
C17616 vdd.n8437 vss 0.00413f
C17617 vdd.n8438 vss 0.0471f
C17618 vdd.n8439 vss 0.00324f
C17619 vdd.n8440 vss 0.0471f
C17620 vdd.n8441 vss 0.00324f
C17621 vdd.n8442 vss 0.0424f
C17622 vdd.t40 vss 0.0471f
C17623 vdd.n8444 vss 0.00425f
C17624 vdd.n8445 vss 0.00925f
C17625 vdd.n8446 vss 0.0132f
C17626 vdd.n8447 vss 0.00324f
C17627 vdd.n8448 vss 0.0128f
C17628 vdd.n8449 vss 0.02f
C17629 vdd.n8450 vss 0.00425f
C17630 vdd.n8451 vss 0.00413f
C17631 vdd.n8452 vss 0.00251f
C17632 vdd.t1420 vss 0.0471f
C17633 vdd.n8453 vss 0.00251f
C17634 vdd.n8454 vss 0.00517f
C17635 vdd.n8455 vss 0.00679f
C17636 vdd.n8456 vss 0.00324f
C17637 vdd.n8457 vss 0.00679f
C17638 vdd.n8458 vss 0.00517f
C17639 vdd.n8459 vss 0.00251f
C17640 vdd.n8460 vss 0.00413f
C17641 vdd.n8461 vss 0.0471f
C17642 vdd.t1149 vss 0.0471f
C17643 vdd.n8462 vss 0.00425f
C17644 vdd.n8463 vss 0.0424f
C17645 vdd.n8464 vss 0.0132f
C17646 vdd.n8465 vss 0.02f
C17647 vdd.n8466 vss 0.00425f
C17648 vdd.n8467 vss 0.00413f
C17649 vdd.n8468 vss 0.00251f
C17650 vdd.n8469 vss 0.0112f
C17651 vdd.n8470 vss 0.0707f
C17652 vdd.n8471 vss 0.0393f
C17653 vdd.n8472 vss 0.032f
C17654 vdd.n8473 vss 0.0608f
C17655 vdd.t1065 vss 0.00134f
C17656 vdd.t212 vss 0.0013f
C17657 vdd.n8474 vss 0.032f
C17658 vdd.n8475 vss 0.0393f
C17659 vdd.n8476 vss 0.00324f
C17660 vdd.n8477 vss 0.0112f
C17661 vdd.n8478 vss 0.0128f
C17662 vdd.n8479 vss 0.00413f
C17663 vdd.t1063 vss 0.0471f
C17664 vdd.n8480 vss 0.00324f
C17665 vdd.n8482 vss 0.00925f
C17666 vdd.n8483 vss 0.00413f
C17667 vdd.n8484 vss 0.00679f
C17668 vdd.n8485 vss 0.00413f
C17669 vdd.n8486 vss 0.0471f
C17670 vdd.n8487 vss 0.00324f
C17671 vdd.n8488 vss 0.0471f
C17672 vdd.n8489 vss 0.00324f
C17673 vdd.n8490 vss 0.0424f
C17674 vdd.t211 vss 0.0471f
C17675 vdd.n8492 vss 0.00425f
C17676 vdd.n8493 vss 0.00925f
C17677 vdd.n8494 vss 0.0132f
C17678 vdd.n8495 vss 0.00324f
C17679 vdd.n8496 vss 0.0128f
C17680 vdd.n8497 vss 0.02f
C17681 vdd.n8498 vss 0.00425f
C17682 vdd.n8499 vss 0.00413f
C17683 vdd.n8500 vss 0.00251f
C17684 vdd.t1064 vss 0.0471f
C17685 vdd.n8501 vss 0.00251f
C17686 vdd.n8502 vss 0.00517f
C17687 vdd.n8503 vss 0.00679f
C17688 vdd.n8504 vss 0.00324f
C17689 vdd.n8505 vss 0.00679f
C17690 vdd.n8506 vss 0.00517f
C17691 vdd.n8507 vss 0.00251f
C17692 vdd.n8508 vss 0.00413f
C17693 vdd.n8509 vss 0.0471f
C17694 vdd.t1066 vss 0.0471f
C17695 vdd.n8510 vss 0.00425f
C17696 vdd.n8511 vss 0.0424f
C17697 vdd.n8512 vss 0.0132f
C17698 vdd.n8513 vss 0.02f
C17699 vdd.n8514 vss 0.00425f
C17700 vdd.n8515 vss 0.00413f
C17701 vdd.n8516 vss 0.00251f
C17702 vdd.n8517 vss 0.0112f
C17703 vdd.n8518 vss 0.0128f
C17704 vdd.n8519 vss 0.0418f
C17705 vdd.n8520 vss 0.299f
C17706 vdd.n8521 vss 0.00324f
C17707 vdd.n8522 vss 0.0112f
C17708 vdd.n8523 vss 0.0128f
C17709 vdd.n8524 vss 0.00413f
C17710 vdd.n8525 vss 0.00413f
C17711 vdd.n8526 vss 0.0471f
C17712 vdd.n8527 vss 0.00251f
C17713 vdd.t482 vss 0.0471f
C17714 vdd.n8528 vss 0.00324f
C17715 vdd.n8530 vss 0.00679f
C17716 vdd.n8531 vss 0.00413f
C17717 vdd.n8532 vss 0.00324f
C17718 vdd.n8533 vss 0.00413f
C17719 vdd.n8534 vss 0.0471f
C17720 vdd.n8535 vss 0.00324f
C17721 vdd.n8537 vss 0.00925f
C17722 vdd.t634 vss 0.0471f
C17723 vdd.n8538 vss 0.00425f
C17724 vdd.n8539 vss 0.0424f
C17725 vdd.n8540 vss 0.0132f
C17726 vdd.n8541 vss 0.00324f
C17727 vdd.n8542 vss 0.0128f
C17728 vdd.n8543 vss 0.02f
C17729 vdd.n8544 vss 0.00425f
C17730 vdd.n8545 vss 0.00413f
C17731 vdd.n8546 vss 0.00251f
C17732 vdd.t1451 vss 0.0471f
C17733 vdd.n8547 vss 0.00251f
C17734 vdd.n8548 vss 0.00517f
C17735 vdd.n8549 vss 0.00679f
C17736 vdd.n8550 vss 0.00517f
C17737 vdd.n8551 vss 0.00679f
C17738 vdd.n8552 vss 0.02f
C17739 vdd.n8553 vss 0.00425f
C17740 vdd.n8554 vss 0.0424f
C17741 vdd.n8555 vss 0.0132f
C17742 vdd.n8556 vss 0.00925f
C17743 vdd.n8557 vss 0.00425f
C17744 vdd.n8558 vss 0.00413f
C17745 vdd.n8559 vss 0.00324f
C17746 vdd.n8560 vss 0.0471f
C17747 vdd.t1452 vss 0.0471f
C17748 vdd.n8561 vss 0.00251f
C17749 vdd.n8562 vss 0.0112f
C17750 vdd.n8563 vss 0.0128f
C17751 vdd.t1453 vss 0.00134f
C17752 vdd.t483 vss 0.0013f
C17753 vdd.n8564 vss 0.0332f
C17754 vdd.n8565 vss 0.0393f
C17755 vdd.n8566 vss 0.0345f
C17756 vdd.n8567 vss 0.262f
C17757 vdd.t849 vss 0.0013f
C17758 vdd.t1081 vss 0.00134f
C17759 vdd.n8568 vss 0.00324f
C17760 vdd.n8569 vss 0.0112f
C17761 vdd.n8570 vss 0.0128f
C17762 vdd.n8571 vss 0.00413f
C17763 vdd.n8572 vss 0.00413f
C17764 vdd.n8573 vss 0.0471f
C17765 vdd.n8574 vss 0.00251f
C17766 vdd.t773 vss 0.0471f
C17767 vdd.n8575 vss 0.00324f
C17768 vdd.n8577 vss 0.00679f
C17769 vdd.n8578 vss 0.00413f
C17770 vdd.n8579 vss 0.00324f
C17771 vdd.n8580 vss 0.00413f
C17772 vdd.n8581 vss 0.0471f
C17773 vdd.n8582 vss 0.00324f
C17774 vdd.n8584 vss 0.00925f
C17775 vdd.t412 vss 0.0471f
C17776 vdd.n8585 vss 0.00425f
C17777 vdd.n8586 vss 0.0424f
C17778 vdd.n8587 vss 0.0132f
C17779 vdd.n8588 vss 0.00324f
C17780 vdd.n8589 vss 0.0128f
C17781 vdd.n8590 vss 0.02f
C17782 vdd.n8591 vss 0.00425f
C17783 vdd.n8592 vss 0.00413f
C17784 vdd.n8593 vss 0.00251f
C17785 vdd.t764 vss 0.0471f
C17786 vdd.n8594 vss 0.00251f
C17787 vdd.n8595 vss 0.00517f
C17788 vdd.n8596 vss 0.00679f
C17789 vdd.n8597 vss 0.00517f
C17790 vdd.n8598 vss 0.00679f
C17791 vdd.n8599 vss 0.02f
C17792 vdd.n8600 vss 0.00425f
C17793 vdd.n8601 vss 0.0424f
C17794 vdd.n8602 vss 0.0132f
C17795 vdd.n8603 vss 0.00925f
C17796 vdd.n8604 vss 0.00425f
C17797 vdd.n8605 vss 0.00413f
C17798 vdd.n8606 vss 0.00324f
C17799 vdd.n8607 vss 0.0471f
C17800 vdd.t762 vss 0.0471f
C17801 vdd.n8608 vss 0.00251f
C17802 vdd.n8609 vss 0.0112f
C17803 vdd.n8610 vss 0.0128f
C17804 vdd.t763 vss 0.00134f
C17805 vdd.t774 vss 0.0013f
C17806 vdd.n8611 vss 0.0332f
C17807 vdd.n8612 vss 0.0393f
C17808 vdd.n8613 vss 0.119f
C17809 vdd.n8614 vss 0.00324f
C17810 vdd.n8615 vss 0.0112f
C17811 vdd.n8616 vss 0.0128f
C17812 vdd.n8617 vss 0.00413f
C17813 vdd.n8618 vss 0.00413f
C17814 vdd.n8619 vss 0.0471f
C17815 vdd.n8620 vss 0.00251f
C17816 vdd.t848 vss 0.0471f
C17817 vdd.n8621 vss 0.00324f
C17818 vdd.n8623 vss 0.00679f
C17819 vdd.n8624 vss 0.00413f
C17820 vdd.n8625 vss 0.00324f
C17821 vdd.n8626 vss 0.00413f
C17822 vdd.n8627 vss 0.0471f
C17823 vdd.n8628 vss 0.00324f
C17824 vdd.n8630 vss 0.00925f
C17825 vdd.t284 vss 0.0471f
C17826 vdd.n8631 vss 0.00425f
C17827 vdd.n8632 vss 0.0424f
C17828 vdd.n8633 vss 0.0132f
C17829 vdd.n8634 vss 0.00324f
C17830 vdd.n8635 vss 0.0128f
C17831 vdd.n8636 vss 0.02f
C17832 vdd.n8637 vss 0.00425f
C17833 vdd.n8638 vss 0.00413f
C17834 vdd.n8639 vss 0.00251f
C17835 vdd.t1079 vss 0.0471f
C17836 vdd.n8640 vss 0.00251f
C17837 vdd.n8641 vss 0.00517f
C17838 vdd.n8642 vss 0.00679f
C17839 vdd.n8643 vss 0.00517f
C17840 vdd.n8644 vss 0.00679f
C17841 vdd.n8645 vss 0.02f
C17842 vdd.n8646 vss 0.00425f
C17843 vdd.n8647 vss 0.0424f
C17844 vdd.n8648 vss 0.0132f
C17845 vdd.n8649 vss 0.00925f
C17846 vdd.n8650 vss 0.00425f
C17847 vdd.n8651 vss 0.00413f
C17848 vdd.n8652 vss 0.00324f
C17849 vdd.n8653 vss 0.0471f
C17850 vdd.t1080 vss 0.0471f
C17851 vdd.n8654 vss 0.00251f
C17852 vdd.n8655 vss 0.0112f
C17853 vdd.n8656 vss 0.0128f
C17854 vdd.n8657 vss 0.118f
C17855 vdd.n8658 vss 0.0393f
C17856 vdd.n8659 vss 0.0332f
C17857 vdd.n8660 vss 0.0596f
C17858 vdd.n8661 vss 0.00324f
C17859 vdd.n8662 vss 0.0112f
C17860 vdd.n8663 vss 0.0128f
C17861 vdd.n8664 vss 0.00413f
C17862 vdd.n8665 vss 0.00413f
C17863 vdd.n8666 vss 0.0471f
C17864 vdd.n8667 vss 0.00251f
C17865 vdd.t1314 vss 0.0471f
C17866 vdd.n8668 vss 0.00324f
C17867 vdd.n8670 vss 0.00679f
C17868 vdd.n8671 vss 0.00413f
C17869 vdd.n8672 vss 0.00324f
C17870 vdd.n8673 vss 0.00413f
C17871 vdd.n8674 vss 0.0471f
C17872 vdd.n8675 vss 0.00324f
C17873 vdd.n8677 vss 0.00925f
C17874 vdd.t1143 vss 0.0471f
C17875 vdd.n8678 vss 0.00425f
C17876 vdd.n8679 vss 0.0424f
C17877 vdd.n8680 vss 0.0132f
C17878 vdd.n8681 vss 0.00324f
C17879 vdd.n8682 vss 0.0128f
C17880 vdd.n8683 vss 0.02f
C17881 vdd.n8684 vss 0.00425f
C17882 vdd.n8685 vss 0.00413f
C17883 vdd.n8686 vss 0.00251f
C17884 vdd.t254 vss 0.0471f
C17885 vdd.n8687 vss 0.00251f
C17886 vdd.n8688 vss 0.00517f
C17887 vdd.n8689 vss 0.00679f
C17888 vdd.n8690 vss 0.00517f
C17889 vdd.n8691 vss 0.00679f
C17890 vdd.n8692 vss 0.02f
C17891 vdd.n8693 vss 0.00425f
C17892 vdd.n8694 vss 0.0424f
C17893 vdd.n8695 vss 0.0132f
C17894 vdd.n8696 vss 0.00925f
C17895 vdd.n8697 vss 0.00425f
C17896 vdd.n8698 vss 0.00413f
C17897 vdd.n8699 vss 0.00324f
C17898 vdd.n8700 vss 0.0471f
C17899 vdd.t255 vss 0.0471f
C17900 vdd.n8701 vss 0.00251f
C17901 vdd.n8702 vss 0.0112f
C17902 vdd.n8703 vss 0.0128f
C17903 vdd.t256 vss 0.00134f
C17904 vdd.t1315 vss 0.0013f
C17905 vdd.n8704 vss 0.0332f
C17906 vdd.n8705 vss 0.0393f
C17907 vdd.n8706 vss 0.0418f
C17908 vdd.n8707 vss 0.118f
C17909 vdd.n8708 vss 0.121f
C17910 vdd.t857 vss 0.0013f
C17911 vdd.t935 vss 0.00134f
C17912 vdd.n8709 vss 0.00324f
C17913 vdd.n8710 vss 0.0112f
C17914 vdd.n8711 vss 0.0128f
C17915 vdd.n8712 vss 0.00413f
C17916 vdd.n8713 vss 0.00413f
C17917 vdd.n8714 vss 0.0471f
C17918 vdd.n8715 vss 0.00251f
C17919 vdd.t856 vss 0.0471f
C17920 vdd.n8716 vss 0.00324f
C17921 vdd.n8718 vss 0.00679f
C17922 vdd.n8719 vss 0.00413f
C17923 vdd.n8720 vss 0.00324f
C17924 vdd.n8721 vss 0.00413f
C17925 vdd.n8722 vss 0.0471f
C17926 vdd.n8723 vss 0.00324f
C17927 vdd.n8725 vss 0.00925f
C17928 vdd.t658 vss 0.0471f
C17929 vdd.n8726 vss 0.00425f
C17930 vdd.n8727 vss 0.0424f
C17931 vdd.n8728 vss 0.0132f
C17932 vdd.n8729 vss 0.00324f
C17933 vdd.n8730 vss 0.0128f
C17934 vdd.n8731 vss 0.02f
C17935 vdd.n8732 vss 0.00425f
C17936 vdd.n8733 vss 0.00413f
C17937 vdd.n8734 vss 0.00251f
C17938 vdd.t933 vss 0.0471f
C17939 vdd.n8735 vss 0.00251f
C17940 vdd.n8736 vss 0.00517f
C17941 vdd.n8737 vss 0.00679f
C17942 vdd.n8738 vss 0.00517f
C17943 vdd.n8739 vss 0.00679f
C17944 vdd.n8740 vss 0.02f
C17945 vdd.n8741 vss 0.00425f
C17946 vdd.n8742 vss 0.0424f
C17947 vdd.n8743 vss 0.0132f
C17948 vdd.n8744 vss 0.00925f
C17949 vdd.n8745 vss 0.00425f
C17950 vdd.n8746 vss 0.00413f
C17951 vdd.n8747 vss 0.00324f
C17952 vdd.n8748 vss 0.0471f
C17953 vdd.t934 vss 0.0471f
C17954 vdd.n8749 vss 0.00251f
C17955 vdd.n8750 vss 0.0112f
C17956 vdd.n8751 vss 0.0707f
C17957 vdd.n8752 vss 0.0393f
C17958 vdd.n8753 vss 0.0332f
C17959 vdd.n8754 vss 0.0596f
C17960 vdd.n8755 vss 0.00324f
C17961 vdd.n8756 vss 0.0112f
C17962 vdd.n8757 vss 0.0128f
C17963 vdd.n8758 vss 0.00413f
C17964 vdd.n8759 vss 0.00413f
C17965 vdd.n8760 vss 0.0471f
C17966 vdd.n8761 vss 0.00251f
C17967 vdd.t1467 vss 0.0471f
C17968 vdd.n8762 vss 0.00324f
C17969 vdd.n8764 vss 0.00679f
C17970 vdd.n8765 vss 0.00413f
C17971 vdd.n8766 vss 0.00324f
C17972 vdd.n8767 vss 0.00413f
C17973 vdd.n8768 vss 0.0471f
C17974 vdd.n8769 vss 0.00324f
C17975 vdd.n8771 vss 0.00925f
C17976 vdd.t1507 vss 0.0471f
C17977 vdd.n8772 vss 0.00425f
C17978 vdd.n8773 vss 0.0424f
C17979 vdd.n8774 vss 0.0132f
C17980 vdd.n8775 vss 0.00324f
C17981 vdd.n8776 vss 0.0128f
C17982 vdd.n8777 vss 0.02f
C17983 vdd.n8778 vss 0.00425f
C17984 vdd.n8779 vss 0.00413f
C17985 vdd.n8780 vss 0.00251f
C17986 vdd.t190 vss 0.0471f
C17987 vdd.n8781 vss 0.00251f
C17988 vdd.n8782 vss 0.00517f
C17989 vdd.n8783 vss 0.00679f
C17990 vdd.n8784 vss 0.00517f
C17991 vdd.n8785 vss 0.00679f
C17992 vdd.n8786 vss 0.02f
C17993 vdd.n8787 vss 0.00425f
C17994 vdd.n8788 vss 0.0424f
C17995 vdd.n8789 vss 0.0132f
C17996 vdd.n8790 vss 0.00925f
C17997 vdd.n8791 vss 0.00425f
C17998 vdd.n8792 vss 0.00413f
C17999 vdd.n8793 vss 0.00324f
C18000 vdd.n8794 vss 0.0471f
C18001 vdd.t188 vss 0.0471f
C18002 vdd.n8795 vss 0.00251f
C18003 vdd.n8796 vss 0.0112f
C18004 vdd.n8797 vss 0.0128f
C18005 vdd.t189 vss 0.00134f
C18006 vdd.t1468 vss 0.0013f
C18007 vdd.n8798 vss 0.0332f
C18008 vdd.n8799 vss 0.0393f
C18009 vdd.n8800 vss 0.0418f
C18010 vdd.n8801 vss 0.0912f
C18011 vdd.n8802 vss 0.0824f
C18012 vdd.n8803 vss 0.059f
C18013 vdd.t826 vss 0.0013f
C18014 vdd.t138 vss 0.00134f
C18015 vdd.n8804 vss 0.00324f
C18016 vdd.n8805 vss 0.0112f
C18017 vdd.n8806 vss 0.0128f
C18018 vdd.n8807 vss 0.00413f
C18019 vdd.n8808 vss 0.00413f
C18020 vdd.n8809 vss 0.0471f
C18021 vdd.n8810 vss 0.00251f
C18022 vdd.t1129 vss 0.0471f
C18023 vdd.n8811 vss 0.00324f
C18024 vdd.n8813 vss 0.00679f
C18025 vdd.n8814 vss 0.00413f
C18026 vdd.n8815 vss 0.00324f
C18027 vdd.n8816 vss 0.00413f
C18028 vdd.n8817 vss 0.0471f
C18029 vdd.n8818 vss 0.00324f
C18030 vdd.n8820 vss 0.00925f
C18031 vdd.t264 vss 0.0471f
C18032 vdd.n8821 vss 0.00425f
C18033 vdd.n8822 vss 0.0424f
C18034 vdd.n8823 vss 0.0132f
C18035 vdd.n8824 vss 0.00324f
C18036 vdd.n8825 vss 0.0128f
C18037 vdd.n8826 vss 0.02f
C18038 vdd.n8827 vss 0.00425f
C18039 vdd.n8828 vss 0.00413f
C18040 vdd.n8829 vss 0.00251f
C18041 vdd.t1201 vss 0.0471f
C18042 vdd.n8830 vss 0.00251f
C18043 vdd.n8831 vss 0.00517f
C18044 vdd.n8832 vss 0.00679f
C18045 vdd.n8833 vss 0.00517f
C18046 vdd.n8834 vss 0.00679f
C18047 vdd.n8835 vss 0.02f
C18048 vdd.n8836 vss 0.00425f
C18049 vdd.n8837 vss 0.0424f
C18050 vdd.n8838 vss 0.0132f
C18051 vdd.n8839 vss 0.00925f
C18052 vdd.n8840 vss 0.00425f
C18053 vdd.n8841 vss 0.00413f
C18054 vdd.n8842 vss 0.00324f
C18055 vdd.n8843 vss 0.0471f
C18056 vdd.t1199 vss 0.0471f
C18057 vdd.n8844 vss 0.00251f
C18058 vdd.n8845 vss 0.0112f
C18059 vdd.n8846 vss 0.0128f
C18060 vdd.t1200 vss 0.00134f
C18061 vdd.t1130 vss 0.0013f
C18062 vdd.n8847 vss 0.0332f
C18063 vdd.n8848 vss 0.0393f
C18064 vdd.n8849 vss 0.158f
C18065 vdd.n8850 vss 0.00324f
C18066 vdd.n8851 vss 0.0112f
C18067 vdd.n8852 vss 0.0128f
C18068 vdd.n8853 vss 0.00413f
C18069 vdd.n8854 vss 0.00413f
C18070 vdd.n8855 vss 0.0471f
C18071 vdd.n8856 vss 0.00251f
C18072 vdd.t765 vss 0.0471f
C18073 vdd.n8857 vss 0.00324f
C18074 vdd.n8859 vss 0.00679f
C18075 vdd.n8860 vss 0.00413f
C18076 vdd.n8861 vss 0.00324f
C18077 vdd.n8862 vss 0.00413f
C18078 vdd.n8863 vss 0.0471f
C18079 vdd.n8864 vss 0.00324f
C18080 vdd.n8866 vss 0.00925f
C18081 vdd.t1195 vss 0.0471f
C18082 vdd.n8867 vss 0.00425f
C18083 vdd.n8868 vss 0.0424f
C18084 vdd.n8869 vss 0.0132f
C18085 vdd.n8870 vss 0.00324f
C18086 vdd.n8871 vss 0.0128f
C18087 vdd.n8872 vss 0.02f
C18088 vdd.n8873 vss 0.00425f
C18089 vdd.n8874 vss 0.00413f
C18090 vdd.n8875 vss 0.00251f
C18091 vdd.t584 vss 0.0471f
C18092 vdd.n8876 vss 0.00251f
C18093 vdd.n8877 vss 0.00517f
C18094 vdd.n8878 vss 0.00679f
C18095 vdd.n8879 vss 0.00517f
C18096 vdd.n8880 vss 0.00679f
C18097 vdd.n8881 vss 0.02f
C18098 vdd.n8882 vss 0.00425f
C18099 vdd.n8883 vss 0.0424f
C18100 vdd.n8884 vss 0.0132f
C18101 vdd.n8885 vss 0.00925f
C18102 vdd.n8886 vss 0.00425f
C18103 vdd.n8887 vss 0.00413f
C18104 vdd.n8888 vss 0.00324f
C18105 vdd.n8889 vss 0.0471f
C18106 vdd.t585 vss 0.0471f
C18107 vdd.n8890 vss 0.00251f
C18108 vdd.n8891 vss 0.0112f
C18109 vdd.n8892 vss 0.0128f
C18110 vdd.t586 vss 0.00134f
C18111 vdd.t766 vss 0.0013f
C18112 vdd.n8893 vss 0.0332f
C18113 vdd.n8894 vss 0.0393f
C18114 vdd.n8895 vss 0.0316f
C18115 vdd.n8896 vss 0.256f
C18116 vdd.n8897 vss 0.00324f
C18117 vdd.n8898 vss 0.0112f
C18118 vdd.n8899 vss 0.0128f
C18119 vdd.n8900 vss 0.00413f
C18120 vdd.n8901 vss 0.00413f
C18121 vdd.n8902 vss 0.0471f
C18122 vdd.n8903 vss 0.00251f
C18123 vdd.t825 vss 0.0471f
C18124 vdd.n8904 vss 0.00324f
C18125 vdd.n8906 vss 0.00679f
C18126 vdd.n8907 vss 0.00413f
C18127 vdd.n8908 vss 0.00324f
C18128 vdd.n8909 vss 0.00413f
C18129 vdd.n8910 vss 0.0471f
C18130 vdd.n8911 vss 0.00324f
C18131 vdd.n8913 vss 0.00925f
C18132 vdd.t66 vss 0.0471f
C18133 vdd.n8914 vss 0.00425f
C18134 vdd.n8915 vss 0.0424f
C18135 vdd.n8916 vss 0.0132f
C18136 vdd.n8917 vss 0.00324f
C18137 vdd.n8918 vss 0.0128f
C18138 vdd.n8919 vss 0.02f
C18139 vdd.n8920 vss 0.00425f
C18140 vdd.n8921 vss 0.00413f
C18141 vdd.n8922 vss 0.00251f
C18142 vdd.t139 vss 0.0471f
C18143 vdd.n8923 vss 0.00251f
C18144 vdd.n8924 vss 0.00517f
C18145 vdd.n8925 vss 0.00679f
C18146 vdd.n8926 vss 0.00517f
C18147 vdd.n8927 vss 0.00679f
C18148 vdd.n8928 vss 0.02f
C18149 vdd.n8929 vss 0.00425f
C18150 vdd.n8930 vss 0.0424f
C18151 vdd.n8931 vss 0.0132f
C18152 vdd.n8932 vss 0.00925f
C18153 vdd.n8933 vss 0.00425f
C18154 vdd.n8934 vss 0.00413f
C18155 vdd.n8935 vss 0.00324f
C18156 vdd.n8936 vss 0.0471f
C18157 vdd.t137 vss 0.0471f
C18158 vdd.n8937 vss 0.00251f
C18159 vdd.n8938 vss 0.0112f
C18160 vdd.n8939 vss 0.0128f
C18161 vdd.n8940 vss 0.0953f
C18162 vdd.n8941 vss 0.0393f
C18163 vdd.n8942 vss 0.0332f
C18164 vdd.n8943 vss 0.0596f
C18165 vdd.n8944 vss 0.00324f
C18166 vdd.n8945 vss 0.0112f
C18167 vdd.n8946 vss 0.0128f
C18168 vdd.n8947 vss 0.00413f
C18169 vdd.n8948 vss 0.00413f
C18170 vdd.n8949 vss 0.0471f
C18171 vdd.n8950 vss 0.00251f
C18172 vdd.t458 vss 0.0471f
C18173 vdd.n8951 vss 0.00324f
C18174 vdd.n8953 vss 0.00679f
C18175 vdd.n8954 vss 0.00413f
C18176 vdd.n8955 vss 0.00324f
C18177 vdd.n8956 vss 0.00413f
C18178 vdd.n8957 vss 0.0471f
C18179 vdd.n8958 vss 0.00324f
C18180 vdd.n8960 vss 0.00925f
C18181 vdd.t758 vss 0.0471f
C18182 vdd.n8961 vss 0.00425f
C18183 vdd.n8962 vss 0.0424f
C18184 vdd.n8963 vss 0.0132f
C18185 vdd.n8964 vss 0.00324f
C18186 vdd.n8965 vss 0.0128f
C18187 vdd.n8966 vss 0.02f
C18188 vdd.n8967 vss 0.00425f
C18189 vdd.n8968 vss 0.00413f
C18190 vdd.n8969 vss 0.00251f
C18191 vdd.t755 vss 0.0471f
C18192 vdd.n8970 vss 0.00251f
C18193 vdd.n8971 vss 0.00517f
C18194 vdd.n8972 vss 0.00679f
C18195 vdd.n8973 vss 0.00517f
C18196 vdd.n8974 vss 0.00679f
C18197 vdd.n8975 vss 0.02f
C18198 vdd.n8976 vss 0.00425f
C18199 vdd.n8977 vss 0.0424f
C18200 vdd.n8978 vss 0.0132f
C18201 vdd.n8979 vss 0.00925f
C18202 vdd.n8980 vss 0.00425f
C18203 vdd.n8981 vss 0.00413f
C18204 vdd.n8982 vss 0.00324f
C18205 vdd.n8983 vss 0.0471f
C18206 vdd.t756 vss 0.0471f
C18207 vdd.n8984 vss 0.00251f
C18208 vdd.n8985 vss 0.0112f
C18209 vdd.n8986 vss 0.0128f
C18210 vdd.t757 vss 0.00134f
C18211 vdd.t459 vss 0.0013f
C18212 vdd.n8987 vss 0.0332f
C18213 vdd.n8988 vss 0.0393f
C18214 vdd.n8989 vss 0.0418f
C18215 vdd.n8990 vss 0.118f
C18216 vdd.n8991 vss 0.121f
C18217 vdd.t865 vss 0.0013f
C18218 vdd.t639 vss 0.00134f
C18219 vdd.n8992 vss 0.00324f
C18220 vdd.n8993 vss 0.0112f
C18221 vdd.n8994 vss 0.0128f
C18222 vdd.n8995 vss 0.00413f
C18223 vdd.n8996 vss 0.00413f
C18224 vdd.n8997 vss 0.0471f
C18225 vdd.n8998 vss 0.00251f
C18226 vdd.t864 vss 0.0471f
C18227 vdd.n8999 vss 0.00324f
C18228 vdd.n9001 vss 0.00679f
C18229 vdd.n9002 vss 0.00413f
C18230 vdd.n9003 vss 0.00324f
C18231 vdd.n9004 vss 0.00413f
C18232 vdd.n9005 vss 0.0471f
C18233 vdd.n9006 vss 0.00324f
C18234 vdd.n9008 vss 0.00925f
C18235 vdd.t1062 vss 0.0471f
C18236 vdd.n9009 vss 0.00425f
C18237 vdd.n9010 vss 0.0424f
C18238 vdd.n9011 vss 0.0132f
C18239 vdd.n9012 vss 0.00324f
C18240 vdd.n9013 vss 0.0128f
C18241 vdd.n9014 vss 0.02f
C18242 vdd.n9015 vss 0.00425f
C18243 vdd.n9016 vss 0.00413f
C18244 vdd.n9017 vss 0.00251f
C18245 vdd.t640 vss 0.0471f
C18246 vdd.n9018 vss 0.00251f
C18247 vdd.n9019 vss 0.00517f
C18248 vdd.n9020 vss 0.00679f
C18249 vdd.n9021 vss 0.00517f
C18250 vdd.n9022 vss 0.00679f
C18251 vdd.n9023 vss 0.02f
C18252 vdd.n9024 vss 0.00425f
C18253 vdd.n9025 vss 0.0424f
C18254 vdd.n9026 vss 0.0132f
C18255 vdd.n9027 vss 0.00925f
C18256 vdd.n9028 vss 0.00425f
C18257 vdd.n9029 vss 0.00413f
C18258 vdd.n9030 vss 0.00324f
C18259 vdd.n9031 vss 0.0471f
C18260 vdd.t638 vss 0.0471f
C18261 vdd.n9032 vss 0.00251f
C18262 vdd.n9033 vss 0.0112f
C18263 vdd.n9034 vss 0.0707f
C18264 vdd.n9035 vss 0.0393f
C18265 vdd.n9036 vss 0.0332f
C18266 vdd.n9037 vss 0.0596f
C18267 vdd.n9038 vss 0.00324f
C18268 vdd.n9039 vss 0.0112f
C18269 vdd.n9040 vss 0.0128f
C18270 vdd.n9041 vss 0.00413f
C18271 vdd.n9042 vss 0.00413f
C18272 vdd.n9043 vss 0.0471f
C18273 vdd.n9044 vss 0.00251f
C18274 vdd.t1477 vss 0.0471f
C18275 vdd.n9045 vss 0.00324f
C18276 vdd.n9047 vss 0.00679f
C18277 vdd.n9048 vss 0.00413f
C18278 vdd.n9049 vss 0.00324f
C18279 vdd.n9050 vss 0.00413f
C18280 vdd.n9051 vss 0.0471f
C18281 vdd.n9052 vss 0.00324f
C18282 vdd.n9054 vss 0.00925f
C18283 vdd.t1108 vss 0.0471f
C18284 vdd.n9055 vss 0.00425f
C18285 vdd.n9056 vss 0.0424f
C18286 vdd.n9057 vss 0.0132f
C18287 vdd.n9058 vss 0.00324f
C18288 vdd.n9059 vss 0.0128f
C18289 vdd.n9060 vss 0.02f
C18290 vdd.n9061 vss 0.00425f
C18291 vdd.n9062 vss 0.00413f
C18292 vdd.n9063 vss 0.00251f
C18293 vdd.t1526 vss 0.0471f
C18294 vdd.n9064 vss 0.00251f
C18295 vdd.n9065 vss 0.00517f
C18296 vdd.n9066 vss 0.00679f
C18297 vdd.n9067 vss 0.00517f
C18298 vdd.n9068 vss 0.00679f
C18299 vdd.n9069 vss 0.02f
C18300 vdd.n9070 vss 0.00425f
C18301 vdd.n9071 vss 0.0424f
C18302 vdd.n9072 vss 0.0132f
C18303 vdd.n9073 vss 0.00925f
C18304 vdd.n9074 vss 0.00425f
C18305 vdd.n9075 vss 0.00413f
C18306 vdd.n9076 vss 0.00324f
C18307 vdd.n9077 vss 0.0471f
C18308 vdd.t1524 vss 0.0471f
C18309 vdd.n9078 vss 0.00251f
C18310 vdd.n9079 vss 0.0112f
C18311 vdd.n9080 vss 0.0128f
C18312 vdd.t1525 vss 0.00134f
C18313 vdd.t1478 vss 0.0013f
C18314 vdd.n9081 vss 0.0332f
C18315 vdd.n9082 vss 0.0393f
C18316 vdd.n9083 vss 0.0418f
C18317 vdd.n9084 vss 0.118f
C18318 vdd.n9085 vss 0.0951f
C18319 vdd.t1007 vss 0.0013f
C18320 vdd.t79 vss 0.00134f
C18321 vdd.n9086 vss 0.00324f
C18322 vdd.n9087 vss 0.0112f
C18323 vdd.n9088 vss 0.0128f
C18324 vdd.n9089 vss 0.00413f
C18325 vdd.n9090 vss 0.00413f
C18326 vdd.n9091 vss 0.0471f
C18327 vdd.n9092 vss 0.00251f
C18328 vdd.t430 vss 0.0471f
C18329 vdd.n9093 vss 0.00324f
C18330 vdd.n9095 vss 0.00679f
C18331 vdd.n9096 vss 0.00413f
C18332 vdd.n9097 vss 0.00324f
C18333 vdd.n9098 vss 0.00413f
C18334 vdd.n9099 vss 0.0471f
C18335 vdd.n9100 vss 0.00324f
C18336 vdd.n9102 vss 0.00925f
C18337 vdd.t1024 vss 0.0471f
C18338 vdd.n9103 vss 0.00425f
C18339 vdd.n9104 vss 0.0424f
C18340 vdd.n9105 vss 0.0132f
C18341 vdd.n9106 vss 0.00324f
C18342 vdd.n9107 vss 0.0128f
C18343 vdd.n9108 vss 0.02f
C18344 vdd.n9109 vss 0.00425f
C18345 vdd.n9110 vss 0.00413f
C18346 vdd.n9111 vss 0.00251f
C18347 vdd.t785 vss 0.0471f
C18348 vdd.n9112 vss 0.00251f
C18349 vdd.n9113 vss 0.00517f
C18350 vdd.n9114 vss 0.00679f
C18351 vdd.n9115 vss 0.00517f
C18352 vdd.n9116 vss 0.00679f
C18353 vdd.n9117 vss 0.02f
C18354 vdd.n9118 vss 0.00425f
C18355 vdd.n9119 vss 0.0424f
C18356 vdd.n9120 vss 0.0132f
C18357 vdd.n9121 vss 0.00925f
C18358 vdd.n9122 vss 0.00425f
C18359 vdd.n9123 vss 0.00413f
C18360 vdd.n9124 vss 0.00324f
C18361 vdd.n9125 vss 0.0471f
C18362 vdd.t783 vss 0.0471f
C18363 vdd.n9126 vss 0.00251f
C18364 vdd.n9127 vss 0.0112f
C18365 vdd.n9128 vss 0.0128f
C18366 vdd.t784 vss 0.00134f
C18367 vdd.t431 vss 0.0013f
C18368 vdd.n9129 vss 0.0332f
C18369 vdd.n9130 vss 0.0393f
C18370 vdd.n9131 vss 0.119f
C18371 vdd.n9132 vss 0.00324f
C18372 vdd.n9133 vss 0.0112f
C18373 vdd.n9134 vss 0.0128f
C18374 vdd.n9135 vss 0.00413f
C18375 vdd.n9136 vss 0.00413f
C18376 vdd.n9137 vss 0.0471f
C18377 vdd.n9138 vss 0.00251f
C18378 vdd.t1006 vss 0.0471f
C18379 vdd.n9139 vss 0.00324f
C18380 vdd.n9141 vss 0.00679f
C18381 vdd.n9142 vss 0.00413f
C18382 vdd.n9143 vss 0.00324f
C18383 vdd.n9144 vss 0.00413f
C18384 vdd.n9145 vss 0.0471f
C18385 vdd.n9146 vss 0.00324f
C18386 vdd.n9148 vss 0.00925f
C18387 vdd.t64 vss 0.0471f
C18388 vdd.n9149 vss 0.00425f
C18389 vdd.n9150 vss 0.0424f
C18390 vdd.n9151 vss 0.0132f
C18391 vdd.n9152 vss 0.00324f
C18392 vdd.n9153 vss 0.0128f
C18393 vdd.n9154 vss 0.02f
C18394 vdd.n9155 vss 0.00425f
C18395 vdd.n9156 vss 0.00413f
C18396 vdd.n9157 vss 0.00251f
C18397 vdd.t77 vss 0.0471f
C18398 vdd.n9158 vss 0.00251f
C18399 vdd.n9159 vss 0.00517f
C18400 vdd.n9160 vss 0.00679f
C18401 vdd.n9161 vss 0.00517f
C18402 vdd.n9162 vss 0.00679f
C18403 vdd.n9163 vss 0.02f
C18404 vdd.n9164 vss 0.00425f
C18405 vdd.n9165 vss 0.0424f
C18406 vdd.n9166 vss 0.0132f
C18407 vdd.n9167 vss 0.00925f
C18408 vdd.n9168 vss 0.00425f
C18409 vdd.n9169 vss 0.00413f
C18410 vdd.n9170 vss 0.00324f
C18411 vdd.n9171 vss 0.0471f
C18412 vdd.t78 vss 0.0471f
C18413 vdd.n9172 vss 0.00251f
C18414 vdd.n9173 vss 0.0112f
C18415 vdd.n9174 vss 0.0128f
C18416 vdd.n9175 vss 0.118f
C18417 vdd.n9176 vss 0.0393f
C18418 vdd.n9177 vss 0.0332f
C18419 vdd.n9178 vss 0.0596f
C18420 vdd.n9179 vss 0.00324f
C18421 vdd.n9180 vss 0.0112f
C18422 vdd.n9181 vss 0.0128f
C18423 vdd.n9182 vss 0.00413f
C18424 vdd.n9183 vss 0.00413f
C18425 vdd.n9184 vss 0.0471f
C18426 vdd.n9185 vss 0.00251f
C18427 vdd.t566 vss 0.0471f
C18428 vdd.n9186 vss 0.00324f
C18429 vdd.n9188 vss 0.00679f
C18430 vdd.n9189 vss 0.00413f
C18431 vdd.n9190 vss 0.00324f
C18432 vdd.n9191 vss 0.00413f
C18433 vdd.n9192 vss 0.0471f
C18434 vdd.n9193 vss 0.00324f
C18435 vdd.n9195 vss 0.00925f
C18436 vdd.t1270 vss 0.0471f
C18437 vdd.n9196 vss 0.00425f
C18438 vdd.n9197 vss 0.0424f
C18439 vdd.n9198 vss 0.0132f
C18440 vdd.n9199 vss 0.00324f
C18441 vdd.n9200 vss 0.0128f
C18442 vdd.n9201 vss 0.02f
C18443 vdd.n9202 vss 0.00425f
C18444 vdd.n9203 vss 0.00413f
C18445 vdd.n9204 vss 0.00251f
C18446 vdd.t1267 vss 0.0471f
C18447 vdd.n9205 vss 0.00251f
C18448 vdd.n9206 vss 0.00517f
C18449 vdd.n9207 vss 0.00679f
C18450 vdd.n9208 vss 0.00517f
C18451 vdd.n9209 vss 0.00679f
C18452 vdd.n9210 vss 0.02f
C18453 vdd.n9211 vss 0.00425f
C18454 vdd.n9212 vss 0.0424f
C18455 vdd.n9213 vss 0.0132f
C18456 vdd.n9214 vss 0.00925f
C18457 vdd.n9215 vss 0.00425f
C18458 vdd.n9216 vss 0.00413f
C18459 vdd.n9217 vss 0.00324f
C18460 vdd.n9218 vss 0.0471f
C18461 vdd.t1268 vss 0.0471f
C18462 vdd.n9219 vss 0.00251f
C18463 vdd.n9220 vss 0.0112f
C18464 vdd.n9221 vss 0.0128f
C18465 vdd.t1269 vss 0.00134f
C18466 vdd.t567 vss 0.0013f
C18467 vdd.n9222 vss 0.0332f
C18468 vdd.n9223 vss 0.0393f
C18469 vdd.n9224 vss 0.0418f
C18470 vdd.n9225 vss 0.118f
C18471 vdd.n9226 vss 0.121f
C18472 vdd.t43 vss 0.0013f
C18473 vdd.t746 vss 0.00134f
C18474 vdd.n9227 vss 0.00324f
C18475 vdd.n9228 vss 0.0112f
C18476 vdd.n9229 vss 0.0128f
C18477 vdd.n9230 vss 0.00413f
C18478 vdd.n9231 vss 0.00413f
C18479 vdd.n9232 vss 0.0471f
C18480 vdd.n9233 vss 0.00251f
C18481 vdd.t42 vss 0.0471f
C18482 vdd.n9234 vss 0.00324f
C18483 vdd.n9236 vss 0.00679f
C18484 vdd.n9237 vss 0.00413f
C18485 vdd.n9238 vss 0.00324f
C18486 vdd.n9239 vss 0.00413f
C18487 vdd.n9240 vss 0.0471f
C18488 vdd.n9241 vss 0.00324f
C18489 vdd.n9243 vss 0.00925f
C18490 vdd.t675 vss 0.0471f
C18491 vdd.n9244 vss 0.00425f
C18492 vdd.n9245 vss 0.0424f
C18493 vdd.n9246 vss 0.0132f
C18494 vdd.n9247 vss 0.00324f
C18495 vdd.n9248 vss 0.0128f
C18496 vdd.n9249 vss 0.02f
C18497 vdd.n9250 vss 0.00425f
C18498 vdd.n9251 vss 0.00413f
C18499 vdd.n9252 vss 0.00251f
C18500 vdd.t744 vss 0.0471f
C18501 vdd.n9253 vss 0.00251f
C18502 vdd.n9254 vss 0.00517f
C18503 vdd.n9255 vss 0.00679f
C18504 vdd.n9256 vss 0.00517f
C18505 vdd.n9257 vss 0.00679f
C18506 vdd.n9258 vss 0.02f
C18507 vdd.n9259 vss 0.00425f
C18508 vdd.n9260 vss 0.0424f
C18509 vdd.n9261 vss 0.0132f
C18510 vdd.n9262 vss 0.00925f
C18511 vdd.n9263 vss 0.00425f
C18512 vdd.n9264 vss 0.00413f
C18513 vdd.n9265 vss 0.00324f
C18514 vdd.n9266 vss 0.0471f
C18515 vdd.t745 vss 0.0471f
C18516 vdd.n9267 vss 0.00251f
C18517 vdd.n9268 vss 0.0112f
C18518 vdd.n9269 vss 0.0707f
C18519 vdd.n9270 vss 0.0393f
C18520 vdd.n9271 vss 0.0332f
C18521 vdd.n9272 vss 0.0596f
C18522 vdd.n9273 vss 0.00324f
C18523 vdd.n9274 vss 0.0112f
C18524 vdd.n9275 vss 0.0128f
C18525 vdd.n9276 vss 0.00413f
C18526 vdd.n9277 vss 0.00413f
C18527 vdd.n9278 vss 0.0471f
C18528 vdd.n9279 vss 0.00251f
C18529 vdd.t1302 vss 0.0471f
C18530 vdd.n9280 vss 0.00324f
C18531 vdd.n9282 vss 0.00679f
C18532 vdd.n9283 vss 0.00413f
C18533 vdd.n9284 vss 0.00324f
C18534 vdd.n9285 vss 0.00413f
C18535 vdd.n9286 vss 0.0471f
C18536 vdd.n9287 vss 0.00324f
C18537 vdd.n9289 vss 0.00925f
C18538 vdd.t547 vss 0.0471f
C18539 vdd.n9290 vss 0.00425f
C18540 vdd.n9291 vss 0.0424f
C18541 vdd.n9292 vss 0.0132f
C18542 vdd.n9293 vss 0.00324f
C18543 vdd.n9294 vss 0.0128f
C18544 vdd.n9295 vss 0.02f
C18545 vdd.n9296 vss 0.00425f
C18546 vdd.n9297 vss 0.00413f
C18547 vdd.n9298 vss 0.00251f
C18548 vdd.t401 vss 0.0471f
C18549 vdd.n9299 vss 0.00251f
C18550 vdd.n9300 vss 0.00517f
C18551 vdd.n9301 vss 0.00679f
C18552 vdd.n9302 vss 0.00517f
C18553 vdd.n9303 vss 0.00679f
C18554 vdd.n9304 vss 0.02f
C18555 vdd.n9305 vss 0.00425f
C18556 vdd.n9306 vss 0.0424f
C18557 vdd.n9307 vss 0.0132f
C18558 vdd.n9308 vss 0.00925f
C18559 vdd.n9309 vss 0.00425f
C18560 vdd.n9310 vss 0.00413f
C18561 vdd.n9311 vss 0.00324f
C18562 vdd.n9312 vss 0.0471f
C18563 vdd.t399 vss 0.0471f
C18564 vdd.n9313 vss 0.00251f
C18565 vdd.n9314 vss 0.0112f
C18566 vdd.n9315 vss 0.0128f
C18567 vdd.t400 vss 0.00134f
C18568 vdd.t1303 vss 0.0013f
C18569 vdd.n9316 vss 0.0332f
C18570 vdd.n9317 vss 0.0393f
C18571 vdd.n9318 vss 0.0418f
C18572 vdd.n9319 vss 0.0912f
C18573 vdd.n9320 vss 0.0824f
C18574 vdd.n9321 vss 0.059f
C18575 vdd.t989 vss 0.0013f
C18576 vdd.t178 vss 0.00134f
C18577 vdd.n9322 vss 0.00324f
C18578 vdd.n9323 vss 0.0112f
C18579 vdd.n9324 vss 0.0128f
C18580 vdd.n9325 vss 0.00413f
C18581 vdd.n9326 vss 0.00413f
C18582 vdd.n9327 vss 0.0471f
C18583 vdd.n9328 vss 0.00251f
C18584 vdd.t627 vss 0.0471f
C18585 vdd.n9329 vss 0.00324f
C18586 vdd.n9331 vss 0.00679f
C18587 vdd.n9332 vss 0.00413f
C18588 vdd.n9333 vss 0.00324f
C18589 vdd.n9334 vss 0.00413f
C18590 vdd.n9335 vss 0.0471f
C18591 vdd.n9336 vss 0.00324f
C18592 vdd.n9338 vss 0.00925f
C18593 vdd.t1031 vss 0.0471f
C18594 vdd.n9339 vss 0.00425f
C18595 vdd.n9340 vss 0.0424f
C18596 vdd.n9341 vss 0.0132f
C18597 vdd.n9342 vss 0.00324f
C18598 vdd.n9343 vss 0.0128f
C18599 vdd.n9344 vss 0.02f
C18600 vdd.n9345 vss 0.00425f
C18601 vdd.n9346 vss 0.00413f
C18602 vdd.n9347 vss 0.00251f
C18603 vdd.t1028 vss 0.0471f
C18604 vdd.n9348 vss 0.00251f
C18605 vdd.n9349 vss 0.00517f
C18606 vdd.n9350 vss 0.00679f
C18607 vdd.n9351 vss 0.00517f
C18608 vdd.n9352 vss 0.00679f
C18609 vdd.n9353 vss 0.02f
C18610 vdd.n9354 vss 0.00425f
C18611 vdd.n9355 vss 0.0424f
C18612 vdd.n9356 vss 0.0132f
C18613 vdd.n9357 vss 0.00925f
C18614 vdd.n9358 vss 0.00425f
C18615 vdd.n9359 vss 0.00413f
C18616 vdd.n9360 vss 0.00324f
C18617 vdd.n9361 vss 0.0471f
C18618 vdd.t1029 vss 0.0471f
C18619 vdd.n9362 vss 0.00251f
C18620 vdd.n9363 vss 0.0112f
C18621 vdd.n9364 vss 0.0128f
C18622 vdd.t1030 vss 0.00134f
C18623 vdd.t628 vss 0.0013f
C18624 vdd.n9365 vss 0.0332f
C18625 vdd.n9366 vss 0.0393f
C18626 vdd.n9367 vss 0.119f
C18627 vdd.n9368 vss 0.00324f
C18628 vdd.n9369 vss 0.0112f
C18629 vdd.n9370 vss 0.0128f
C18630 vdd.n9371 vss 0.00413f
C18631 vdd.n9372 vss 0.00413f
C18632 vdd.n9373 vss 0.0471f
C18633 vdd.n9374 vss 0.00251f
C18634 vdd.t988 vss 0.0471f
C18635 vdd.n9375 vss 0.00324f
C18636 vdd.n9377 vss 0.00679f
C18637 vdd.n9378 vss 0.00413f
C18638 vdd.n9379 vss 0.00324f
C18639 vdd.n9380 vss 0.00413f
C18640 vdd.n9381 vss 0.0471f
C18641 vdd.n9382 vss 0.00324f
C18642 vdd.n9384 vss 0.00925f
C18643 vdd.t523 vss 0.0471f
C18644 vdd.n9385 vss 0.00425f
C18645 vdd.n9386 vss 0.0424f
C18646 vdd.n9387 vss 0.0132f
C18647 vdd.n9388 vss 0.00324f
C18648 vdd.n9389 vss 0.0128f
C18649 vdd.n9390 vss 0.02f
C18650 vdd.n9391 vss 0.00425f
C18651 vdd.n9392 vss 0.00413f
C18652 vdd.n9393 vss 0.00251f
C18653 vdd.t176 vss 0.0471f
C18654 vdd.n9394 vss 0.00251f
C18655 vdd.n9395 vss 0.00517f
C18656 vdd.n9396 vss 0.00679f
C18657 vdd.n9397 vss 0.00517f
C18658 vdd.n9398 vss 0.00679f
C18659 vdd.n9399 vss 0.02f
C18660 vdd.n9400 vss 0.00425f
C18661 vdd.n9401 vss 0.0424f
C18662 vdd.n9402 vss 0.0132f
C18663 vdd.n9403 vss 0.00925f
C18664 vdd.n9404 vss 0.00425f
C18665 vdd.n9405 vss 0.00413f
C18666 vdd.n9406 vss 0.00324f
C18667 vdd.n9407 vss 0.0471f
C18668 vdd.t177 vss 0.0471f
C18669 vdd.n9408 vss 0.00251f
C18670 vdd.n9409 vss 0.0112f
C18671 vdd.n9410 vss 0.0128f
C18672 vdd.n9411 vss 0.118f
C18673 vdd.n9412 vss 0.0393f
C18674 vdd.n9413 vss 0.0332f
C18675 vdd.n9414 vss 0.0596f
C18676 vdd.n9415 vss 0.00324f
C18677 vdd.n9416 vss 0.0112f
C18678 vdd.n9417 vss 0.0128f
C18679 vdd.n9418 vss 0.00413f
C18680 vdd.n9419 vss 0.00413f
C18681 vdd.n9420 vss 0.0471f
C18682 vdd.n9421 vss 0.00251f
C18683 vdd.t601 vss 0.0471f
C18684 vdd.n9422 vss 0.00324f
C18685 vdd.n9424 vss 0.00679f
C18686 vdd.n9425 vss 0.00413f
C18687 vdd.n9426 vss 0.00324f
C18688 vdd.n9427 vss 0.00413f
C18689 vdd.n9428 vss 0.0471f
C18690 vdd.n9429 vss 0.00324f
C18691 vdd.n9431 vss 0.00925f
C18692 vdd.t428 vss 0.0471f
C18693 vdd.n9432 vss 0.00425f
C18694 vdd.n9433 vss 0.0424f
C18695 vdd.n9434 vss 0.0132f
C18696 vdd.n9435 vss 0.00324f
C18697 vdd.n9436 vss 0.0128f
C18698 vdd.n9437 vss 0.02f
C18699 vdd.n9438 vss 0.00425f
C18700 vdd.n9439 vss 0.00413f
C18701 vdd.n9440 vss 0.00251f
C18702 vdd.t546 vss 0.0471f
C18703 vdd.n9441 vss 0.00251f
C18704 vdd.n9442 vss 0.00517f
C18705 vdd.n9443 vss 0.00679f
C18706 vdd.n9444 vss 0.00517f
C18707 vdd.n9445 vss 0.00679f
C18708 vdd.n9446 vss 0.02f
C18709 vdd.n9447 vss 0.00425f
C18710 vdd.n9448 vss 0.0424f
C18711 vdd.n9449 vss 0.0132f
C18712 vdd.n9450 vss 0.00925f
C18713 vdd.n9451 vss 0.00425f
C18714 vdd.n9452 vss 0.00413f
C18715 vdd.n9453 vss 0.00324f
C18716 vdd.n9454 vss 0.0471f
C18717 vdd.t544 vss 0.0471f
C18718 vdd.n9455 vss 0.00251f
C18719 vdd.n9456 vss 0.0112f
C18720 vdd.n9457 vss 0.0128f
C18721 vdd.t545 vss 0.00134f
C18722 vdd.t602 vss 0.0013f
C18723 vdd.n9458 vss 0.0332f
C18724 vdd.n9459 vss 0.0393f
C18725 vdd.n9460 vss 0.0418f
C18726 vdd.n9461 vss 0.118f
C18727 vdd.n9462 vss 0.121f
C18728 vdd.t861 vss 0.0013f
C18729 vdd.t663 vss 0.00134f
C18730 vdd.n9463 vss 0.00324f
C18731 vdd.n9464 vss 0.0112f
C18732 vdd.n9465 vss 0.0128f
C18733 vdd.n9466 vss 0.00413f
C18734 vdd.n9467 vss 0.00413f
C18735 vdd.n9468 vss 0.0471f
C18736 vdd.n9469 vss 0.00251f
C18737 vdd.t860 vss 0.0471f
C18738 vdd.n9470 vss 0.00324f
C18739 vdd.n9472 vss 0.00679f
C18740 vdd.n9473 vss 0.00413f
C18741 vdd.n9474 vss 0.00324f
C18742 vdd.n9475 vss 0.00413f
C18743 vdd.n9476 vss 0.0471f
C18744 vdd.n9477 vss 0.00324f
C18745 vdd.n9479 vss 0.00925f
C18746 vdd.t1191 vss 0.0471f
C18747 vdd.n9480 vss 0.00425f
C18748 vdd.n9481 vss 0.0424f
C18749 vdd.n9482 vss 0.0132f
C18750 vdd.n9483 vss 0.00324f
C18751 vdd.n9484 vss 0.0128f
C18752 vdd.n9485 vss 0.02f
C18753 vdd.n9486 vss 0.00425f
C18754 vdd.n9487 vss 0.00413f
C18755 vdd.n9488 vss 0.00251f
C18756 vdd.t661 vss 0.0471f
C18757 vdd.n9489 vss 0.00251f
C18758 vdd.n9490 vss 0.00517f
C18759 vdd.n9491 vss 0.00679f
C18760 vdd.n9492 vss 0.00517f
C18761 vdd.n9493 vss 0.00679f
C18762 vdd.n9494 vss 0.02f
C18763 vdd.n9495 vss 0.00425f
C18764 vdd.n9496 vss 0.0424f
C18765 vdd.n9497 vss 0.0132f
C18766 vdd.n9498 vss 0.00925f
C18767 vdd.n9499 vss 0.00425f
C18768 vdd.n9500 vss 0.00413f
C18769 vdd.n9501 vss 0.00324f
C18770 vdd.n9502 vss 0.0471f
C18771 vdd.t662 vss 0.0471f
C18772 vdd.n9503 vss 0.00251f
C18773 vdd.n9504 vss 0.0112f
C18774 vdd.n9505 vss 0.0707f
C18775 vdd.n9506 vss 0.0393f
C18776 vdd.n9507 vss 0.0332f
C18777 vdd.n9508 vss 0.0596f
C18778 vdd.n9509 vss 0.00324f
C18779 vdd.n9510 vss 0.0112f
C18780 vdd.n9511 vss 0.0128f
C18781 vdd.n9512 vss 0.00413f
C18782 vdd.n9513 vss 0.00413f
C18783 vdd.n9514 vss 0.0471f
C18784 vdd.n9515 vss 0.00251f
C18785 vdd.t1041 vss 0.0471f
C18786 vdd.n9516 vss 0.00324f
C18787 vdd.n9518 vss 0.00679f
C18788 vdd.n9519 vss 0.00413f
C18789 vdd.n9520 vss 0.00324f
C18790 vdd.n9521 vss 0.00413f
C18791 vdd.n9522 vss 0.0471f
C18792 vdd.n9523 vss 0.00324f
C18793 vdd.n9525 vss 0.00925f
C18794 vdd.t76 vss 0.0471f
C18795 vdd.n9526 vss 0.00425f
C18796 vdd.n9527 vss 0.0424f
C18797 vdd.n9528 vss 0.0132f
C18798 vdd.n9529 vss 0.00324f
C18799 vdd.n9530 vss 0.0128f
C18800 vdd.n9531 vss 0.02f
C18801 vdd.n9532 vss 0.00425f
C18802 vdd.n9533 vss 0.00413f
C18803 vdd.n9534 vss 0.00251f
C18804 vdd.t1518 vss 0.0471f
C18805 vdd.n9535 vss 0.00251f
C18806 vdd.n9536 vss 0.00517f
C18807 vdd.n9537 vss 0.00679f
C18808 vdd.n9538 vss 0.00517f
C18809 vdd.n9539 vss 0.00679f
C18810 vdd.n9540 vss 0.02f
C18811 vdd.n9541 vss 0.00425f
C18812 vdd.n9542 vss 0.0424f
C18813 vdd.n9543 vss 0.0132f
C18814 vdd.n9544 vss 0.00925f
C18815 vdd.n9545 vss 0.00425f
C18816 vdd.n9546 vss 0.00413f
C18817 vdd.n9547 vss 0.00324f
C18818 vdd.n9548 vss 0.0471f
C18819 vdd.t1519 vss 0.0471f
C18820 vdd.n9549 vss 0.00251f
C18821 vdd.n9550 vss 0.0112f
C18822 vdd.n9551 vss 0.0128f
C18823 vdd.t1520 vss 0.00134f
C18824 vdd.t1042 vss 0.0013f
C18825 vdd.n9552 vss 0.0332f
C18826 vdd.n9553 vss 0.0393f
C18827 vdd.n9554 vss 0.0418f
C18828 vdd.n9555 vss 0.121f
C18829 vdd.n9556 vss 0.291f
C18830 vdd.n9557 vss 0.227f
C18831 vdd.n9558 vss 0.00324f
C18832 vdd.n9559 vss 0.0112f
C18833 vdd.n9560 vss 0.0128f
C18834 vdd.n9561 vss 0.00413f
C18835 vdd.n9562 vss 0.00413f
C18836 vdd.n9563 vss 0.0471f
C18837 vdd.n9564 vss 0.00251f
C18838 vdd.t984 vss 0.0471f
C18839 vdd.n9565 vss 0.00324f
C18840 vdd.n9567 vss 0.00679f
C18841 vdd.n9568 vss 0.00413f
C18842 vdd.n9569 vss 0.00324f
C18843 vdd.n9570 vss 0.00413f
C18844 vdd.n9571 vss 0.0471f
C18845 vdd.n9572 vss 0.00324f
C18846 vdd.n9574 vss 0.00925f
C18847 vdd.t237 vss 0.0471f
C18848 vdd.n9575 vss 0.00425f
C18849 vdd.n9576 vss 0.0424f
C18850 vdd.n9577 vss 0.0132f
C18851 vdd.n9578 vss 0.00324f
C18852 vdd.n9579 vss 0.0128f
C18853 vdd.n9580 vss 0.02f
C18854 vdd.n9581 vss 0.00425f
C18855 vdd.n9582 vss 0.00413f
C18856 vdd.n9583 vss 0.00251f
C18857 vdd.t1113 vss 0.0471f
C18858 vdd.n9584 vss 0.00251f
C18859 vdd.n9585 vss 0.00517f
C18860 vdd.n9586 vss 0.00679f
C18861 vdd.n9587 vss 0.00517f
C18862 vdd.n9588 vss 0.00679f
C18863 vdd.n9589 vss 0.02f
C18864 vdd.n9590 vss 0.00425f
C18865 vdd.n9591 vss 0.0424f
C18866 vdd.n9592 vss 0.0132f
C18867 vdd.n9593 vss 0.00925f
C18868 vdd.n9594 vss 0.00425f
C18869 vdd.n9595 vss 0.00413f
C18870 vdd.n9596 vss 0.00324f
C18871 vdd.n9597 vss 0.0471f
C18872 vdd.t1114 vss 0.0471f
C18873 vdd.n9598 vss 0.00251f
C18874 vdd.n9599 vss 0.0112f
C18875 vdd.n9600 vss 0.0128f
C18876 vdd.n9601 vss 0.152f
C18877 vdd.n9602 vss 0.0393f
C18878 vdd.n9603 vss 0.0332f
C18879 vdd.n9604 vss 0.00324f
C18880 vdd.n9605 vss 0.0112f
C18881 vdd.n9606 vss 0.0128f
C18882 vdd.n9607 vss 0.00413f
C18883 vdd.n9608 vss 0.00413f
C18884 vdd.n9609 vss 0.0471f
C18885 vdd.n9610 vss 0.00251f
C18886 vdd.t26 vss 0.0471f
C18887 vdd.n9611 vss 0.00324f
C18888 vdd.n9613 vss 0.00679f
C18889 vdd.n9614 vss 0.00413f
C18890 vdd.n9615 vss 0.00324f
C18891 vdd.n9616 vss 0.00413f
C18892 vdd.n9617 vss 0.0471f
C18893 vdd.n9618 vss 0.00324f
C18894 vdd.n9620 vss 0.00925f
C18895 vdd.t706 vss 0.0471f
C18896 vdd.n9621 vss 0.00425f
C18897 vdd.n9622 vss 0.0424f
C18898 vdd.n9623 vss 0.0132f
C18899 vdd.n9624 vss 0.00324f
C18900 vdd.n9625 vss 0.0128f
C18901 vdd.n9626 vss 0.02f
C18902 vdd.n9627 vss 0.00425f
C18903 vdd.n9628 vss 0.00413f
C18904 vdd.n9629 vss 0.00251f
C18905 vdd.t912 vss 0.0471f
C18906 vdd.n9630 vss 0.00251f
C18907 vdd.n9631 vss 0.00517f
C18908 vdd.n9632 vss 0.00679f
C18909 vdd.n9633 vss 0.00517f
C18910 vdd.n9634 vss 0.00679f
C18911 vdd.n9635 vss 0.02f
C18912 vdd.n9636 vss 0.00425f
C18913 vdd.n9637 vss 0.0424f
C18914 vdd.n9638 vss 0.0132f
C18915 vdd.n9639 vss 0.00925f
C18916 vdd.n9640 vss 0.00425f
C18917 vdd.n9641 vss 0.00413f
C18918 vdd.n9642 vss 0.00324f
C18919 vdd.n9643 vss 0.0471f
C18920 vdd.t910 vss 0.0471f
C18921 vdd.n9644 vss 0.00251f
C18922 vdd.n9645 vss 0.0112f
C18923 vdd.n9646 vss 0.0128f
C18924 vdd.n9647 vss 0.221f
C18925 vdd.n9648 vss 0.0393f
C18926 vdd.n9649 vss 0.0332f
C18927 vdd.n9650 vss 0.00324f
C18928 vdd.n9651 vss 0.0112f
C18929 vdd.n9652 vss 0.0128f
C18930 vdd.n9653 vss 0.00413f
C18931 vdd.n9654 vss 0.00413f
C18932 vdd.n9655 vss 0.0471f
C18933 vdd.n9656 vss 0.00251f
C18934 vdd.t1354 vss 0.0471f
C18935 vdd.n9657 vss 0.00324f
C18936 vdd.n9659 vss 0.00679f
C18937 vdd.n9660 vss 0.00413f
C18938 vdd.n9661 vss 0.00324f
C18939 vdd.n9662 vss 0.00413f
C18940 vdd.n9663 vss 0.0471f
C18941 vdd.n9664 vss 0.00324f
C18942 vdd.n9666 vss 0.00925f
C18943 vdd.t1514 vss 0.0471f
C18944 vdd.n9667 vss 0.00425f
C18945 vdd.n9668 vss 0.0424f
C18946 vdd.n9669 vss 0.0132f
C18947 vdd.n9670 vss 0.00324f
C18948 vdd.n9671 vss 0.0128f
C18949 vdd.n9672 vss 0.02f
C18950 vdd.n9673 vss 0.00425f
C18951 vdd.n9674 vss 0.00413f
C18952 vdd.n9675 vss 0.00251f
C18953 vdd.t1511 vss 0.0471f
C18954 vdd.n9676 vss 0.00251f
C18955 vdd.n9677 vss 0.00517f
C18956 vdd.n9678 vss 0.00679f
C18957 vdd.n9679 vss 0.00517f
C18958 vdd.n9680 vss 0.00679f
C18959 vdd.n9681 vss 0.02f
C18960 vdd.n9682 vss 0.00425f
C18961 vdd.n9683 vss 0.0424f
C18962 vdd.n9684 vss 0.0132f
C18963 vdd.n9685 vss 0.00925f
C18964 vdd.n9686 vss 0.00425f
C18965 vdd.n9687 vss 0.00413f
C18966 vdd.n9688 vss 0.00324f
C18967 vdd.n9689 vss 0.0471f
C18968 vdd.t1512 vss 0.0471f
C18969 vdd.n9690 vss 0.00251f
C18970 vdd.n9691 vss 0.0112f
C18971 vdd.n9692 vss 0.0128f
C18972 vdd.t1513 vss 0.00134f
C18973 vdd.t1355 vss 0.0013f
C18974 vdd.n9693 vss 0.0332f
C18975 vdd.n9694 vss 0.0393f
C18976 vdd.n9695 vss 0.0418f
C18977 vdd.n9696 vss 0.00324f
C18978 vdd.n9697 vss 0.0112f
C18979 vdd.n9698 vss 0.0128f
C18980 vdd.n9699 vss 0.00413f
C18981 vdd.n9700 vss 0.00413f
C18982 vdd.n9701 vss 0.0471f
C18983 vdd.n9702 vss 0.00251f
C18984 vdd.t1322 vss 0.0471f
C18985 vdd.n9703 vss 0.00324f
C18986 vdd.n9705 vss 0.00679f
C18987 vdd.n9706 vss 0.00413f
C18988 vdd.n9707 vss 0.00324f
C18989 vdd.n9708 vss 0.00413f
C18990 vdd.n9709 vss 0.0471f
C18991 vdd.n9710 vss 0.00324f
C18992 vdd.n9712 vss 0.00925f
C18993 vdd.t71 vss 0.0471f
C18994 vdd.n9713 vss 0.00425f
C18995 vdd.n9714 vss 0.0424f
C18996 vdd.n9715 vss 0.0132f
C18997 vdd.n9716 vss 0.00324f
C18998 vdd.n9717 vss 0.0128f
C18999 vdd.n9718 vss 0.02f
C19000 vdd.n9719 vss 0.00425f
C19001 vdd.n9720 vss 0.00413f
C19002 vdd.n9721 vss 0.00251f
C19003 vdd.t1387 vss 0.0471f
C19004 vdd.n9722 vss 0.00251f
C19005 vdd.n9723 vss 0.00517f
C19006 vdd.n9724 vss 0.00679f
C19007 vdd.n9725 vss 0.00517f
C19008 vdd.n9726 vss 0.00679f
C19009 vdd.n9727 vss 0.02f
C19010 vdd.n9728 vss 0.00425f
C19011 vdd.n9729 vss 0.0424f
C19012 vdd.n9730 vss 0.0132f
C19013 vdd.n9731 vss 0.00925f
C19014 vdd.n9732 vss 0.00425f
C19015 vdd.n9733 vss 0.00413f
C19016 vdd.n9734 vss 0.00324f
C19017 vdd.n9735 vss 0.0471f
C19018 vdd.t1388 vss 0.0471f
C19019 vdd.n9736 vss 0.00251f
C19020 vdd.n9737 vss 0.0112f
C19021 vdd.n9738 vss 0.0128f
C19022 vdd.t1389 vss 0.00134f
C19023 vdd.t1323 vss 0.0013f
C19024 vdd.n9739 vss 0.0332f
C19025 vdd.n9740 vss 0.0393f
C19026 vdd.n9741 vss 0.0345f
C19027 vdd.n9742 vss 0.00335f
C19028 vdd.t1462 vss 0.0013f
C19029 vdd.n9743 vss 0.0309f
C19030 vdd.n9744 vss 0.00991f
C19031 vdd.n9745 vss 0.0424f
C19032 vdd.n9746 vss 0.00679f
C19033 vdd.n9747 vss 0.00413f
C19034 vdd.n9748 vss 0.0471f
C19035 vdd.n9749 vss 0.00251f
C19036 vdd.n9750 vss 0.00324f
C19037 vdd.n9751 vss 0.0128f
C19038 vdd.n9752 vss 0.00413f
C19039 vdd.n9753 vss 0.00413f
C19040 vdd.n9754 vss 0.0471f
C19041 vdd.n9755 vss 0.00251f
C19042 vdd.n9756 vss 0.00324f
C19043 vdd.n9757 vss 0.00413f
C19044 vdd.n9758 vss 0.00324f
C19045 vdd.n9759 vss 0.0132f
C19046 vdd.n9760 vss 0.0424f
C19047 vdd.n9761 vss 0.00324f
C19048 vdd.n9762 vss 0.00413f
C19049 vdd.n9763 vss 0.02f
C19050 vdd.n9764 vss 0.00425f
C19051 vdd.t964 vss 0.0471f
C19052 vdd.n9766 vss 0.00425f
C19053 vdd.n9767 vss 0.00925f
C19054 vdd.n9768 vss 0.00679f
C19055 vdd.n9769 vss 0.00517f
C19056 vdd.n9770 vss 0.00679f
C19057 vdd.n9771 vss 0.00517f
C19058 vdd.n9772 vss 0.00251f
C19059 vdd.t1364 vss 0.0471f
C19060 vdd.n9773 vss 0.0471f
C19061 vdd.t1363 vss 0.0471f
C19062 vdd.n9774 vss 0.00251f
C19063 vdd.n9775 vss 0.0105f
C19064 vdd.t1365 vss 0.00134f
C19065 vdd.n9776 vss 0.0393f
C19066 vdd.n9777 vss 0.0633f
C19067 vdd.n9778 vss 0.00805f
C19068 vdd.n9779 vss 0.0112f
C19069 vdd.n9780 vss 0.0128f
C19070 vdd.n9781 vss 0.00324f
C19071 vdd.n9782 vss 0.00324f
C19072 vdd.n9783 vss 0.00413f
C19073 vdd.n9784 vss 0.00425f
C19074 vdd.t1461 vss 0.0471f
C19075 vdd.n9786 vss 0.00425f
C19076 vdd.n9787 vss 0.00925f
C19077 vdd.n9788 vss 0.0107f
C19078 vdd.n9789 vss 0.0126f
C19079 vdd.n9790 vss 9.89e-19
C19080 vdd.n9791 vss 0.00163f
C19081 vdd.n9792 vss 0.00145f
C19082 vdd.n9793 vss 0.0271f
C19083 vdd.n9794 vss 0.00324f
C19084 vdd.n9795 vss 0.0112f
C19085 vdd.n9796 vss 0.0128f
C19086 vdd.n9797 vss 0.00413f
C19087 vdd.n9798 vss 0.00413f
C19088 vdd.n9799 vss 0.0471f
C19089 vdd.n9800 vss 0.00251f
C19090 vdd.t478 vss 0.0471f
C19091 vdd.n9801 vss 0.00324f
C19092 vdd.n9803 vss 0.00679f
C19093 vdd.n9804 vss 0.00413f
C19094 vdd.n9805 vss 0.00324f
C19095 vdd.n9806 vss 0.00413f
C19096 vdd.n9807 vss 0.0471f
C19097 vdd.n9808 vss 0.00324f
C19098 vdd.n9810 vss 0.00925f
C19099 vdd.t360 vss 0.0471f
C19100 vdd.n9811 vss 0.00425f
C19101 vdd.n9812 vss 0.0424f
C19102 vdd.n9813 vss 0.0132f
C19103 vdd.n9814 vss 0.00324f
C19104 vdd.n9815 vss 0.0128f
C19105 vdd.n9816 vss 0.02f
C19106 vdd.n9817 vss 0.00425f
C19107 vdd.n9818 vss 0.00413f
C19108 vdd.n9819 vss 0.00251f
C19109 vdd.t727 vss 0.0471f
C19110 vdd.n9820 vss 0.00251f
C19111 vdd.n9821 vss 0.00517f
C19112 vdd.n9822 vss 0.00679f
C19113 vdd.n9823 vss 0.00517f
C19114 vdd.n9824 vss 0.00679f
C19115 vdd.n9825 vss 0.02f
C19116 vdd.n9826 vss 0.00425f
C19117 vdd.n9827 vss 0.0424f
C19118 vdd.n9828 vss 0.0132f
C19119 vdd.n9829 vss 0.00925f
C19120 vdd.n9830 vss 0.00425f
C19121 vdd.n9831 vss 0.00413f
C19122 vdd.n9832 vss 0.00324f
C19123 vdd.n9833 vss 0.0471f
C19124 vdd.t725 vss 0.0471f
C19125 vdd.n9834 vss 0.00251f
C19126 vdd.n9835 vss 0.0112f
C19127 vdd.n9836 vss 0.0128f
C19128 vdd.t726 vss 0.00134f
C19129 vdd.t479 vss 0.0013f
C19130 vdd.n9837 vss 0.0332f
C19131 vdd.n9838 vss 0.0393f
C19132 vdd.n9839 vss 0.0418f
C19133 vdd.n9840 vss 0.00324f
C19134 vdd.n9841 vss 0.0112f
C19135 vdd.n9842 vss 0.0128f
C19136 vdd.n9843 vss 0.00413f
C19137 vdd.n9844 vss 0.00413f
C19138 vdd.n9845 vss 0.0471f
C19139 vdd.n9846 vss 0.00251f
C19140 vdd.t1059 vss 0.0471f
C19141 vdd.n9847 vss 0.00324f
C19142 vdd.n9849 vss 0.00679f
C19143 vdd.n9850 vss 0.00413f
C19144 vdd.n9851 vss 0.00324f
C19145 vdd.n9852 vss 0.00413f
C19146 vdd.n9853 vss 0.0471f
C19147 vdd.n9854 vss 0.00324f
C19148 vdd.n9856 vss 0.00925f
C19149 vdd.t1284 vss 0.0471f
C19150 vdd.n9857 vss 0.00425f
C19151 vdd.n9858 vss 0.0424f
C19152 vdd.n9859 vss 0.0132f
C19153 vdd.n9860 vss 0.00324f
C19154 vdd.n9861 vss 0.0128f
C19155 vdd.n9862 vss 0.02f
C19156 vdd.n9863 vss 0.00425f
C19157 vdd.n9864 vss 0.00413f
C19158 vdd.n9865 vss 0.00251f
C19159 vdd.t1179 vss 0.0471f
C19160 vdd.n9866 vss 0.00251f
C19161 vdd.n9867 vss 0.00517f
C19162 vdd.n9868 vss 0.00679f
C19163 vdd.n9869 vss 0.00517f
C19164 vdd.n9870 vss 0.00679f
C19165 vdd.n9871 vss 0.02f
C19166 vdd.n9872 vss 0.00425f
C19167 vdd.n9873 vss 0.0424f
C19168 vdd.n9874 vss 0.0132f
C19169 vdd.n9875 vss 0.00925f
C19170 vdd.n9876 vss 0.00425f
C19171 vdd.n9877 vss 0.00413f
C19172 vdd.n9878 vss 0.00324f
C19173 vdd.n9879 vss 0.0471f
C19174 vdd.t1180 vss 0.0471f
C19175 vdd.n9880 vss 0.00251f
C19176 vdd.n9881 vss 0.0112f
C19177 vdd.n9882 vss 0.0128f
C19178 vdd.t1181 vss 0.00134f
C19179 vdd.t1060 vss 0.0013f
C19180 vdd.n9883 vss 0.0332f
C19181 vdd.n9884 vss 0.0393f
C19182 vdd.n9885 vss 0.0345f
C19183 vdd.n9886 vss 0.00324f
C19184 vdd.n9887 vss 0.0112f
C19185 vdd.n9888 vss 0.0128f
C19186 vdd.n9889 vss 0.00413f
C19187 vdd.n9890 vss 0.00413f
C19188 vdd.n9891 vss 0.0471f
C19189 vdd.n9892 vss 0.00251f
C19190 vdd.t15 vss 0.0471f
C19191 vdd.n9893 vss 0.00324f
C19192 vdd.n9895 vss 0.00679f
C19193 vdd.n9896 vss 0.00413f
C19194 vdd.n9897 vss 0.00324f
C19195 vdd.n9898 vss 0.00413f
C19196 vdd.n9899 vss 0.0471f
C19197 vdd.n9900 vss 0.00324f
C19198 vdd.n9902 vss 0.00925f
C19199 vdd.t1023 vss 0.0471f
C19200 vdd.n9903 vss 0.00425f
C19201 vdd.n9904 vss 0.0424f
C19202 vdd.n9905 vss 0.0132f
C19203 vdd.n9906 vss 0.00324f
C19204 vdd.n9907 vss 0.0128f
C19205 vdd.n9908 vss 0.02f
C19206 vdd.n9909 vss 0.00425f
C19207 vdd.n9910 vss 0.00413f
C19208 vdd.n9911 vss 0.00251f
C19209 vdd.t259 vss 0.0471f
C19210 vdd.n9912 vss 0.00251f
C19211 vdd.n9913 vss 0.00517f
C19212 vdd.n9914 vss 0.00679f
C19213 vdd.n9915 vss 0.00517f
C19214 vdd.n9916 vss 0.00679f
C19215 vdd.n9917 vss 0.02f
C19216 vdd.n9918 vss 0.00425f
C19217 vdd.n9919 vss 0.0424f
C19218 vdd.n9920 vss 0.0132f
C19219 vdd.n9921 vss 0.00925f
C19220 vdd.n9922 vss 0.00425f
C19221 vdd.n9923 vss 0.00413f
C19222 vdd.n9924 vss 0.00324f
C19223 vdd.n9925 vss 0.0471f
C19224 vdd.t257 vss 0.0471f
C19225 vdd.n9926 vss 0.00251f
C19226 vdd.n9927 vss 0.0112f
C19227 vdd.n9928 vss 0.0128f
C19228 vdd.t258 vss 0.00134f
C19229 vdd.t16 vss 0.0013f
C19230 vdd.n9929 vss 0.0332f
C19231 vdd.n9930 vss 0.0393f
C19232 vdd.n9931 vss 0.0418f
C19233 vdd.n9932 vss 0.00324f
C19234 vdd.n9933 vss 0.0112f
C19235 vdd.n9934 vss 0.0128f
C19236 vdd.n9935 vss 0.00413f
C19237 vdd.n9936 vss 0.00413f
C19238 vdd.n9937 vss 0.0471f
C19239 vdd.n9938 vss 0.00251f
C19240 vdd.t490 vss 0.0471f
C19241 vdd.n9939 vss 0.00324f
C19242 vdd.n9941 vss 0.00679f
C19243 vdd.n9942 vss 0.00413f
C19244 vdd.n9943 vss 0.00324f
C19245 vdd.n9944 vss 0.00413f
C19246 vdd.n9945 vss 0.0471f
C19247 vdd.n9946 vss 0.00324f
C19248 vdd.n9948 vss 0.00925f
C19249 vdd.t960 vss 0.0471f
C19250 vdd.n9949 vss 0.00425f
C19251 vdd.n9950 vss 0.0424f
C19252 vdd.n9951 vss 0.0132f
C19253 vdd.n9952 vss 0.00324f
C19254 vdd.n9953 vss 0.0128f
C19255 vdd.n9954 vss 0.02f
C19256 vdd.n9955 vss 0.00425f
C19257 vdd.n9956 vss 0.00413f
C19258 vdd.n9957 vss 0.00251f
C19259 vdd.t62 vss 0.0471f
C19260 vdd.n9958 vss 0.00251f
C19261 vdd.n9959 vss 0.00517f
C19262 vdd.n9960 vss 0.00679f
C19263 vdd.n9961 vss 0.00517f
C19264 vdd.n9962 vss 0.00679f
C19265 vdd.n9963 vss 0.02f
C19266 vdd.n9964 vss 0.00425f
C19267 vdd.n9965 vss 0.0424f
C19268 vdd.n9966 vss 0.0132f
C19269 vdd.n9967 vss 0.00925f
C19270 vdd.n9968 vss 0.00425f
C19271 vdd.n9969 vss 0.00413f
C19272 vdd.n9970 vss 0.00324f
C19273 vdd.n9971 vss 0.0471f
C19274 vdd.t60 vss 0.0471f
C19275 vdd.n9972 vss 0.00251f
C19276 vdd.n9973 vss 0.0112f
C19277 vdd.n9974 vss 0.0128f
C19278 vdd.t61 vss 0.00134f
C19279 vdd.t491 vss 0.0013f
C19280 vdd.n9975 vss 0.0332f
C19281 vdd.n9976 vss 0.0393f
C19282 vdd.n9977 vss 0.0345f
C19283 vdd.n9978 vss 0.00335f
C19284 vdd.t576 vss 0.0013f
C19285 vdd.n9979 vss 0.0309f
C19286 vdd.n9980 vss 0.00991f
C19287 vdd.n9981 vss 0.0424f
C19288 vdd.n9982 vss 0.00679f
C19289 vdd.n9983 vss 0.00413f
C19290 vdd.n9984 vss 0.0471f
C19291 vdd.n9985 vss 0.00251f
C19292 vdd.n9986 vss 0.00324f
C19293 vdd.n9987 vss 0.0128f
C19294 vdd.n9988 vss 0.00413f
C19295 vdd.n9989 vss 0.00413f
C19296 vdd.n9990 vss 0.0471f
C19297 vdd.n9991 vss 0.00251f
C19298 vdd.n9992 vss 0.00324f
C19299 vdd.n9993 vss 0.00413f
C19300 vdd.n9994 vss 0.00324f
C19301 vdd.n9995 vss 0.0132f
C19302 vdd.n9996 vss 0.0424f
C19303 vdd.n9997 vss 0.00324f
C19304 vdd.n9998 vss 0.00413f
C19305 vdd.n9999 vss 0.02f
C19306 vdd.n10000 vss 0.00425f
C19307 vdd.t694 vss 0.0471f
C19308 vdd.n10002 vss 0.00425f
C19309 vdd.n10003 vss 0.00925f
C19310 vdd.n10004 vss 0.00679f
C19311 vdd.n10005 vss 0.00517f
C19312 vdd.n10006 vss 0.00679f
C19313 vdd.n10007 vss 0.00517f
C19314 vdd.n10008 vss 0.00251f
C19315 vdd.t1398 vss 0.0471f
C19316 vdd.n10009 vss 0.0471f
C19317 vdd.t1397 vss 0.0471f
C19318 vdd.n10010 vss 0.00251f
C19319 vdd.n10011 vss 0.0105f
C19320 vdd.t1399 vss 0.00134f
C19321 vdd.n10012 vss 0.0393f
C19322 vdd.n10013 vss 0.0633f
C19323 vdd.n10014 vss 0.00805f
C19324 vdd.n10015 vss 0.0112f
C19325 vdd.n10016 vss 0.0128f
C19326 vdd.n10017 vss 0.00324f
C19327 vdd.n10018 vss 0.00324f
C19328 vdd.n10019 vss 0.00413f
C19329 vdd.n10020 vss 0.00425f
C19330 vdd.t575 vss 0.0471f
C19331 vdd.n10022 vss 0.00425f
C19332 vdd.n10023 vss 0.00925f
C19333 vdd.n10024 vss 0.0107f
C19334 vdd.n10025 vss 0.0126f
C19335 vdd.n10026 vss 9.89e-19
C19336 vdd.n10027 vss 0.00163f
C19337 vdd.n10028 vss 0.00145f
C19338 vdd.n10029 vss 0.0271f
C19339 vdd.n10030 vss 0.00324f
C19340 vdd.n10031 vss 0.0112f
C19341 vdd.n10032 vss 0.0128f
C19342 vdd.n10033 vss 0.00413f
C19343 vdd.n10034 vss 0.00413f
C19344 vdd.n10035 vss 0.0471f
C19345 vdd.n10036 vss 0.00251f
C19346 vdd.t1334 vss 0.0471f
C19347 vdd.n10037 vss 0.00324f
C19348 vdd.n10039 vss 0.00679f
C19349 vdd.n10040 vss 0.00413f
C19350 vdd.n10041 vss 0.00324f
C19351 vdd.n10042 vss 0.00413f
C19352 vdd.n10043 vss 0.0471f
C19353 vdd.n10044 vss 0.00324f
C19354 vdd.n10046 vss 0.00925f
C19355 vdd.t548 vss 0.0471f
C19356 vdd.n10047 vss 0.00425f
C19357 vdd.n10048 vss 0.0424f
C19358 vdd.n10049 vss 0.0132f
C19359 vdd.n10050 vss 0.00324f
C19360 vdd.n10051 vss 0.0128f
C19361 vdd.n10052 vss 0.02f
C19362 vdd.n10053 vss 0.00425f
C19363 vdd.n10054 vss 0.00413f
C19364 vdd.n10055 vss 0.00251f
C19365 vdd.t337 vss 0.0471f
C19366 vdd.n10056 vss 0.00251f
C19367 vdd.n10057 vss 0.00517f
C19368 vdd.n10058 vss 0.00679f
C19369 vdd.n10059 vss 0.00517f
C19370 vdd.n10060 vss 0.00679f
C19371 vdd.n10061 vss 0.02f
C19372 vdd.n10062 vss 0.00425f
C19373 vdd.n10063 vss 0.0424f
C19374 vdd.n10064 vss 0.0132f
C19375 vdd.n10065 vss 0.00925f
C19376 vdd.n10066 vss 0.00425f
C19377 vdd.n10067 vss 0.00413f
C19378 vdd.n10068 vss 0.00324f
C19379 vdd.n10069 vss 0.0471f
C19380 vdd.t338 vss 0.0471f
C19381 vdd.n10070 vss 0.00251f
C19382 vdd.n10071 vss 0.0112f
C19383 vdd.n10072 vss 0.0128f
C19384 vdd.t339 vss 0.00134f
C19385 vdd.t1335 vss 0.0013f
C19386 vdd.n10073 vss 0.0332f
C19387 vdd.n10074 vss 0.0393f
C19388 vdd.n10075 vss 0.0418f
C19389 vdd.n10076 vss 0.00324f
C19390 vdd.n10077 vss 0.0112f
C19391 vdd.n10078 vss 0.0128f
C19392 vdd.n10079 vss 0.00413f
C19393 vdd.n10080 vss 0.00413f
C19394 vdd.n10081 vss 0.0471f
C19395 vdd.n10082 vss 0.00251f
C19396 vdd.t568 vss 0.0471f
C19397 vdd.n10083 vss 0.00324f
C19398 vdd.n10085 vss 0.00679f
C19399 vdd.n10086 vss 0.00413f
C19400 vdd.n10087 vss 0.00324f
C19401 vdd.n10088 vss 0.00413f
C19402 vdd.n10089 vss 0.0471f
C19403 vdd.n10090 vss 0.00324f
C19404 vdd.n10092 vss 0.00925f
C19405 vdd.t1164 vss 0.0471f
C19406 vdd.n10093 vss 0.00425f
C19407 vdd.n10094 vss 0.0424f
C19408 vdd.n10095 vss 0.0132f
C19409 vdd.n10096 vss 0.00324f
C19410 vdd.n10097 vss 0.0128f
C19411 vdd.n10098 vss 0.02f
C19412 vdd.n10099 vss 0.00425f
C19413 vdd.n10100 vss 0.00413f
C19414 vdd.n10101 vss 0.00251f
C19415 vdd.t1087 vss 0.0471f
C19416 vdd.n10102 vss 0.00251f
C19417 vdd.n10103 vss 0.00517f
C19418 vdd.n10104 vss 0.00679f
C19419 vdd.n10105 vss 0.00517f
C19420 vdd.n10106 vss 0.00679f
C19421 vdd.n10107 vss 0.02f
C19422 vdd.n10108 vss 0.00425f
C19423 vdd.n10109 vss 0.0424f
C19424 vdd.n10110 vss 0.0132f
C19425 vdd.n10111 vss 0.00925f
C19426 vdd.n10112 vss 0.00425f
C19427 vdd.n10113 vss 0.00413f
C19428 vdd.n10114 vss 0.00324f
C19429 vdd.n10115 vss 0.0471f
C19430 vdd.t1085 vss 0.0471f
C19431 vdd.n10116 vss 0.00251f
C19432 vdd.n10117 vss 0.0112f
C19433 vdd.n10118 vss 0.0128f
C19434 vdd.t1086 vss 0.00134f
C19435 vdd.t569 vss 0.0013f
C19436 vdd.n10119 vss 0.0332f
C19437 vdd.n10120 vss 0.0393f
C19438 vdd.n10121 vss 0.0418f
C19439 vdd.n10122 vss 0.118f
C19440 vdd.n10123 vss 0.121f
C19441 vdd.t909 vss 0.0013f
C19442 vdd.t782 vss 0.00134f
C19443 vdd.n10124 vss 0.00324f
C19444 vdd.n10125 vss 0.0112f
C19445 vdd.n10126 vss 0.0128f
C19446 vdd.n10127 vss 0.00413f
C19447 vdd.n10128 vss 0.00413f
C19448 vdd.n10129 vss 0.0471f
C19449 vdd.n10130 vss 0.00251f
C19450 vdd.t908 vss 0.0471f
C19451 vdd.n10131 vss 0.00324f
C19452 vdd.n10133 vss 0.00679f
C19453 vdd.n10134 vss 0.00413f
C19454 vdd.n10135 vss 0.00324f
C19455 vdd.n10136 vss 0.00413f
C19456 vdd.n10137 vss 0.0471f
C19457 vdd.n10138 vss 0.00324f
C19458 vdd.n10140 vss 0.00925f
C19459 vdd.t1438 vss 0.0471f
C19460 vdd.n10141 vss 0.00425f
C19461 vdd.n10142 vss 0.0424f
C19462 vdd.n10143 vss 0.0132f
C19463 vdd.n10144 vss 0.00324f
C19464 vdd.n10145 vss 0.0128f
C19465 vdd.n10146 vss 0.02f
C19466 vdd.n10147 vss 0.00425f
C19467 vdd.n10148 vss 0.00413f
C19468 vdd.n10149 vss 0.00251f
C19469 vdd.t780 vss 0.0471f
C19470 vdd.n10150 vss 0.00251f
C19471 vdd.n10151 vss 0.00517f
C19472 vdd.n10152 vss 0.00679f
C19473 vdd.n10153 vss 0.00517f
C19474 vdd.n10154 vss 0.00679f
C19475 vdd.n10155 vss 0.02f
C19476 vdd.n10156 vss 0.00425f
C19477 vdd.n10157 vss 0.0424f
C19478 vdd.n10158 vss 0.0132f
C19479 vdd.n10159 vss 0.00925f
C19480 vdd.n10160 vss 0.00425f
C19481 vdd.n10161 vss 0.00413f
C19482 vdd.n10162 vss 0.00324f
C19483 vdd.n10163 vss 0.0471f
C19484 vdd.t781 vss 0.0471f
C19485 vdd.n10164 vss 0.00251f
C19486 vdd.n10165 vss 0.0112f
C19487 vdd.n10166 vss 0.0707f
C19488 vdd.n10167 vss 0.0393f
C19489 vdd.n10168 vss 0.0332f
C19490 vdd.n10169 vss 0.0596f
C19491 vdd.n10170 vss 0.00324f
C19492 vdd.n10171 vss 0.0112f
C19493 vdd.n10172 vss 0.0128f
C19494 vdd.n10173 vss 0.00413f
C19495 vdd.n10174 vss 0.00413f
C19496 vdd.n10175 vss 0.0471f
C19497 vdd.n10176 vss 0.00251f
C19498 vdd.t597 vss 0.0471f
C19499 vdd.n10177 vss 0.00324f
C19500 vdd.n10179 vss 0.00679f
C19501 vdd.n10180 vss 0.00413f
C19502 vdd.n10181 vss 0.00324f
C19503 vdd.n10182 vss 0.00413f
C19504 vdd.n10183 vss 0.0471f
C19505 vdd.n10184 vss 0.00324f
C19506 vdd.n10186 vss 0.00925f
C19507 vdd.t418 vss 0.0471f
C19508 vdd.n10187 vss 0.00425f
C19509 vdd.n10188 vss 0.0424f
C19510 vdd.n10189 vss 0.0132f
C19511 vdd.n10190 vss 0.00324f
C19512 vdd.n10191 vss 0.0128f
C19513 vdd.n10192 vss 0.02f
C19514 vdd.n10193 vss 0.00425f
C19515 vdd.n10194 vss 0.00413f
C19516 vdd.n10195 vss 0.00251f
C19517 vdd.t1020 vss 0.0471f
C19518 vdd.n10196 vss 0.00251f
C19519 vdd.n10197 vss 0.00517f
C19520 vdd.n10198 vss 0.00679f
C19521 vdd.n10199 vss 0.00517f
C19522 vdd.n10200 vss 0.00679f
C19523 vdd.n10201 vss 0.02f
C19524 vdd.n10202 vss 0.00425f
C19525 vdd.n10203 vss 0.0424f
C19526 vdd.n10204 vss 0.0132f
C19527 vdd.n10205 vss 0.00925f
C19528 vdd.n10206 vss 0.00425f
C19529 vdd.n10207 vss 0.00413f
C19530 vdd.n10208 vss 0.00324f
C19531 vdd.n10209 vss 0.0471f
C19532 vdd.t1021 vss 0.0471f
C19533 vdd.n10210 vss 0.00251f
C19534 vdd.n10211 vss 0.0112f
C19535 vdd.n10212 vss 0.0128f
C19536 vdd.t1022 vss 0.00134f
C19537 vdd.t598 vss 0.0013f
C19538 vdd.n10213 vss 0.0332f
C19539 vdd.n10214 vss 0.0393f
C19540 vdd.n10215 vss 0.0418f
C19541 vdd.n10216 vss 0.0912f
C19542 vdd.n10217 vss 0.0824f
C19543 vdd.n10218 vss 0.059f
C19544 vdd.t939 vss 0.0013f
C19545 vdd.t689 vss 0.00134f
C19546 vdd.n10219 vss 0.00324f
C19547 vdd.n10220 vss 0.0112f
C19548 vdd.n10221 vss 0.0128f
C19549 vdd.n10222 vss 0.00413f
C19550 vdd.n10223 vss 0.00413f
C19551 vdd.n10224 vss 0.0471f
C19552 vdd.n10225 vss 0.00251f
C19553 vdd.t1379 vss 0.0471f
C19554 vdd.n10226 vss 0.00324f
C19555 vdd.n10228 vss 0.00679f
C19556 vdd.n10229 vss 0.00413f
C19557 vdd.n10230 vss 0.00324f
C19558 vdd.n10231 vss 0.00413f
C19559 vdd.n10232 vss 0.0471f
C19560 vdd.n10233 vss 0.00324f
C19561 vdd.n10235 vss 0.00925f
C19562 vdd.t659 vss 0.0471f
C19563 vdd.n10236 vss 0.00425f
C19564 vdd.n10237 vss 0.0424f
C19565 vdd.n10238 vss 0.0132f
C19566 vdd.n10239 vss 0.00324f
C19567 vdd.n10240 vss 0.0128f
C19568 vdd.n10241 vss 0.02f
C19569 vdd.n10242 vss 0.00425f
C19570 vdd.n10243 vss 0.00413f
C19571 vdd.n10244 vss 0.00251f
C19572 vdd.t1416 vss 0.0471f
C19573 vdd.n10245 vss 0.00251f
C19574 vdd.n10246 vss 0.00517f
C19575 vdd.n10247 vss 0.00679f
C19576 vdd.n10248 vss 0.00517f
C19577 vdd.n10249 vss 0.00679f
C19578 vdd.n10250 vss 0.02f
C19579 vdd.n10251 vss 0.00425f
C19580 vdd.n10252 vss 0.0424f
C19581 vdd.n10253 vss 0.0132f
C19582 vdd.n10254 vss 0.00925f
C19583 vdd.n10255 vss 0.00425f
C19584 vdd.n10256 vss 0.00413f
C19585 vdd.n10257 vss 0.00324f
C19586 vdd.n10258 vss 0.0471f
C19587 vdd.t1417 vss 0.0471f
C19588 vdd.n10259 vss 0.00251f
C19589 vdd.n10260 vss 0.0112f
C19590 vdd.n10261 vss 0.0128f
C19591 vdd.t1418 vss 0.00134f
C19592 vdd.t1380 vss 0.0013f
C19593 vdd.n10262 vss 0.0332f
C19594 vdd.n10263 vss 0.0393f
C19595 vdd.n10264 vss 0.158f
C19596 vdd.n10265 vss 0.00324f
C19597 vdd.n10266 vss 0.0112f
C19598 vdd.n10267 vss 0.0128f
C19599 vdd.n10268 vss 0.00413f
C19600 vdd.n10269 vss 0.00413f
C19601 vdd.n10270 vss 0.0471f
C19602 vdd.n10271 vss 0.00251f
C19603 vdd.t54 vss 0.0471f
C19604 vdd.n10272 vss 0.00324f
C19605 vdd.n10274 vss 0.00679f
C19606 vdd.n10275 vss 0.00413f
C19607 vdd.n10276 vss 0.00324f
C19608 vdd.n10277 vss 0.00413f
C19609 vdd.n10278 vss 0.0471f
C19610 vdd.n10279 vss 0.00324f
C19611 vdd.n10281 vss 0.00925f
C19612 vdd.t502 vss 0.0471f
C19613 vdd.n10282 vss 0.00425f
C19614 vdd.n10283 vss 0.0424f
C19615 vdd.n10284 vss 0.0132f
C19616 vdd.n10285 vss 0.00324f
C19617 vdd.n10286 vss 0.0128f
C19618 vdd.n10287 vss 0.02f
C19619 vdd.n10288 vss 0.00425f
C19620 vdd.n10289 vss 0.00413f
C19621 vdd.n10290 vss 0.00251f
C19622 vdd.t299 vss 0.0471f
C19623 vdd.n10291 vss 0.00251f
C19624 vdd.n10292 vss 0.00517f
C19625 vdd.n10293 vss 0.00679f
C19626 vdd.n10294 vss 0.00517f
C19627 vdd.n10295 vss 0.00679f
C19628 vdd.n10296 vss 0.02f
C19629 vdd.n10297 vss 0.00425f
C19630 vdd.n10298 vss 0.0424f
C19631 vdd.n10299 vss 0.0132f
C19632 vdd.n10300 vss 0.00925f
C19633 vdd.n10301 vss 0.00425f
C19634 vdd.n10302 vss 0.00413f
C19635 vdd.n10303 vss 0.00324f
C19636 vdd.n10304 vss 0.0471f
C19637 vdd.t300 vss 0.0471f
C19638 vdd.n10305 vss 0.00251f
C19639 vdd.n10306 vss 0.0112f
C19640 vdd.n10307 vss 0.0128f
C19641 vdd.t301 vss 0.00134f
C19642 vdd.t55 vss 0.0013f
C19643 vdd.n10308 vss 0.0332f
C19644 vdd.n10309 vss 0.0393f
C19645 vdd.n10310 vss 0.0316f
C19646 vdd.n10311 vss 0.256f
C19647 vdd.n10312 vss 0.00324f
C19648 vdd.n10313 vss 0.0112f
C19649 vdd.n10314 vss 0.0128f
C19650 vdd.n10315 vss 0.00413f
C19651 vdd.n10316 vss 0.00413f
C19652 vdd.n10317 vss 0.0471f
C19653 vdd.n10318 vss 0.00251f
C19654 vdd.t938 vss 0.0471f
C19655 vdd.n10319 vss 0.00324f
C19656 vdd.n10321 vss 0.00679f
C19657 vdd.n10322 vss 0.00413f
C19658 vdd.n10323 vss 0.00324f
C19659 vdd.n10324 vss 0.00413f
C19660 vdd.n10325 vss 0.0471f
C19661 vdd.n10326 vss 0.00324f
C19662 vdd.n10328 vss 0.00925f
C19663 vdd.t702 vss 0.0471f
C19664 vdd.n10329 vss 0.00425f
C19665 vdd.n10330 vss 0.0424f
C19666 vdd.n10331 vss 0.0132f
C19667 vdd.n10332 vss 0.00324f
C19668 vdd.n10333 vss 0.0128f
C19669 vdd.n10334 vss 0.02f
C19670 vdd.n10335 vss 0.00425f
C19671 vdd.n10336 vss 0.00413f
C19672 vdd.n10337 vss 0.00251f
C19673 vdd.t687 vss 0.0471f
C19674 vdd.n10338 vss 0.00251f
C19675 vdd.n10339 vss 0.00517f
C19676 vdd.n10340 vss 0.00679f
C19677 vdd.n10341 vss 0.00517f
C19678 vdd.n10342 vss 0.00679f
C19679 vdd.n10343 vss 0.02f
C19680 vdd.n10344 vss 0.00425f
C19681 vdd.n10345 vss 0.0424f
C19682 vdd.n10346 vss 0.0132f
C19683 vdd.n10347 vss 0.00925f
C19684 vdd.n10348 vss 0.00425f
C19685 vdd.n10349 vss 0.00413f
C19686 vdd.n10350 vss 0.00324f
C19687 vdd.n10351 vss 0.0471f
C19688 vdd.t688 vss 0.0471f
C19689 vdd.n10352 vss 0.00251f
C19690 vdd.n10353 vss 0.0112f
C19691 vdd.n10354 vss 0.0128f
C19692 vdd.n10355 vss 0.0953f
C19693 vdd.n10356 vss 0.0393f
C19694 vdd.n10357 vss 0.0332f
C19695 vdd.n10358 vss 0.0596f
C19696 vdd.n10359 vss 0.00324f
C19697 vdd.n10360 vss 0.0112f
C19698 vdd.n10361 vss 0.0128f
C19699 vdd.n10362 vss 0.00413f
C19700 vdd.n10363 vss 0.00413f
C19701 vdd.n10364 vss 0.0471f
C19702 vdd.n10365 vss 0.00251f
C19703 vdd.t383 vss 0.0471f
C19704 vdd.n10366 vss 0.00324f
C19705 vdd.n10368 vss 0.00679f
C19706 vdd.n10369 vss 0.00413f
C19707 vdd.n10370 vss 0.00324f
C19708 vdd.n10371 vss 0.00413f
C19709 vdd.n10372 vss 0.0471f
C19710 vdd.n10373 vss 0.00324f
C19711 vdd.n10375 vss 0.00925f
C19712 vdd.t1138 vss 0.0471f
C19713 vdd.n10376 vss 0.00425f
C19714 vdd.n10377 vss 0.0424f
C19715 vdd.n10378 vss 0.0132f
C19716 vdd.n10379 vss 0.00324f
C19717 vdd.n10380 vss 0.0128f
C19718 vdd.n10381 vss 0.02f
C19719 vdd.n10382 vss 0.00425f
C19720 vdd.n10383 vss 0.00413f
C19721 vdd.n10384 vss 0.00251f
C19722 vdd.t354 vss 0.0471f
C19723 vdd.n10385 vss 0.00251f
C19724 vdd.n10386 vss 0.00517f
C19725 vdd.n10387 vss 0.00679f
C19726 vdd.n10388 vss 0.00517f
C19727 vdd.n10389 vss 0.00679f
C19728 vdd.n10390 vss 0.02f
C19729 vdd.n10391 vss 0.00425f
C19730 vdd.n10392 vss 0.0424f
C19731 vdd.n10393 vss 0.0132f
C19732 vdd.n10394 vss 0.00925f
C19733 vdd.n10395 vss 0.00425f
C19734 vdd.n10396 vss 0.00413f
C19735 vdd.n10397 vss 0.00324f
C19736 vdd.n10398 vss 0.0471f
C19737 vdd.t355 vss 0.0471f
C19738 vdd.n10399 vss 0.00251f
C19739 vdd.n10400 vss 0.0112f
C19740 vdd.n10401 vss 0.0128f
C19741 vdd.t356 vss 0.00134f
C19742 vdd.t384 vss 0.0013f
C19743 vdd.n10402 vss 0.0332f
C19744 vdd.n10403 vss 0.0393f
C19745 vdd.n10404 vss 0.0418f
C19746 vdd.n10405 vss 0.118f
C19747 vdd.n10406 vss 0.121f
C19748 vdd.t847 vss 0.0013f
C19749 vdd.t1402 vss 0.00134f
C19750 vdd.n10407 vss 0.00324f
C19751 vdd.n10408 vss 0.0112f
C19752 vdd.n10409 vss 0.0128f
C19753 vdd.n10410 vss 0.00413f
C19754 vdd.n10411 vss 0.00413f
C19755 vdd.n10412 vss 0.0471f
C19756 vdd.n10413 vss 0.00251f
C19757 vdd.t846 vss 0.0471f
C19758 vdd.n10414 vss 0.00324f
C19759 vdd.n10416 vss 0.00679f
C19760 vdd.n10417 vss 0.00413f
C19761 vdd.n10418 vss 0.00324f
C19762 vdd.n10419 vss 0.00413f
C19763 vdd.n10420 vss 0.0471f
C19764 vdd.n10421 vss 0.00324f
C19765 vdd.n10423 vss 0.00925f
C19766 vdd.t1454 vss 0.0471f
C19767 vdd.n10424 vss 0.00425f
C19768 vdd.n10425 vss 0.0424f
C19769 vdd.n10426 vss 0.0132f
C19770 vdd.n10427 vss 0.00324f
C19771 vdd.n10428 vss 0.0128f
C19772 vdd.n10429 vss 0.02f
C19773 vdd.n10430 vss 0.00425f
C19774 vdd.n10431 vss 0.00413f
C19775 vdd.n10432 vss 0.00251f
C19776 vdd.t1400 vss 0.0471f
C19777 vdd.n10433 vss 0.00251f
C19778 vdd.n10434 vss 0.00517f
C19779 vdd.n10435 vss 0.00679f
C19780 vdd.n10436 vss 0.00517f
C19781 vdd.n10437 vss 0.00679f
C19782 vdd.n10438 vss 0.02f
C19783 vdd.n10439 vss 0.00425f
C19784 vdd.n10440 vss 0.0424f
C19785 vdd.n10441 vss 0.0132f
C19786 vdd.n10442 vss 0.00925f
C19787 vdd.n10443 vss 0.00425f
C19788 vdd.n10444 vss 0.00413f
C19789 vdd.n10445 vss 0.00324f
C19790 vdd.n10446 vss 0.0471f
C19791 vdd.t1401 vss 0.0471f
C19792 vdd.n10447 vss 0.00251f
C19793 vdd.n10448 vss 0.0112f
C19794 vdd.n10449 vss 0.0707f
C19795 vdd.n10450 vss 0.0393f
C19796 vdd.n10451 vss 0.0332f
C19797 vdd.n10452 vss 0.0596f
C19798 vdd.n10453 vss 0.00324f
C19799 vdd.n10454 vss 0.0112f
C19800 vdd.n10455 vss 0.0128f
C19801 vdd.n10456 vss 0.00413f
C19802 vdd.n10457 vss 0.00413f
C19803 vdd.n10458 vss 0.0471f
C19804 vdd.n10459 vss 0.00251f
C19805 vdd.t1306 vss 0.0471f
C19806 vdd.n10460 vss 0.00324f
C19807 vdd.n10462 vss 0.00679f
C19808 vdd.n10463 vss 0.00413f
C19809 vdd.n10464 vss 0.00324f
C19810 vdd.n10465 vss 0.00413f
C19811 vdd.n10466 vss 0.0471f
C19812 vdd.n10467 vss 0.00324f
C19813 vdd.n10469 vss 0.00925f
C19814 vdd.t1257 vss 0.0471f
C19815 vdd.n10470 vss 0.00425f
C19816 vdd.n10471 vss 0.0424f
C19817 vdd.n10472 vss 0.0132f
C19818 vdd.n10473 vss 0.00324f
C19819 vdd.n10474 vss 0.0128f
C19820 vdd.n10475 vss 0.02f
C19821 vdd.n10476 vss 0.00425f
C19822 vdd.n10477 vss 0.00413f
C19823 vdd.n10478 vss 0.00251f
C19824 vdd.t803 vss 0.0471f
C19825 vdd.n10479 vss 0.00251f
C19826 vdd.n10480 vss 0.00517f
C19827 vdd.n10481 vss 0.00679f
C19828 vdd.n10482 vss 0.00517f
C19829 vdd.n10483 vss 0.00679f
C19830 vdd.n10484 vss 0.02f
C19831 vdd.n10485 vss 0.00425f
C19832 vdd.n10486 vss 0.0424f
C19833 vdd.n10487 vss 0.0132f
C19834 vdd.n10488 vss 0.00925f
C19835 vdd.n10489 vss 0.00425f
C19836 vdd.n10490 vss 0.00413f
C19837 vdd.n10491 vss 0.00324f
C19838 vdd.n10492 vss 0.0471f
C19839 vdd.t804 vss 0.0471f
C19840 vdd.n10493 vss 0.00251f
C19841 vdd.n10494 vss 0.0112f
C19842 vdd.n10495 vss 0.0128f
C19843 vdd.t805 vss 0.00134f
C19844 vdd.t1307 vss 0.0013f
C19845 vdd.n10496 vss 0.0332f
C19846 vdd.n10497 vss 0.0393f
C19847 vdd.n10498 vss 0.0418f
C19848 vdd.n10499 vss 0.118f
C19849 vdd.n10500 vss 0.0951f
C19850 vdd.t1005 vss 0.0013f
C19851 vdd.t1262 vss 0.00134f
C19852 vdd.n10501 vss 0.00324f
C19853 vdd.n10502 vss 0.0112f
C19854 vdd.n10503 vss 0.0128f
C19855 vdd.n10504 vss 0.00413f
C19856 vdd.n10505 vss 0.00413f
C19857 vdd.n10506 vss 0.0471f
C19858 vdd.n10507 vss 0.00251f
C19859 vdd.t775 vss 0.0471f
C19860 vdd.n10508 vss 0.00324f
C19861 vdd.n10510 vss 0.00679f
C19862 vdd.n10511 vss 0.00413f
C19863 vdd.n10512 vss 0.00324f
C19864 vdd.n10513 vss 0.00413f
C19865 vdd.n10514 vss 0.0471f
C19866 vdd.n10515 vss 0.00324f
C19867 vdd.n10517 vss 0.00925f
C19868 vdd.t1102 vss 0.0471f
C19869 vdd.n10518 vss 0.00425f
C19870 vdd.n10519 vss 0.0424f
C19871 vdd.n10520 vss 0.0132f
C19872 vdd.n10521 vss 0.00324f
C19873 vdd.n10522 vss 0.0128f
C19874 vdd.n10523 vss 0.02f
C19875 vdd.n10524 vss 0.00425f
C19876 vdd.n10525 vss 0.00413f
C19877 vdd.n10526 vss 0.00251f
C19878 vdd.t261 vss 0.0471f
C19879 vdd.n10527 vss 0.00251f
C19880 vdd.n10528 vss 0.00517f
C19881 vdd.n10529 vss 0.00679f
C19882 vdd.n10530 vss 0.00517f
C19883 vdd.n10531 vss 0.00679f
C19884 vdd.n10532 vss 0.02f
C19885 vdd.n10533 vss 0.00425f
C19886 vdd.n10534 vss 0.0424f
C19887 vdd.n10535 vss 0.0132f
C19888 vdd.n10536 vss 0.00925f
C19889 vdd.n10537 vss 0.00425f
C19890 vdd.n10538 vss 0.00413f
C19891 vdd.n10539 vss 0.00324f
C19892 vdd.n10540 vss 0.0471f
C19893 vdd.t262 vss 0.0471f
C19894 vdd.n10541 vss 0.00251f
C19895 vdd.n10542 vss 0.0112f
C19896 vdd.n10543 vss 0.0128f
C19897 vdd.t263 vss 0.00134f
C19898 vdd.t776 vss 0.0013f
C19899 vdd.n10544 vss 0.0332f
C19900 vdd.n10545 vss 0.0393f
C19901 vdd.n10546 vss 0.119f
C19902 vdd.n10547 vss 0.00324f
C19903 vdd.n10548 vss 0.0112f
C19904 vdd.n10549 vss 0.0128f
C19905 vdd.n10550 vss 0.00413f
C19906 vdd.n10551 vss 0.00413f
C19907 vdd.n10552 vss 0.0471f
C19908 vdd.n10553 vss 0.00251f
C19909 vdd.t1004 vss 0.0471f
C19910 vdd.n10554 vss 0.00324f
C19911 vdd.n10556 vss 0.00679f
C19912 vdd.n10557 vss 0.00413f
C19913 vdd.n10558 vss 0.00324f
C19914 vdd.n10559 vss 0.00413f
C19915 vdd.n10560 vss 0.0471f
C19916 vdd.n10561 vss 0.00324f
C19917 vdd.n10563 vss 0.00925f
C19918 vdd.t1366 vss 0.0471f
C19919 vdd.n10564 vss 0.00425f
C19920 vdd.n10565 vss 0.0424f
C19921 vdd.n10566 vss 0.0132f
C19922 vdd.n10567 vss 0.00324f
C19923 vdd.n10568 vss 0.0128f
C19924 vdd.n10569 vss 0.02f
C19925 vdd.n10570 vss 0.00425f
C19926 vdd.n10571 vss 0.00413f
C19927 vdd.n10572 vss 0.00251f
C19928 vdd.t1260 vss 0.0471f
C19929 vdd.n10573 vss 0.00251f
C19930 vdd.n10574 vss 0.00517f
C19931 vdd.n10575 vss 0.00679f
C19932 vdd.n10576 vss 0.00517f
C19933 vdd.n10577 vss 0.00679f
C19934 vdd.n10578 vss 0.02f
C19935 vdd.n10579 vss 0.00425f
C19936 vdd.n10580 vss 0.0424f
C19937 vdd.n10581 vss 0.0132f
C19938 vdd.n10582 vss 0.00925f
C19939 vdd.n10583 vss 0.00425f
C19940 vdd.n10584 vss 0.00413f
C19941 vdd.n10585 vss 0.00324f
C19942 vdd.n10586 vss 0.0471f
C19943 vdd.t1261 vss 0.0471f
C19944 vdd.n10587 vss 0.00251f
C19945 vdd.n10588 vss 0.0112f
C19946 vdd.n10589 vss 0.0128f
C19947 vdd.n10590 vss 0.118f
C19948 vdd.n10591 vss 0.0393f
C19949 vdd.n10592 vss 0.0332f
C19950 vdd.n10593 vss 0.0596f
C19951 vdd.n10594 vss 0.00324f
C19952 vdd.n10595 vss 0.0112f
C19953 vdd.n10596 vss 0.0128f
C19954 vdd.n10597 vss 0.00413f
C19955 vdd.n10598 vss 0.00413f
C19956 vdd.n10599 vss 0.0471f
C19957 vdd.n10600 vss 0.00251f
C19958 vdd.t1491 vss 0.0471f
C19959 vdd.n10601 vss 0.00324f
C19960 vdd.n10603 vss 0.00679f
C19961 vdd.n10604 vss 0.00413f
C19962 vdd.n10605 vss 0.00324f
C19963 vdd.n10606 vss 0.00413f
C19964 vdd.n10607 vss 0.0471f
C19965 vdd.n10608 vss 0.00324f
C19966 vdd.n10610 vss 0.00925f
C19967 vdd.t1019 vss 0.0471f
C19968 vdd.n10611 vss 0.00425f
C19969 vdd.n10612 vss 0.0424f
C19970 vdd.n10613 vss 0.0132f
C19971 vdd.n10614 vss 0.00324f
C19972 vdd.n10615 vss 0.0128f
C19973 vdd.n10616 vss 0.02f
C19974 vdd.n10617 vss 0.00425f
C19975 vdd.n10618 vss 0.00413f
C19976 vdd.n10619 vss 0.00251f
C19977 vdd.t1077 vss 0.0471f
C19978 vdd.n10620 vss 0.00251f
C19979 vdd.n10621 vss 0.00517f
C19980 vdd.n10622 vss 0.00679f
C19981 vdd.n10623 vss 0.00517f
C19982 vdd.n10624 vss 0.00679f
C19983 vdd.n10625 vss 0.02f
C19984 vdd.n10626 vss 0.00425f
C19985 vdd.n10627 vss 0.0424f
C19986 vdd.n10628 vss 0.0132f
C19987 vdd.n10629 vss 0.00925f
C19988 vdd.n10630 vss 0.00425f
C19989 vdd.n10631 vss 0.00413f
C19990 vdd.n10632 vss 0.00324f
C19991 vdd.n10633 vss 0.0471f
C19992 vdd.t1075 vss 0.0471f
C19993 vdd.n10634 vss 0.00251f
C19994 vdd.n10635 vss 0.0112f
C19995 vdd.n10636 vss 0.0128f
C19996 vdd.t1076 vss 0.00134f
C19997 vdd.t1492 vss 0.0013f
C19998 vdd.n10637 vss 0.0332f
C19999 vdd.n10638 vss 0.0393f
C20000 vdd.n10639 vss 0.0418f
C20001 vdd.n10640 vss 0.118f
C20002 vdd.n10641 vss 0.121f
C20003 vdd.t818 vss 0.0013f
C20004 vdd.t609 vss 0.00134f
C20005 vdd.n10642 vss 0.00324f
C20006 vdd.n10643 vss 0.0112f
C20007 vdd.n10644 vss 0.0128f
C20008 vdd.n10645 vss 0.00413f
C20009 vdd.n10646 vss 0.00413f
C20010 vdd.n10647 vss 0.0471f
C20011 vdd.n10648 vss 0.00251f
C20012 vdd.t817 vss 0.0471f
C20013 vdd.n10649 vss 0.00324f
C20014 vdd.n10651 vss 0.00679f
C20015 vdd.n10652 vss 0.00413f
C20016 vdd.n10653 vss 0.00324f
C20017 vdd.n10654 vss 0.00413f
C20018 vdd.n10655 vss 0.0471f
C20019 vdd.n10656 vss 0.00324f
C20020 vdd.n10658 vss 0.00925f
C20021 vdd.t253 vss 0.0471f
C20022 vdd.n10659 vss 0.00425f
C20023 vdd.n10660 vss 0.0424f
C20024 vdd.n10661 vss 0.0132f
C20025 vdd.n10662 vss 0.00324f
C20026 vdd.n10663 vss 0.0128f
C20027 vdd.n10664 vss 0.02f
C20028 vdd.n10665 vss 0.00425f
C20029 vdd.n10666 vss 0.00413f
C20030 vdd.n10667 vss 0.00251f
C20031 vdd.t610 vss 0.0471f
C20032 vdd.n10668 vss 0.00251f
C20033 vdd.n10669 vss 0.00517f
C20034 vdd.n10670 vss 0.00679f
C20035 vdd.n10671 vss 0.00517f
C20036 vdd.n10672 vss 0.00679f
C20037 vdd.n10673 vss 0.02f
C20038 vdd.n10674 vss 0.00425f
C20039 vdd.n10675 vss 0.0424f
C20040 vdd.n10676 vss 0.0132f
C20041 vdd.n10677 vss 0.00925f
C20042 vdd.n10678 vss 0.00425f
C20043 vdd.n10679 vss 0.00413f
C20044 vdd.n10680 vss 0.00324f
C20045 vdd.n10681 vss 0.0471f
C20046 vdd.t608 vss 0.0471f
C20047 vdd.n10682 vss 0.00251f
C20048 vdd.n10683 vss 0.0112f
C20049 vdd.n10684 vss 0.0707f
C20050 vdd.n10685 vss 0.0393f
C20051 vdd.n10686 vss 0.0332f
C20052 vdd.n10687 vss 0.0596f
C20053 vdd.n10688 vss 0.00324f
C20054 vdd.n10689 vss 0.0112f
C20055 vdd.n10690 vss 0.0128f
C20056 vdd.n10691 vss 0.00413f
C20057 vdd.n10692 vss 0.00413f
C20058 vdd.n10693 vss 0.0471f
C20059 vdd.n10694 vss 0.00251f
C20060 vdd.t1352 vss 0.0471f
C20061 vdd.n10695 vss 0.00324f
C20062 vdd.n10697 vss 0.00679f
C20063 vdd.n10698 vss 0.00413f
C20064 vdd.n10699 vss 0.00324f
C20065 vdd.n10700 vss 0.00413f
C20066 vdd.n10701 vss 0.0471f
C20067 vdd.n10702 vss 0.00324f
C20068 vdd.n10704 vss 0.00925f
C20069 vdd.t292 vss 0.0471f
C20070 vdd.n10705 vss 0.00425f
C20071 vdd.n10706 vss 0.0424f
C20072 vdd.n10707 vss 0.0132f
C20073 vdd.n10708 vss 0.00324f
C20074 vdd.n10709 vss 0.0128f
C20075 vdd.n10710 vss 0.02f
C20076 vdd.n10711 vss 0.00425f
C20077 vdd.n10712 vss 0.00413f
C20078 vdd.n10713 vss 0.00251f
C20079 vdd.t146 vss 0.0471f
C20080 vdd.n10714 vss 0.00251f
C20081 vdd.n10715 vss 0.00517f
C20082 vdd.n10716 vss 0.00679f
C20083 vdd.n10717 vss 0.00517f
C20084 vdd.n10718 vss 0.00679f
C20085 vdd.n10719 vss 0.02f
C20086 vdd.n10720 vss 0.00425f
C20087 vdd.n10721 vss 0.0424f
C20088 vdd.n10722 vss 0.0132f
C20089 vdd.n10723 vss 0.00925f
C20090 vdd.n10724 vss 0.00425f
C20091 vdd.n10725 vss 0.00413f
C20092 vdd.n10726 vss 0.00324f
C20093 vdd.n10727 vss 0.0471f
C20094 vdd.t147 vss 0.0471f
C20095 vdd.n10728 vss 0.00251f
C20096 vdd.n10729 vss 0.0112f
C20097 vdd.n10730 vss 0.0128f
C20098 vdd.t148 vss 0.00134f
C20099 vdd.t1353 vss 0.0013f
C20100 vdd.n10731 vss 0.0332f
C20101 vdd.n10732 vss 0.0393f
C20102 vdd.n10733 vss 0.0418f
C20103 vdd.n10734 vss 0.0912f
C20104 vdd.n10735 vss 0.0824f
C20105 vdd.n10736 vss 0.059f
C20106 vdd.t903 vss 0.0013f
C20107 vdd.t1236 vss 0.00134f
C20108 vdd.n10737 vss 0.00324f
C20109 vdd.n10738 vss 0.0112f
C20110 vdd.n10739 vss 0.0128f
C20111 vdd.n10740 vss 0.00413f
C20112 vdd.n10741 vss 0.00413f
C20113 vdd.n10742 vss 0.0471f
C20114 vdd.n10743 vss 0.00251f
C20115 vdd.t629 vss 0.0471f
C20116 vdd.n10744 vss 0.00324f
C20117 vdd.n10746 vss 0.00679f
C20118 vdd.n10747 vss 0.00413f
C20119 vdd.n10748 vss 0.00324f
C20120 vdd.n10749 vss 0.00413f
C20121 vdd.n10750 vss 0.0471f
C20122 vdd.n10751 vss 0.00324f
C20123 vdd.n10753 vss 0.00925f
C20124 vdd.t1247 vss 0.0471f
C20125 vdd.n10754 vss 0.00425f
C20126 vdd.n10755 vss 0.0424f
C20127 vdd.n10756 vss 0.0132f
C20128 vdd.n10757 vss 0.00324f
C20129 vdd.n10758 vss 0.0128f
C20130 vdd.n10759 vss 0.02f
C20131 vdd.n10760 vss 0.00425f
C20132 vdd.n10761 vss 0.00413f
C20133 vdd.n10762 vss 0.00251f
C20134 vdd.t1244 vss 0.0471f
C20135 vdd.n10763 vss 0.00251f
C20136 vdd.n10764 vss 0.00517f
C20137 vdd.n10765 vss 0.00679f
C20138 vdd.n10766 vss 0.00517f
C20139 vdd.n10767 vss 0.00679f
C20140 vdd.n10768 vss 0.02f
C20141 vdd.n10769 vss 0.00425f
C20142 vdd.n10770 vss 0.0424f
C20143 vdd.n10771 vss 0.0132f
C20144 vdd.n10772 vss 0.00925f
C20145 vdd.n10773 vss 0.00425f
C20146 vdd.n10774 vss 0.00413f
C20147 vdd.n10775 vss 0.00324f
C20148 vdd.n10776 vss 0.0471f
C20149 vdd.t1245 vss 0.0471f
C20150 vdd.n10777 vss 0.00251f
C20151 vdd.n10778 vss 0.0112f
C20152 vdd.n10779 vss 0.0128f
C20153 vdd.t1246 vss 0.00134f
C20154 vdd.t630 vss 0.0013f
C20155 vdd.n10780 vss 0.0332f
C20156 vdd.n10781 vss 0.0393f
C20157 vdd.n10782 vss 0.119f
C20158 vdd.n10783 vss 0.00324f
C20159 vdd.n10784 vss 0.0112f
C20160 vdd.n10785 vss 0.0128f
C20161 vdd.n10786 vss 0.00413f
C20162 vdd.n10787 vss 0.00413f
C20163 vdd.n10788 vss 0.0471f
C20164 vdd.n10789 vss 0.00251f
C20165 vdd.t902 vss 0.0471f
C20166 vdd.n10790 vss 0.00324f
C20167 vdd.n10792 vss 0.00679f
C20168 vdd.n10793 vss 0.00413f
C20169 vdd.n10794 vss 0.00324f
C20170 vdd.n10795 vss 0.00413f
C20171 vdd.n10796 vss 0.0471f
C20172 vdd.n10797 vss 0.00324f
C20173 vdd.n10799 vss 0.00925f
C20174 vdd.t742 vss 0.0471f
C20175 vdd.n10800 vss 0.00425f
C20176 vdd.n10801 vss 0.0424f
C20177 vdd.n10802 vss 0.0132f
C20178 vdd.n10803 vss 0.00324f
C20179 vdd.n10804 vss 0.0128f
C20180 vdd.n10805 vss 0.02f
C20181 vdd.n10806 vss 0.00425f
C20182 vdd.n10807 vss 0.00413f
C20183 vdd.n10808 vss 0.00251f
C20184 vdd.t1234 vss 0.0471f
C20185 vdd.n10809 vss 0.00251f
C20186 vdd.n10810 vss 0.00517f
C20187 vdd.n10811 vss 0.00679f
C20188 vdd.n10812 vss 0.00517f
C20189 vdd.n10813 vss 0.00679f
C20190 vdd.n10814 vss 0.02f
C20191 vdd.n10815 vss 0.00425f
C20192 vdd.n10816 vss 0.0424f
C20193 vdd.n10817 vss 0.0132f
C20194 vdd.n10818 vss 0.00925f
C20195 vdd.n10819 vss 0.00425f
C20196 vdd.n10820 vss 0.00413f
C20197 vdd.n10821 vss 0.00324f
C20198 vdd.n10822 vss 0.0471f
C20199 vdd.t1235 vss 0.0471f
C20200 vdd.n10823 vss 0.00251f
C20201 vdd.n10824 vss 0.0112f
C20202 vdd.n10825 vss 0.0128f
C20203 vdd.n10826 vss 0.118f
C20204 vdd.n10827 vss 0.0393f
C20205 vdd.n10828 vss 0.0332f
C20206 vdd.n10829 vss 0.0596f
C20207 vdd.n10830 vss 0.00324f
C20208 vdd.n10831 vss 0.0112f
C20209 vdd.n10832 vss 0.0128f
C20210 vdd.n10833 vss 0.00413f
C20211 vdd.n10834 vss 0.00413f
C20212 vdd.n10835 vss 0.0471f
C20213 vdd.n10836 vss 0.00251f
C20214 vdd.t480 vss 0.0471f
C20215 vdd.n10837 vss 0.00324f
C20216 vdd.n10839 vss 0.00679f
C20217 vdd.n10840 vss 0.00413f
C20218 vdd.n10841 vss 0.00324f
C20219 vdd.n10842 vss 0.00413f
C20220 vdd.n10843 vss 0.0471f
C20221 vdd.n10844 vss 0.00324f
C20222 vdd.n10846 vss 0.00925f
C20223 vdd.t417 vss 0.0471f
C20224 vdd.n10847 vss 0.00425f
C20225 vdd.n10848 vss 0.0424f
C20226 vdd.n10849 vss 0.0132f
C20227 vdd.n10850 vss 0.00324f
C20228 vdd.n10851 vss 0.0128f
C20229 vdd.n10852 vss 0.02f
C20230 vdd.n10853 vss 0.00425f
C20231 vdd.n10854 vss 0.00413f
C20232 vdd.n10855 vss 0.00251f
C20233 vdd.t1162 vss 0.0471f
C20234 vdd.n10856 vss 0.00251f
C20235 vdd.n10857 vss 0.00517f
C20236 vdd.n10858 vss 0.00679f
C20237 vdd.n10859 vss 0.00517f
C20238 vdd.n10860 vss 0.00679f
C20239 vdd.n10861 vss 0.02f
C20240 vdd.n10862 vss 0.00425f
C20241 vdd.n10863 vss 0.0424f
C20242 vdd.n10864 vss 0.0132f
C20243 vdd.n10865 vss 0.00925f
C20244 vdd.n10866 vss 0.00425f
C20245 vdd.n10867 vss 0.00413f
C20246 vdd.n10868 vss 0.00324f
C20247 vdd.n10869 vss 0.0471f
C20248 vdd.t1160 vss 0.0471f
C20249 vdd.n10870 vss 0.00251f
C20250 vdd.n10871 vss 0.0112f
C20251 vdd.n10872 vss 0.0128f
C20252 vdd.t1161 vss 0.00134f
C20253 vdd.t481 vss 0.0013f
C20254 vdd.n10873 vss 0.0332f
C20255 vdd.n10874 vss 0.0393f
C20256 vdd.n10875 vss 0.0418f
C20257 vdd.n10876 vss 0.118f
C20258 vdd.n10877 vss 0.121f
C20259 vdd.t937 vss 0.0013f
C20260 vdd.t950 vss 0.00134f
C20261 vdd.n10878 vss 0.00324f
C20262 vdd.n10879 vss 0.0112f
C20263 vdd.n10880 vss 0.0128f
C20264 vdd.n10881 vss 0.00413f
C20265 vdd.n10882 vss 0.00413f
C20266 vdd.n10883 vss 0.0471f
C20267 vdd.n10884 vss 0.00251f
C20268 vdd.t936 vss 0.0471f
C20269 vdd.n10885 vss 0.00324f
C20270 vdd.n10887 vss 0.00679f
C20271 vdd.n10888 vss 0.00413f
C20272 vdd.n10889 vss 0.00324f
C20273 vdd.n10890 vss 0.00413f
C20274 vdd.n10891 vss 0.0471f
C20275 vdd.n10892 vss 0.00324f
C20276 vdd.n10894 vss 0.00925f
C20277 vdd.t285 vss 0.0471f
C20278 vdd.n10895 vss 0.00425f
C20279 vdd.n10896 vss 0.0424f
C20280 vdd.n10897 vss 0.0132f
C20281 vdd.n10898 vss 0.00324f
C20282 vdd.n10899 vss 0.0128f
C20283 vdd.n10900 vss 0.02f
C20284 vdd.n10901 vss 0.00425f
C20285 vdd.n10902 vss 0.00413f
C20286 vdd.n10903 vss 0.00251f
C20287 vdd.t948 vss 0.0471f
C20288 vdd.n10904 vss 0.00251f
C20289 vdd.n10905 vss 0.00517f
C20290 vdd.n10906 vss 0.00679f
C20291 vdd.n10907 vss 0.00517f
C20292 vdd.n10908 vss 0.00679f
C20293 vdd.n10909 vss 0.02f
C20294 vdd.n10910 vss 0.00425f
C20295 vdd.n10911 vss 0.0424f
C20296 vdd.n10912 vss 0.0132f
C20297 vdd.n10913 vss 0.00925f
C20298 vdd.n10914 vss 0.00425f
C20299 vdd.n10915 vss 0.00413f
C20300 vdd.n10916 vss 0.00324f
C20301 vdd.n10917 vss 0.0471f
C20302 vdd.t949 vss 0.0471f
C20303 vdd.n10918 vss 0.00251f
C20304 vdd.n10919 vss 0.0112f
C20305 vdd.n10920 vss 0.0707f
C20306 vdd.n10921 vss 0.0393f
C20307 vdd.n10922 vss 0.0332f
C20308 vdd.n10923 vss 0.0596f
C20309 vdd.n10924 vss 0.00324f
C20310 vdd.n10925 vss 0.0112f
C20311 vdd.n10926 vss 0.0128f
C20312 vdd.n10927 vss 0.00413f
C20313 vdd.n10928 vss 0.00413f
C20314 vdd.n10929 vss 0.0471f
C20315 vdd.n10930 vss 0.00251f
C20316 vdd.t5 vss 0.0471f
C20317 vdd.n10931 vss 0.00324f
C20318 vdd.n10933 vss 0.00679f
C20319 vdd.n10934 vss 0.00413f
C20320 vdd.n10935 vss 0.00324f
C20321 vdd.n10936 vss 0.00413f
C20322 vdd.n10937 vss 0.0471f
C20323 vdd.n10938 vss 0.00324f
C20324 vdd.n10940 vss 0.00925f
C20325 vdd.t690 vss 0.0471f
C20326 vdd.n10941 vss 0.00425f
C20327 vdd.n10942 vss 0.0424f
C20328 vdd.n10943 vss 0.0132f
C20329 vdd.n10944 vss 0.00324f
C20330 vdd.n10945 vss 0.0128f
C20331 vdd.n10946 vss 0.02f
C20332 vdd.n10947 vss 0.00425f
C20333 vdd.n10948 vss 0.00413f
C20334 vdd.n10949 vss 0.00251f
C20335 vdd.t1196 vss 0.0471f
C20336 vdd.n10950 vss 0.00251f
C20337 vdd.n10951 vss 0.00517f
C20338 vdd.n10952 vss 0.00679f
C20339 vdd.n10953 vss 0.00517f
C20340 vdd.n10954 vss 0.00679f
C20341 vdd.n10955 vss 0.02f
C20342 vdd.n10956 vss 0.00425f
C20343 vdd.n10957 vss 0.0424f
C20344 vdd.n10958 vss 0.0132f
C20345 vdd.n10959 vss 0.00925f
C20346 vdd.n10960 vss 0.00425f
C20347 vdd.n10961 vss 0.00413f
C20348 vdd.n10962 vss 0.00324f
C20349 vdd.n10963 vss 0.0471f
C20350 vdd.t1197 vss 0.0471f
C20351 vdd.n10964 vss 0.00251f
C20352 vdd.n10965 vss 0.0112f
C20353 vdd.n10966 vss 0.0128f
C20354 vdd.t1198 vss 0.00134f
C20355 vdd.t6 vss 0.0013f
C20356 vdd.n10967 vss 0.0332f
C20357 vdd.n10968 vss 0.0393f
C20358 vdd.n10969 vss 0.0418f
C20359 vdd.n10970 vss 0.121f
C20360 vdd.n10971 vss 0.32f
C20361 vdd.n10972 vss 0.202f
C20362 vdd.t822 vss 0.0013f
C20363 vdd.t287 vss 0.00134f
C20364 vdd.n10973 vss 0.00324f
C20365 vdd.n10974 vss 0.0112f
C20366 vdd.n10975 vss 0.0128f
C20367 vdd.n10976 vss 0.00413f
C20368 vdd.t288 vss 0.0471f
C20369 vdd.n10977 vss 0.00324f
C20370 vdd.n10979 vss 0.00925f
C20371 vdd.n10980 vss 0.00413f
C20372 vdd.n10981 vss 0.00679f
C20373 vdd.n10982 vss 0.00413f
C20374 vdd.n10983 vss 0.0471f
C20375 vdd.n10984 vss 0.00324f
C20376 vdd.n10985 vss 0.0471f
C20377 vdd.n10986 vss 0.00324f
C20378 vdd.n10987 vss 0.0424f
C20379 vdd.t821 vss 0.0471f
C20380 vdd.n10989 vss 0.00425f
C20381 vdd.n10990 vss 0.00925f
C20382 vdd.n10991 vss 0.0132f
C20383 vdd.n10992 vss 0.00324f
C20384 vdd.n10993 vss 0.0128f
C20385 vdd.n10994 vss 0.02f
C20386 vdd.n10995 vss 0.00425f
C20387 vdd.n10996 vss 0.00413f
C20388 vdd.n10997 vss 0.00251f
C20389 vdd.t286 vss 0.0471f
C20390 vdd.n10998 vss 0.00251f
C20391 vdd.n10999 vss 0.00517f
C20392 vdd.n11000 vss 0.00679f
C20393 vdd.n11001 vss 0.00324f
C20394 vdd.n11002 vss 0.00679f
C20395 vdd.n11003 vss 0.00517f
C20396 vdd.n11004 vss 0.00251f
C20397 vdd.n11005 vss 0.00413f
C20398 vdd.n11006 vss 0.0471f
C20399 vdd.t498 vss 0.0471f
C20400 vdd.n11007 vss 0.00425f
C20401 vdd.n11008 vss 0.0424f
C20402 vdd.n11009 vss 0.0132f
C20403 vdd.n11010 vss 0.02f
C20404 vdd.n11011 vss 0.00425f
C20405 vdd.n11012 vss 0.00413f
C20406 vdd.n11013 vss 0.00251f
C20407 vdd.n11014 vss 0.0112f
C20408 vdd.n11015 vss 0.0128f
C20409 vdd.t646 vss 0.00134f
C20410 vdd.t59 vss 0.0013f
C20411 vdd.n11016 vss 0.032f
C20412 vdd.n11017 vss 0.0393f
C20413 vdd.n11018 vss 0.00324f
C20414 vdd.n11019 vss 0.0112f
C20415 vdd.n11020 vss 0.0128f
C20416 vdd.n11021 vss 0.00413f
C20417 vdd.t647 vss 0.0471f
C20418 vdd.n11022 vss 0.00324f
C20419 vdd.n11024 vss 0.00925f
C20420 vdd.n11025 vss 0.00413f
C20421 vdd.n11026 vss 0.00679f
C20422 vdd.n11027 vss 0.00413f
C20423 vdd.n11028 vss 0.0471f
C20424 vdd.n11029 vss 0.00324f
C20425 vdd.n11030 vss 0.0471f
C20426 vdd.n11031 vss 0.00324f
C20427 vdd.n11032 vss 0.0424f
C20428 vdd.t58 vss 0.0471f
C20429 vdd.n11034 vss 0.00425f
C20430 vdd.n11035 vss 0.00925f
C20431 vdd.n11036 vss 0.0132f
C20432 vdd.n11037 vss 0.00324f
C20433 vdd.n11038 vss 0.0128f
C20434 vdd.n11039 vss 0.02f
C20435 vdd.n11040 vss 0.00425f
C20436 vdd.n11041 vss 0.00413f
C20437 vdd.n11042 vss 0.00251f
C20438 vdd.t645 vss 0.0471f
C20439 vdd.n11043 vss 0.00251f
C20440 vdd.n11044 vss 0.00517f
C20441 vdd.n11045 vss 0.00679f
C20442 vdd.n11046 vss 0.00324f
C20443 vdd.n11047 vss 0.00679f
C20444 vdd.n11048 vss 0.00517f
C20445 vdd.n11049 vss 0.00251f
C20446 vdd.n11050 vss 0.00413f
C20447 vdd.n11051 vss 0.0471f
C20448 vdd.t1251 vss 0.0471f
C20449 vdd.n11052 vss 0.00425f
C20450 vdd.n11053 vss 0.0424f
C20451 vdd.n11054 vss 0.0132f
C20452 vdd.n11055 vss 0.02f
C20453 vdd.n11056 vss 0.00425f
C20454 vdd.n11057 vss 0.00413f
C20455 vdd.n11058 vss 0.00251f
C20456 vdd.n11059 vss 0.0112f
C20457 vdd.n11060 vss 0.0128f
C20458 vdd.n11061 vss 0.119f
C20459 vdd.n11062 vss 0.118f
C20460 vdd.n11063 vss 0.0393f
C20461 vdd.n11064 vss 0.032f
C20462 vdd.n11065 vss 0.0608f
C20463 vdd.t734 vss 0.00134f
C20464 vdd.t1500 vss 0.0013f
C20465 vdd.n11066 vss 0.032f
C20466 vdd.n11067 vss 0.0393f
C20467 vdd.n11068 vss 0.00324f
C20468 vdd.n11069 vss 0.0112f
C20469 vdd.n11070 vss 0.0128f
C20470 vdd.n11071 vss 0.00413f
C20471 vdd.t735 vss 0.0471f
C20472 vdd.n11072 vss 0.00324f
C20473 vdd.n11074 vss 0.00925f
C20474 vdd.n11075 vss 0.00413f
C20475 vdd.n11076 vss 0.00679f
C20476 vdd.n11077 vss 0.00413f
C20477 vdd.n11078 vss 0.0471f
C20478 vdd.n11079 vss 0.00324f
C20479 vdd.n11080 vss 0.0471f
C20480 vdd.n11081 vss 0.00324f
C20481 vdd.n11082 vss 0.0424f
C20482 vdd.t1499 vss 0.0471f
C20483 vdd.n11084 vss 0.00425f
C20484 vdd.n11085 vss 0.00925f
C20485 vdd.n11086 vss 0.0132f
C20486 vdd.n11087 vss 0.00324f
C20487 vdd.n11088 vss 0.0128f
C20488 vdd.n11089 vss 0.02f
C20489 vdd.n11090 vss 0.00425f
C20490 vdd.n11091 vss 0.00413f
C20491 vdd.n11092 vss 0.00251f
C20492 vdd.t733 vss 0.0471f
C20493 vdd.n11093 vss 0.00251f
C20494 vdd.n11094 vss 0.00517f
C20495 vdd.n11095 vss 0.00679f
C20496 vdd.n11096 vss 0.00324f
C20497 vdd.n11097 vss 0.00679f
C20498 vdd.n11098 vss 0.00517f
C20499 vdd.n11099 vss 0.00251f
C20500 vdd.n11100 vss 0.00413f
C20501 vdd.n11101 vss 0.0471f
C20502 vdd.t538 vss 0.0471f
C20503 vdd.n11102 vss 0.00425f
C20504 vdd.n11103 vss 0.0424f
C20505 vdd.n11104 vss 0.0132f
C20506 vdd.n11105 vss 0.02f
C20507 vdd.n11106 vss 0.00425f
C20508 vdd.n11107 vss 0.00413f
C20509 vdd.n11108 vss 0.00251f
C20510 vdd.n11109 vss 0.0112f
C20511 vdd.n11110 vss 0.0128f
C20512 vdd.n11111 vss 0.0418f
C20513 vdd.n11112 vss 0.118f
C20514 vdd.n11113 vss 0.121f
C20515 vdd.t997 vss 0.0013f
C20516 vdd.t295 vss 0.00134f
C20517 vdd.n11114 vss 0.00324f
C20518 vdd.n11115 vss 0.0112f
C20519 vdd.n11116 vss 0.0128f
C20520 vdd.n11117 vss 0.00413f
C20521 vdd.t293 vss 0.0471f
C20522 vdd.n11118 vss 0.00324f
C20523 vdd.n11120 vss 0.00925f
C20524 vdd.n11121 vss 0.00413f
C20525 vdd.n11122 vss 0.00679f
C20526 vdd.n11123 vss 0.00413f
C20527 vdd.n11124 vss 0.0471f
C20528 vdd.n11125 vss 0.00324f
C20529 vdd.n11126 vss 0.0471f
C20530 vdd.n11127 vss 0.00324f
C20531 vdd.n11128 vss 0.0424f
C20532 vdd.t996 vss 0.0471f
C20533 vdd.n11130 vss 0.00425f
C20534 vdd.n11131 vss 0.00925f
C20535 vdd.n11132 vss 0.0132f
C20536 vdd.n11133 vss 0.00324f
C20537 vdd.n11134 vss 0.0128f
C20538 vdd.n11135 vss 0.02f
C20539 vdd.n11136 vss 0.00425f
C20540 vdd.n11137 vss 0.00413f
C20541 vdd.n11138 vss 0.00251f
C20542 vdd.t294 vss 0.0471f
C20543 vdd.n11139 vss 0.00251f
C20544 vdd.n11140 vss 0.00517f
C20545 vdd.n11141 vss 0.00679f
C20546 vdd.n11142 vss 0.00324f
C20547 vdd.n11143 vss 0.00679f
C20548 vdd.n11144 vss 0.00517f
C20549 vdd.n11145 vss 0.00251f
C20550 vdd.n11146 vss 0.00413f
C20551 vdd.n11147 vss 0.0471f
C20552 vdd.t539 vss 0.0471f
C20553 vdd.n11148 vss 0.00425f
C20554 vdd.n11149 vss 0.0424f
C20555 vdd.n11150 vss 0.0132f
C20556 vdd.n11151 vss 0.02f
C20557 vdd.n11152 vss 0.00425f
C20558 vdd.n11153 vss 0.00413f
C20559 vdd.n11154 vss 0.00251f
C20560 vdd.n11155 vss 0.0112f
C20561 vdd.n11156 vss 0.0707f
C20562 vdd.n11157 vss 0.0393f
C20563 vdd.n11158 vss 0.032f
C20564 vdd.n11159 vss 0.0608f
C20565 vdd.t351 vss 0.00134f
C20566 vdd.t1295 vss 0.0013f
C20567 vdd.n11160 vss 0.032f
C20568 vdd.n11161 vss 0.0393f
C20569 vdd.n11162 vss 0.00324f
C20570 vdd.n11163 vss 0.0112f
C20571 vdd.n11164 vss 0.0128f
C20572 vdd.n11165 vss 0.00413f
C20573 vdd.t352 vss 0.0471f
C20574 vdd.n11166 vss 0.00324f
C20575 vdd.n11168 vss 0.00925f
C20576 vdd.n11169 vss 0.00413f
C20577 vdd.n11170 vss 0.00679f
C20578 vdd.n11171 vss 0.00413f
C20579 vdd.n11172 vss 0.0471f
C20580 vdd.n11173 vss 0.00324f
C20581 vdd.n11174 vss 0.0471f
C20582 vdd.n11175 vss 0.00324f
C20583 vdd.n11176 vss 0.0424f
C20584 vdd.t1294 vss 0.0471f
C20585 vdd.n11178 vss 0.00425f
C20586 vdd.n11179 vss 0.00925f
C20587 vdd.n11180 vss 0.0132f
C20588 vdd.n11181 vss 0.00324f
C20589 vdd.n11182 vss 0.0128f
C20590 vdd.n11183 vss 0.02f
C20591 vdd.n11184 vss 0.00425f
C20592 vdd.n11185 vss 0.00413f
C20593 vdd.n11186 vss 0.00251f
C20594 vdd.t350 vss 0.0471f
C20595 vdd.n11187 vss 0.00251f
C20596 vdd.n11188 vss 0.00517f
C20597 vdd.n11189 vss 0.00679f
C20598 vdd.n11190 vss 0.00324f
C20599 vdd.n11191 vss 0.00679f
C20600 vdd.n11192 vss 0.00517f
C20601 vdd.n11193 vss 0.00251f
C20602 vdd.n11194 vss 0.00413f
C20603 vdd.n11195 vss 0.0471f
C20604 vdd.t216 vss 0.0471f
C20605 vdd.n11196 vss 0.00425f
C20606 vdd.n11197 vss 0.0424f
C20607 vdd.n11198 vss 0.0132f
C20608 vdd.n11199 vss 0.02f
C20609 vdd.n11200 vss 0.00425f
C20610 vdd.n11201 vss 0.00413f
C20611 vdd.n11202 vss 0.00251f
C20612 vdd.n11203 vss 0.0112f
C20613 vdd.n11204 vss 0.0128f
C20614 vdd.n11205 vss 0.0418f
C20615 vdd.n11206 vss 0.0912f
C20616 vdd.n11207 vss 0.0824f
C20617 vdd.n11208 vss 0.0567f
C20618 vdd.t966 vss 0.0013f
C20619 vdd.t515 vss 0.00134f
C20620 vdd.n11209 vss 0.00324f
C20621 vdd.n11210 vss 0.0112f
C20622 vdd.n11211 vss 0.0128f
C20623 vdd.n11212 vss 0.00413f
C20624 vdd.t513 vss 0.0471f
C20625 vdd.n11213 vss 0.00324f
C20626 vdd.n11215 vss 0.00925f
C20627 vdd.n11216 vss 0.00413f
C20628 vdd.n11217 vss 0.00679f
C20629 vdd.n11218 vss 0.00413f
C20630 vdd.n11219 vss 0.0471f
C20631 vdd.n11220 vss 0.00324f
C20632 vdd.n11221 vss 0.0471f
C20633 vdd.n11222 vss 0.00324f
C20634 vdd.n11223 vss 0.0424f
C20635 vdd.t965 vss 0.0471f
C20636 vdd.n11225 vss 0.00425f
C20637 vdd.n11226 vss 0.00925f
C20638 vdd.n11227 vss 0.0132f
C20639 vdd.n11228 vss 0.00324f
C20640 vdd.n11229 vss 0.0128f
C20641 vdd.n11230 vss 0.02f
C20642 vdd.n11231 vss 0.00425f
C20643 vdd.n11232 vss 0.00413f
C20644 vdd.n11233 vss 0.00251f
C20645 vdd.t514 vss 0.0471f
C20646 vdd.n11234 vss 0.00251f
C20647 vdd.n11235 vss 0.00517f
C20648 vdd.n11236 vss 0.00679f
C20649 vdd.n11237 vss 0.00324f
C20650 vdd.n11238 vss 0.00679f
C20651 vdd.n11239 vss 0.00517f
C20652 vdd.n11240 vss 0.00251f
C20653 vdd.n11241 vss 0.00413f
C20654 vdd.n11242 vss 0.0471f
C20655 vdd.t115 vss 0.0471f
C20656 vdd.n11243 vss 0.00425f
C20657 vdd.n11244 vss 0.0424f
C20658 vdd.n11245 vss 0.0132f
C20659 vdd.n11246 vss 0.02f
C20660 vdd.n11247 vss 0.00425f
C20661 vdd.n11248 vss 0.00413f
C20662 vdd.n11249 vss 0.00251f
C20663 vdd.n11250 vss 0.0112f
C20664 vdd.n11251 vss 0.0128f
C20665 vdd.t890 vss 0.00134f
C20666 vdd.t797 vss 0.0013f
C20667 vdd.n11252 vss 0.032f
C20668 vdd.n11253 vss 0.0393f
C20669 vdd.n11254 vss 0.00324f
C20670 vdd.n11255 vss 0.0112f
C20671 vdd.n11256 vss 0.0128f
C20672 vdd.n11257 vss 0.00413f
C20673 vdd.t891 vss 0.0471f
C20674 vdd.n11258 vss 0.00324f
C20675 vdd.n11260 vss 0.00925f
C20676 vdd.n11261 vss 0.00413f
C20677 vdd.n11262 vss 0.00679f
C20678 vdd.n11263 vss 0.00413f
C20679 vdd.n11264 vss 0.0471f
C20680 vdd.n11265 vss 0.00324f
C20681 vdd.n11266 vss 0.0471f
C20682 vdd.n11267 vss 0.00324f
C20683 vdd.n11268 vss 0.0424f
C20684 vdd.t796 vss 0.0471f
C20685 vdd.n11270 vss 0.00425f
C20686 vdd.n11271 vss 0.00925f
C20687 vdd.n11272 vss 0.0132f
C20688 vdd.n11273 vss 0.00324f
C20689 vdd.n11274 vss 0.0128f
C20690 vdd.n11275 vss 0.02f
C20691 vdd.n11276 vss 0.00425f
C20692 vdd.n11277 vss 0.00413f
C20693 vdd.n11278 vss 0.00251f
C20694 vdd.t889 vss 0.0471f
C20695 vdd.n11279 vss 0.00251f
C20696 vdd.n11280 vss 0.00517f
C20697 vdd.n11281 vss 0.00679f
C20698 vdd.n11282 vss 0.00324f
C20699 vdd.n11283 vss 0.00679f
C20700 vdd.n11284 vss 0.00517f
C20701 vdd.n11285 vss 0.00251f
C20702 vdd.n11286 vss 0.00413f
C20703 vdd.n11287 vss 0.0471f
C20704 vdd.t531 vss 0.0471f
C20705 vdd.n11288 vss 0.00425f
C20706 vdd.n11289 vss 0.0424f
C20707 vdd.n11290 vss 0.0132f
C20708 vdd.n11291 vss 0.02f
C20709 vdd.n11292 vss 0.00425f
C20710 vdd.n11293 vss 0.00413f
C20711 vdd.n11294 vss 0.00251f
C20712 vdd.n11295 vss 0.0112f
C20713 vdd.n11296 vss 0.0128f
C20714 vdd.n11297 vss 0.0316f
C20715 vdd.t406 vss 0.00134f
C20716 vdd.t1378 vss 0.0013f
C20717 vdd.n11298 vss 0.032f
C20718 vdd.n11299 vss 0.0393f
C20719 vdd.n11300 vss 0.00324f
C20720 vdd.n11301 vss 0.0112f
C20721 vdd.n11302 vss 0.0128f
C20722 vdd.n11303 vss 0.00413f
C20723 vdd.t407 vss 0.0471f
C20724 vdd.n11304 vss 0.00324f
C20725 vdd.n11306 vss 0.00925f
C20726 vdd.n11307 vss 0.00413f
C20727 vdd.n11308 vss 0.00679f
C20728 vdd.n11309 vss 0.00413f
C20729 vdd.n11310 vss 0.0471f
C20730 vdd.n11311 vss 0.00324f
C20731 vdd.n11312 vss 0.0471f
C20732 vdd.n11313 vss 0.00324f
C20733 vdd.n11314 vss 0.0424f
C20734 vdd.t1377 vss 0.0471f
C20735 vdd.n11316 vss 0.00425f
C20736 vdd.n11317 vss 0.00925f
C20737 vdd.n11318 vss 0.0132f
C20738 vdd.n11319 vss 0.00324f
C20739 vdd.n11320 vss 0.0128f
C20740 vdd.n11321 vss 0.02f
C20741 vdd.n11322 vss 0.00425f
C20742 vdd.n11323 vss 0.00413f
C20743 vdd.n11324 vss 0.00251f
C20744 vdd.t405 vss 0.0471f
C20745 vdd.n11325 vss 0.00251f
C20746 vdd.n11326 vss 0.00517f
C20747 vdd.n11327 vss 0.00679f
C20748 vdd.n11328 vss 0.00324f
C20749 vdd.n11329 vss 0.00679f
C20750 vdd.n11330 vss 0.00517f
C20751 vdd.n11331 vss 0.00251f
C20752 vdd.n11332 vss 0.00413f
C20753 vdd.n11333 vss 0.0471f
C20754 vdd.t1037 vss 0.0471f
C20755 vdd.n11334 vss 0.00425f
C20756 vdd.n11335 vss 0.0424f
C20757 vdd.n11336 vss 0.0132f
C20758 vdd.n11337 vss 0.02f
C20759 vdd.n11338 vss 0.00425f
C20760 vdd.n11339 vss 0.00413f
C20761 vdd.n11340 vss 0.00251f
C20762 vdd.n11341 vss 0.0112f
C20763 vdd.n11342 vss 0.0128f
C20764 vdd.n11343 vss 0.158f
C20765 vdd.n11344 vss 0.256f
C20766 vdd.n11345 vss 0.0953f
C20767 vdd.n11346 vss 0.0393f
C20768 vdd.n11347 vss 0.032f
C20769 vdd.n11348 vss 0.0608f
C20770 vdd.t1146 vss 0.00134f
C20771 vdd.t200 vss 0.0013f
C20772 vdd.n11349 vss 0.032f
C20773 vdd.n11350 vss 0.0393f
C20774 vdd.n11351 vss 0.00324f
C20775 vdd.n11352 vss 0.0112f
C20776 vdd.n11353 vss 0.0128f
C20777 vdd.n11354 vss 0.00413f
C20778 vdd.t1144 vss 0.0471f
C20779 vdd.n11355 vss 0.00324f
C20780 vdd.n11357 vss 0.00925f
C20781 vdd.n11358 vss 0.00413f
C20782 vdd.n11359 vss 0.00679f
C20783 vdd.n11360 vss 0.00413f
C20784 vdd.n11361 vss 0.0471f
C20785 vdd.n11362 vss 0.00324f
C20786 vdd.n11363 vss 0.0471f
C20787 vdd.n11364 vss 0.00324f
C20788 vdd.n11365 vss 0.0424f
C20789 vdd.t199 vss 0.0471f
C20790 vdd.n11367 vss 0.00425f
C20791 vdd.n11368 vss 0.00925f
C20792 vdd.n11369 vss 0.0132f
C20793 vdd.n11370 vss 0.00324f
C20794 vdd.n11371 vss 0.0128f
C20795 vdd.n11372 vss 0.02f
C20796 vdd.n11373 vss 0.00425f
C20797 vdd.n11374 vss 0.00413f
C20798 vdd.n11375 vss 0.00251f
C20799 vdd.t1145 vss 0.0471f
C20800 vdd.n11376 vss 0.00251f
C20801 vdd.n11377 vss 0.00517f
C20802 vdd.n11378 vss 0.00679f
C20803 vdd.n11379 vss 0.00324f
C20804 vdd.n11380 vss 0.00679f
C20805 vdd.n11381 vss 0.00517f
C20806 vdd.n11382 vss 0.00251f
C20807 vdd.n11383 vss 0.00413f
C20808 vdd.n11384 vss 0.0471f
C20809 vdd.t1147 vss 0.0471f
C20810 vdd.n11385 vss 0.00425f
C20811 vdd.n11386 vss 0.0424f
C20812 vdd.n11387 vss 0.0132f
C20813 vdd.n11388 vss 0.02f
C20814 vdd.n11389 vss 0.00425f
C20815 vdd.n11390 vss 0.00413f
C20816 vdd.n11391 vss 0.00251f
C20817 vdd.n11392 vss 0.0112f
C20818 vdd.n11393 vss 0.0128f
C20819 vdd.n11394 vss 0.0418f
C20820 vdd.n11395 vss 0.118f
C20821 vdd.n11396 vss 0.121f
C20822 vdd.t851 vss 0.0013f
C20823 vdd.t283 vss 0.00134f
C20824 vdd.n11397 vss 0.00324f
C20825 vdd.n11398 vss 0.0112f
C20826 vdd.n11399 vss 0.0128f
C20827 vdd.n11400 vss 0.00413f
C20828 vdd.t281 vss 0.0471f
C20829 vdd.n11401 vss 0.00324f
C20830 vdd.n11403 vss 0.00925f
C20831 vdd.n11404 vss 0.00413f
C20832 vdd.n11405 vss 0.00679f
C20833 vdd.n11406 vss 0.00413f
C20834 vdd.n11407 vss 0.0471f
C20835 vdd.n11408 vss 0.00324f
C20836 vdd.n11409 vss 0.0471f
C20837 vdd.n11410 vss 0.00324f
C20838 vdd.n11411 vss 0.0424f
C20839 vdd.t850 vss 0.0471f
C20840 vdd.n11413 vss 0.00425f
C20841 vdd.n11414 vss 0.00925f
C20842 vdd.n11415 vss 0.0132f
C20843 vdd.n11416 vss 0.00324f
C20844 vdd.n11417 vss 0.0128f
C20845 vdd.n11418 vss 0.02f
C20846 vdd.n11419 vss 0.00425f
C20847 vdd.n11420 vss 0.00413f
C20848 vdd.n11421 vss 0.00251f
C20849 vdd.t282 vss 0.0471f
C20850 vdd.n11422 vss 0.00251f
C20851 vdd.n11423 vss 0.00517f
C20852 vdd.n11424 vss 0.00679f
C20853 vdd.n11425 vss 0.00324f
C20854 vdd.n11426 vss 0.00679f
C20855 vdd.n11427 vss 0.00517f
C20856 vdd.n11428 vss 0.00251f
C20857 vdd.n11429 vss 0.00413f
C20858 vdd.n11430 vss 0.0471f
C20859 vdd.t958 vss 0.0471f
C20860 vdd.n11431 vss 0.00425f
C20861 vdd.n11432 vss 0.0424f
C20862 vdd.n11433 vss 0.0132f
C20863 vdd.n11434 vss 0.02f
C20864 vdd.n11435 vss 0.00425f
C20865 vdd.n11436 vss 0.00413f
C20866 vdd.n11437 vss 0.00251f
C20867 vdd.n11438 vss 0.0112f
C20868 vdd.n11439 vss 0.0707f
C20869 vdd.n11440 vss 0.0393f
C20870 vdd.n11441 vss 0.032f
C20871 vdd.n11442 vss 0.0608f
C20872 vdd.t1522 vss 0.00134f
C20873 vdd.t1341 vss 0.0013f
C20874 vdd.n11443 vss 0.032f
C20875 vdd.n11444 vss 0.0393f
C20876 vdd.n11445 vss 0.00324f
C20877 vdd.n11446 vss 0.0112f
C20878 vdd.n11447 vss 0.0128f
C20879 vdd.n11448 vss 0.00413f
C20880 vdd.t1523 vss 0.0471f
C20881 vdd.n11449 vss 0.00324f
C20882 vdd.n11451 vss 0.00925f
C20883 vdd.n11452 vss 0.00413f
C20884 vdd.n11453 vss 0.00679f
C20885 vdd.n11454 vss 0.00413f
C20886 vdd.n11455 vss 0.0471f
C20887 vdd.n11456 vss 0.00324f
C20888 vdd.n11457 vss 0.0471f
C20889 vdd.n11458 vss 0.00324f
C20890 vdd.n11459 vss 0.0424f
C20891 vdd.t1340 vss 0.0471f
C20892 vdd.n11461 vss 0.00425f
C20893 vdd.n11462 vss 0.00925f
C20894 vdd.n11463 vss 0.0132f
C20895 vdd.n11464 vss 0.00324f
C20896 vdd.n11465 vss 0.0128f
C20897 vdd.n11466 vss 0.02f
C20898 vdd.n11467 vss 0.00425f
C20899 vdd.n11468 vss 0.00413f
C20900 vdd.n11469 vss 0.00251f
C20901 vdd.t1521 vss 0.0471f
C20902 vdd.n11470 vss 0.00251f
C20903 vdd.n11471 vss 0.00517f
C20904 vdd.n11472 vss 0.00679f
C20905 vdd.n11473 vss 0.00324f
C20906 vdd.n11474 vss 0.00679f
C20907 vdd.n11475 vss 0.00517f
C20908 vdd.n11476 vss 0.00251f
C20909 vdd.n11477 vss 0.00413f
C20910 vdd.n11478 vss 0.0471f
C20911 vdd.t1242 vss 0.0471f
C20912 vdd.n11479 vss 0.00425f
C20913 vdd.n11480 vss 0.0424f
C20914 vdd.n11481 vss 0.0132f
C20915 vdd.n11482 vss 0.02f
C20916 vdd.n11483 vss 0.00425f
C20917 vdd.n11484 vss 0.00413f
C20918 vdd.n11485 vss 0.00251f
C20919 vdd.n11486 vss 0.0112f
C20920 vdd.n11487 vss 0.0128f
C20921 vdd.n11488 vss 0.0418f
C20922 vdd.n11489 vss 0.118f
C20923 vdd.n11490 vss 0.0935f
C20924 vdd.t812 vss 0.0013f
C20925 vdd.t271 vss 0.00134f
C20926 vdd.n11491 vss 0.00324f
C20927 vdd.n11492 vss 0.0112f
C20928 vdd.n11493 vss 0.0128f
C20929 vdd.n11494 vss 0.00413f
C20930 vdd.t272 vss 0.0471f
C20931 vdd.n11495 vss 0.00324f
C20932 vdd.n11497 vss 0.00925f
C20933 vdd.n11498 vss 0.00413f
C20934 vdd.n11499 vss 0.00679f
C20935 vdd.n11500 vss 0.00413f
C20936 vdd.n11501 vss 0.0471f
C20937 vdd.n11502 vss 0.00324f
C20938 vdd.n11503 vss 0.0471f
C20939 vdd.n11504 vss 0.00324f
C20940 vdd.n11505 vss 0.0424f
C20941 vdd.t811 vss 0.0471f
C20942 vdd.n11507 vss 0.00425f
C20943 vdd.n11508 vss 0.00925f
C20944 vdd.n11509 vss 0.0132f
C20945 vdd.n11510 vss 0.00324f
C20946 vdd.n11511 vss 0.0128f
C20947 vdd.n11512 vss 0.02f
C20948 vdd.n11513 vss 0.00425f
C20949 vdd.n11514 vss 0.00413f
C20950 vdd.n11515 vss 0.00251f
C20951 vdd.t270 vss 0.0471f
C20952 vdd.n11516 vss 0.00251f
C20953 vdd.n11517 vss 0.00517f
C20954 vdd.n11518 vss 0.00679f
C20955 vdd.n11519 vss 0.00324f
C20956 vdd.n11520 vss 0.00679f
C20957 vdd.n11521 vss 0.00517f
C20958 vdd.n11522 vss 0.00251f
C20959 vdd.n11523 vss 0.00413f
C20960 vdd.n11524 vss 0.0471f
C20961 vdd.t273 vss 0.0471f
C20962 vdd.n11525 vss 0.00425f
C20963 vdd.n11526 vss 0.0424f
C20964 vdd.n11527 vss 0.0132f
C20965 vdd.n11528 vss 0.02f
C20966 vdd.n11529 vss 0.00425f
C20967 vdd.n11530 vss 0.00413f
C20968 vdd.n11531 vss 0.00251f
C20969 vdd.n11532 vss 0.0112f
C20970 vdd.n11533 vss 0.0128f
C20971 vdd.t1440 vss 0.00134f
C20972 vdd.t795 vss 0.0013f
C20973 vdd.n11534 vss 0.032f
C20974 vdd.n11535 vss 0.0393f
C20975 vdd.n11536 vss 0.00324f
C20976 vdd.n11537 vss 0.0112f
C20977 vdd.n11538 vss 0.0128f
C20978 vdd.n11539 vss 0.00413f
C20979 vdd.t1441 vss 0.0471f
C20980 vdd.n11540 vss 0.00324f
C20981 vdd.n11542 vss 0.00925f
C20982 vdd.n11543 vss 0.00413f
C20983 vdd.n11544 vss 0.00679f
C20984 vdd.n11545 vss 0.00413f
C20985 vdd.n11546 vss 0.0471f
C20986 vdd.n11547 vss 0.00324f
C20987 vdd.n11548 vss 0.0471f
C20988 vdd.n11549 vss 0.00324f
C20989 vdd.n11550 vss 0.0424f
C20990 vdd.t794 vss 0.0471f
C20991 vdd.n11552 vss 0.00425f
C20992 vdd.n11553 vss 0.00925f
C20993 vdd.n11554 vss 0.0132f
C20994 vdd.n11555 vss 0.00324f
C20995 vdd.n11556 vss 0.0128f
C20996 vdd.n11557 vss 0.02f
C20997 vdd.n11558 vss 0.00425f
C20998 vdd.n11559 vss 0.00413f
C20999 vdd.n11560 vss 0.00251f
C21000 vdd.t1439 vss 0.0471f
C21001 vdd.n11561 vss 0.00251f
C21002 vdd.n11562 vss 0.00517f
C21003 vdd.n11563 vss 0.00679f
C21004 vdd.n11564 vss 0.00324f
C21005 vdd.n11565 vss 0.00679f
C21006 vdd.n11566 vss 0.00517f
C21007 vdd.n11567 vss 0.00251f
C21008 vdd.n11568 vss 0.00413f
C21009 vdd.n11569 vss 0.0471f
C21010 vdd.t307 vss 0.0471f
C21011 vdd.n11570 vss 0.00425f
C21012 vdd.n11571 vss 0.0424f
C21013 vdd.n11572 vss 0.0132f
C21014 vdd.n11573 vss 0.02f
C21015 vdd.n11574 vss 0.00425f
C21016 vdd.n11575 vss 0.00413f
C21017 vdd.n11576 vss 0.00251f
C21018 vdd.n11577 vss 0.0112f
C21019 vdd.n11578 vss 0.0128f
C21020 vdd.n11579 vss 0.119f
C21021 vdd.n11580 vss 0.118f
C21022 vdd.n11581 vss 0.0393f
C21023 vdd.n11582 vss 0.032f
C21024 vdd.n11583 vss 0.0608f
C21025 vdd.t1391 vss 0.00134f
C21026 vdd.t1287 vss 0.0013f
C21027 vdd.n11584 vss 0.032f
C21028 vdd.n11585 vss 0.0393f
C21029 vdd.n11586 vss 0.00324f
C21030 vdd.n11587 vss 0.0112f
C21031 vdd.n11588 vss 0.0128f
C21032 vdd.n11589 vss 0.00413f
C21033 vdd.t1392 vss 0.0471f
C21034 vdd.n11590 vss 0.00324f
C21035 vdd.n11592 vss 0.00925f
C21036 vdd.n11593 vss 0.00413f
C21037 vdd.n11594 vss 0.00679f
C21038 vdd.n11595 vss 0.00413f
C21039 vdd.n11596 vss 0.0471f
C21040 vdd.n11597 vss 0.00324f
C21041 vdd.n11598 vss 0.0471f
C21042 vdd.n11599 vss 0.00324f
C21043 vdd.n11600 vss 0.0424f
C21044 vdd.t1286 vss 0.0471f
C21045 vdd.n11602 vss 0.00425f
C21046 vdd.n11603 vss 0.00925f
C21047 vdd.n11604 vss 0.0132f
C21048 vdd.n11605 vss 0.00324f
C21049 vdd.n11606 vss 0.0128f
C21050 vdd.n11607 vss 0.02f
C21051 vdd.n11608 vss 0.00425f
C21052 vdd.n11609 vss 0.00413f
C21053 vdd.n11610 vss 0.00251f
C21054 vdd.t1390 vss 0.0471f
C21055 vdd.n11611 vss 0.00251f
C21056 vdd.n11612 vss 0.00517f
C21057 vdd.n11613 vss 0.00679f
C21058 vdd.n11614 vss 0.00324f
C21059 vdd.n11615 vss 0.00679f
C21060 vdd.n11616 vss 0.00517f
C21061 vdd.n11617 vss 0.00251f
C21062 vdd.n11618 vss 0.00413f
C21063 vdd.n11619 vss 0.0471f
C21064 vdd.t535 vss 0.0471f
C21065 vdd.n11620 vss 0.00425f
C21066 vdd.n11621 vss 0.0424f
C21067 vdd.n11622 vss 0.0132f
C21068 vdd.n11623 vss 0.02f
C21069 vdd.n11624 vss 0.00425f
C21070 vdd.n11625 vss 0.00413f
C21071 vdd.n11626 vss 0.00251f
C21072 vdd.n11627 vss 0.0112f
C21073 vdd.n11628 vss 0.0128f
C21074 vdd.n11629 vss 0.0418f
C21075 vdd.n11630 vss 0.118f
C21076 vdd.n11631 vss 0.121f
C21077 vdd.t995 vss 0.0013f
C21078 vdd.t1249 vss 0.00134f
C21079 vdd.n11632 vss 0.00324f
C21080 vdd.n11633 vss 0.0112f
C21081 vdd.n11634 vss 0.0128f
C21082 vdd.n11635 vss 0.00413f
C21083 vdd.t1250 vss 0.0471f
C21084 vdd.n11636 vss 0.00324f
C21085 vdd.n11638 vss 0.00925f
C21086 vdd.n11639 vss 0.00413f
C21087 vdd.n11640 vss 0.00679f
C21088 vdd.n11641 vss 0.00413f
C21089 vdd.n11642 vss 0.0471f
C21090 vdd.n11643 vss 0.00324f
C21091 vdd.n11644 vss 0.0471f
C21092 vdd.n11645 vss 0.00324f
C21093 vdd.n11646 vss 0.0424f
C21094 vdd.t994 vss 0.0471f
C21095 vdd.n11648 vss 0.00425f
C21096 vdd.n11649 vss 0.00925f
C21097 vdd.n11650 vss 0.0132f
C21098 vdd.n11651 vss 0.00324f
C21099 vdd.n11652 vss 0.0128f
C21100 vdd.n11653 vss 0.02f
C21101 vdd.n11654 vss 0.00425f
C21102 vdd.n11655 vss 0.00413f
C21103 vdd.n11656 vss 0.00251f
C21104 vdd.t1248 vss 0.0471f
C21105 vdd.n11657 vss 0.00251f
C21106 vdd.n11658 vss 0.00517f
C21107 vdd.n11659 vss 0.00679f
C21108 vdd.n11660 vss 0.00324f
C21109 vdd.n11661 vss 0.00679f
C21110 vdd.n11662 vss 0.00517f
C21111 vdd.n11663 vss 0.00251f
C21112 vdd.n11664 vss 0.00413f
C21113 vdd.n11665 vss 0.0471f
C21114 vdd.t641 vss 0.0471f
C21115 vdd.n11666 vss 0.00425f
C21116 vdd.n11667 vss 0.0424f
C21117 vdd.n11668 vss 0.0132f
C21118 vdd.n11669 vss 0.02f
C21119 vdd.n11670 vss 0.00425f
C21120 vdd.n11671 vss 0.00413f
C21121 vdd.n11672 vss 0.00251f
C21122 vdd.n11673 vss 0.0112f
C21123 vdd.n11674 vss 0.0707f
C21124 vdd.n11675 vss 0.0393f
C21125 vdd.n11676 vss 0.032f
C21126 vdd.n11677 vss 0.0608f
C21127 vdd.t529 vss 0.00134f
C21128 vdd.t1339 vss 0.0013f
C21129 vdd.n11678 vss 0.032f
C21130 vdd.n11679 vss 0.0393f
C21131 vdd.n11680 vss 0.00324f
C21132 vdd.n11681 vss 0.0112f
C21133 vdd.n11682 vss 0.0128f
C21134 vdd.n11683 vss 0.00413f
C21135 vdd.t530 vss 0.0471f
C21136 vdd.n11684 vss 0.00324f
C21137 vdd.n11686 vss 0.00925f
C21138 vdd.n11687 vss 0.00413f
C21139 vdd.n11688 vss 0.00679f
C21140 vdd.n11689 vss 0.00413f
C21141 vdd.n11690 vss 0.0471f
C21142 vdd.n11691 vss 0.00324f
C21143 vdd.n11692 vss 0.0471f
C21144 vdd.n11693 vss 0.00324f
C21145 vdd.n11694 vss 0.0424f
C21146 vdd.t1338 vss 0.0471f
C21147 vdd.n11696 vss 0.00425f
C21148 vdd.n11697 vss 0.00925f
C21149 vdd.n11698 vss 0.0132f
C21150 vdd.n11699 vss 0.00324f
C21151 vdd.n11700 vss 0.0128f
C21152 vdd.n11701 vss 0.02f
C21153 vdd.n11702 vss 0.00425f
C21154 vdd.n11703 vss 0.00413f
C21155 vdd.n11704 vss 0.00251f
C21156 vdd.t528 vss 0.0471f
C21157 vdd.n11705 vss 0.00251f
C21158 vdd.n11706 vss 0.00517f
C21159 vdd.n11707 vss 0.00679f
C21160 vdd.n11708 vss 0.00324f
C21161 vdd.n11709 vss 0.00679f
C21162 vdd.n11710 vss 0.00517f
C21163 vdd.n11711 vss 0.00251f
C21164 vdd.n11712 vss 0.00413f
C21165 vdd.n11713 vss 0.0471f
C21166 vdd.t1120 vss 0.0471f
C21167 vdd.n11714 vss 0.00425f
C21168 vdd.n11715 vss 0.0424f
C21169 vdd.n11716 vss 0.0132f
C21170 vdd.n11717 vss 0.02f
C21171 vdd.n11718 vss 0.00425f
C21172 vdd.n11719 vss 0.00413f
C21173 vdd.n11720 vss 0.00251f
C21174 vdd.n11721 vss 0.0112f
C21175 vdd.n11722 vss 0.0128f
C21176 vdd.n11723 vss 0.0418f
C21177 vdd.n11724 vss 0.0912f
C21178 vdd.n11725 vss 0.0824f
C21179 vdd.n11726 vss 0.0567f
C21180 vdd.t1015 vss 0.0013f
C21181 vdd.t358 vss 0.00134f
C21182 vdd.n11727 vss 0.00324f
C21183 vdd.n11728 vss 0.0112f
C21184 vdd.n11729 vss 0.0128f
C21185 vdd.n11730 vss 0.00413f
C21186 vdd.t359 vss 0.0471f
C21187 vdd.n11731 vss 0.00324f
C21188 vdd.n11733 vss 0.00925f
C21189 vdd.n11734 vss 0.00413f
C21190 vdd.n11735 vss 0.00679f
C21191 vdd.n11736 vss 0.00413f
C21192 vdd.n11737 vss 0.0471f
C21193 vdd.n11738 vss 0.00324f
C21194 vdd.n11739 vss 0.0471f
C21195 vdd.n11740 vss 0.00324f
C21196 vdd.n11741 vss 0.0424f
C21197 vdd.t1014 vss 0.0471f
C21198 vdd.n11743 vss 0.00425f
C21199 vdd.n11744 vss 0.00925f
C21200 vdd.n11745 vss 0.0132f
C21201 vdd.n11746 vss 0.00324f
C21202 vdd.n11747 vss 0.0128f
C21203 vdd.n11748 vss 0.02f
C21204 vdd.n11749 vss 0.00425f
C21205 vdd.n11750 vss 0.00413f
C21206 vdd.n11751 vss 0.00251f
C21207 vdd.t357 vss 0.0471f
C21208 vdd.n11752 vss 0.00251f
C21209 vdd.n11753 vss 0.00517f
C21210 vdd.n11754 vss 0.00679f
C21211 vdd.n11755 vss 0.00324f
C21212 vdd.n11756 vss 0.00679f
C21213 vdd.n11757 vss 0.00517f
C21214 vdd.n11758 vss 0.00251f
C21215 vdd.n11759 vss 0.00413f
C21216 vdd.n11760 vss 0.0471f
C21217 vdd.t49 vss 0.0471f
C21218 vdd.n11761 vss 0.00425f
C21219 vdd.n11762 vss 0.0424f
C21220 vdd.n11763 vss 0.0132f
C21221 vdd.n11764 vss 0.02f
C21222 vdd.n11765 vss 0.00425f
C21223 vdd.n11766 vss 0.00413f
C21224 vdd.n11767 vss 0.00251f
C21225 vdd.n11768 vss 0.0112f
C21226 vdd.n11769 vss 0.0128f
C21227 vdd.t105 vss 0.00134f
C21228 vdd.t793 vss 0.0013f
C21229 vdd.n11770 vss 0.032f
C21230 vdd.n11771 vss 0.0393f
C21231 vdd.n11772 vss 0.00324f
C21232 vdd.n11773 vss 0.0112f
C21233 vdd.n11774 vss 0.0128f
C21234 vdd.n11775 vss 0.00413f
C21235 vdd.t106 vss 0.0471f
C21236 vdd.n11776 vss 0.00324f
C21237 vdd.n11778 vss 0.00925f
C21238 vdd.n11779 vss 0.00413f
C21239 vdd.n11780 vss 0.00679f
C21240 vdd.n11781 vss 0.00413f
C21241 vdd.n11782 vss 0.0471f
C21242 vdd.n11783 vss 0.00324f
C21243 vdd.n11784 vss 0.0471f
C21244 vdd.n11785 vss 0.00324f
C21245 vdd.n11786 vss 0.0424f
C21246 vdd.t792 vss 0.0471f
C21247 vdd.n11788 vss 0.00425f
C21248 vdd.n11789 vss 0.00925f
C21249 vdd.n11790 vss 0.0132f
C21250 vdd.n11791 vss 0.00324f
C21251 vdd.n11792 vss 0.0128f
C21252 vdd.n11793 vss 0.02f
C21253 vdd.n11794 vss 0.00425f
C21254 vdd.n11795 vss 0.00413f
C21255 vdd.n11796 vss 0.00251f
C21256 vdd.t104 vss 0.0471f
C21257 vdd.n11797 vss 0.00251f
C21258 vdd.n11798 vss 0.00517f
C21259 vdd.n11799 vss 0.00679f
C21260 vdd.n11800 vss 0.00324f
C21261 vdd.n11801 vss 0.00679f
C21262 vdd.n11802 vss 0.00517f
C21263 vdd.n11803 vss 0.00251f
C21264 vdd.n11804 vss 0.00413f
C21265 vdd.n11805 vss 0.0471f
C21266 vdd.t1396 vss 0.0471f
C21267 vdd.n11806 vss 0.00425f
C21268 vdd.n11807 vss 0.0424f
C21269 vdd.n11808 vss 0.0132f
C21270 vdd.n11809 vss 0.02f
C21271 vdd.n11810 vss 0.00425f
C21272 vdd.n11811 vss 0.00413f
C21273 vdd.n11812 vss 0.00251f
C21274 vdd.n11813 vss 0.0112f
C21275 vdd.n11814 vss 0.0128f
C21276 vdd.n11815 vss 0.119f
C21277 vdd.n11816 vss 0.118f
C21278 vdd.n11817 vss 0.0393f
C21279 vdd.n11818 vss 0.032f
C21280 vdd.n11819 vss 0.0608f
C21281 vdd.t317 vss 0.00134f
C21282 vdd.t1321 vss 0.0013f
C21283 vdd.n11820 vss 0.032f
C21284 vdd.n11821 vss 0.0393f
C21285 vdd.n11822 vss 0.00324f
C21286 vdd.n11823 vss 0.0112f
C21287 vdd.n11824 vss 0.0128f
C21288 vdd.n11825 vss 0.00413f
C21289 vdd.t315 vss 0.0471f
C21290 vdd.n11826 vss 0.00324f
C21291 vdd.n11828 vss 0.00925f
C21292 vdd.n11829 vss 0.00413f
C21293 vdd.n11830 vss 0.00679f
C21294 vdd.n11831 vss 0.00413f
C21295 vdd.n11832 vss 0.0471f
C21296 vdd.n11833 vss 0.00324f
C21297 vdd.n11834 vss 0.0471f
C21298 vdd.n11835 vss 0.00324f
C21299 vdd.n11836 vss 0.0424f
C21300 vdd.t1320 vss 0.0471f
C21301 vdd.n11838 vss 0.00425f
C21302 vdd.n11839 vss 0.00925f
C21303 vdd.n11840 vss 0.0132f
C21304 vdd.n11841 vss 0.00324f
C21305 vdd.n11842 vss 0.0128f
C21306 vdd.n11843 vss 0.02f
C21307 vdd.n11844 vss 0.00425f
C21308 vdd.n11845 vss 0.00413f
C21309 vdd.n11846 vss 0.00251f
C21310 vdd.t316 vss 0.0471f
C21311 vdd.n11847 vss 0.00251f
C21312 vdd.n11848 vss 0.00517f
C21313 vdd.n11849 vss 0.00679f
C21314 vdd.n11850 vss 0.00324f
C21315 vdd.n11851 vss 0.00679f
C21316 vdd.n11852 vss 0.00517f
C21317 vdd.n11853 vss 0.00251f
C21318 vdd.n11854 vss 0.00413f
C21319 vdd.n11855 vss 0.0471f
C21320 vdd.t1271 vss 0.0471f
C21321 vdd.n11856 vss 0.00425f
C21322 vdd.n11857 vss 0.0424f
C21323 vdd.n11858 vss 0.0132f
C21324 vdd.n11859 vss 0.02f
C21325 vdd.n11860 vss 0.00425f
C21326 vdd.n11861 vss 0.00413f
C21327 vdd.n11862 vss 0.00251f
C21328 vdd.n11863 vss 0.0112f
C21329 vdd.n11864 vss 0.0128f
C21330 vdd.n11865 vss 0.0418f
C21331 vdd.n11866 vss 0.118f
C21332 vdd.n11867 vss 0.121f
C21333 vdd.t814 vss 0.0013f
C21334 vdd.t753 vss 0.00134f
C21335 vdd.n11868 vss 0.00324f
C21336 vdd.n11869 vss 0.0112f
C21337 vdd.n11870 vss 0.0128f
C21338 vdd.n11871 vss 0.00413f
C21339 vdd.t754 vss 0.0471f
C21340 vdd.n11872 vss 0.00324f
C21341 vdd.n11874 vss 0.00925f
C21342 vdd.n11875 vss 0.00413f
C21343 vdd.n11876 vss 0.00679f
C21344 vdd.n11877 vss 0.00413f
C21345 vdd.n11878 vss 0.0471f
C21346 vdd.n11879 vss 0.00324f
C21347 vdd.n11880 vss 0.0471f
C21348 vdd.n11881 vss 0.00324f
C21349 vdd.n11882 vss 0.0424f
C21350 vdd.t813 vss 0.0471f
C21351 vdd.n11884 vss 0.00425f
C21352 vdd.n11885 vss 0.00925f
C21353 vdd.n11886 vss 0.0132f
C21354 vdd.n11887 vss 0.00324f
C21355 vdd.n11888 vss 0.0128f
C21356 vdd.n11889 vss 0.02f
C21357 vdd.n11890 vss 0.00425f
C21358 vdd.n11891 vss 0.00413f
C21359 vdd.n11892 vss 0.00251f
C21360 vdd.t752 vss 0.0471f
C21361 vdd.n11893 vss 0.00251f
C21362 vdd.n11894 vss 0.00517f
C21363 vdd.n11895 vss 0.00679f
C21364 vdd.n11896 vss 0.00324f
C21365 vdd.n11897 vss 0.00679f
C21366 vdd.n11898 vss 0.00517f
C21367 vdd.n11899 vss 0.00251f
C21368 vdd.n11900 vss 0.00413f
C21369 vdd.n11901 vss 0.0471f
C21370 vdd.t619 vss 0.0471f
C21371 vdd.n11902 vss 0.00425f
C21372 vdd.n11903 vss 0.0424f
C21373 vdd.n11904 vss 0.0132f
C21374 vdd.n11905 vss 0.02f
C21375 vdd.n11906 vss 0.00425f
C21376 vdd.n11907 vss 0.00413f
C21377 vdd.n11908 vss 0.00251f
C21378 vdd.n11909 vss 0.0112f
C21379 vdd.n11910 vss 0.0707f
C21380 vdd.n11911 vss 0.0393f
C21381 vdd.n11912 vss 0.032f
C21382 vdd.n11913 vss 0.0608f
C21383 vdd.t341 vss 0.00134f
C21384 vdd.t1293 vss 0.0013f
C21385 vdd.n11914 vss 0.032f
C21386 vdd.n11915 vss 0.0393f
C21387 vdd.n11916 vss 0.00324f
C21388 vdd.n11917 vss 0.0112f
C21389 vdd.n11918 vss 0.0128f
C21390 vdd.n11919 vss 0.00413f
C21391 vdd.t342 vss 0.0471f
C21392 vdd.n11920 vss 0.00324f
C21393 vdd.n11922 vss 0.00925f
C21394 vdd.n11923 vss 0.00413f
C21395 vdd.n11924 vss 0.00679f
C21396 vdd.n11925 vss 0.00413f
C21397 vdd.n11926 vss 0.0471f
C21398 vdd.n11927 vss 0.00324f
C21399 vdd.n11928 vss 0.0471f
C21400 vdd.n11929 vss 0.00324f
C21401 vdd.n11930 vss 0.0424f
C21402 vdd.t1292 vss 0.0471f
C21403 vdd.n11932 vss 0.00425f
C21404 vdd.n11933 vss 0.00925f
C21405 vdd.n11934 vss 0.0132f
C21406 vdd.n11935 vss 0.00324f
C21407 vdd.n11936 vss 0.0128f
C21408 vdd.n11937 vss 0.02f
C21409 vdd.n11938 vss 0.00425f
C21410 vdd.n11939 vss 0.00413f
C21411 vdd.n11940 vss 0.00251f
C21412 vdd.t340 vss 0.0471f
C21413 vdd.n11941 vss 0.00251f
C21414 vdd.n11942 vss 0.00517f
C21415 vdd.n11943 vss 0.00679f
C21416 vdd.n11944 vss 0.00324f
C21417 vdd.n11945 vss 0.00679f
C21418 vdd.n11946 vss 0.00517f
C21419 vdd.n11947 vss 0.00251f
C21420 vdd.n11948 vss 0.00413f
C21421 vdd.n11949 vss 0.0471f
C21422 vdd.t1071 vss 0.0471f
C21423 vdd.n11950 vss 0.00425f
C21424 vdd.n11951 vss 0.0424f
C21425 vdd.n11952 vss 0.0132f
C21426 vdd.n11953 vss 0.02f
C21427 vdd.n11954 vss 0.00425f
C21428 vdd.n11955 vss 0.00413f
C21429 vdd.n11956 vss 0.00251f
C21430 vdd.n11957 vss 0.0112f
C21431 vdd.n11958 vss 0.0128f
C21432 vdd.n11959 vss 0.0418f
C21433 vdd.n11960 vss 0.299f
C21434 vdd.n11961 vss 0.262f
C21435 vdd.n11962 vss 0.0471f
C21436 vdd.n11963 vss 0.00324f
C21437 vdd.n11964 vss 0.00324f
C21438 vdd.n11965 vss 0.0471f
C21439 vdd.n11966 vss 0.00324f
C21440 vdd.n11967 vss 0.00324f
C21441 vdd.n11968 vss 0.0424f
C21442 vdd.n11969 vss 0.0132f
C21443 vdd.n11970 vss 0.00925f
C21444 vdd.n11971 vss 0.00425f
C21445 vdd.t829 vss 0.0471f
C21446 vdd.n11973 vss 0.00425f
C21447 vdd.n11974 vss 0.02f
C21448 vdd.n11975 vss 0.0128f
C21449 vdd.n11976 vss 0.00413f
C21450 vdd.n11977 vss 0.00413f
C21451 vdd.n11978 vss 0.00413f
C21452 vdd.n11979 vss 0.00679f
C21453 vdd.n11980 vss 0.00517f
C21454 vdd.n11981 vss 0.00251f
C21455 vdd.t1082 vss 0.0471f
C21456 vdd.n11982 vss 0.00251f
C21457 vdd.n11983 vss 0.0112f
C21458 vdd.n11984 vss 0.0471f
C21459 vdd.n11985 vss 0.00324f
C21460 vdd.n11986 vss 0.00324f
C21461 vdd.n11987 vss 0.0424f
C21462 vdd.n11988 vss 0.0132f
C21463 vdd.n11989 vss 0.00925f
C21464 vdd.n11990 vss 0.00425f
C21465 vdd.t1471 vss 0.0471f
C21466 vdd.n11992 vss 0.00425f
C21467 vdd.n11993 vss 0.02f
C21468 vdd.n11994 vss 0.0128f
C21469 vdd.n11995 vss 0.00413f
C21470 vdd.n11996 vss 0.00413f
C21471 vdd.n11997 vss 0.00413f
C21472 vdd.n11998 vss 0.00679f
C21473 vdd.n11999 vss 0.00679f
C21474 vdd.n12000 vss 0.00517f
C21475 vdd.n12001 vss 0.00251f
C21476 vdd.t1083 vss 0.0471f
C21477 vdd.n12002 vss 0.00251f
C21478 vdd.n12003 vss 0.0112f
C21479 vdd.n12004 vss 0.0128f
C21480 vdd.t1084 vss 0.00134f
C21481 vdd.t1472 vss 0.0013f
C21482 vdd.n12005 vss 0.0332f
C21483 vdd.n12006 vss 0.0393f
C21484 vdd.n12007 vss 0.035f
.ends

