MACRO INV
  ORIGIN 0 0 ;
  FOREIGN INV 0 0 ;
  SIZE 5.16 BY 7.56 ;
  PIN N_BODY
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 2.84 6.58 4.04 6.86 ;
    END
  END N_BODY
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
      LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
      LAYER M2 ;
        RECT 2.15 0.28 3.01 0.56 ;
    END
  END OUT
  PIN IN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
      LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
      LAYER M2 ;
        RECT 2.15 4.48 3.01 4.76 ;
    END
  END IN
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
    END
  END VSS
  PIN P_BODY
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
    END
  END P_BODY
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
    END
  END VDD
  OBS 
  LAYER M1 ;
        RECT 3.745 0.335 3.995 3.865 ;
  LAYER M1 ;
        RECT 3.745 4.115 3.995 5.125 ;
  LAYER M1 ;
        RECT 3.745 6.215 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 3.865 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 3.865 ;
  LAYER M2 ;
        RECT 2.84 6.58 4.04 6.86 ;
  LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
  LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 3.865 ;
  LAYER M1 ;
        RECT 1.165 4.115 1.415 5.125 ;
  LAYER M1 ;
        RECT 1.165 6.215 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.595 0.335 1.845 3.865 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
  LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  END 
END INV
