magic
tech sky130B
magscale 1 2
timestamp 1688377021
<< metal1 >>
rect 2600 7740 2640 7780
rect 1480 7540 1680 7740
rect 4800 7720 4840 7760
rect 3100 6984 3140 7024
rect 5300 6078 5340 6118
rect 5600 4132 5640 4172
rect 5806 4122 5816 4182
rect 5876 4122 5886 4182
rect 6770 3842 6780 3902
rect 6840 3842 6850 3902
rect 7350 3462 7430 3472
rect 7350 3402 7360 3462
rect 7420 3402 7430 3462
rect 4964 1074 5084 1174
rect 5616 1074 5626 1174
rect 5726 1074 5736 1174
rect 7350 1070 7430 3402
rect 7350 1010 7360 1070
rect 7420 1010 7430 1070
rect 7350 1000 7430 1010
rect 1366 200 1798 600
rect 2560 200 2712 600
rect 5300 -154 5452 600
rect 5600 360 5640 400
rect 6780 360 6820 400
rect 7350 -116 7430 -106
rect 5300 -306 5600 -154
rect 7350 -176 7360 -116
rect 7420 -176 7430 -116
rect 7350 -2362 7430 -176
rect 7350 -2422 7360 -2362
rect 7420 -2422 7430 -2362
rect 7350 -2436 7430 -2422
rect 6770 -3100 6780 -3040
rect 6840 -3100 6850 -3040
rect 5806 -3502 5816 -3442
rect 5876 -3502 5886 -3442
rect 1480 -6940 1680 -6740
<< via1 >>
rect 5816 4122 5876 4182
rect 6780 3842 6840 3902
rect 7360 3402 7420 3462
rect 5626 1074 5726 1174
rect 7360 1010 7420 1070
rect 7360 -176 7420 -116
rect 7360 -2422 7420 -2362
rect 6780 -3100 6840 -3040
rect 5816 -3502 5876 -3442
<< metal2 >>
rect 5590 4186 5892 4196
rect 5590 4118 5600 4186
rect 5668 4182 5892 4186
rect 5668 4122 5816 4182
rect 5876 4122 5892 4182
rect 5668 4118 5892 4122
rect 5590 4108 5892 4118
rect 6770 3902 6852 3912
rect 6770 3842 6780 3902
rect 6840 3842 6852 3902
rect 6770 3838 6852 3842
rect 6770 3770 6776 3838
rect 6844 3770 6852 3838
rect 6770 3758 6852 3770
rect 4990 3648 5070 3660
rect 4990 3580 4996 3648
rect 5064 3580 5070 3648
rect 1580 1246 3180 1326
rect 4990 1268 5070 3580
rect 6760 3468 7440 3484
rect 6760 3400 6776 3468
rect 6844 3462 7440 3468
rect 6844 3402 7360 3462
rect 7420 3402 7440 3462
rect 6844 3400 7440 3402
rect 6760 3384 7440 3400
rect 1580 -200 1660 1246
rect 4990 1200 4996 1268
rect 5064 1200 5070 1268
rect 4990 1190 5070 1200
rect 5300 1194 5380 2246
rect 5300 1126 5306 1194
rect 5374 1126 5380 1194
rect 5300 1116 5380 1126
rect 5600 1174 5746 1200
rect 5600 1074 5626 1174
rect 5726 1074 5746 1174
rect 5600 998 5746 1074
rect 7180 1070 7430 1080
rect 7180 1010 7360 1070
rect 7420 1010 7430 1070
rect 7180 1000 7430 1010
rect 4948 846 5746 998
rect 5300 648 5380 660
rect 4948 200 5100 600
rect 5300 580 5306 648
rect 5374 580 5380 648
rect 4990 -126 5070 -112
rect 4990 -194 4996 -126
rect 5064 -194 5070 -126
rect 1580 -280 3180 -200
rect 3100 -660 3180 -280
rect 4990 -2612 5070 -194
rect 5300 -1486 5380 580
rect 7310 -116 7430 -106
rect 7310 -176 7360 -116
rect 7420 -176 7430 -116
rect 7310 -186 7430 -176
rect 4990 -2680 4996 -2612
rect 5064 -2680 5070 -2612
rect 6766 -2362 7430 -2348
rect 6766 -2422 7360 -2362
rect 7420 -2422 7430 -2362
rect 6766 -2436 7430 -2422
rect 6766 -2572 6854 -2436
rect 6766 -2640 6776 -2572
rect 6844 -2640 6854 -2572
rect 6766 -2650 6854 -2640
rect 4990 -2690 5070 -2680
rect 6770 -2964 6852 -2952
rect 6770 -3032 6776 -2964
rect 6844 -3032 6852 -2964
rect 6770 -3040 6852 -3032
rect 6770 -3100 6780 -3040
rect 6840 -3100 6852 -3040
rect 6770 -3110 6852 -3100
rect 5594 -3438 5892 -3428
rect 5594 -3506 5600 -3438
rect 5668 -3442 5892 -3438
rect 5668 -3502 5816 -3442
rect 5876 -3502 5892 -3442
rect 5668 -3506 5892 -3502
rect 5594 -3516 5892 -3506
<< via2 >>
rect 5600 4118 5668 4186
rect 6776 3770 6844 3838
rect 4996 3580 5064 3648
rect 6776 3400 6844 3468
rect 4996 1200 5064 1268
rect 5306 1126 5374 1194
rect 5306 580 5374 648
rect 4996 -194 5064 -126
rect 4996 -2680 5064 -2612
rect 6776 -2640 6844 -2572
rect 6776 -3032 6844 -2964
rect 5600 -3506 5668 -3438
<< metal3 >>
rect 4986 4186 5680 4196
rect 4986 4118 5600 4186
rect 5668 4118 5680 4186
rect 4986 4108 5680 4118
rect 4986 3648 5074 4108
rect 4986 3580 4996 3648
rect 5064 3580 5074 3648
rect 4986 3570 5074 3580
rect 6760 3838 6860 3848
rect 6760 3770 6776 3838
rect 6844 3770 6860 3838
rect 6760 3468 6860 3770
rect 6760 3400 6776 3468
rect 6844 3400 6860 3468
rect 6760 3384 6860 3400
rect 4986 1268 5074 1278
rect 4986 1200 4996 1268
rect 5064 1200 5074 1268
rect 4986 -126 5074 1200
rect 5290 1194 5390 1200
rect 5290 1126 5306 1194
rect 5374 1126 5390 1194
rect 5290 648 5390 1126
rect 5290 580 5306 648
rect 5374 580 5390 648
rect 5290 570 5390 580
rect 4986 -194 4996 -126
rect 5064 -194 5074 -126
rect 4986 -199 5074 -194
rect 6760 -2572 6860 -2556
rect 4986 -2612 5074 -2607
rect 4986 -2680 4996 -2612
rect 5064 -2680 5074 -2612
rect 4986 -3428 5074 -2680
rect 6760 -2640 6776 -2572
rect 6844 -2640 6860 -2572
rect 6760 -2964 6860 -2640
rect 6760 -3032 6776 -2964
rect 6844 -3032 6860 -2964
rect 6760 -3048 6860 -3032
rect 4986 -3438 5680 -3428
rect 4986 -3506 5600 -3438
rect 5668 -3506 5680 -3438
rect 4986 -3516 5680 -3506
use 3bit_dac  X1
timestamp 1688376520
transform 1 0 400 0 1 3812
box 800 -3212 6920 4012
use 3bit_dac  X2
timestamp 1688376520
transform 1 0 400 0 1 -3812
box 800 -3212 6920 4012
use sw  X3
timestamp 1687966408
transform 1 0 5600 0 1 480
box 0 -786 1720 720
<< labels >>
flabel metal1 1480 7540 1680 7740 0 FreeSans 256 0 0 0 vrefh
port 2 nsew
flabel metal1 1480 -6940 1680 -6740 0 FreeSans 256 0 0 0 vrefl
port 3 nsew
flabel metal1 4800 7720 4840 7760 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 2600 7740 2640 7780 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 3100 6984 3140 7024 0 FreeSans 256 0 0 0 d0
port 4 nsew
flabel metal1 5300 6078 5340 6118 0 FreeSans 256 0 0 0 d1
port 5 nsew
flabel metal1 5600 4132 5640 4172 0 FreeSans 256 0 0 0 d2
port 6 nsew
flabel metal1 5600 360 5640 400 0 FreeSans 256 0 0 0 d3
port 7 nsew
flabel metal1 6780 360 6820 400 0 FreeSans 256 0 0 0 vout
port 8 nsew
<< end >>
