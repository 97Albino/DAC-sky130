* NGSPICE file created from 2bit_dac.ext - technology: sky130B

.subckt sky130_fd_pr__res_high_po_0p35_2NY7PZ a_n35_109# a_n165_n671# a_n35_n541#
X0 a_n35_n541# a_n35_109# a_n165_n671# sky130_fd_pr__res_high_po_0p35 l=1.09
.ends

.subckt sky130_fd_pr__pfet_01v8_XPYSY6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 a_n50_n197# w_n246_n319# 0.119f
C1 a_n108_n100# w_n246_n319# 0.0852f
C2 a_50_n100# w_n246_n319# 0.0852f
C3 a_n50_n197# a_n108_n100# 0.0163f
C4 a_n50_n197# a_50_n100# 0.0163f
C5 a_n108_n100# a_50_n100# 0.0906f
C6 a_50_n100# VSUBS 0.0558f
C7 a_n108_n100# VSUBS 0.0558f
C8 a_n50_n197# VSUBS 0.179f
C9 w_n246_n319# VSUBS 1.41f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFH27D a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt sw vdd din vin1 vin2 vout vss
XXM1 vdd din m1_994_178# vdd vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM2 vdd m1_994_178# m1_688_n494# vdd vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM3 vdd m1_994_178# vout vin1 vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM4 vdd m1_688_n494# vin2 vout vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM5 m1_994_178# vss vss din sky130_fd_pr__nfet_01v8_ZFH27D
XXM6 m1_688_n494# vss vss m1_994_178# sky130_fd_pr__nfet_01v8_ZFH27D
XXM7 vout vss vin2 m1_994_178# sky130_fd_pr__nfet_01v8_ZFH27D
XXM8 vin1 vss vout m1_688_n494# sky130_fd_pr__nfet_01v8_ZFH27D
C0 vdd vin2 0.147f
C1 vdd vin1 0.259f
C2 din m1_994_178# 0.477f
C3 vdd vout 0.192f
C4 vdd m1_688_n494# 0.182f
C5 m1_994_178# vin2 0.0836f
C6 vin1 m1_994_178# 0.154f
C7 m1_994_178# vout 0.323f
C8 din vin2 4.93e-19
C9 din vin1 5.3e-19
C10 m1_994_178# m1_688_n494# 0.393f
C11 din m1_688_n494# 0.00777f
C12 vin1 vin2 0.514f
C13 vin2 vout -0.0571f
C14 vin1 vout -0.0258f
C15 vin2 m1_688_n494# 0.247f
C16 vin1 m1_688_n494# 0.382f
C17 vdd m1_994_178# 0.619f
C18 vout m1_688_n494# 0.374f
C19 din vdd 0.31f
C20 m1_688_n494# vss 0.491f
C21 m1_994_178# vss 0.662f
C22 din vss 0.416f
C23 vin1 vss 0.246f
C24 vout vss 0.195f
C25 vin2 vss 0.679f
C26 vdd vss 4.95f
.ends

.subckt x2bit_dac vdd vss vrefh vrefl d0 d1 vout
XXR1 vrefh vss X1/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XXR2 X1/vin2 vss X1/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XXR3 X1/vin2 vss X2/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XXR4 vrefl vss X2/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XX1 vdd d0 X1/vin1 X1/vin2 X3/vin1 vss sw
XX2 vdd d0 X2/vin1 vrefl X3/vin2 vss sw
XX3 vdd d1 X3/vin1 X3/vin2 vout vss sw
C0 X3/m1_688_n494# vss 0.339f
C1 X3/m1_994_178# vss 0.188f
C2 d1 vss 0.174f
C3 vout vss 0.0395f
C4 X2/m1_688_n494# vss 0.339f
C5 X2/m1_994_178# vss 0.188f
C6 d0 vss 0.348f
C7 X2/vin1 vss 0.186f
C8 X3/vin2 vss 0.517f
C9 vrefl vss 0.477f
C10 vdd vss 14.3f
C11 X1/m1_688_n494# vss 0.339f
C12 X1/m1_994_178# vss 0.188f
C13 X1/vin1 vss 0.186f
C14 X3/vin1 vss 0.226f
C15 X1/vin2 vss 0.477f
.ends

