* NGSPICE file created from sw.ext - technology: sky130B

.subckt sky130_fd_pr__pfet_01v8_XHX9Y6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_XPYSY6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFH27D a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_HEL24J a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt sw vdd vss din vin1 vin2 vout
XXM2 XM4/w_n246_n319# m1_800_578# m1_488_106# vdd sky130_fd_pr__pfet_01v8_XHX9Y6
XXM3 XM4/w_n246_n319# m1_800_578# vout vin1 sky130_fd_pr__pfet_01v8_XHX9Y6
XXM4 XM4/w_n246_n319# m1_488_106# vin2 vout sky130_fd_pr__pfet_01v8_XPYSY6
XXM5 m1_800_578# VSUBS vss din sky130_fd_pr__nfet_01v8_ZFH27D
XXM6 m1_488_106# VSUBS vss m1_800_578# sky130_fd_pr__nfet_01v8_HEL24J
Xsky130_fd_pr__pfet_01v8_XPYSY6_0 XM4/w_n246_n319# din m1_800_578# vdd sky130_fd_pr__pfet_01v8_XPYSY6
XXM7 vout VSUBS vin2 m1_800_578# sky130_fd_pr__nfet_01v8_HEL24J
XXM8 vin1 VSUBS vout m1_488_106# sky130_fd_pr__nfet_01v8_ZFH27D
.ends

