magic
tech sky130B
magscale 1 2
timestamp 1687214096
<< checkpaint >>
rect 3773 10526 6763 10579
rect 3773 8211 7180 10526
rect 2179 6473 7180 8211
rect 2179 4139 7597 6473
rect -235 2585 7597 4139
rect -1313 -713 7597 2585
rect -1260 -925 7597 -713
rect -1260 -2860 1460 -925
rect 1640 -978 7597 -925
rect 2179 -1031 7597 -978
rect 2976 -1084 7597 -1031
rect 3773 -1137 7597 -1084
rect 4190 -1190 7597 -1137
rect 4607 -1243 7597 -1190
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__nfet_01v8_34YWRA  xm1
timestamp 0
transform 1 0 243 0 1 936
box -296 -389 296 389
use sky130_fd_pr__nfet_01v8_34YWRA  xm2
timestamp 0
transform 1 0 782 0 1 883
box -296 -389 296 389
use sky130_fd_pr__pfet_01v8_GGAEPD  xm3
timestamp 0
transform 1 0 1321 0 1 1660
box -296 -1219 296 1219
use sky130_fd_pr__pfet_01v8_GGAEPD  xm4
timestamp 0
transform 1 0 1860 0 1 1607
box -296 -1219 296 1219
use sky130_fd_pr__nfet_01v8_EF4BLE  xm5
timestamp 0
transform 1 0 2528 0 1 1545
box -425 -1210 425 1210
use sky130_fd_pr__nfet_01v8_6WXQK8  xm6
timestamp 0
transform 1 0 3196 0 1 1492
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_RLGYC7  xm7
timestamp 0
transform 1 0 3864 0 1 3590
box -425 -3361 425 3361
use sky130_fd_pr__nfet_01v8_6WGMFU  xm8
timestamp 0
transform 1 0 4661 0 1 3528
box -425 -3352 425 3352
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR1
timestamp 0
transform 1 0 5268 0 1 4721
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_NKSDAM  xR2
timestamp 0
transform 1 0 5685 0 1 4668
box -235 -4598 235 4598
use sky130_fd_pr__res_high_po_0p69_YVB7ZU  xR3
timestamp 0
transform 1 0 6102 0 1 2615
box -235 -2598 235 2598
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 in1
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 in2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 out2
port 4 nsew
<< end >>
