* SPICE3 file created from 8bit_dac_flat.ext - technology: sky130B

.subckt x8bit_dac_flat vrefh vrefl d0 d1 d2 d3 d4 d5 d6 d7 vout vss vdd
X0 X1.X2.X1.X2.X3.vin2 a_19722_10916# X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 X1.X1.X1.X2.X1.X2.X1.vin2 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X3 X2.X2.X1.X2.X1.X1.X3.vin2 a_46116_15634# X2.X2.X1.X2.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X4 X2.X2.X1.X3.vin1 a_49002_18540# X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X5 vdd a_11072_4110# a_10686_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X6 a_46502_9916# a_46116_9916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X7 X2.X1.X1.X1.X1.X2.X3.vin1 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X8 vss a_52492_18358# a_52106_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X9 X1.X2.X2.X2.X1.X1.X3.vin2 a_23512_20264# X1.X2.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X10 a_35312_892# a_34926_892# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 a_2582_13728# a_2196_13728# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X12 a_16836_25164# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X13 vdd a_8872_16452# a_8486_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 a_33676_12822# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X15 X1.X1.X2.X1.X2.X1.X1.vin2 a_11072_11734# X1.X1.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X16 X2.X2.X1.X1.X1.X2.X3.vin1 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X17 a_46502_4198# a_46116_4198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X19 X2.X2.X2.X1.X1.X2.X3.vin1 a_54606_7922# X2.X2.X2.X1.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X20 X2.X1.X1.X1.X2.X2.X3.vin2 a_34062_20446# X2.X1.X1.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 X2.X2.X2.X2.X1.X2.X1.vin1 a_54992_23170# X2.X2.X2.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X22 X2.X1.X2.X2.X1.X1.vout a_37766_20264# X2.X1.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X23 a_16836_4198# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X24 X1.X2.X2.X1.X1.X1.vout a_23126_5016# X1.X2.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X25 X2.X2.X1.X2.X3.vin1 a_49002_10916# X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X26 X1.X1.X1.X2.X1.X1.X3.vin2 a_4782_16634# X1.X1.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X27 X1.X1.X2.X1.X1.X1.X1.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X28 vss d0 a_54992_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X29 vdd a_23212_6962# a_22826_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 a_46502_15634# a_46116_15634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X31 vss d0 a_25712_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X32 X1.X1.X2.X3.vin2 a_8186_25982# X1.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X33 a_17222_19446# a_16836_19446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X34 X2.X1.X1.X1.X2.X1.vout a_34362_22312# X2.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X35 X1.X2.X1.X1.X1.X2.X3.vin2 a_19422_28070# X1.X2.X1.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X36 vdd d0 a_11072_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X37 X2.X1.X1.X2.X2.X2.X1.vin2 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X38 X1.X1.X1.X1.X1.X1.X3.vin2 a_2196_30882# X1.X1.X1.X1.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X39 X1.X2.X2.X2.X1.X2.X1.vin2 a_25712_23170# X1.X2.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X40 a_19422_31882# a_19036_31882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X41 X2.X2.X2.X2.X2.X1.vout a_52492_29834# X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X42 X2.X2.vrefh X2.X2.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X43 X2.X2.X1.X1.X2.X2.vout a_49002_22312# X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X44 a_46502_28976# a_46116_28976# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X45 vdd d1 a_38152_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X46 a_4782_31882# a_4396_31882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X47 vdd d0 a_25712_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X48 X1.X1.X1.X2.X1.X2.X2.vin1 a_2582_11822# X1.X1.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X49 vss a_25712_28888# a_25326_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X50 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X51 X1.X2.X1.X2.vrefh a_17222_19446# X1.X2.X1.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X52 a_2582_32788# a_2196_32788# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X53 X2.X2.X2.X2.X2.X2.X3.vin1 a_52792_31700# X2.X2.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X54 X1.X2.X1.X1.X2.X2.vout a_19036_20446# X1.X2.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X55 X2.X1.X2.X2.X1.X2.X3.vin1 a_39966_23170# X2.X1.X2.X2.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X56 X2.X2.X2.X2.X2.X2.X3.vin2 a_54606_32700# vrefl vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X57 X2.X2.X2.X2.X2.X2.X3.vin1 a_54606_30794# X2.X2.X2.X2.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X58 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X59 a_5082_18540# a_4696_18540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X60 X1.X1.X1.X1.X3.vin1 a_4696_29936# X1.X1.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X61 vdd d0 a_54992_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X62 vdd d0 a_25712_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X63 a_4782_5198# a_4396_5198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X64 vdd d3 a_23212_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X65 X1.X1.X1.X1.X2.X1.X1.vin2 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X66 vss a_40352_15546# a_39966_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X67 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X68 X2.X1.X1.X1.X2.X1.vout a_33676_24258# X2.X1.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X69 a_5646_892# d5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X70 a_4396_20446# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X71 X2.X1.X1.X3.vin1 a_33976_26164# X2.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X72 X2.X1.X2.X2.X3.vin2 a_37466_29834# X2.X1.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X73 a_5082_10916# a_4696_10916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X74 X2.X1.X2.X2.X1.X1.X1.vin1 a_40352_19358# X2.X1.X2.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X75 a_17222_6104# a_16836_6104# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X76 X1.X2.X1.X1.X2.X1.X1.vin1 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X77 X2.X1.X1.X2.X2.X1.vout a_34362_7064# X2.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X78 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X79 vrefl a_54992_32700# X2.X2.X2.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X80 X2.X1.X2.X2.X2.X2.vout a_37766_31700# X2.X1.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X81 vdd a_23512_8828# a_23126_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X82 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X83 X1.X1.X2.X1.X1.X1.X3.vin1 a_8872_5016# X1.X1.X2.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X84 X1.X1.X1.X2.X1.X2.X3.vin1 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X85 X2.X1.X1.X2.X2.X2.X3.vin2 a_34062_5198# X2.X1.X1.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X86 a_31862_19446# a_31476_19446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X87 X1.X1.X2.X2.X2.X1.vout a_8486_27888# X1.X1.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X88 X2.X2.X2.X1.X1.X1.X3.vin1 a_52792_5016# X2.X2.X2.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X89 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X90 X2.X2.X2.vrefh a_46502_4198# X2.X2.X1.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X91 vdd a_54992_7922# a_54606_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X92 vss a_11072_6016# a_10686_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X93 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X94 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X95 a_34062_31882# a_33676_31882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X96 X1.X2.X1.X1.X3.vin1 a_19336_29936# X1.X2.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X97 vss d0 a_11072_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X98 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X99 X1.X1.X2.X2.X2.X2.X1.vin1 a_11072_30794# X1.X1.X2.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X100 X2.X1.X1.X2.X2.vrefh a_31862_11822# X2.X1.X1.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X101 X1.X1.X2.X1.X2.X1.X3.vin1 a_10686_11734# X1.X1.X2.X1.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X102 X2.X2.X2.X1.X2.X2.X3.vin1 a_54606_15546# X2.X2.X2.X1.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X103 X1.X2.X2.X2.X1.X1.X3.vin1 a_25326_19358# X1.X2.X2.X2.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X104 vss a_25712_19358# a_25326_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X105 a_4782_28070# a_4396_28070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X106 vss a_52792_16452# a_52406_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X107 X2.X1.X2.X2.X2.X2.X3.vin2 a_39966_32700# X2.X1.X2.X2.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X108 a_48316_28070# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X109 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X110 vdd d0 a_54992_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X111 X1.X3.vin2 a_20286_892# X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X112 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X113 a_46116_30882# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X114 vss d0 a_54992_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X115 a_49002_18540# a_48616_18540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X116 X2.X1.X1.X1.X3.vin2 a_33976_22312# X2.X1.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X117 a_17222_23258# a_16836_23258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X118 a_16836_19446# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X119 X1.X2.X1.X2.X2.X1.X3.vin2 a_16836_8010# X1.X2.X1.X2.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X120 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X121 a_19036_31882# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X122 X2.X1.X1.X2.X1.X1.X1.vin1 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X123 X2.X2.X2.X1.X2.X2.X2.vin1 a_54992_17452# X2.X2.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X124 X1.X2.X1.X2.X1.X2.X3.vin2 a_16836_11822# X1.X2.X1.X2.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X125 X1.X1.X1.X3.vin1 a_4696_26164# X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X126 vss d4 a_37852_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X127 a_48316_20446# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X128 X2.X1.X2.X2.X2.X2.vrefh a_40352_28888# X2.X1.X2.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X129 X1.X2.X2.X2.X2.X1.vout a_23126_27888# X1.X2.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X130 vdd a_52792_24076# a_52406_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X131 X1.X1.X1.X2.X1.X2.X3.vin2 a_2196_11822# X1.X1.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X132 a_19422_12822# a_19036_12822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X133 a_49002_10916# a_48616_10916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X134 vss d2 a_8572_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X135 vss d0 a_54992_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X136 vdd a_37852_6962# a_37466_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X137 a_2582_6104# a_2196_6104# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X138 vss d1 a_8872_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X139 vss d2 a_52492_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X140 a_2196_11822# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X141 X1.X1.X1.X1.X2.X1.X3.vin1 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X142 X1.X2.X2.X2.vrefh a_25712_17452# X1.X2.X2.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X143 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X144 X2.X2.X1.X2.X2.X1.X3.vin1 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X145 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X146 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X147 a_19722_7064# a_19336_7064# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X148 X1.X1.X2.X2.X1.X2.vout a_8572_22210# X1.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X149 X1.X2.X1.X2.X1.X1.X3.vin1 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X150 X2.X2.X2.X2.X2.X2.vout a_52492_29834# X2.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X151 a_2196_6104# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X152 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X153 X2.X1.X2.X1.X2.X2.X3.vin2 a_39966_17452# X2.X1.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X154 a_49002_22312# a_48616_22312# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X155 X1.X1.X1.X2.X2.X1.X3.vin2 a_4782_9010# X1.X1.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X156 X1.X1.X2.X1.X1.X2.X3.vin1 a_10686_7922# X1.X1.X2.X1.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X157 vdd a_54992_26982# a_54606_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X158 a_31476_21352# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X159 X1.X2.X2.X2.X2.X1.X3.vin2 a_25326_28888# X1.X2.X2.X2.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X160 vdd d0 a_54992_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X161 vss a_54992_25076# a_54606_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X162 a_46116_13728# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X163 vdd d0 a_25712_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X164 vdd d0 a_40352_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X165 vss a_23212_22210# a_22826_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X166 X2.X1.X2.X1.X3.vin2 a_37852_10734# X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X167 a_19336_7064# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X168 X1.X2.X1.X1.X2.X2.X3.vin2 a_19422_20446# X1.X2.X1.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X169 X1.X2.X2.X2.X1.X2.X2.vin1 a_25712_25076# X1.X2.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X170 a_2196_17540# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X171 X2.X1.X2.X1.X1.X2.X3.vin1 a_39966_7922# X2.X1.X2.X1.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X172 X1.X2.X1.X3.vin1 a_19336_26164# X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X173 a_31862_23258# a_31476_23258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X174 X2.X2.X1.X1.X1.X2.X3.vin1 a_48702_28070# X2.X2.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X175 X2.X2.X2.X1.X1.X2.X1.vin2 a_54992_7922# X2.X2.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X176 X2.X2.X2.X2.X1.X1.vout a_52492_22210# X2.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X177 X1.X1.X3.vin2 a_8186_18358# X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X178 X2.X2.X1.X1.X1.X2.vrefh a_46502_30882# X2.X2.X1.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X179 X1.X2.X1.X1.X2.X2.X2.vin1 a_17222_19446# X1.X2.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X180 X1.X1.X2.X2.X2.X2.X3.vin1 a_10686_30794# X1.X1.X2.X2.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X181 X2.X1.X1.X1.X1.X2.X1.vin1 a_31862_28976# X2.X1.X1.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X182 X2.X1.X2.X2.X3.vin2 a_37466_29834# X2.X1.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X183 X2.X2.X2.X2.X2.X1.X1.vin2 a_54992_26982# X2.X2.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X184 X2.X1.X2.X2.X1.X1.X1.vin2 a_40352_19358# X2.X1.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X185 X1.X1.X1.X1.X3.vin1 a_4696_29936# X1.X1.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X186 vdd a_38152_8828# a_37766_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X187 X1.X1.X2.X2.X1.X2.X1.vin2 a_11072_23170# X1.X1.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X188 a_33676_24258# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X189 X1.X2.X1.X2.X2.X2.X1.vin2 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X190 X1.X1.X1.X2.X2.X1.X3.vin2 a_2196_8010# X1.X1.X1.X2.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X191 a_34062_12822# a_33676_12822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X192 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X193 vdd d1 a_8872_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X194 a_48316_16634# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X195 vdd d1 a_23512_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X196 X2.X2.X1.X1.X2.X2.X3.vin1 a_48702_20446# X2.X2.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X197 X1.X2.X2.X2.X1.X2.vout a_23212_22210# X1.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X198 a_13696_892# d6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X199 X1.X2.X1.X2.X2.X2.vout a_19036_5198# X1.X2.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X200 X2.X2.X2.X1.X2.X1.vout a_52492_14586# X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X201 a_16836_23258# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X202 X2.X1.X2.X2.X3.vin1 a_37466_22210# X2.X1.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X203 a_4396_5198# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X204 X1.X1.X1.X2.X1.X2.vout a_4396_12822# X1.X1.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X205 vss a_54992_9828# a_54606_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X206 X1.X1.X2.X2.X3.vin2 a_8572_25982# X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X207 a_46116_11822# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X208 X3.vin1 a_28482_892# vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X209 vss a_25712_13640# a_25326_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X210 X2.X2.X1.X2.vrefh X2.X2.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X211 X1.X2.X1.X1.X1.X2.X3.vin1 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X212 vdd a_11072_13640# a_10686_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X213 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X214 X2.X1.X2.X2.X2.X1.X3.vin1 a_39966_26982# X2.X1.X2.X2.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X215 X1.X2.X2.X2.X1.X1.X3.vin1 a_25326_19358# X1.X2.X2.X2.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X216 a_31476_32788# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X217 X2.X1.X2.X2.X1.X2.X3.vin2 a_38152_24076# X2.X1.X2.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X218 a_5082_7064# a_4696_7064# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X219 a_19036_12822# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X220 X2.X1.X2.X1.X1.X2.vout a_37852_6962# X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X221 X2.X2.X2.X1.X2.X2.vout a_52406_16452# X2.X2.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X222 a_31476_17540# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X223 X1.X1.X1.X1.X2.X1.X2.vin1 a_2582_23258# X1.X1.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X224 a_46116_25164# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X225 vss a_23212_25982# a_22826_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X226 vss d0 a_25712_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X227 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X228 X2.X2.X1.X2.X1.X2.X1.vin2 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X229 X1.X1.X1.X1.X1.X2.vout a_5082_29936# X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X230 a_2196_28976# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X231 a_31476_8010# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X232 X1.X2.X1.X1.X3.vin1 a_19336_29936# X1.X2.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X233 vss d1 a_38152_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X234 vss d0 a_40352_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X235 X2.X1.X2.X1.X3.vin2 a_37466_14586# X2.X1.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X236 vdd a_25712_21264# a_25326_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X237 a_4696_7064# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X238 X2.X1.X1.X1.X2.X1.X3.vin2 a_34062_24258# X2.X1.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X239 a_34062_9010# a_33676_9010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X240 a_31476_9916# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X241 a_4782_20446# a_4396_20446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X242 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X243 X2.X1.X1.X2.X2.X1.X3.vin1 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X244 X2.X2.X2.X2.X1.X2.vout a_52406_24076# X2.X2.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X245 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X246 X2.X1.X2.X2.X2.X1.vout a_37852_29834# X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X247 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X248 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X249 vdd a_40352_28888# a_39966_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X250 X1.X2.X2.X2.X3.vin2 a_23212_25982# X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X251 X2.X1.X1.X1.X1.X1.X3.vin2 a_31476_30882# X2.X1.X1.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X252 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X253 X2.X2.X1.X2.X1.X1.X3.vin2 a_48702_16634# X2.X2.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X254 X2.X2.X1.X1.X1.X2.vout a_48316_28070# X2.X2.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X255 a_49566_892# d5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X256 X2.X2.X1.X1.X1.X1.X3.vin2 a_46116_30882# X2.X2.X1.X1.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X257 a_17222_4198# a_16836_4198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X258 X1.X1.X2.X2.X2.X1.X3.vin1 a_8872_27888# X1.X1.X2.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X259 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X260 X1.X2.X2.X1.X1.X2.X3.vin1 a_25326_7922# X1.X2.X2.X1.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X261 X1.X2.X1.X1.X2.X2.vrefh a_17222_23258# X1.X2.X1.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X262 a_31476_15634# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X263 a_34362_18540# a_33976_18540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X264 X1.X2.X1.X1.X2.X1.vout a_19036_24258# X1.X2.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X265 vdd d0 a_54992_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X266 X2.X1.X2.X1.X1.X2.X1.vin2 a_40352_7922# X2.X1.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X267 X2.X2.X1.X2.X1.X2.X2.vin1 a_46502_11822# X2.X2.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X268 X2.X2.X2.X2.X2.X1.X3.vin1 a_54606_26982# X2.X2.X2.X2.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X269 X2.X2.X2.X2.X1.X2.X3.vin2 a_52792_24076# X2.X2.X2.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X270 X1.X1.X2.X2.X1.X2.X3.vin1 a_10686_23170# X1.X1.X2.X2.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X271 X2.X2.X2.X2.X1.X2.X3.vin2 a_54606_25076# X2.X2.X2.X2.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X272 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X273 X1.X2.X2.X2.X1.X1.X1.vin1 a_25712_19358# X1.X2.X2.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X274 X2.X2.X1.X1.X2.X2.vout a_48316_20446# X2.X2.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X275 vss d0 a_25712_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X276 X2.X2.X1.X1.X3.vin1 a_48616_29936# X2.X2.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X277 a_31476_28976# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X278 vdd a_23512_27888# a_23126_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X279 X1.X2.X2.X2.X3.vin1 a_22826_22210# X1.X2.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X280 a_17222_21352# a_16836_21352# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X281 X1.X2.X1.X2.X2.X2.X3.vin1 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X282 a_14082_892# a_13696_892# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X283 vss d1 a_52792_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X284 a_4396_24258# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X285 X2.X2.X1.X1.X2.X1.X1.vin2 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X286 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X287 a_34362_10916# a_33976_10916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X288 a_48702_28070# a_48316_28070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X289 a_4696_26164# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X290 a_46502_30882# a_46116_30882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X291 vdd a_25712_32700# a_25326_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X292 X2.X1.X2.X1.X2.X2.vrefh a_40352_13640# X2.X1.X2.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X293 vss a_25712_30794# a_25326_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X294 vss d2 a_8572_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X295 X1.X1.X2.X2.vrefh a_11072_17452# X1.X1.X2.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X296 a_19336_18540# d4 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X297 vss a_52792_27888# a_52406_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X298 vss d1 a_8872_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X299 X2.X1.X2.X2.X1.X2.vout a_37766_24076# X2.X1.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X300 X2.X2.X2.X1.X1.X2.X2.vin1 a_54992_9828# X2.X2.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X301 vss d1 a_52792_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X302 a_34362_22312# a_33976_22312# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X303 X1.X1.X1.X1.X2.X1.X3.vin2 a_2196_23258# X1.X1.X1.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X304 X1.X2.X2.X2.X2.X1.X3.vin1 a_23512_27888# X1.X2.X2.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X305 X1.X1.X1.X1.X3.vin1 a_5082_26164# X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X306 a_48702_20446# a_48316_20446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X307 vdd d1 a_52792_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X308 a_19422_24258# a_19036_24258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X309 vss a_11072_21264# a_10686_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X310 X1.X2.X2.X1.X1.X1.X1.vin2 a_25712_4110# X1.X2.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X311 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X312 X2.X2.X1.X2.X1.X2.X3.vin1 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X313 X2.X2.X1.X2.X2.X1.vout a_48316_9010# X2.X2.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X314 vss a_38152_16452# a_37766_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X315 X2.X1.X1.X1.X1.X2.X3.vin2 a_31476_27070# X2.X1.X1.X1.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X316 X1.X2.X2.X1.X1.X2.vout a_23212_6962# X1.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X317 a_19336_10916# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X318 X2.X1.X2.X2.X1.X1.X2.vin1 a_40352_21264# X2.X1.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X319 a_2582_11822# a_2196_11822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X320 X1.X1.X2.X2.X1.X2.X2.vin1 a_11072_25076# X1.X1.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X321 a_16836_9916# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X322 X2.X2.X2.X1.X1.X2.X3.vin2 a_54606_9828# X2.X2.X2.X1.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X323 X1.X2.X2.X1.X2.X1.X3.vin2 a_25326_13640# X1.X2.X2.X1.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X324 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X325 vss d0 a_40352_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X326 X2.X1.X1.X2.X1.X1.vout a_33676_16634# X2.X1.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X327 a_2582_4198# a_2196_4198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X328 a_31862_21352# a_31476_21352# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X329 X1.X2.X2.X3.vin2 a_22826_25982# X1.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X330 vdd d0 a_54992_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X331 a_19336_22312# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X332 X1.X2.X2.X2.X2.X2.vrefh a_25712_28888# X1.X2.X2.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X333 vss d0 a_54992_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X334 vdd a_38152_24076# a_37766_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X335 a_46116_8010# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X336 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X337 a_17222_32788# a_16836_32788# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X338 vdd a_54992_11734# a_54606_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X339 a_46502_13728# a_46116_13728# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X340 X2.X2.X1.X2.X1.X1.vout a_48316_16634# X2.X2.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X341 a_4696_22312# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X342 vdd a_25712_7922# a_25326_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X343 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X344 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X345 vdd a_25712_15546# a_25326_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X346 a_17222_17540# a_16836_17540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X347 vss d2 a_23212_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X348 a_2582_17540# a_2196_17540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X349 X1.X2.X2.X2.X1.X1.X3.vin2 a_25326_21264# X1.X2.X2.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X350 a_48702_9010# a_48316_9010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X351 X1.X1.X1.X2.X3.vin1 a_4696_14688# X1.X1.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X352 X1.X1.X1.X2.X2.X2.X3.vin1 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X353 X1.X1.X2.X1.X1.X1.vout a_8486_5016# X1.X1.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X354 X1.X1.X2.X3.vin2 a_8572_18358# X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X355 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X356 a_33976_18540# d4 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X357 X2.X2.X1.X3.vin1 a_48616_26164# X2.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X358 X2.X2.X1.X2.X1.X2.X3.vin2 a_46116_11822# X2.X2.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X359 vdd d3 a_8572_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X360 a_17222_9916# a_16836_9916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X361 X2.X1.X2.X2.X2.X2.vout a_37852_29834# X2.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X362 X1.X1.X1.X1.X1.X1.vout a_5082_29936# X1.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X363 vdd d0 a_40352_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X364 a_34062_24258# a_33676_24258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X365 a_16836_21352# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X366 vdd a_8872_12640# a_8486_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X367 vss a_23212_18358# a_22826_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X368 a_48702_16634# a_48316_16634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X369 X2.X2.X1.X1.X2.X1.X3.vin1 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X370 a_33976_10916# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X371 X2.X2.X2.X1.X1.X1.X3.vin1 a_54606_4110# X2.X2.X2.X1.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X372 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X373 X2.X2.X2.X3.vin1 a_52492_18358# X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X374 X2.X1.X2.X2.X2.X2.X2.vin1 a_40352_32700# X2.X1.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X375 X2.X1.X2.X2.X2.X2.X1.vin2 a_40352_30794# X2.X1.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X376 vss a_8572_14586# a_8186_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X377 X1.X1.X2.X1.X2.X2.X3.vin2 a_10686_17452# X1.X1.X2.X1.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X378 X2.X1.X2.X2.X1.X1.vout a_37852_22210# X2.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X379 vss d0 a_54992_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X380 X1.X1.X1.X2.X1.X2.X3.vin2 a_4782_12822# X1.X1.X1.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X381 a_46116_23258# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X382 vss d0 a_25712_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X383 a_46502_11822# a_46116_11822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X384 vss d0 a_25712_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X385 X1.X2.X1.X1.X2.X1.X3.vin2 a_19422_24258# X1.X2.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X386 a_17222_15634# a_16836_15634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X387 vdd d0 a_11072_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X388 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X389 a_33976_22312# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X390 X1.X2.X1.X2.X3.vin1 a_19336_14688# X1.X2.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X391 a_48616_29936# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X392 X1.X2.X1.X1.X3.vin2 a_19722_26164# X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X393 X1.X2.X2.X2.X1.X1.X1.vin2 a_25712_19358# X1.X2.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X394 a_31862_32788# a_31476_32788# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X395 a_19036_24258# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X396 X1.X2.X2.X3.vin2 a_23212_18358# X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X397 X1.X2.vrefh X1.X2.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X398 a_31862_17540# a_31476_17540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X399 a_46502_25164# a_46116_25164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X400 vss d3 a_23212_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X401 a_17222_28976# a_16836_28976# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X402 X2.X1.X2.X1.X1.X2.X2.vin1 a_40352_9828# X2.X1.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X403 a_2582_28976# a_2196_28976# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X404 X1.X1.X2.X2.X1.X2.X3.vin2 a_10686_25076# X1.X1.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X405 X2.X1.X3.vin2 a_37466_18358# X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X406 X1.X2.X2.X2.X2.X2.X3.vin2 a_25326_32700# X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X407 X2.X1.X1.X2.X2.X1.vout a_33676_9010# X2.X1.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X408 X1.X2.X2.X2.X2.X2.X3.vin1 a_25326_30794# X1.X2.X2.X2.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X409 X1.X2.X1.X2.X2.X1.X3.vin2 a_19422_9010# X1.X2.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X410 X2.X1.X2.X1.X2.X1.vout a_37852_14586# X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X411 vdd d0 a_25712_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X412 vdd d0 a_40352_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X413 X2.X2.X2.X2.X2.X1.vout a_52406_27888# X2.X2.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X414 X2.X2.X1.X1.X3.vin1 a_48616_29936# X2.X2.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X415 vss a_40352_11734# a_39966_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X416 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X417 a_31862_9916# a_31476_9916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X418 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X419 vss a_11072_15546# a_10686_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X420 X2.X2.X1.X2.X2.X1.X3.vin2 a_48702_9010# X2.X2.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X421 a_16836_32788# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X422 X2.X1.X2.X1.X2.X2.X1.vin1 a_40352_15546# X2.X1.X2.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X423 a_16836_17540# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X424 X1.X1.X2.X2.X1.X1.X1.vin1 a_11072_19358# X1.X1.X2.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X425 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X426 X1.X2.X1.X1.X2.X2.X1.vin1 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X427 X2.X1.X1.X1.X1.X1.X2.vin1 a_31862_30882# X2.X1.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X428 X1.X2.X2.X1.X1.X1.X2.vin1 a_25712_6016# X1.X2.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X429 a_31862_15634# a_31476_15634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X430 vdd a_8572_25982# a_8186_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X431 X1.X2.X1.X1.X2.X1.vout a_19722_22312# X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X432 X2.X1.X2.X1.X1.X1.X3.vin1 a_38152_5016# X2.X1.X2.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X433 a_16836_9916# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X434 vdd a_54992_4110# a_54606_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X435 X2.X2.X1.X1.X2.X1.X2.vin1 a_46502_23258# X2.X2.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X436 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X437 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X438 a_31476_4198# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X439 X2.X1.X1.X2.X1.X2.vout a_34362_14688# X2.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X440 X2.X1.X1.X1.X2.X2.X3.vin2 a_31476_19446# X2.X1.X1.X1.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X441 X2.X2.X2.X1.X2.X1.X3.vin1 a_54606_11734# X2.X2.X2.X1.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X442 X2.X2.X1.X1.X1.X2.vout a_49002_29936# X2.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X443 a_31862_28976# a_31476_28976# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X444 X2.X2.X1.X2.X2.X1.X3.vin2 a_46116_8010# X2.X2.X1.X2.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X445 X1.X2.X2.X1.X2.X2.X3.vin1 a_25326_15546# X1.X2.X2.X1.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X446 X3.vin2 a_28482_892# vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X447 a_4782_24258# a_4396_24258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X448 X1.X2.X1.X1.X1.X1.X3.vin2 a_16836_30882# X1.X2.X1.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X449 X1.X1.X1.X2.X2.X2.X1.vin2 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X450 X2.X2.X2.X1.X1.X1.X3.vin2 a_54606_6016# X2.X2.X2.X1.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X451 vss a_52792_12640# a_52406_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X452 vdd d0 a_11072_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X453 vss a_8872_20264# a_8486_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X454 a_5082_26164# a_4696_26164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X455 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X456 vdd d0 a_25712_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X457 a_48616_26164# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X458 vss d0 a_25712_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X459 X2.X2.X2.X1.X1.X1.X1.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X460 a_16836_15634# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X461 a_19722_18540# a_19336_18540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X462 a_2196_30882# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X463 vss d1 a_52792_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X464 X1.X2.X1.X2.X2.X2.X3.vin2 a_16836_4198# X1.X2.X1.X2.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X465 X2.X1.X1.X1.X2.X1.X3.vin1 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X466 X1.X2.X2.X1.X1.X2.X3.vin2 a_23512_8828# X1.X2.X2.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X467 X2.X2.X2.X1.X2.X1.X2.vin1 a_54992_13640# X2.X2.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X468 X1.X2.X3.vin2 a_22826_18358# X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X469 vss a_40352_7922# a_39966_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X470 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X471 a_16836_28976# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X472 vdd a_52792_20264# a_52406_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X473 vss d0 a_11072_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X474 X1.X2.X1.X1.X1.X1.X1.vin1 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X475 a_19036_9010# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X476 X1.X1.X2.X2.X2.X2.vrefh a_11072_28888# X1.X1.X2.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X477 vss d1 a_38152_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X478 X1.X2.X1.X2.X1.X1.X1.vin2 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X479 X2.X1.X1.X1.X2.vrefh a_31862_27070# X2.X1.X1.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X480 a_20672_892# a_20286_892# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X481 a_19722_10916# a_19336_10916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X482 X2.X2.X2.X1.X3.vin1 a_52106_6962# X2.X2.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X483 X2.X1.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X484 vdd a_40352_30794# a_39966_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X485 X1.X2.X2.X1.X2.X2.vrefh a_25712_13640# X1.X2.X2.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X486 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X487 X1.X3.vin2 a_14082_892# X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X488 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X489 vss d0 a_40352_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X490 vss a_38152_27888# a_37766_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X491 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X492 X2.X1.X1.X2.X1.X1.X3.vin1 a_34062_16634# X2.X1.X1.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X493 X1.X2.X1.X2.X2.X1.X1.vin2 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X494 X2.X1.X2.X1.X2.X1.X3.vin2 a_39966_13640# X2.X1.X2.X1.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X495 X1.X1.X1.X2.X2.X2.X3.vin2 a_4782_5198# X1.X1.X1.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X496 a_19722_22312# a_19336_22312# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X497 X1.X1.X2.X1.X1.X1.X3.vin1 a_10686_4110# X1.X1.X2.X1.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X498 X1.X1.X2.X2.X1.X1.X3.vin1 a_10686_19358# X1.X1.X2.X2.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X499 vdd d1 a_38152_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X500 vdd a_54992_23170# a_54606_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X501 vdd a_25712_26982# a_25326_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X502 vdd d0 a_25712_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X503 vdd d0 a_54992_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X504 a_5082_22312# a_4696_22312# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X505 X1.X1.X2.X1.X1.X2.X1.vin2 a_11072_7922# X1.X1.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X506 vss a_25712_25076# a_25326_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X507 vdd d0 a_25712_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X508 X1.X2.X1.X1.X1.X2.X3.vin2 a_16836_27070# X1.X2.X1.X1.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X509 a_33676_28070# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X510 X1.X2.X2.X2.X1.X1.X2.vin1 a_25712_21264# X1.X2.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X511 a_31476_30882# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X512 a_48616_29936# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X513 X2.X1.X2.X1.X1.X1.X3.vin1 a_39966_4110# X2.X1.X2.X1.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X514 X1.X1.X1.X2.X1.X1.vout a_5082_14688# X1.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X515 X1.X1.X1.X1.X2.X2.X1.vin2 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X516 X2.X2.X1.X1.X2.X1.X3.vin2 a_46116_23258# X2.X2.X1.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X517 X2.X2.X1.X1.X3.vin1 a_49002_26164# X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X518 X2.X1.X1.X2.X2.X1.X2.vin1 a_31862_8010# X2.X1.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X519 X2.X2.X1.X2.X2.X2.vout a_48316_5198# X2.X2.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X520 X2.X1.X1.X2.X3.vin1 a_33976_14688# X2.X1.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X521 vss a_54992_6016# a_54606_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X522 X1.X2.X1.X2.X1.X1.X2.vin1 a_17222_15634# X1.X2.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X523 X1.X1.X2.X1.X2.X2.vout a_8486_16452# X1.X1.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X524 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X525 a_2196_27070# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X526 X1.X2.X1.X2.X1.X1.vout a_19036_16634# X1.X2.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X527 vdd d3 a_8572_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X528 X1.X1.X1.X1.X1.X1.vout a_4396_31882# X1.X1.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X529 X1.X1.X1.X2.X2.X2.vout a_5082_7064# X1.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X530 X2.X2.X2.X1.X1.X2.vout a_52406_8828# X2.X2.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X531 vss d4 a_23212_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X532 a_33676_20446# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X533 a_31862_6104# a_31476_6104# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X534 X1.X1.X1.X2.X2.X2.X3.vin2 a_2196_4198# X1.X1.X1.X2.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X535 vdd d1 a_8872_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X536 X1.X1.X2.X2.X1.X1.X1.vin2 a_11072_19358# X1.X1.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X537 vdd a_52792_31700# a_52406_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X538 a_48316_12822# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X539 X1.X1.X3.vin1 a_4696_18540# X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X540 X1.X2.X1.X1.X1.X2.X1.vin2 a_17222_28976# X1.X2.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X541 vdd a_23512_5016# a_23126_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X542 X2.X1.X1.X2.X2.X1.X3.vin2 a_31476_8010# X2.X1.X1.X2.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X543 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X544 vss d1 a_23512_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X545 a_4396_16634# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X546 X1.X1.X1.X1.X1.X2.X2.vin1 a_2582_27070# X1.X1.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X547 a_46116_4198# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X548 X1.X1.X2.X2.X1.X2.vout a_8486_24076# X1.X1.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X549 a_46502_23258# a_46116_23258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X550 vss a_25712_9828# a_25326_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X551 X1.X1.X1.X3.vin2 a_4696_10916# X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X552 a_49002_29936# a_48616_29936# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X553 a_34926_892# d5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X554 X1.X2.X1.X2.vrefh X1.X2.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X555 X2.X2.X2.X3.vin1 a_52106_10734# X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X556 X1.X1.X2.X2.X2.X1.X3.vin2 a_10686_28888# X1.X1.X2.X2.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X557 vss a_54992_32700# a_54606_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X558 X2.X2.X2.X1.X2.X1.vout a_52406_12640# X2.X2.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X559 a_31476_13728# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X560 X2.X2.X1.X2.X3.vin1 a_48616_14688# X2.X2.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X561 X2.X2.X2.X2.X1.X2.vrefh a_54992_21264# X2.X2.X2.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X562 X1.X2.X2.X1.X2.X2.vout a_23126_16452# X1.X2.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X563 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X564 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X565 X2.X1.X2.X3.vin1 a_37852_18358# X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X566 a_34362_7064# a_33976_7064# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X567 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X568 X1.X2.X2.X2.X2.X2.X2.vin1 a_25712_32700# X1.X2.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X569 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X570 X1.X2.X2.X2.X2.X2.X1.vin2 a_25712_30794# X1.X2.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X571 X2.X1.X1.X1.X2.X2.X3.vin2 a_31476_19446# X2.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X572 vss a_40352_23170# a_39966_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X573 X1.X2.X3.vin1 a_19336_18540# X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X574 X2.X2.X1.X1.X1.X1.vout a_49002_29936# X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X575 X2.X1.X1.X1.X1.X1.vout a_33676_31882# X2.X1.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X576 vss d0 a_11072_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X577 a_34062_5198# a_33676_5198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X578 X3.vin1 a_13696_892# X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X579 a_19422_9010# a_19036_9010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X580 X2.X2.X2.X2.X1.X1.vout a_52406_20264# X2.X2.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X581 X2.X1.X2.X2.X2.X1.X1.vin1 a_40352_26982# X2.X1.X2.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X582 X1.X1.X2.X1.X1.X1.X3.vin2 a_10686_6016# X1.X1.X2.X1.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X583 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X584 X1.X1.X1.X1.X1.X2.vout a_4396_28070# X1.X1.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X585 X2.X1.X2.X2.X2.vrefh a_40352_25076# X2.X1.X2.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X586 X1.X2.X2.X2.X1.X2.vout a_23126_24076# X1.X2.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X587 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X588 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X1.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X589 a_33676_16634# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X590 vdd a_11072_28888# a_10686_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X591 X2.X1.X2.X2.X1.X1.X3.vin2 a_39966_21264# X2.X1.X2.X2.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X592 X1.X2.X1.X3.vin2 a_19336_10916# X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X593 X2.X2.X1.X2.X1.X2.X3.vin2 a_48702_12822# X2.X2.X1.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X594 vdd a_8872_8828# a_8486_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X595 vss d0 a_40352_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X596 vdd a_40352_9828# a_39966_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X597 X2.X1.X2.X1.X1.X1.X3.vin2 a_39966_6016# X2.X1.X2.X1.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X598 X1.X1.X1.X1.X2.X2.X3.vin1 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X599 vdd a_52792_8828# a_52406_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X600 X2.X2.X1.X2.X2.X2.X3.vin1 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X601 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X602 X1.X2.X2.X1.X1.X1.X3.vin1 a_25326_4110# X1.X2.X2.X1.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X603 a_31476_11822# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X604 vdd a_54992_17452# a_54606_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X605 vdd a_8572_10734# a_8186_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X606 X2.X1.X1.X2.vrefh a_31862_19446# X2.X1.X1.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X607 a_16836_8010# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X608 X1.X1.X2.X2.X1.X1.X3.vin1 a_10686_19358# X1.X1.X2.X2.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X609 X2.X2.X2.X2.X1.X2.X3.vin1 a_54606_23170# X2.X2.X2.X2.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X610 X1.X2.X2.X2.X2.X1.X3.vin1 a_25326_26982# X1.X2.X2.X2.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X611 X2.X1.X1.X2.X2.X2.vout a_33676_5198# X2.X1.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X612 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X613 X2.X1.X2.X2.X2.X2.X3.vin2 a_38152_31700# X2.X1.X2.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X614 X1.X2.X2.X2.X1.X2.X3.vin2 a_25326_25076# X1.X2.X2.X2.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X615 X1.X2.X2.X1.X2.X2.X1.vin1 a_25712_15546# X1.X2.X2.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X616 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X617 a_31476_25164# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X618 vss d3 a_52492_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X619 vdd d0 a_40352_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X620 vss d1 a_52792_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X621 X1.X1.X1.X2.X1.X2.vrefh a_2582_15634# X1.X1.X1.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X622 vss d1 a_23512_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X623 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X624 vss d1 a_8872_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X625 X1.X1.X1.X1.X1.X2.X3.vin2 a_2196_27070# X1.X1.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X626 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X627 X2.X2.X3.vin1 a_49952_892# X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X628 a_19422_28070# a_19036_28070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X629 X1.X1.X2.X1.X1.X2.vout a_8572_6962# X1.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X630 X2.X2.X2.X1.X1.X1.X1.vin2 a_54992_4110# X2.X2.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X631 a_49002_26164# a_48616_26164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X632 X2.X1.X2.X1.X3.vin1 a_37466_6962# X2.X1.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X633 X1.X3.vin1 a_5646_892# X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X634 a_17222_30882# a_16836_30882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X635 X2.X1.X2.X1.X2.vrefh a_40352_9828# X2.X1.X2.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X636 X1.X1.X2.X1.X1.X2.X2.vin1 a_11072_9828# X1.X1.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X637 X2.X2.X2.X2.X3.vin2 a_52106_29834# X2.X2.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X638 X2.X2.X2.X1.X1.X2.vout a_52492_6962# X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X639 X1.X1.X2.X1.X2.X2.vrefh a_11072_13640# X1.X1.X2.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X640 a_2582_30882# a_2196_30882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X641 X2.X3.vin2 a_49566_892# X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X642 X2.X1.X1.X1.X2.X1.X1.vin1 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X643 a_2196_8010# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X644 a_46502_6104# a_46116_6104# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X645 vss d1 a_8872_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X646 X1.X2.X1.X1.X2.X2.X3.vin2 a_16836_19446# X1.X2.X1.X1.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X647 X2.X2.X2.X2.X2.X2.vout a_52406_31700# X2.X2.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X648 vdd a_38152_5016# a_37766_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X649 X1.X2.X1.X2.X1.X1.X3.vin1 a_19422_16634# X1.X2.X1.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X650 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X651 vss d1 a_52792_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X652 vdd d1 a_52792_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X653 vss a_37852_10734# a_37466_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X654 a_19422_20446# a_19036_20446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X655 vdd d1 a_23512_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X656 a_4782_9010# a_4396_9010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X657 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X658 vss a_38152_12640# a_37766_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X659 X2.X1.X1.X1.X2.X1.X3.vin2 a_31476_23258# X2.X1.X1.X1.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X660 a_2196_19446# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X661 X1.X1.X2.X2.X1.X1.X2.vin1 a_11072_21264# X1.X1.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X662 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X663 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X664 X1.X2.X2.X1.X1.X2.X3.vin2 a_25326_9828# X1.X2.X2.X1.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X665 X2.X1.X2.X1.X2.X2.X3.vin1 a_38152_16452# X2.X1.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X666 vss d1 a_38152_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X667 vss a_54992_26982# a_54606_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X668 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X669 X1.X1.X1.X2.X1.X2.X1.vin1 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X670 X1.X2.X1.X1.X2.X1.X3.vin1 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X671 X2.X2.X2.X1.X2.X2.X1.vin2 a_54992_15546# X2.X2.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X672 X1.X2.X1.X2.X2.X1.X2.vin1 a_17222_8010# X1.X2.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X673 X2.X1.X1.X2.X1.X2.vout a_33676_12822# X2.X1.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X674 X2.X2.X2.X2.X2.X2.X3.vin2 a_52792_31700# X2.X2.X2.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X675 X2.X2.X2.X2.X2.X2.X3.vin2 a_54606_32700# X2.X2.X2.X2.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X676 a_48616_14688# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X677 vdd d0 a_54992_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X678 vdd d0 a_25712_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X679 vdd a_38152_20264# a_37766_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X680 a_46116_21352# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X681 vss d0 a_25712_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X682 vdd a_25712_4110# a_25326_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X683 X2.X1.X2.X1.X1.X2.vout a_37766_8828# X2.X1.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X684 X2.X2.X1.X2.X1.X2.vout a_48316_12822# X2.X2.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X685 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X686 a_17222_13728# a_16836_13728# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X687 vss a_40352_17452# a_39966_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X688 vdd a_25712_11734# a_25326_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X689 a_34062_28070# a_33676_28070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X690 a_2196_25164# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X691 a_31862_30882# a_31476_30882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X692 a_49002_29936# a_48616_29936# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X693 a_48702_5198# a_48316_5198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X694 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X695 a_19036_5198# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X696 X1.X2.X2.X1.X1.X1.X3.vin2 a_25326_6016# X1.X2.X2.X1.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X697 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X698 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X699 X1.X1.X2.X1.X2.X2.X3.vin2 a_8872_16452# X1.X1.X2.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X700 vdd d2 a_52492_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X701 X2.X1.X1.X2.X2.X2.X3.vin1 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X702 a_2582_27070# a_2196_27070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X703 X2.X1.X2.X1.X2.X2.X3.vin1 a_39966_15546# X2.X1.X2.X1.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X704 X1.X1.X1.X1.X1.X1.X3.vin1 a_4782_31882# X1.X1.X1.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X705 X2.X1.X2.X2.X2.X2.vout a_37766_31700# X2.X1.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X706 a_34362_29936# a_33976_29936# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X707 vss a_52492_10734# a_52106_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X708 a_34062_20446# a_33676_20446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X709 a_46116_27070# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X710 X1.X1.X1.X1.X1.X1.X1.vin2 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X711 vdd d1 a_52792_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X712 vdd a_40352_25076# a_39966_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X713 a_48702_12822# a_48316_12822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X714 X1.X1.X1.X2.X1.X1.X3.vin2 a_2196_15634# X1.X1.X1.X2.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X715 X1.X1.X1.X3.vin2 a_5082_18540# X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X716 a_19422_16634# a_19036_16634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X717 vss a_23512_16452# a_23126_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X718 X1.X1.X2.X2.X2.X1.vout a_8486_27888# X1.X1.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X719 X2.X2.X1.X2.X2.X2.X1.vin2 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X720 vss a_11072_7922# a_10686_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X721 a_4782_16634# a_4396_16634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X722 a_19036_28070# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X723 a_34926_892# d5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X724 X1.X1.X2.X2.X2.X2.X2.vin1 a_11072_32700# X1.X1.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X725 a_16836_30882# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X726 a_49002_7064# a_48616_7064# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X727 X2.X2.X2.X1.X2.X2.X3.vin1 a_52792_16452# X2.X2.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X728 X1.X1.X2.X2.X2.X2.X1.vin2 a_11072_30794# X1.X1.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X729 X2.X2.X2.X1.X2.X2.X3.vin2 a_54606_17452# X2.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X730 X1.X1.X2.X2.X1.X2.X3.vin1 a_8872_24076# X1.X1.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X731 X1.X1.X2.X1.X2.X1.X3.vin2 a_10686_13640# X1.X1.X2.X1.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X732 X1.X1.X1.X1.X2.X2.vout a_4396_20446# X1.X1.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X733 X2.X1.X2.X1.X1.X1.X1.vin2 a_40352_4110# X2.X1.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X734 vss d0 a_25712_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X735 vdd a_37852_29834# a_37466_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X736 a_17222_11822# a_16836_11822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X737 X1.X1.X1.X2.X3.vin2 a_5082_10916# X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X738 vdd d0 a_40352_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X739 a_19336_29936# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X740 vdd a_23512_24076# a_23126_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X741 a_31476_9916# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X742 a_19036_20446# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X743 vss d0 a_54992_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X744 vdd a_38152_31700# a_37766_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X745 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X746 X2.X2.X1.X2.X1.X1.vout a_49002_14688# X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X747 a_31862_13728# a_31476_13728# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X748 X1.X2.X2.X1.X2.X2.X3.vin2 a_23512_16452# X1.X2.X2.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X749 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X750 a_17222_25164# a_16836_25164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X751 X2.X1.X1.X2.X2.X2.X2.vin1 a_31862_4198# X2.X1.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X752 X2.X2.X1.X1.X2.X2.X1.vin2 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X753 a_4696_14688# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X754 X1.X1.X2.X2.X1.X1.X3.vin2 a_10686_21264# X1.X1.X2.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X755 X2.X1.X1.X1.X2.X2.X2.vin1 a_31862_19446# X2.X1.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X756 vdd a_8872_27888# a_8486_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X757 X1.X2.X1.X2.X2.X2.X3.vin2 a_19422_5198# X1.X2.X1.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X758 X2.X1.X2.X1.X2.X2.vout a_37766_16452# X2.X1.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X759 X2.X2.X2.X2.X3.vin2 a_52106_29834# X2.X2.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X760 X2.X1.X1.X1.X1.X1.X3.vin2 a_34062_31882# X2.X1.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X761 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X762 X1.X1.X1.X2.X1.X2.X3.vin1 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X763 X1.X2.X2.X2.X2.X1.vout a_23126_27888# X1.X2.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X764 vss a_52792_24076# a_52406_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X765 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X766 vss a_11072_11734# a_10686_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X767 X2.X2.X3.vin1 a_48616_18540# X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X768 X2.X2.X2.X1.X1.X1.X2.vin1 a_54992_6016# X2.X2.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X769 X1.X1.X1.X1.X1.X2.X3.vin2 a_4782_28070# X1.X1.X1.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X770 X1.X2.X2.X2.X1.X2.X3.vin1 a_23512_24076# X1.X2.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X771 X2.X2.X1.X2.X2.X2.X3.vin2 a_48702_5198# X2.X2.X1.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X772 X2.X1.X2.X1.X2.X1.X1.vin1 a_40352_11734# X2.X1.X2.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X773 a_34062_16634# a_33676_16634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X774 X2.X2.X1.X1.X1.X2.X2.vin1 a_46502_27070# X2.X2.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X775 a_16836_13728# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X776 X1.X1.X2.X1.X2.X2.X1.vin1 a_11072_15546# X1.X1.X2.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X777 vdd d0 a_11072_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X778 vss a_25712_6016# a_25326_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X779 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X780 X2.X2.X2.X2.X3.vin1 a_52106_22210# X2.X2.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X781 a_35312_892# a_34926_892# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X782 a_16836_6104# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X783 X1.X2.X2.X1.X1.X2.vout a_23126_8828# X1.X2.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X784 X1.X2.X1.X1.X2.X2.X3.vin2 a_16836_19446# X1.X2.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X785 X2.X2.X1.X3.vin2 a_48616_10916# X2.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X786 X2.X1.X1.X2.X3.vin2 a_33976_7064# X2.X1.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X787 X1.X2.X1.X2.X2.X2.vout a_19722_7064# X1.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X788 X1.X2.X1.X1.X1.X2.vrefh a_17222_30882# X1.X2.X1.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X789 X2.X2.X2.X2.X2.X1.X3.vin1 a_54606_26982# X2.X2.X2.X2.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X790 a_31476_23258# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X791 a_34362_26164# a_33976_26164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X792 X1.X2.X1.X1.X1.X1.vout a_19036_31882# X1.X2.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X793 vdd a_52492_29834# a_52106_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X794 a_31862_11822# a_31476_11822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X795 vdd d0 a_54992_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X796 a_46116_15634# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X797 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X798 vss d0 a_40352_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X799 X2.X3.vin1 a_34926_892# X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X800 a_33976_29936# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X801 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X802 X1.X2.X2.X2.X2.X1.X1.vin1 a_25712_26982# X1.X2.X2.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X803 a_2196_19446# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X804 X1.X1.X1.X1.X1.X1.X3.vin1 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X805 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X806 X1.X2.X2.X2.X2.vrefh a_25712_25076# X1.X2.X2.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X807 X2.X2.X1.X2.X2.X2.vout a_49002_7064# X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X808 X1.X2.X1.X2.X2.X1.vout a_19036_9010# X1.X2.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X809 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X810 X2.X2.X1.X2.X2.X2.X3.vin2 a_46116_4198# X2.X2.X1.X2.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X811 X1.X1.X2.X1.X1.X2.X3.vin2 a_8872_8828# X1.X1.X2.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X812 a_31862_25164# a_31476_25164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X813 X1.X2.X2.X1.X2.X1.X3.vin1 a_25326_11734# X1.X2.X2.X1.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X814 a_19036_16634# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X815 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X816 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X817 a_4396_31882# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X818 X2.X2.X2.X1.X3.vin2 a_52106_14586# X2.X2.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X819 X2.X2.X2.X1.X1.X2.X3.vin2 a_52792_8828# X2.X2.X2.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X820 vdd d0 a_11072_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X821 X1.X1.X2.X2.X2.X2.X3.vin2 a_10686_32700# X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X822 X1.X1.X2.X2.X2.X2.X3.vin1 a_10686_30794# X1.X1.X2.X2.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X823 vss d2 a_8572_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X824 vss d2 a_52492_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X825 a_19336_26164# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X826 a_16836_11822# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X827 vdd a_40352_19358# a_39966_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X828 vss d1 a_23512_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X829 X1.X1.X1.X2.X2.X1.vout a_4396_9010# X1.X1.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X830 X2.X1.X1.X1.X2.X2.X3.vin1 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X831 X1.X2.X2.X1.X1.X1.X3.vin2 a_23512_5016# X1.X2.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X832 a_42976_892# d6 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X833 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X834 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X835 vss d3 a_37852_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X836 a_16836_25164# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X837 X2.X2.X2.X1.X2.X2.vout a_52492_14586# X2.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X838 X2.X2.X1.X1.X2.X2.X3.vin1 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X839 vdd d2 a_23212_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X840 vss d1 a_38152_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X841 X1.X2.X1.X2.X1.X2.X1.vin2 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X842 X2.X1.X1.X1.X2.X2.vrefh a_31862_23258# X2.X1.X1.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X843 a_46116_13728# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X844 a_2582_19446# a_2196_19446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X845 vdd d2 a_52492_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X846 a_34362_29936# a_33976_29936# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X847 vdd a_11072_30794# a_10686_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X848 X1.X2.X2.X1.X2.vrefh a_25712_9828# X1.X2.X2.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X849 vss a_8572_6962# a_8186_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X850 vss a_37852_29834# a_37466_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X851 vss d0 a_54992_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X852 a_46116_9916# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X853 vss d0 a_40352_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X854 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X855 X2.X1.X1.X1.X2.X1.vout a_33676_24258# X2.X1.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X856 vdd a_11072_9828# a_10686_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X857 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X858 vss a_52492_6962# a_52106_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X859 X2.X1.X1.X2.X1.X2.X3.vin1 a_34062_12822# X2.X1.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X860 X1.X2.X1.X2.X1.X2.vout a_19722_14688# X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X861 X2.X2.X1.X2.X1.X2.vrefh a_46502_15634# X2.X2.X1.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X862 a_6032_892# a_5646_892# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X863 a_49002_14688# a_48616_14688# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X864 X1.X1.X2.X1.X2.X2.X3.vin1 a_10686_15546# X1.X1.X2.X1.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X865 X2.X2.X1.X1.X1.X2.X3.vin2 a_46116_27070# X2.X2.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X866 vdd d1 a_38152_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X867 a_46502_21352# a_46116_21352# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X868 X2.X1.X2.X1.X1.X1.X2.vin1 a_40352_6016# X2.X1.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X869 X2.X1.X2.X1.X3.vin2 a_37466_14586# X2.X1.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X870 vdd a_25712_23170# a_25326_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X871 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X872 vdd d0 a_25712_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X873 X2.X2.X2.X2.X2.X1.X2.vin1 a_54992_28888# X2.X2.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X874 a_2196_4198# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X875 a_2582_25164# a_2196_25164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X876 vdd d2 a_52492_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X877 X1.X2.X1.X1.X2.X1.X3.vin2 a_16836_23258# X1.X2.X1.X1.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X878 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X879 vdd a_37852_22210# a_37466_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X880 a_48316_31882# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X881 vss d3 a_8572_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X882 a_33976_26164# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X883 a_19336_29936# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X884 X2.X2.X2.X2.X1.X2.vout a_52406_24076# X2.X2.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X885 a_46116_32788# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X886 X1.X1.X2.X3.vin1 a_8186_10734# X1.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X887 a_48616_18540# d4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X888 vss a_40352_28888# a_39966_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X889 X1.X2.X1.X2.X3.vin2 a_19336_7064# X1.X2.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X890 X1.X1.X2.X1.X2.X1.vout a_8486_12640# X1.X1.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X891 X2.X1.X1.X1.X1.X1.X3.vin1 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X892 X1.X2.X1.X2.X1.X2.X2.vin1 a_17222_11822# X1.X2.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X893 a_2196_23258# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X894 X1.X2.X1.X2.X1.X2.vout a_19036_12822# X1.X2.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X895 X2.X1.X1.X2.X1.X1.X3.vin1 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X896 a_46502_27070# a_46116_27070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X897 a_17222_6104# a_16836_6104# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X898 X1.X1.X2.X2.X2.X1.X3.vin2 a_8872_27888# X1.X1.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X899 X1.X2.X1.X1.X2.X1.X1.vin2 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X900 X2.X1.X1.X2.X2.X2.vout a_34362_7064# X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X901 X2.X1.X2.X2.X2.X1.X3.vin2 a_39966_28888# X2.X1.X2.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X902 X2.X2.X2.X2.X3.vin1 a_52492_25982# X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X903 X2.X1.X1.X2.X2.X2.X3.vin2 a_31476_4198# X2.X1.X1.X2.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X904 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X905 vdd d0 a_54992_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X906 vss d0 a_11072_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X907 a_48616_10916# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X908 vdd a_37852_14586# a_37466_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X909 X1.X2.X1.X2.X2.X2.X2.vin1 a_17222_4198# X1.X2.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X910 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X1.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X911 a_4396_12822# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X912 vss d1 a_23512_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X913 X2.X2.X1.X2.X1.X2.X1.vin1 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X914 vss a_8572_22210# a_8186_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X915 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X916 X2.X1.X1.X2.X2.X1.X3.vin1 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X917 X1.X1.X1.X1.X2.X2.X3.vin2 a_4782_20446# X1.X1.X1.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X918 vss a_52492_29834# a_52106_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X919 X1.X1.X2.X2.X1.X1.vout a_8486_20264# X1.X1.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X920 a_33676_9010# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X921 vss a_23512_27888# a_23126_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X922 a_17222_23258# a_16836_23258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X923 X1.X2.X1.X1.X1.X1.X3.vin2 a_19422_31882# X1.X2.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X924 vdd d2 a_37852_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X925 a_19722_29936# a_19336_29936# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X926 vdd d1 a_38152_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X927 vss a_25712_32700# a_25326_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X928 X1.X2.X2.X1.X2.X1.vout a_23126_12640# X1.X2.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X929 a_5082_14688# a_4696_14688# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X930 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X931 vdd a_52492_22210# a_52106_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X932 X2.X1.X2.X3.vin2 a_37466_25982# X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X933 vdd d1 a_8872_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X934 a_33976_29936# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X935 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X936 X2.X1.X1.X2.X1.X1.X3.vin2 a_31476_15634# X2.X1.X1.X2.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X937 X2.X1.X1.X3.vin1 a_34362_18540# X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X938 a_48316_28070# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X939 X2.X2.X1.X1.X1.X1.X3.vin1 a_48702_31882# X2.X2.X1.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X940 vss a_40352_19358# a_39966_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X941 X1.X2.X2.X2.X2.X1.X3.vin2 a_23512_27888# X1.X2.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X942 vss d1 a_52792_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X943 vss a_11072_23170# a_10686_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X944 X2.X2.X1.X1.X1.X1.X1.vin2 a_46502_32788# X2.X2.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X945 vss d0 a_11072_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X946 X2.X2.X1.X2.X1.X1.X3.vin2 a_46116_15634# X2.X2.X1.X2.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X947 X2.X2.X1.X3.vin2 a_49002_18540# X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X948 a_19422_5198# a_19036_5198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X949 X2.X1.X1.X1.X1.X2.X3.vin1 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X950 vdd d2 a_37852_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X951 vss a_40352_4110# a_39966_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X952 X2.X1.X2.X2.X1.X2.X1.vin1 a_40352_23170# X2.X1.X2.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X953 X1.X1.X2.X2.X2.X1.X1.vin1 a_11072_26982# X1.X1.X2.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X954 X1.X1.X1.X1.X2.X1.vout a_4396_24258# X1.X1.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X955 X1.X2.X2.X2.X1.X1.vout a_23126_20264# X1.X2.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X956 X1.X1.X1.X2.X2.X1.X2.vin1 a_2582_8010# X1.X1.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X957 X1.X1.X2.X2.X2.vrefh a_11072_25076# X1.X1.X2.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X958 X2.X1.X1.X2.X3.vin1 a_34362_10916# X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X959 a_33676_12822# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X960 X1.X1.X1.X3.vin1 a_4696_26164# X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X961 vdd a_52492_14586# a_52106_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X962 X1.X1.X2.X2.X3.vin2 a_8186_29834# X1.X1.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X963 a_28482_892# a_28096_892# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X964 vss d0 a_40352_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X965 vss a_8572_25982# a_8186_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X966 a_2582_6104# a_2196_6104# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X967 X2.X2.X1.X2.X3.vin2 a_49002_10916# X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X968 X1.X1.X2.X2.X2.X2.vout a_8486_31700# X1.X1.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X969 a_31862_23258# a_31476_23258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X970 vss a_38152_24076# a_37766_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X971 a_46502_15634# a_46116_15634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X972 vdd a_54992_13640# a_54606_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X973 X2.X1.X1.X1.X2.X2.vout a_34362_22312# X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X974 vdd a_25712_17452# a_25326_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X975 a_19722_7064# a_19336_7064# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X976 a_2582_19446# a_2196_19446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X977 a_16836_4198# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X978 X2.X2.X3.vin2 a_52106_18358# X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X979 X1.X2.X2.X2.X1.X2.X3.vin1 a_25326_23170# X1.X2.X2.X2.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X980 X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X981 X1.X2.X2.X1.X2.X1.X1.vin1 a_25712_11734# X1.X2.X2.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X982 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X983 X1.X1.X2.X1.X1.X1.X1.vin2 a_11072_4110# X1.X1.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X984 a_4782_31882# a_4396_31882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X985 vdd d0 a_40352_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X986 X1.X1.X1.X2.X2.vrefh a_2582_11822# X1.X1.X1.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X987 X2.X2.X1.X2.X1.X2.X3.vin1 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X988 vss d1 a_23512_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X989 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X990 vdd d1 a_38152_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X991 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X992 vdd d0 a_40352_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X993 X1.X2.X1.X3.vin1 a_19336_26164# X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X994 a_19722_26164# a_19336_26164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X995 a_16836_23258# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X996 X2.X2.X1.X1.X1.X2.X3.vin2 a_48702_28070# X2.X2.X1.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X997 X1.X1.X2.X1.X2.vrefh a_11072_9828# X1.X1.X2.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X998 X2.X1.X1.X1.X2.X2.X1.vin1 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X999 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1000 X2.X1.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1001 a_14082_892# a_13696_892# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1002 X1.X2.X1.X2.X1.X2.X3.vin1 a_19422_12822# X1.X2.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1003 X1.X1.X1.X1.X3.vin2 a_4696_22312# X1.X1.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1004 X2.X2.X2.X1.X1.X1.vout a_52406_5016# X2.X2.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1005 X2.X2.vrefh a_40352_32700# X2.X1.X2.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1006 X2.X1.X2.X1.X1.X1.X1.vin1 X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1007 X1.X2.X2.X2.X2.X2.vout a_23126_31700# X1.X2.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1008 a_34362_14688# a_33976_14688# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1009 a_4782_5198# a_4396_5198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1010 X1.X1.X1.X2.X1.X1.X1.vin1 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1011 vdd d1 a_23512_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1012 a_46502_13728# a_46116_13728# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1013 a_48316_9010# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1014 vss d4 a_8572_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1015 X2.X1.X3.vin1 a_33976_18540# X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1016 X2.X2.X1.X1.X1.X1.vout a_48316_31882# X2.X2.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1017 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1018 vdd d0 a_11072_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1019 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1020 X2.X2.X1.X1.X1.X1.X3.vin1 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1021 X2.X1.X2.X1.X2.X1.X3.vin1 a_38152_12640# X2.X1.X2.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1022 vss d2 a_37852_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1023 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1024 X1.X2.X2.X1.X3.vin1 a_22826_6962# X1.X2.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1025 X2.X1.X1.X1.X2.X1.X3.vin1 a_34062_24258# X2.X1.X1.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1026 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1027 X2.X2.X2.X1.X2.X1.X1.vin2 a_54992_11734# X2.X2.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1028 X1.X2.X1.X1.X2.X2.X3.vin1 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1029 vss a_25712_26982# a_25326_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1030 X2.X3.vin2 a_43362_892# X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1031 a_31862_8010# a_31476_8010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1032 X1.X1.X2.X2.X2.X1.X3.vin1 a_10686_26982# X1.X1.X2.X2.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1033 X1.X1.X2.X2.X1.X2.X3.vin2 a_10686_25076# X1.X1.X2.X2.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1034 X1.X2.X2.X2.X2.X2.X3.vin2 a_25326_32700# X1.X2.X2.X2.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1035 X2.X1.X1.X3.vin2 a_33976_10916# X2.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1036 a_19336_14688# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1037 X2.X1.X2.X1.X2.X2.vout a_37852_14586# X2.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1038 vdd d4 a_52492_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1039 vdd d0 a_25712_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1040 vdd d0 a_40352_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1041 a_5082_7064# a_4696_7064# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1042 vss d0 a_40352_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1043 vss a_40352_13640# a_39966_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1044 X1.X1.X1.X2.X2.X2.vout a_4396_5198# X1.X1.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1045 X2.X1.X1.X2.X2.X1.X1.vin1 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1046 vss a_11072_17452# a_10686_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1047 a_2196_21352# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1048 vdd d2 a_37852_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1049 a_48702_31882# a_48316_31882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1050 a_43362_892# a_42976_892# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1051 X1.X2.X1.X1.X3.vin2 a_19336_22312# X1.X2.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1052 a_31476_8010# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1053 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1054 a_19722_29936# a_19336_29936# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1055 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1056 a_46502_32788# a_46116_32788# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1057 a_49952_892# a_49566_892# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1058 X1.X1.X2.X1.X3.vin2 a_8572_10734# X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1059 X2.X1.X2.X1.X2.X2.X2.vin1 a_40352_17452# X2.X1.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1060 a_49002_18540# a_48616_18540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1061 X2.X1.X1.X1.X3.vin2 a_33976_22312# X2.X1.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1062 X1.X2.X1.X1.X2.X1.X2.vin1 a_17222_23258# X1.X2.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1063 X2.X1.X1.X1.X1.X1.X1.vin1 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1064 X1.X2.X1.X1.X2.X1.vout a_19036_24258# X1.X2.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1065 X1.X1.X2.X1.X2.X1.X3.vin2 a_8872_12640# X1.X1.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1066 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1067 a_2582_23258# a_2196_23258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1068 X2.X1.X2.X1.X2.X1.X3.vin1 a_39966_11734# X2.X1.X2.X1.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1069 X2.X1.X1.X2.X1.X1.X1.vin2 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1070 X1.X1.X2.X1.X3.vin1 a_8186_6962# X1.X1.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1071 vss a_54992_21264# a_54606_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1072 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1073 a_48316_20446# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1074 vdd a_40352_21264# a_39966_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1075 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1076 vss a_23212_10734# a_22826_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1077 X1.X1.X1.X2.X1.X2.X3.vin2 a_2196_11822# X1.X1.X1.X2.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1078 vdd d1 a_23512_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1079 X1.X1.X1.X1.X1.X2.X1.vin1 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1080 vdd a_11072_25076# a_10686_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1081 vdd a_37852_18358# a_37466_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1082 X1.X2.X2.X1.X1.X2.X1.vin1 a_25712_7922# X1.X2.X2.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1083 X2.X3.vin1 a_34926_892# X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1084 X1.X1.X2.X2.X3.vin2 a_8186_29834# X1.X1.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1085 vss a_23512_12640# a_23126_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1086 a_19422_12822# a_19036_12822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1087 a_49002_10916# a_48616_10916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1088 vdd d2 a_37852_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1089 a_4396_24258# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1090 vdd a_8872_5016# a_8486_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1091 vdd a_40352_6016# a_39966_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1092 a_4782_12822# a_4396_12822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1093 X2.X2.X2.X1.X3.vin1 a_52492_10734# X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1094 vdd a_52792_5016# a_52406_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1095 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1096 X2.X2.X2.X1.X2.X1.X3.vin1 a_52792_12640# X2.X2.X2.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1097 X2.X2.X1.X1.X1.X2.vout a_48316_28070# X2.X2.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1098 X2.X1.X1.X2.X2.X1.X1.vin2 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1099 X1.X1.X2.X1.X1.X2.X3.vin2 a_10686_9828# X1.X1.X2.X1.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1100 X2.X2.X2.X1.X2.X1.X3.vin2 a_54606_13640# X2.X2.X2.X1.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1101 X1.X1.X2.X2.X1.X1.X3.vin1 a_8872_20264# X1.X1.X2.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1102 X1.X2.X2.X1.X2.X2.X3.vin2 a_25326_17452# X1.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1103 X1.X2.X1.X1.X1.X1.X3.vin1 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1104 X2.X2.X2.X1.X1.X2.X3.vin1 a_54606_7922# X2.X2.X2.X1.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1105 vdd d0 a_40352_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1106 X1.X2.X1.X2.X1.X1.X3.vin1 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1107 X1.X1.X2.X2.X3.vin1 a_8186_22210# X1.X1.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1108 a_33976_14688# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1109 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1110 X1.X2.X2.X1.X3.vin2 a_23212_10734# X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1111 X1.X1.X1.X2.X1.X1.X3.vin1 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1112 vdd a_23512_20264# a_23126_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1113 a_31476_21352# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1114 X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1115 vss d0 a_25712_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1116 X1.X2.X2.X1.X2.X1.X3.vin2 a_23512_12640# X1.X2.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1117 vss a_23212_6962# a_22826_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1118 X2.X1.X2.X2.X3.vin1 a_37852_25982# X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1119 X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1120 vss a_8572_18358# a_8186_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1121 a_2196_32788# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1122 X1.X2.X1.X2.X2.X2.X3.vin1 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1123 X2.X1.X2.X3.vin1 a_37466_10734# X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1124 X2.X1.X1.X2.X1.X1.X2.vin1 a_31862_15634# X2.X1.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1125 a_2196_17540# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1126 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1127 a_48702_28070# a_48316_28070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1128 X1.X2.X1.X2.X2.X1.X3.vin1 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1129 X2.X1.X2.X1.X2.X1.vout a_37766_12640# X2.X1.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1130 X1.X1.X2.X1.X1.X1.X2.vin1 a_11072_6016# X1.X1.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1131 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1132 X1.X1.X2.X1.X1.X2.vout a_8486_8828# X1.X1.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1133 X2.X2.X2.X2.X2.X2.X1.vin1 a_54992_30794# X2.X2.X2.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1134 X2.X1.X2.X2.X2.X1.X1.vin2 a_40352_26982# X2.X1.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1135 vss d0 a_11072_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1136 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1137 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1138 X1.X1.X2.X1.X3.vin2 a_8186_14586# X1.X1.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1139 X2.X1.X1.X1.X1.X2.X1.vin2 a_31862_28976# X2.X1.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1140 X2.X1.X2.X2.X1.X1.X3.vin2 a_38152_20264# X2.X1.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1141 a_31476_27070# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1142 X1.X1.X1.X1.X2.X1.X3.vin2 a_4782_24258# X1.X1.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1143 X1.X2.X2.X2.X1.X1.X3.vin1 a_23512_20264# X1.X2.X2.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1144 vdd a_52492_18358# a_52106_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1145 vdd a_40352_32700# a_39966_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1146 a_2196_9916# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1147 a_34062_12822# a_33676_12822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1148 vss a_40352_30794# a_39966_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1149 X1.X1.X1.X1.X3.vin2 a_5082_26164# X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1150 a_33676_5198# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1151 X1.X1.X2.X1.X2.X1.X1.vin1 a_11072_11734# X1.X1.X2.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1152 X2.X2.X2.X2.X2.X2.X2.vin1 vrefl vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1153 X2.X2.X1.X1.X2.X2.X3.vin2 a_48702_20446# X2.X2.X1.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1154 X1.X1.X2.X2.X2.X1.vout a_8572_29834# X1.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1155 X2.X2.X1.X2.X2.X1.vout a_48316_9010# X2.X2.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1156 X1.X2.X1.X2.X1.X1.X3.vin2 a_16836_15634# X1.X2.X1.X2.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1157 X1.X1.X2.X2.X2.X2.X3.vin1 a_8872_31700# X1.X1.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1158 a_46502_8010# a_46116_8010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1159 X2.X1.X2.X2.X2.X2.X3.vin1 a_39966_30794# X2.X1.X2.X2.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1160 X1.X2.X2.X2.X2.X1.X3.vin1 a_25326_26982# X1.X2.X2.X2.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1161 vss d1 a_38152_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1162 vdd d0 a_54992_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1163 vdd d0 a_25712_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1164 vdd a_23212_29834# a_22826_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1165 a_5646_892# d5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1166 a_46116_11822# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1167 vdd d0 a_25712_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1168 X1.X2.X1.X1.X1.X2.X3.vin1 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1169 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1170 X1.X2.X2.X2.X1.X2.X1.vin1 a_25712_23170# X1.X2.X2.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1171 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1172 a_2196_15634# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1173 vdd a_23512_31700# a_23126_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1174 X1.X1.X1.X1.X1.X2.X3.vin1 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1175 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1176 X1.X2.X1.X2.X2.X2.vout a_19036_5198# X1.X2.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1177 X1.X1.X2.X1.X1.X1.X3.vin2 a_8872_5016# X1.X1.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1178 a_19036_12822# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1179 X2.X1.X2.X1.X1.X1.vout a_37766_5016# X2.X1.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1180 X1.X2.X2.X1.X1.X1.X1.vin1 X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1181 a_46116_8010# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1182 X2.X2.X2.X1.X1.X1.X3.vin2 a_52792_5016# X2.X2.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1183 X2.X1.X2.X1.X1.X2.X3.vin2 a_38152_8828# X2.X1.X2.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1184 vss a_54992_7922# a_54606_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1185 a_2196_28976# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1186 a_2196_9916# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1187 X1.X3.vin1 a_5646_892# X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1188 vout a_28096_892# X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1189 X1.X1.X1.X2.X2.X2.X3.vin1 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1190 X1.X1.X1.X2.X2.X2.X2.vin1 a_2582_4198# X1.X1.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1191 vss a_54992_15546# a_54606_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1192 a_46116_17540# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1193 vss a_52792_31700# a_52406_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1194 X1.X2.X2.X2.X2.X1.vout a_23212_29834# X1.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1195 vdd a_40352_15546# a_39966_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1196 vdd a_11072_19358# a_10686_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1197 X2.X2.X2.X2.X1.X1.X3.vin2 a_52792_20264# X2.X2.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1198 X2.X2.X1.X3.vin1 a_48616_26164# X2.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1199 X2.X2.X2.X2.X1.X1.X3.vin2 a_54606_21264# X2.X2.X2.X2.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1200 X1.X2.X1.X1.X2.X1.X3.vin1 a_19422_24258# X1.X2.X1.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1201 X1.X1.X1.X1.X2.X1.vout a_5082_22312# X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1202 X1.X2.X2.X3.vin1 a_22826_10734# X1.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1203 X1.X2.X2.X2.X2.X2.X3.vin1 a_23512_31700# X1.X2.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1204 X2.X1.X1.X1.X1.X2.vout a_33676_28070# X2.X1.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1205 X1.X1.X2.X2.X1.X2.vout a_8486_24076# X1.X1.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1206 a_28096_892# d7 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1207 X2.X1.X1.X1.X1.X1.X3.vin2 a_31476_30882# X2.X1.X1.X1.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1208 vss a_11072_4110# a_10686_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1209 X1.X2.X1.X2.X2.X1.X1.vin1 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1210 vss a_8872_16452# a_8486_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1211 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1212 a_31476_15634# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1213 a_34362_18540# a_33976_18540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1214 X2.X2.X2.X2.X1.X2.X1.vin2 a_54992_23170# X2.X2.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1215 vss d0 a_25712_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1216 X2.X1.X1.X1.X2.X2.vout a_33676_20446# X2.X1.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1217 X2.X1.X2.X2.X1.X1.vout a_37766_20264# X2.X1.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1218 vss a_37852_6962# a_37466_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1219 X1.X1.X1.X2.X3.vin2 a_4696_7064# X1.X1.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1220 X2.X2.X1.X2.X2.vrefh a_46502_11822# X2.X2.X1.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1221 a_31476_6104# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1222 X2.X1.X1.X2.X2.X1.X3.vin1 a_34062_9010# X2.X1.X1.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1223 X2.vrefh a_25712_32700# X1.X2.X2.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1224 X1.X1.X2.X1.X2.X1.X3.vin1 a_10686_11734# X1.X1.X2.X1.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1225 a_19722_14688# a_19336_14688# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1226 X2.X2.X1.X2.X2.X1.X2.vin1 a_46502_8010# X2.X2.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1227 X2.X2.X1.X1.X2.X2.vout a_48316_20446# X2.X2.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1228 X1.X1.X1.X2.X1.X1.vout a_4396_16634# X1.X1.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1229 a_17222_21352# a_16836_21352# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1230 X2.X2.X2.X1.X1.X2.X3.vin2 a_54606_9828# X2.X2.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1231 vss d0 a_11072_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1232 a_2582_21352# a_2196_21352# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1233 vdd a_52792_16452# a_52406_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1234 vdd a_8872_24076# a_8486_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1235 a_34362_10916# a_33976_10916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1236 X2.X1.X1.X2.X2.X1.vout a_33676_9010# X2.X1.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1237 X1.X1.X2.X1.X1.X2.X3.vin1 a_10686_7922# X1.X1.X2.X1.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1238 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1239 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1240 X2.X2.X1.X1.X3.vin2 a_48616_22312# X2.X2.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1241 X1.X2.X2.X2.X1.X2.vout a_23126_24076# X1.X2.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1242 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1243 a_46116_28976# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1244 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1245 X2.X1.X2.X2.X1.X2.X3.vin1 a_39966_23170# X2.X1.X2.X2.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1246 a_19336_18540# d4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1247 X2.X2.X1.X2.X1.X1.X1.vin1 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1248 vss a_11072_28888# a_10686_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1249 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1250 a_48316_5198# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1251 a_4696_18540# d4 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1252 X2.X1.X1.X2.X1.X2.X3.vin1 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1253 vss d0 a_54992_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1254 X2.X1.X2.X1.X1.X2.X3.vin1 a_39966_7922# X2.X1.X2.X1.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1255 a_17222_27070# a_16836_27070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1256 vss d3 a_23212_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1257 a_48702_20446# a_48316_20446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1258 vdd d4 a_37852_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1259 vdd d0 a_11072_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1260 X1.X1.X2.X2.X2.X2.vout a_8572_29834# X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1261 a_4782_24258# a_4396_24258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1262 X2.X1.X2.vrefh X2.X1.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1263 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1264 a_31476_13728# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1265 vdd d0 a_54992_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1266 X1.X2.X2.X1.X1.X1.vout a_23126_5016# X1.X2.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1267 X1.X1.X2.X1.X1.X1.X1.vin1 X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1268 a_31862_4198# a_31476_4198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1269 a_19336_10916# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1270 a_4696_10916# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1271 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1272 X1.X2.X2.X2.X3.vin2 a_22826_29834# X1.X2.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1273 X1.X2.X2.X1.X2.X2.X2.vin1 a_25712_17452# X1.X2.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1274 vss a_23212_29834# a_22826_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1275 vdd d0 a_40352_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1276 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1277 vss d0 a_40352_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1278 vss a_23512_8828# a_23126_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1279 X1.X1.X2.X2.X1.X1.vout a_8572_22210# X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1280 X2.X1.X1.X2.X1.X1.vout a_33676_16634# X2.X1.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1281 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1282 a_31862_21352# a_31476_21352# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1283 a_4696_22312# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1284 a_2582_32788# a_2196_32788# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1285 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1286 vdd a_23212_22210# a_22826_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1287 X2.X1.X2.X1.X3.vin1 a_37852_10734# X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1288 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1289 a_33676_31882# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1290 a_2582_17540# a_2196_17540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1291 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1292 X2.X1.X1.X2.X1.X2.X3.vin2 a_31476_11822# X2.X1.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1293 X2.X2.X2.X1.X2.X2.X3.vin1 a_54606_15546# X2.X2.X2.X1.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1294 X2.X2.X2.X2.X2.X2.vout a_52406_31700# X2.X2.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1295 a_48316_24258# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1296 a_31476_32788# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1297 X1.X2.X2.X2.X2.X2.vout a_23212_29834# X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1298 a_33976_18540# d4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1299 a_48616_26164# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1300 X1.X1.X3.vin2 a_8186_18358# X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1301 a_33976_7064# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1302 vss a_11072_19358# a_10686_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1303 X2.X2.X1.X1.X1.X2.X1.vin1 a_46502_28976# X2.X2.X1.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1304 vss d1 a_23512_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1305 X2.X2.X1.X2.X1.X2.X3.vin2 a_46116_11822# X2.X2.X1.X2.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1306 X1.X1.X2.X1.X2.X1.vout a_8572_14586# X1.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1307 vdd a_54992_9828# a_54606_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1308 X2.X1.X1.X1.X2.X1.X3.vin1 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1309 a_31862_27070# a_31476_27070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1310 a_2582_9916# a_2196_9916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1311 a_16836_21352# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1312 X1.X1.X2.X2.X1.X2.X1.vin1 a_11072_23170# X1.X1.X2.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1313 a_19036_9010# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1314 a_33976_10916# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1315 vdd a_23212_14586# a_22826_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1316 X1.X2.X2.X2.X1.X1.vout a_23212_22210# X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1317 vss d0 a_40352_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1318 X2.X2.X2.X2.vrefh a_54992_17452# X2.X2.X2.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1319 X1.X1.X1.X1.X1.X1.X2.vin1 a_2582_30882# X1.X1.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1320 X1.X2.X2.X2.X2.X2.X1.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1321 X1.X2.X2.X2.X2.X1.X1.vin2 a_25712_26982# X1.X2.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1322 a_46116_6104# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1323 X2.X2.X1.X2.X1.X1.X3.vin1 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1324 vdd d2 a_23212_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1325 vdd a_11072_6016# a_10686_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1326 a_46502_11822# a_46116_11822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1327 vdd a_25712_13640# a_25326_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1328 a_17222_15634# a_16836_15634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1329 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1330 a_2582_15634# a_2196_15634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1331 a_16836_27070# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1332 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1333 a_4396_9010# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1334 X2.X2.X2.X1.X2.X2.vout a_52406_16452# X2.X2.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1335 X2.X2.X2.X2.X1.X2.X2.vin1 a_54992_25076# X2.X2.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1336 X1.X2.X2.X1.X2.X1.vout a_23212_14586# X1.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1337 X1.X2.X2.X1.X1.X2.X3.vin1 a_25326_7922# X1.X2.X2.X1.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1338 vss d0 a_54992_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1339 a_2582_28976# a_2196_28976# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1340 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1341 X2.X1.X2.X1.X2.X2.X3.vin2 a_39966_17452# X2.X1.X2.X1.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1342 X1.X2.X1.X3.vin1 a_19722_18540# X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1343 a_48616_22312# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1344 a_33676_28070# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1345 X1.X2.X2.vrefh X1.X2.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1346 vdd d0 a_40352_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1347 vss d0 a_54992_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1348 vdd a_40352_26982# a_39966_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1349 a_46502_17540# a_46116_17540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1350 X2.X2.X1.X1.X2.X1.X3.vin2 a_48702_24258# X2.X2.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1351 vss d1 a_52792_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1352 vss a_40352_25076# a_39966_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1353 X2.X2.X1.X1.X3.vin2 a_49002_26164# X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1354 vdd d0 a_11072_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1355 X2.X1.X1.X2.X2.X2.vrefh a_31862_8010# X2.X1.X1.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1356 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1357 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1358 X1.X1.X2.X1.X1.X2.X3.vin2 a_10686_9828# X1.X1.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1359 X2.X2.X2.X2.X1.X2.vout a_52492_22210# X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1360 vdd a_54992_28888# a_54606_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1361 a_46502_4198# a_46116_4198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1362 X1.X2.X1.X2.X3.vin1 a_19722_10916# X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1363 X1.X2.vrefh a_11072_32700# X1.X1.X2.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1364 X2.X1.X1.X1.X1.X2.X3.vin1 a_34062_28070# X2.X1.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1365 X1.X1.X2.X2.X1.X2.X3.vin2 a_8872_24076# X1.X1.X2.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1366 X1.X2.X1.X1.X2.X2.X1.vin2 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1367 X2.X1.X1.X1.X1.X2.vrefh a_31862_30882# X2.X1.X1.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1368 X2.X1.X2.X2.X1.X2.X3.vin2 a_39966_25076# X2.X1.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1369 vdd d2 a_8572_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1370 a_17222_13728# a_16836_13728# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1371 vdd d2 a_52492_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1372 X2.X1.X2.X1.X1.X2.X3.vin2 a_39966_9828# X2.X1.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1373 vss a_38152_8828# a_37766_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1374 X1.X2.X2.X2.X3.vin2 a_22826_29834# X1.X2.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1375 vss d1 a_8872_16452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1376 X1.X1.X1.X1.X2.vrefh a_2582_27070# X1.X1.X1.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1377 X1.X3.vin2 a_20286_892# X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1378 vss a_23512_24076# a_23126_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1379 a_31862_15634# a_31476_15634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1380 vss a_38152_31700# a_37766_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1381 X2.X2.X1.X1.X1.X1.X1.vin2 X2.X2.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1382 X2.X2.X1.X1.X1.X2.X3.vin1 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1383 X1.X2.X1.X1.X2.X2.vout a_19722_22312# X1.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1384 X2.X1.X1.X1.X1.X2.vout a_34362_29936# X2.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1385 X2.X1.X1.X1.X2.X2.X3.vin1 a_34062_20446# X2.X1.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1386 X1.X3.vin1 a_14082_892# X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1387 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1388 X1.X1.X2.X2.X1.X2.X3.vin1 a_10686_23170# X1.X1.X2.X2.X1.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1389 a_17222_8010# a_16836_8010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1390 vss a_8872_27888# a_8486_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1391 X1.X2.X1.X1.X1.X2.X2.vin1 a_17222_27070# X1.X2.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1392 X2.X1.X2.X2.X3.vin1 a_37466_22210# X2.X1.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1393 X1.X1.X1.X2.X1.X1.X3.vin1 a_4782_16634# X1.X1.X1.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1394 X1.X2.X1.X1.X1.X2.vout a_19036_28070# X1.X2.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1395 X1.X2.X2.X2.X3.vin1 a_22826_22210# X1.X2.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1396 X1.X2.X1.X1.X1.X1.X3.vin2 a_16836_30882# X1.X2.X1.X1.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1397 vss a_40352_9828# a_39966_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1398 vdd d1 a_52792_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1399 a_20286_892# d5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1400 vdd d1 a_8872_24076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1401 vss a_11072_13640# a_10686_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1402 X1.X1.X1.X1.X1.X1.X3.vin2 a_2196_30882# X1.X1.X1.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1403 a_48616_7064# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1404 a_34362_7064# a_33976_7064# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1405 a_19422_31882# a_19036_31882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1406 a_31476_4198# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1407 X2.X2.X2.X1.X1.X2.X1.vin1 a_54992_7922# X2.X2.X2.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1408 X2.X2.X1.X1.X2.X1.vout a_49002_22312# X2.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1409 a_46502_28976# a_46116_28976# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1410 X1.X2.X2.X2.X1.X2.X3.vin2 a_23512_24076# X1.X2.X2.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1411 X2.X1.X2.X1.X2.X1.X2.vin1 a_40352_13640# X2.X1.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1412 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1413 a_4396_28070# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1414 a_28482_892# a_28096_892# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1415 a_17222_32788# a_16836_32788# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1416 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1417 a_16836_15634# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1418 X1.X1.X2.X1.X2.X2.X2.vin1 a_11072_17452# X1.X1.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1419 vss a_25712_7922# a_25326_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1420 a_19722_18540# a_19336_18540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1421 a_49566_892# d5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1422 a_2196_30882# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1423 vss d0 a_11072_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1424 X1.X2.X1.X1.X2.X2.vout a_19036_20446# X1.X2.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1425 a_5082_18540# a_4696_18540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1426 vdd d1 a_8872_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1427 X2.X1.X1.X2.X1.X2.X1.vin2 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1428 X2.X2.X2.X2.X3.vin2 a_52492_25982# X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1429 X2.X1.X2.X2.X2.X1.X3.vin1 a_38152_27888# X2.X1.X2.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1430 vdd d1 a_52792_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1431 X1.X1.X1.X2.X3.vin1 a_4696_14688# X1.X1.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1432 vss a_25712_21264# a_25326_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1433 X1.X2.X2.X1.X3.vin2 a_22826_14586# X1.X2.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1434 X1.X2.X1.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1435 vdd a_11072_21264# a_10686_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1436 X1.X2.X2.X1.X1.X1.X1.vin1 a_25712_4110# X1.X2.X2.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1437 a_31862_13728# a_31476_13728# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1438 vdd a_38152_16452# a_37766_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1439 a_4396_20446# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1440 a_19722_10916# a_19336_10916# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1441 X2.X1.X1.X2.X2.X2.X3.vin1 a_34062_5198# X2.X1.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1442 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1443 a_5082_10916# a_4696_10916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1444 X2.X2.X1.X1.X2.X1.vout a_48316_24258# X2.X2.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1445 vss d0 a_40352_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1446 X2.X2.X1.X2.X2.X2.X2.vin1 a_46502_4198# X2.X2.X1.X2.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1447 vss d2 a_23212_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1448 X2.X2.X1.X2.X2.X2.X3.vin1 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1449 X1.X2.X2.X1.X2.X1.X3.vin2 a_25326_13640# X1.X2.X2.X1.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1450 X2.X2.X2.X1.X3.vin2 a_52106_14586# X2.X2.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1451 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1452 vdd d0 a_40352_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1453 X2.X1.X1.X2.X1.X1.X3.vin2 a_34062_16634# X2.X1.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1454 X2.X2.X2.X2.X1.X1.X1.vin1 a_54992_19358# X2.X2.X2.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1455 X1.X2.X1.X2.X1.X2.X3.vin1 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1456 X1.X1.X2.X2.X2.X2.X3.vin2 a_10686_32700# X1.X1.X2.X2.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1457 X2.X1.X2.X3.vin2 a_37466_25982# X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1458 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1459 X2.X1.X2.X1.X1.X1.vout a_37852_6962# X2.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1460 X1.X1.X3.vin2 a_6032_892# X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1461 a_5082_22312# a_4696_22312# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1462 X2.X2.X3.vin2 a_49952_892# X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1463 a_16836_13728# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1464 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1465 a_2582_8010# a_2196_8010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1466 vdd d2 a_23212_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1467 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1468 a_34062_31882# a_33676_31882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1469 X2.X1.X1.X1.X2.X1.X3.vin2 a_31476_23258# X2.X1.X1.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1470 X2.X1.X1.X1.X3.vin1 a_34362_26164# X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1471 vdd d1 a_38152_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1472 X2.X1.X1.X2.X1.X2.X2.vin1 a_31862_11822# X2.X1.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1473 a_2196_13728# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1474 X1.X2.X1.X2.X3.vin1 a_19336_14688# X1.X2.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1475 X1.X1.X1.X1.X1.X2.X3.vin2 a_2196_27070# X1.X1.X1.X1.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1476 a_48702_24258# a_48316_24258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1477 a_31862_32788# a_31476_32788# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1478 a_19422_28070# a_19036_28070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1479 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1480 a_49002_26164# a_48616_26164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1481 X1.X1.X2.X3.vin1 a_8572_18358# X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1482 X2.X1.X1.X1.X3.vin1 a_33976_29936# X2.X1.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1483 X1.X2.X2.X1.X1.X2.X3.vin2 a_25326_9828# X1.X2.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1484 vss d0 a_11072_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1485 X1.X1.X1.X2.X2.X1.X1.vin1 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1486 X1.X1.X2.X2.X2.X1.X1.vin2 a_11072_26982# X1.X1.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1487 X1.X2.X1.X2.X1.X2.vrefh a_17222_15634# X1.X2.X1.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1488 X2.X2.X2.X2.X2.X1.X3.vin1 a_52792_27888# X2.X2.X2.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1489 X2.X1.X1.X1.X2.X1.X1.vin2 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1490 a_2196_8010# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1491 X1.X2.X1.X2.X1.X1.vout a_19036_16634# X1.X2.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1492 X2.X1.X2.X2.X1.X1.X3.vin1 a_39966_19358# X2.X1.X2.X2.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1493 X2.X2.X2.X2.X2.X1.X3.vin2 a_54606_28888# X2.X2.X2.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1494 X2.X2.X1.X2.X3.vin2 a_48616_7064# X2.X2.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1495 X1.X1.X1.X1.X1.X1.vout a_4396_31882# X1.X1.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1496 a_46116_30882# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1497 a_33676_20446# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1498 vdd a_23212_18358# a_22826_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1499 vdd a_11072_32700# a_10686_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1500 vss a_11072_30794# a_10686_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1501 vdd d2 a_23212_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1502 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1503 X2.X2.X1.X2.X2.X2.vout a_48316_5198# X2.X2.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1504 a_19036_31882# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1505 a_4396_16634# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1506 X1.X2.X1.X2.X1.X2.X3.vin2 a_16836_11822# X1.X2.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1507 a_16836_32788# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1508 X1.X1.X2.X1.X2.X2.X3.vin2 a_10686_17452# X1.X1.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1509 vdd d0 a_25712_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1510 X2.X1.X2.X1.X1.X2.X1.vin1 a_40352_7922# X2.X1.X2.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1511 vdd d0 a_25712_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1512 X2.X2.X2.X2.X2.X2.vrefh a_54992_28888# X2.X2.X2.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1513 X2.X1.X2.X2.X2.X1.vout a_37766_27888# X2.X1.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1514 X2.X1.X2.X2.X1.X2.vrefh a_40352_21264# X2.X1.X2.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1515 X1.X2.X1.X1.X2.X1.X3.vin1 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1516 X2.X2.X2.X3.vin2 a_52106_25982# X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1517 vss d2 a_52492_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1518 X1.X2.X1.X2.X2.X2.vrefh a_17222_8010# X1.X2.X1.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1519 a_2196_11822# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1520 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1521 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1522 X1.X2.X2.X3.vin1 a_23212_18358# X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1523 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1524 X1.X2.X2.X1.X1.X2.vrefh a_25712_6016# X1.X2.X2.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1525 a_46116_4198# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1526 X1.X1.X1.X2.vrefh a_2582_19446# X1.X1.X1.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1527 X1.X2.X1.X1.X1.X2.X3.vin1 a_19422_28070# X1.X2.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1528 vrefh X1.X1.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1529 X2.X1.X1.X2.X2.X2.X1.vin1 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1530 X2.X1.X2.X1.X1.X1.X3.vin2 a_38152_5016# X2.X1.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1531 X2.X1.X1.X1.X1.X1.vout a_34362_29936# X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1532 X1.X2.X1.X2.X1.X2.X1.vin1 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1533 a_2196_25164# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1534 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1535 a_49002_22312# a_48616_22312# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1536 a_34062_28070# a_33676_28070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1537 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1538 vss a_54992_11734# a_54606_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1539 vdd a_40352_11734# a_39966_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1540 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1541 vss a_25712_15546# a_25326_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1542 vdd a_11072_15546# a_10686_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1543 X2.X1.X1.X2.X2.X2.X3.vin1 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1544 vss d0 a_11072_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1545 X1.X2.X1.X1.X2.X2.X3.vin1 a_19422_20446# X1.X2.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1546 X2.X1.X2.X2.X2.X1.X3.vin2 a_39966_28888# X2.X1.X2.X2.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1547 X1.X2.X2.X2.X1.X1.X3.vin2 a_25326_21264# X1.X2.X2.X2.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1548 vss a_37852_14586# a_37466_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1549 vdd d0 a_54992_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1550 X1.X1.X1.X1.X2.X1.X1.vin1 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1551 a_46116_27070# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1552 a_43362_892# a_42976_892# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1553 X2.X2.X1.X1.X1.X1.X2.vin1 a_46502_30882# X2.X2.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1554 vdd a_25712_9828# a_25326_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1555 X2.X1.X1.X3.vin1 a_33976_26164# X2.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1556 X1.X2.X2.X1.X1.X1.vout a_23212_6962# X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1557 a_19036_28070# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1558 a_4396_5198# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1559 a_31862_9916# a_31476_9916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1560 vss a_8872_12640# a_8486_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1561 X1.X1.X2.X2.X2.X1.X3.vin1 a_10686_26982# X1.X1.X2.X2.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1562 a_48316_16634# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1563 X1.X2.X1.X1.X1.X1.X1.vin2 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1564 vss d1 a_38152_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1565 a_31476_11822# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1566 X2.X2.X2.X2.X1.X1.X1.vin2 a_54992_19358# X2.X2.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1567 X2.X2.X2.X1.X1.X1.X3.vin1 a_54606_4110# X2.X2.X2.X1.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1568 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1569 X2.X2.X2.X3.vin2 a_52492_18358# X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1570 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1571 X2.X2.X2.X1.X3.vin1 a_52106_6962# X2.X2.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1572 vss d1 a_8872_27888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1573 vdd d3 a_52492_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1574 X2.X1.X2.X2.X1.X2.vout a_37852_22210# X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1575 X1.X1.X1.X2.X1.X2.vout a_4396_12822# X1.X1.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1576 vdd a_52792_12640# a_52406_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1577 vss d0 a_11072_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1578 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1579 vdd a_8872_20264# a_8486_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1580 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1581 X1.X1.X2.X1.X1.X1.vout a_8486_5016# X1.X1.X2.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1582 X2.X1.X1.X2.X2.X2.vout a_33676_5198# X2.X1.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1583 a_4782_28070# a_4396_28070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1584 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1585 a_31476_17540# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1586 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1587 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1588 vss d0 a_25712_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1589 a_2582_30882# a_2196_30882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1590 vss a_52492_14586# a_52106_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1591 X2.X1.X2.X2.X1.X1.X3.vin1 a_39966_19358# X2.X1.X2.X2.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1592 X2.X1.X3.vin2 a_37466_18358# X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1593 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1594 X1.X2.X2.X1.X1.X2.X3.vin1 a_23512_8828# X1.X2.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1595 X1.X2.X1.X2.X1.X1.X3.vin2 a_19422_16634# X1.X2.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1596 X1.X2.X3.vin2 a_22826_18358# X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1597 X1.X2.X3.vin1 a_20672_892# X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1598 X1.X1.X1.X2.X1.X2.vout a_5082_14688# X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1599 X1.X1.X1.X1.X2.X2.X3.vin2 a_2196_19446# X1.X1.X1.X1.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1600 vss d0 a_25712_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1601 vdd a_37852_25982# a_37466_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1602 a_19422_20446# a_19036_20446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1603 vdd d0 a_11072_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1604 X1.X2.X1.X2.X2.X1.X3.vin2 a_16836_8010# X1.X2.X1.X2.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1605 X1.X1.X2.X2.X2.X2.vout a_8486_31700# X1.X1.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1606 X2.X1.X1.X1.X3.vin1 a_33976_29936# X2.X1.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1607 X2.X2.X1.X1.X2.vrefh a_46502_27070# X2.X2.X1.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1608 vdd d1 a_38152_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1609 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1610 a_4782_20446# a_4396_20446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1611 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1612 X2.X1.X3.vin2 a_35312_892# X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1613 vdd a_54992_30794# a_54606_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1614 a_17222_4198# a_16836_4198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1615 a_16836_6104# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1616 X2.X1.X2.X1.X2.X2.X1.vin2 a_40352_15546# X2.X1.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1617 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1618 X2.X1.X1.X2.X3.vin2 a_33976_7064# X2.X1.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1619 X1.X2.X2.X1.X2.X1.X2.vin1 a_25712_13640# X1.X2.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1620 a_34362_26164# a_33976_26164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1621 vdd d0 a_40352_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1622 vss a_23512_5016# a_23126_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1623 X2.X2.X1.X2.X1.X1.X3.vin1 a_48702_16634# X2.X2.X1.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1624 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1625 X2.X1.X1.X2.X1.X2.vout a_33676_12822# X2.X1.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1626 X2.X1.X2.X2.X3.vin2 a_37852_25982# X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1627 X1.X1.X1.X1.X2.X1.X3.vin1 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1628 X2.X2.X1.X1.X1.X1.X3.vin2 a_46116_30882# X2.X2.X1.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1629 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1630 vss a_54992_4110# a_54606_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1631 a_2196_6104# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1632 X1.X1.X1.X2.X2.X1.X3.vin1 a_4782_9010# X1.X1.X1.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1633 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1634 X2.X1.X1.X1.X2.X1.X2.vin1 a_31862_23258# X2.X1.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1635 vdd a_8872_31700# a_8486_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1636 a_2582_13728# a_2196_13728# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1637 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1638 X2.X2.X2.X1.X2.X1.X3.vin1 a_54606_11734# X2.X2.X2.X1.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1639 X1.X2.X2.X1.X2.X2.X3.vin1 a_25326_15546# X1.X2.X2.X1.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1640 a_31476_28976# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1641 X1.X2.X2.X2.X2.X2.vout a_23126_31700# X1.X2.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1642 X2.X2.X1.X2.X3.vin1 a_48616_14688# X2.X2.X1.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1643 X1.X1.X1.X1.X2.X2.X2.vin1 a_2582_19446# X1.X1.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1644 a_19336_26164# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1645 a_19336_7064# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1646 X1.X1.X2.X1.X2.X2.vout a_8486_16452# X1.X1.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1647 X1.X1.X1.X1.X1.X1.X3.vin2 a_4782_31882# X1.X1.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1648 vdd a_52492_25982# a_52106_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1649 X1.X1.X1.X2.X2.X1.vout a_4396_9010# X1.X1.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1650 a_46502_30882# a_46116_30882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1651 a_34062_20446# a_33676_20446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1652 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1653 vdd d4 a_23212_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1654 vdd d0 a_11072_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1655 vss d0 a_11072_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1656 a_19036_5198# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1657 a_46502_9916# a_46116_9916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1658 vdd d0 a_11072_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1659 a_4782_16634# a_4396_16634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1660 X2.X2.X2.X1.X2.X2.vrefh a_54992_13640# X2.X2.X2.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1661 X1.X2.X1.X1.X2.X1.X3.vin2 a_16836_23258# X1.X2.X1.X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1662 vdd d1 a_23512_8828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1663 X1.X1.X1.X2.X2.X1.X3.vin2 a_2196_8010# X1.X1.X1.X2.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1664 X1.X2.X1.X2.X2.X2.X1.vin1 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1665 a_34362_22312# a_33976_22312# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1666 vss a_52792_20264# a_52406_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1667 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1668 a_46116_19446# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1669 a_28096_892# d7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1670 a_2582_4198# a_2196_4198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1671 vss d0 a_40352_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1672 a_17222_11822# a_16836_11822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1673 X2.X1.X1.X2.X1.X1.vout a_34362_14688# X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1674 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1675 a_2196_23258# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1676 a_2582_11822# a_2196_11822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1677 X2.X2.X2.X3.vin1 a_52106_10734# X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1678 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1679 a_19036_20446# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1680 X1.X1.X1.X2.vrefh X1.X1.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1681 X2.X2.X1.X1.X1.X2.X3.vin2 a_46116_27070# X2.X2.X1.X1.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1682 X2.X2.X2.X1.X2.X1.vout a_52406_12640# X2.X2.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1683 a_4696_29936# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1684 X2.X2.X2.X2.X1.X1.X2.vin1 a_54992_21264# X2.X2.X2.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1685 X2.X2.X2.X1.X1.X1.X3.vin2 a_54606_6016# X2.X2.X2.X1.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1686 X1.X2.X2.X1.X2.X2.vout a_23126_16452# X1.X2.X2.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1687 a_2582_25164# a_2196_25164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1688 X2.X2.X2.X1.X1.X1.X1.vin1 X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1689 X2.X1.X2.X1.X2.X1.X3.vin2 a_39966_13640# X2.X1.X2.X1.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1690 X1.X1.X2.X1.X1.X1.X3.vin1 a_10686_4110# X1.X1.X2.X1.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1691 a_33676_24258# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1692 a_19336_22312# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1693 vss a_54992_23170# a_54606_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1694 a_46116_25164# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1695 a_33976_26164# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1696 X1.X2.X3.vin2 a_20672_892# X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1697 vss d0 a_54992_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1698 X2.X2.X1.X2.X1.X1.vout a_48316_16634# X2.X2.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1699 vss d0 a_25712_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1700 vdd a_40352_23170# a_39966_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1701 vdd a_11072_26982# a_10686_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1702 a_17222_17540# a_16836_17540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1703 vss d1 a_23512_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1704 vss a_11072_25076# a_10686_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1705 vdd d0 a_11072_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1706 X2.X1.X2.vrefh a_31862_4198# X2.X1.X1.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1707 X1.X2.X1.X2.X3.vin2 a_19336_7064# X1.X2.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1708 vss d2 a_37852_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1709 X1.X2.X2.X2.X1.X2.vrefh a_25712_21264# X1.X2.X2.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1710 vdd a_40352_7922# a_39966_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1711 X2.X1.X2.X1.X1.X1.X3.vin1 a_39966_4110# X2.X1.X2.X1.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1712 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1713 a_46502_27070# a_46116_27070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1714 a_4696_7064# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1715 X2.X1.X2.X1.X3.vin1 a_37466_6962# X2.X1.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1716 vdd a_25712_28888# a_25326_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1717 a_34062_9010# a_33676_9010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1718 X2.X1.X2.X2.X1.X1.X3.vin2 a_39966_21264# X2.X1.X2.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1719 X2.X2.X2.X2.X2.X2.X3.vin1 a_54606_30794# X2.X2.X2.X2.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1720 vss d3 a_8572_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1721 vdd d0 a_40352_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1722 vss a_38152_5016# a_37766_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1723 X2.X2.X2.X1.X1.X2.vout a_52406_8828# X2.X2.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1724 vss d1 a_8872_12640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1725 X1.X1.X1.X1.X2.X2.vrefh a_2582_23258# X1.X1.X1.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1726 a_48702_16634# a_48316_16634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1727 X1.X1.X1.X1.X2.X2.X3.vin2 a_2196_19446# X1.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1728 a_31862_11822# a_31476_11822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1729 X2.X2.X1.X2.X2.X1.X1.vin1 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1730 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1731 a_33676_9010# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1732 X2.X2.X1.X2.vrefh a_46502_19446# X2.X2.X1.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1733 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1734 X1.X1.X1.X1.X2.X1.vout a_4396_24258# X1.X1.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1735 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1736 X1.X1.X2.X1.X1.X2.X1.vin1 a_11072_7922# X1.X1.X2.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1737 X1.X1.X1.X2.X1.X2.X3.vin1 a_4782_12822# X1.X1.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1738 X1.X2.X2.X2.X2.X2.X2.vin1 X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1739 vdd d3 a_52492_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1740 X2.X2.X2.X2.X2.X2.X2.vin1 a_54992_32700# X2.X2.X2.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1741 X2.X2.X2.X2.X2.X2.X1.vin2 a_54992_30794# X2.X2.X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1742 X3.vin2 a_42976_892# X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1743 vdd d1 a_52792_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1744 vss a_11072_9828# a_10686_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1745 vdd d1 a_23512_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1746 vdd d1 a_8872_20264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1747 a_33976_22312# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1748 X1.X1.X2.X1.X3.vin2 a_8186_14586# X1.X1.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1749 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1750 X2.X2.X2.X1.X1.X1.X1.vin1 a_54992_4110# X2.X2.X2.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1751 a_48616_14688# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1752 a_31862_17540# a_31476_17540# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1753 vss a_40352_32700# a_39966_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1754 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1755 a_17222_28976# a_16836_28976# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1756 X2.X2.X1.X1.X2.X1.X1.vin1 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1757 vdd a_54992_6016# a_54606_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1758 a_16836_11822# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1759 X1.X1.X2.X1.X2.X1.X2.vin1 a_11072_13640# X1.X1.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1760 X2.X1.X1.X2.X3.vin1 a_33976_14688# X2.X1.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1761 a_4696_26164# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1762 X2.X1.X2.X3.vin2 a_37852_18358# X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1763 X2.X1.X1.X1.X2.X2.X3.vin1 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1764 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1765 X2.vrefh X2.X1.X1.X1.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1766 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1767 vdd d3 a_37852_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1768 X1.X1.X2.X2.X2.X2.X3.vin2 a_8872_31700# X1.X1.X2.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1769 X1.X1.X1.X2.X2.X2.vrefh a_2582_8010# X1.X1.X1.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1770 vdd a_37852_10734# a_37466_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1771 X2.X1.X2.X2.X2.X2.X3.vin2 a_39966_32700# X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1772 X2.X1.X2.X2.X2.X2.X3.vin1 a_39966_30794# X2.X1.X2.X2.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1773 vdd a_38152_12640# a_37766_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1774 vdd d0 a_54992_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1775 vss d0 a_40352_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1776 X2.X2.X2.X2.X1.X1.vout a_52406_20264# X2.X2.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1777 X2.X2.X2.X2.X2.X2.X2.vin1 X2.X2.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1778 a_13696_892# d6 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1779 a_16836_17540# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1780 vss a_23512_31700# a_23126_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1781 X1.X2.X1.X1.X1.X2.vout a_19722_29936# X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1782 X2.X1.X1.X1.X1.X2.X3.vin2 a_31476_27070# X2.X1.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1783 vss a_8872_8828# a_8486_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1784 X2.X2.X2.X1.X2.X2.X1.vin1 a_54992_15546# X2.X2.X2.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1785 X2.X1.X1.X2.X1.X2.X3.vin2 a_34062_12822# X2.X1.X1.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1786 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1787 X2.X1.X2.X2.X2.X1.X2.vin1 a_40352_28888# X2.X1.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1788 vss a_52792_8828# a_52406_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1789 vdd d2 a_8572_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1790 X1.X2.X2.X1.X1.X1.X3.vin1 a_25326_4110# X1.X2.X2.X1.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1791 vss a_54992_17452# a_54606_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1792 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1793 a_46116_19446# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1794 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1795 vss a_8572_10734# a_8186_10734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1796 vdd a_40352_17452# a_39966_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1797 vdd d1 a_8872_31700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1798 X2.X2.X2.X2.X1.X2.X3.vin1 a_54606_23170# X2.X2.X2.X2.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1799 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1800 a_48316_31882# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1801 X1.X1.X1.X1.X2.X1.X3.vin2 a_2196_23258# X1.X1.X1.X1.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1802 X1.X2.X2.X1.X2.X2.X1.vin2 a_25712_15546# X1.X2.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1803 a_31862_28976# a_31476_28976# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1804 a_19422_24258# a_19036_24258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1805 X1.X2.X2.X2.X2.X2.X3.vin2 a_23512_31700# X1.X2.X2.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1806 X1.X1.X2.X3.vin2 a_8186_25982# X1.X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1807 X1.X2.X1.X2.X2.X2.X3.vin2 a_16836_4198# X1.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1808 X2.X2.X1.X2.X1.X2.vout a_49002_14688# X2.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1809 a_4696_29936# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1810 a_19722_26164# a_19336_26164# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1811 X2.X2.X1.X1.X2.X2.X3.vin2 a_46116_19446# X2.X2.X1.X1.X2.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1812 X1.X1.X2.X1.X2.X2.X3.vin1 a_8872_16452# X1.X1.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1813 X1.X2.X1.X2.X2.vrefh a_17222_11822# X1.X2.X1.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1814 a_2196_4198# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1815 a_48702_9010# a_48316_9010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1816 X1.X2.X1.X2.X1.X2.vout a_19036_12822# X1.X2.X1.X2.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1817 X2.X1.X2.X1.X2.X2.X3.vin1 a_39966_15546# X2.X1.X2.X1.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1818 X1.X1.X2.X1.X1.X1.X3.vin2 a_10686_6016# X1.X1.X2.X1.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1819 X1.X2.X2.X2.X2.X1.X3.vin2 a_25326_28888# X1.X2.X2.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1820 vdd a_54992_25076# a_54606_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1821 vdd a_52492_10734# a_52106_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1822 vdd a_23512_16452# a_23126_16452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1823 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1824 X2.X1.X2.X1.X1.X1.X3.vin2 a_39966_6016# X2.X1.X2.X1.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1825 a_4396_12822# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1826 a_48316_9010# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1827 X2.X2.X2.X1.X1.X2.vrefh a_54992_6016# X2.X2.X2.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1828 vss d1 a_52792_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1829 a_16836_28976# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1830 X2.X2.X1.X1.X2.X1.X3.vin1 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1831 X1.X1.X2.X1.X2.X1.X3.vin2 a_10686_13640# X1.X1.X2.X1.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1832 a_46502_19446# a_46116_19446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1833 X2.X1.X2.X1.X1.X1.X1.vin1 a_40352_4110# X2.X1.X2.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1834 X1.X2.X1.X2.X1.X1.X1.vin1 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1835 X1.X1.X1.X2.X2.X2.X3.vin1 a_4782_5198# X1.X1.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1836 a_2582_23258# a_2196_23258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1837 vss a_8872_24076# a_8486_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1838 X1.X2.X2.vrefh a_17222_4198# X1.X2.X1.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1839 X1.X1.X2.X2.X1.X2.vrefh a_11072_21264# X1.X1.X2.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1840 a_31862_8010# a_31476_8010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1841 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1842 X2.X1.X2.X1.X2.X2.X3.vin2 a_38152_16452# X2.X1.X2.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1843 a_5082_29936# a_4696_29936# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1844 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1845 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1846 X1.X2.X2.X1.X2.X2.X3.vin1 a_23512_16452# X1.X2.X2.X1.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1847 vss a_40352_26982# a_39966_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1848 X2.X1.X3.vin1 a_35312_892# X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1849 X1.X2.X1.X1.X3.vin1 a_19722_26164# X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1850 X2.X2.X1.X1.X2.X2.X2.vin1 a_46502_19446# X2.X2.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1851 a_34062_24258# a_33676_24258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1852 X1.X1.X2.X1.X1.X1.vout a_8572_6962# X1.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1853 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1854 X2.X1.X1.X2.X1.X1.X3.vin2 a_31476_15634# X2.X1.X1.X2.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1855 a_19722_22312# a_19336_22312# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1856 X2.X1.X1.X3.vin2 a_34362_18540# X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1857 vss d0 a_54992_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1858 X2.X2.X1.X1.X1.X1.X3.vin2 a_48702_31882# X2.X2.X1.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1859 a_46502_25164# a_46116_25164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1860 vss a_38152_20264# a_37766_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1861 X2.X2.X2.X1.X1.X1.vout a_52492_6962# X2.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1862 vdd d0 a_11072_26982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1863 vss a_25712_4110# a_25326_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1864 X2.X1.X2.X1.X1.X2.vout a_37766_8828# X2.X1.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1865 vss a_25712_11734# a_25326_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1866 vss d0 a_11072_25076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1867 vdd d1 a_8872_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1868 vdd a_11072_11734# a_10686_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1869 X1.X2.X1.X2.X2.X1.X3.vin1 a_19422_9010# X1.X2.X1.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1870 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1871 vdd a_8572_29834# a_8186_29834# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1872 X2.X1.X2.X2.X1.X2.X3.vin1 a_38152_24076# X2.X1.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1873 X1.X1.X1.X2.X2.X2.X3.vin2 a_2196_4198# X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1874 a_31476_30882# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1875 vdd d1 a_52792_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1876 X1.X1.X1.X1.X2.X2.X1.vin1 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1877 vdd d0 a_25712_28888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1878 a_46116_23258# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1879 X2.X1.X1.X2.X3.vin2 a_34362_10916# X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1880 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1881 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1882 X2.X2.X1.X2.X2.X1.X3.vin1 a_48702_9010# X2.X2.X1.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1883 a_19036_24258# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1884 X1.X1.X1.X2.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1885 a_17222_9916# a_16836_9916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1886 a_48316_12822# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1887 X1.X1.X3.vin1 a_4696_18540# X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1888 X1.X2.X1.X1.X1.X2.X1.vin1 a_17222_28976# X1.X2.X1.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1889 vss d2 a_23212_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1890 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1891 vss d2 a_8572_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1892 X2.X2.X2.X1.X2.X2.X3.vin2 a_52792_16452# X2.X2.X2.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1893 X2.X2.X2.X1.X2.X2.X3.vin2 a_54606_17452# X2.X2.X2.X1.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1894 X1.X1.X1.X1.X2.X1.X3.vin1 a_4782_24258# X1.X1.X1.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1895 X2.X1.X1.X2.X1.X2.X3.vin1 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1896 X1.X1.X2.X1.X1.X2.X3.vin1 a_8872_8828# X1.X1.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1897 X2.X2.X2.X1.X1.X2.X3.vin1 a_52792_8828# X2.X2.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1898 X1.X2.X1.X1.X1.X1.vout a_19722_29936# X1.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1899 vss d0 a_11072_9828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1900 X1.X1.X1.X3.vin2 a_4696_10916# X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1901 X1.X1.X2.X1.X2.X2.vout a_8572_14586# X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1902 X2.X2.X1.X2.X2.X1.X3.vin2 a_46116_8010# X2.X2.X1.X2.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1903 a_49002_14688# a_48616_14688# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1904 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1905 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1906 X1.X2.X1.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1907 X1.X2.X2.X1.X1.X1.X3.vin2 a_25326_6016# X1.X2.X2.X1.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1908 X3.vin2 a_42976_892# X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1909 vdd a_54992_19358# a_54606_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1910 vdd d2 a_8572_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1911 X1.X1.X1.X2.X2.X2.X1.vin1 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1912 a_34062_5198# a_33676_5198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1913 X2.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1914 X2.X1.X2.X1.X1.X2.vrefh a_40352_6016# X2.X1.X2.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1915 a_5082_26164# a_4696_26164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1916 X2.X2.X2.X2.X1.X2.X3.vin1 a_52792_24076# X2.X2.X2.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1917 X2.X1.X1.X1.X2.X2.X1.vin2 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1918 X2.X2.X2.X2.X1.X2.X3.vin2 a_54606_25076# X2.X2.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1919 X1.X1.X2.X2.X1.X1.X3.vin2 a_10686_21264# X1.X1.X2.X2.X1.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1920 vss a_23212_14586# a_22826_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1921 X1.X2.X1.X2.X1.X2.X3.vin2 a_19422_12822# X1.X2.X1.X2.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1922 X1.X1.X1.X1.X3.vin2 a_4696_22312# X1.X1.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1923 X2.X1.X2.X1.X2.X2.vout a_37766_16452# X2.X1.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1924 X1.X1.X1.X1.X1.X1.X1.vin1 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1925 a_31476_27070# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1926 X1.X2.X3.vin1 a_19336_18540# X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1927 vdd d3 a_37852_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1928 X2.X1.X1.X1.X1.X1.vout a_33676_31882# X2.X1.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1929 X1.X1.X1.X2.X1.X1.X1.vin2 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1930 X2.X2.X1.X1.X2.X2.vrefh a_46502_23258# X2.X2.X1.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1931 X2.X2.X1.X1.X2.X2.X3.vin2 a_46116_19446# X2.X2.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1932 a_6032_892# a_5646_892# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1933 vdd d1 a_38152_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1934 vdd a_11072_7922# a_10686_7922# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1935 X2.X1.X1.X1.X1.X1.X3.vin1 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1936 X2.X1.X3.vin1 a_33976_18540# X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1937 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1938 X2.X2.X1.X1.X1.X1.vout a_48316_31882# X2.X2.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1939 vdd a_25712_30794# a_25326_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1940 X1.X1.X3.vin1 a_6032_892# X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1941 X2.X1.X2.X1.X2.X1.X1.vin2 a_40352_11734# X2.X1.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1942 vdd d2 a_8572_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1943 a_33676_16634# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1944 X1.X1.X2.X1.X2.X2.X1.vin2 a_11072_15546# X1.X1.X2.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1945 vdd a_52792_27888# a_52406_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1946 X2.X1.X1.X1.X1.X2.X2.vin1 a_31862_27070# X2.X1.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1947 a_46502_8010# a_46116_8010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1948 X2.X2.X2.X2.X3.vin1 a_52106_22210# X2.X2.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1949 X2.X2.X2.X2.X2.X1.X1.vin1 a_54992_26982# X2.X2.X2.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1950 X1.X2.X1.X3.vin2 a_19336_10916# X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1951 X2.X2.X1.X2.X1.X2.X3.vin1 a_48702_12822# X2.X2.X1.X2.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1952 X2.X2.X2.X2.X2.vrefh a_54992_25076# X2.X2.X2.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1953 X2.X1.X2.X2.X1.X2.vout a_37766_24076# X2.X1.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1954 X1.X1.X1.X2.X2.X1.X1.vin2 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1955 X1.X2.X2.X1.X2.X2.vout a_23212_14586# X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1956 X1.X2.X1.X1.X2.X2.X3.vin1 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1957 vss d0 a_54992_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1958 X1.X2.X2.X1.X1.X2.vout a_23126_8828# X1.X2.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1959 X1.X2.X2.X2.X2.X2.X1.vin1 X1.X2.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1960 a_2582_9916# a_2196_9916# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1961 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1962 X1.X1.X1.X1.X2.X2.X3.vin1 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1963 X2.X1.X1.X3.vin2 a_33976_10916# X2.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1964 vss d0 a_54992_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1965 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1966 a_46502_19446# a_46116_19446# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1967 a_4696_14688# d2 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1968 a_2196_21352# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1969 X1.X2.X1.X1.X3.vin2 a_19336_22312# X1.X2.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1970 a_48702_31882# a_48316_31882# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1971 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1972 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1973 X1.X1.X2.X2.X3.vin1 a_8572_25982# X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1974 X1.X2.X2.X1.X2.X1.X3.vin1 a_25326_11734# X1.X2.X2.X1.X2.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1975 X3.vin1 a_13696_892# X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1976 a_5082_29936# a_4696_29936# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1977 vss a_54992_28888# a_54606_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1978 X1.X1.X2.X3.vin1 a_8186_10734# X1.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1979 X1.X1.X1.X2.X1.X1.X2.vin1 a_2582_15634# X1.X1.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1980 X1.X2.X1.X1.X1.X2.X3.vin2 a_16836_27070# X1.X2.X1.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1981 a_20286_892# d5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1982 X2.X1.X2.X2.X2.X1.X3.vin1 a_39966_26982# X2.X1.X2.X2.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1983 vss d0 a_11072_4110# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1984 X1.X1.X2.X1.X2.X1.vout a_8486_12640# X1.X1.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1985 vss a_8572_29834# a_8186_29834# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1986 X2.X1.X2.X2.X1.X2.X3.vin2 a_39966_25076# X2.X1.X2.X2.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1987 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1988 X1.X1.X1.X2.X2.X2.vout a_4396_5198# X1.X1.X1.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1989 X1.X2.X2.X2.X2.X1.X2.vin1 a_25712_28888# X1.X2.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1990 vdd d0 a_54992_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1991 vdd a_23212_25982# a_22826_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1992 a_17222_30882# a_16836_30882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1993 vdd a_25712_6016# a_25326_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1994 X1.X1.X1.X1.X1.X2.X1.vin2 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1995 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X1996 X2.X1.X1.X1.X1.X2.vout a_33676_28070# X2.X1.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1997 a_2196_27070# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1998 X2.X2.X2.X1.X2.vrefh a_54992_9828# X2.X2.X2.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X1999 a_4782_12822# a_4396_12822# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2000 vss d2 a_37852_6962# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2001 X1.X1.X1.X2.X2.X1.vout a_5082_7064# X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2002 a_31862_6104# a_31476_6104# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2003 vdd a_8572_22210# a_8186_22210# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2004 X2.X2.X2.X3.vin2 a_52106_25982# X2.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2005 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2006 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2007 X2.X1.X1.X2.X2.X1.X3.vin2 a_31476_8010# X2.X1.X1.X2.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2008 X1.X1.X1.X2.X2.X2.vrefh X1.X1.X1.X2.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2009 vss d2 a_52492_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2010 X1.X1.X1.X1.X1.X1.X3.vin1 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2011 X2.X2.X1.X1.X1.X1.X1.vin2 X2.X2.X1.X1.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2012 X1.X2.X2.X2.X3.vin1 a_23212_25982# X1.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2013 vss d1 a_8872_24076# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2014 X1.X1.X1.X2.X3.vin2 a_4696_7064# X1.X1.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2015 a_31476_6104# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2016 X1.X1.X1.X2.X1.X1.X3.vin1 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2017 X2.X1.X1.X2.X2.X1.X3.vin2 a_34062_9010# X2.X1.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2018 X2.X2.X1.X1.X2.X1.X3.vin2 a_46116_23258# X2.X2.X1.X1.X2.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2019 X2.X2.X1.X2.X2.X2.vrefh a_46502_8010# X2.X2.X1.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2020 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2021 X1.X2.X2.X1.X2.X1.vout a_23126_12640# X1.X2.X2.X1.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2022 X2.X1.X2.X2.X2.X2.X1.vin1 a_40352_30794# X2.X1.X2.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2023 a_48702_5198# a_48316_5198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2024 X2.X1.X2.X1.X1.X2.X3.vin2 a_39966_9828# X2.X1.X2.X1.X1.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2025 vdd a_8572_14586# a_8186_14586# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2026 X2.X1.X1.X2.X1.X2.vrefh a_31862_15634# X2.X1.X1.X2.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2027 X1.X1.X2.X1.X2.X2.X3.vin1 a_10686_15546# X1.X1.X2.X1.X2.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2028 X2.X2.X2.X2.X1.X1.X3.vin1 a_54606_19358# X2.X2.X2.X2.X1.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2029 vss d1 a_38152_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2030 vss a_54992_19358# a_54606_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2031 X2.X1.X2.X2.X2.X1.X3.vin2 a_38152_27888# X2.X1.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2032 a_46116_21352# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2033 vss a_25712_23170# a_25326_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2034 X1.X1.X1.X2.X2.X1.X3.vin1 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2035 X2.X2.X1.X2.X1.X2.vout a_48316_12822# X2.X2.X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2036 vss d0 a_25712_11734# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2037 X1.X2.X2.X1.X3.vin2 a_22826_14586# X1.X2.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2038 vdd a_11072_23170# a_10686_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2039 vdd d0 a_11072_11734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2040 vss a_37852_22210# a_37466_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2041 X1.X2.X2.X1.X1.X1.X3.vin1 a_23512_5016# X1.X2.X2.X1.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2042 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2043 vdd a_40352_4110# a_39966_4110# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2044 a_31862_30882# a_31476_30882# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2045 a_46502_23258# a_46116_23258# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2046 vss d0 a_40352_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2047 a_17222_27070# a_16836_27070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2048 a_19422_9010# a_19036_9010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2049 X1.X2.X2.X2.X2.X2.X3.vin1 a_25326_30794# X1.X2.X2.X2.X2.X2.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2050 vdd d0 a_40352_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2051 X1.X1.X1.X1.X1.X2.vout a_4396_28070# X1.X1.X1.X1.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2052 X1.X2.X1.X2.X1.X1.X3.vin2 a_16836_15634# X1.X2.X1.X2.X1.X1.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2053 X2.X2.X2.X2.X2.X1.vout a_52406_27888# X2.X2.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2054 X2.X2.X2.X1.X1.X1.vout a_52406_5016# X2.X2.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2055 a_48316_24258# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2056 a_34362_14688# a_33976_14688# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2057 vdd a_8572_6962# a_8186_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2058 a_48702_12822# a_48316_12822# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2059 X1.X1.X1.X2.X1.X1.X3.vin2 a_2196_15634# X1.X1.X1.X2.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2060 X1.X1.X1.X3.vin1 a_5082_18540# X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2061 a_31476_19446# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2062 a_19422_16634# a_19036_16634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2063 vss d3 a_52492_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2064 a_33676_5198# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2065 X2.X1.X2.X1.X1.X1.X1.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2066 X1.X2.X1.X2.X1.X1.vout a_19722_14688# X1.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2067 vdd a_52492_6962# a_52106_6962# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2068 a_16836_30882# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2069 X2.X1.X1.X2.X1.X2.X1.vin1 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2070 a_2196_15634# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2071 X1.X1.X1.X1.X1.X2.X3.vin1 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2072 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2073 X1.X1.X2.X2.X1.X1.vout a_8486_20264# X1.X1.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2074 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2075 X1.X1.X1.X1.X2.X2.vout a_4396_20446# X1.X1.X1.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2076 X1.X1.X2.X1.X1.X1.X1.vin1 a_11072_4110# X1.X1.X2.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2077 X1.X1.X1.X2.X3.vin1 a_5082_10916# X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2078 vdd d0 a_54992_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2079 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2080 a_16836_8010# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2081 vdd d1 a_23512_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2082 X1.X2.X1.X2.X2.X2.X3.vin1 a_19422_5198# X1.X2.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2083 X2.X2.X2.X2.X2.X1.X3.vin2 a_52792_27888# X2.X2.X2.X2.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2084 X2.X2.X2.X2.X2.X1.X3.vin2 a_54606_28888# X2.X2.X2.X2.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2085 a_31476_25164# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2086 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2087 a_46116_32788# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2088 a_19336_14688# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2089 vdd d0 a_54992_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2090 a_46116_17540# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2091 X2.X2.X1.X1.X2.X2.X1.vin1 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2092 vss a_52492_22210# a_52106_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2093 vss a_11072_32700# a_10686_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2094 vss a_37852_25982# a_37466_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2095 a_33976_7064# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2096 X1.X2.X1.X2.X2.X1.X3.vin1 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2097 vss d2 a_23212_14586# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2098 X1.X2.X2.X3.vin2 a_22826_25982# X1.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2099 X2.X2.X1.X2.X2.X2.X3.vin1 a_48702_5198# X2.X2.X1.X2.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2100 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2101 X1.X1.X1.X1.X2.X2.vout a_5082_22312# X1.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2102 a_31862_27070# a_31476_27070# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2103 X1.X2.X1.X2.X1.X2.X3.vin1 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2104 X2.X1.X1.X1.X1.X1.X3.vin1 a_34062_31882# X2.X1.X1.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2105 X1.X1.X2.vrefh a_2582_4198# X1.X1.X1.X2.X2.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2106 a_46502_6104# a_46116_6104# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2107 vdd d0 a_11072_6016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2108 X2.X1.X1.X1.X1.X1.X1.vin2 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2109 a_46116_9916# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2110 X2.X2.X3.vin1 a_48616_18540# X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2111 vdd d1 a_23512_5016# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2112 vdd d4 a_8572_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2113 X2.X1.X2.X2.X1.X2.X1.vin2 a_40352_23170# X2.X1.X2.X2.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2114 vdd d0 a_25712_30794# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2115 X2.X1.X2.X2.X2.X1.vout a_37766_27888# X2.X1.X2.X2.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2116 X1.X1.X2.X1.X3.vin1 a_8186_6962# X1.X1.X2.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2117 X1.X2.X2.X2.X1.X1.vout a_23126_20264# X1.X2.X2.X2.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2118 a_4782_9010# a_4396_9010# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2119 a_2196_13728# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2120 a_34062_16634# a_33676_16634# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2121 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2122 vdd d1 a_52792_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2123 X2.X2.X1.X1.X2.X1.X3.vin1 a_48702_24258# X2.X2.X1.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2124 a_46116_6104# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2125 X2.X3.vin2 a_49566_892# X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2126 X1.X2.X2.X1.X1.X2.X1.vin2 a_25712_7922# X1.X2.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2127 vss a_8872_5016# a_8486_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2128 X2.X1.X1.X1.X2.X2.vout a_33676_20446# X2.X1.X1.X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2129 X2.X2.X2.X1.X2.X1.X1.vin1 a_54992_11734# X2.X2.X2.X1.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2130 vss a_40352_6016# a_39966_6016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2131 X2.X2.X1.X2.X2.X2.X3.vin2 a_46116_4198# X2.X2.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2132 X2.X2.X1.X3.vin2 a_48616_10916# X2.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2133 vss a_52792_5016# a_52406_5016# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2134 X1.X1.X2.X2.X2.X1.X2.vin1 a_11072_28888# X1.X1.X2.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2135 a_16836_27070# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2136 X2.X3.vin1 a_43362_892# X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2137 X1.X2.X1.X1.X1.X1.X2.vin1 a_17222_30882# X1.X2.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2138 X1.X2.X1.X1.X1.X1.vout a_19036_31882# X1.X2.X1.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2139 a_4396_9010# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2140 vss a_54992_13640# a_54606_13640# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2141 a_5082_14688# a_4696_14688# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2142 X1.X1.X1.X2.X1.X1.vout a_4396_16634# X1.X1.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2143 a_46116_15634# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2144 vss a_25712_17452# a_25326_17452# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2145 vdd a_40352_13640# a_39966_13640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2146 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2147 X1.X2.X1.X1.X1.X1.X3.vin1 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2148 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X1.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2149 a_2582_21352# a_2196_21352# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2150 vdd a_11072_17452# a_10686_17452# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2151 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2152 X2.X2.X2.X2.X1.X1.X3.vin1 a_54606_19358# X2.X2.X2.X2.X1.X1.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2153 X1.X2.X2.X2.X1.X2.X3.vin1 a_25326_23170# X1.X2.X2.X2.X1.X2.X1.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2154 a_33976_14688# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2155 X2.X2.X3.vin2 a_52106_18358# X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2156 X1.X2.X2.X1.X2.X1.X1.vin2 a_25712_11734# X1.X2.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2157 a_19036_16634# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2158 X2.X2.X1.X1.X3.vin2 a_48616_22312# X2.X2.X1.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2159 vss d0 a_54992_28888# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2160 vdd a_38152_27888# a_37766_27888# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2161 vss a_52492_25982# a_52106_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2162 X1.X1.X2.X1.X3.vin1 a_8572_10734# X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2163 a_4396_31882# d1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2164 a_46116_28976# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2165 vss d0 a_40352_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2166 X2.X2.X1.X1.X1.X1.X1.vin1 a_46502_32788# X2.X2.X1.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2167 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2168 X1.X1.X2.X1.X2.X1.X3.vin1 a_8872_12640# X1.X1.X2.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2169 X2.X2.X1.X2.X1.X1.X1.vin2 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2170 a_2196_32788# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2171 X2.X1.X2.X1.X2.X1.X3.vin1 a_39966_11734# X2.X1.X2.X1.X2.X1.X1.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2172 a_4696_18540# d4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2173 vdd d3 a_23212_25982# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2174 vss d1 a_38152_8828# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2175 vdd a_54992_21264# a_54606_21264# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2176 vdd a_25712_25076# a_25326_25076# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2177 X1.X1.X2.X1.X1.X2.vrefh a_11072_6016# X1.X1.X2.X1.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2178 X1.X1.X1.X2.X2.X1.X3.vin1 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2179 vdd a_23212_10734# a_22826_10734# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2180 X2.X1.X1.X1.X1.X2.X3.vin2 a_34062_28070# X2.X1.X1.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2181 a_2582_27070# a_2196_27070# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2182 vdd a_23512_12640# a_23126_12640# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2183 a_48316_5198# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2184 X2.X2.X1.X2.X2.X1.X1.vin2 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2185 vdd d0 a_40352_9828# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2186 a_4696_10916# d3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2187 X2.X2.X1.X1.X2.X2.X3.vin1 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2188 vss d1 a_23512_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2189 X2.X2.X1.X2.X2.X2.X1.vin1 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2190 a_17222_19446# a_16836_19446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2191 a_20672_892# a_20286_892# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2192 a_49002_7064# a_48616_7064# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2193 a_31862_4198# a_31476_4198# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2194 X1.X2.X2.X1.X3.vin1 a_23212_10734# X1.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2195 a_17222_8010# a_16836_8010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2196 X2.X1.X2.X1.X2.X1.X3.vin2 a_38152_12640# X2.X1.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2197 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2198 X1.X2.X1.X1.X2.vrefh a_17222_27070# X1.X2.X1.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2199 a_31476_19446# d0 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2200 X1.X2.X2.X1.X2.X1.X3.vin1 a_23512_12640# X1.X2.X2.X1.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2201 X1.X2.X1.X1.X1.X2.vout a_19036_28070# X1.X2.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2202 vss d0 a_25712_7922# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2203 a_49952_892# a_49566_892# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2204 vdd a_8572_18358# a_8186_18358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2205 X2.X2.X1.X2.X1.X1.X2.vin1 a_46502_15634# X2.X2.X1.X2.X1.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2206 a_33676_31882# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2207 vss a_11072_26982# a_10686_26982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2208 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X2.vrefh vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2209 a_48616_7064# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2210 X2.X1.X1.X2.X1.X2.X3.vin2 a_31476_11822# X2.X1.X1.X2.X1.X2.X2.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2211 vss d0 a_54992_19358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2212 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2213 a_46502_21352# a_46116_21352# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2214 vss d0 a_25712_23170# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2215 X2.X2.X1.X1.X2.X1.vout a_48316_24258# X2.X2.X1.X1.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2216 vss d4 a_52492_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2217 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2218 a_17222_25164# a_16836_25164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2219 X2.X1.X2.X1.X1.X1.vout a_37766_5016# X2.X1.X2.X1.X1.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2220 vdd d0 a_11072_23170# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2221 a_4396_28070# d1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2222 X2.X2.X1.X1.X1.X2.X1.vin2 a_46502_28976# X2.X2.X1.X1.X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2223 vss d2 a_37852_22210# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2224 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2225 X1.X1.X2.X2.X2.X1.X3.vin2 a_10686_28888# X1.X1.X2.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2226 X1.X2.X2.X1.X1.X1.X1.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2227 X2.X1.X2.X2.X1.X1.X3.vin1 a_38152_20264# X2.X1.X2.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2228 vdd a_54992_32700# a_54606_32700# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2229 vss a_54992_30794# a_54606_30794# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2230 X2.X1.X2.X2.vrefh a_40352_17452# X2.X1.X2.X1.X2.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2231 a_48616_18540# d4 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2232 X2.X1.X1.X2.X2.X2.X3.vin2 a_31476_4198# X2.X1.X2.vrefh vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2233 X1.X2.X2.X2.X2.X2.X1.vin1 a_25712_30794# X1.X2.X2.X2.X2.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2234 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2235 X1.X1.X1.X1.X1.X2.X3.vin1 a_4782_28070# X1.X1.X1.X1.X1.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2236 X2.X1.X1.X2.X1.X1.X3.vin1 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2237 a_42976_892# d6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2238 X1.X1.X1.X1.X1.X2.vrefh a_2582_30882# X1.X1.X1.X1.X1.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2239 a_48702_24258# a_48316_24258# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2240 X1.X1.X2.vrefh X1.X1.X1.X2.X2.X2.X2.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2241 vss a_40352_21264# a_39966_21264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2242 a_31862_19446# a_31476_19446# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2243 X2.X2.X1.X1.X1.X1.X3.vin1 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2244 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2245 vss a_37852_18358# a_37466_18358# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2246 X1.X2.X2.X1.X3.vin1 a_22826_6962# X1.X2.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2247 X2.X2.X1.X2.X1.X1.X3.vin1 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2248 a_48616_10916# d3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2249 X2.X2.X2.X1.X3.vin2 a_52492_10734# X2.X2.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2250 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2251 X2.X1.X2.X2.X1.X2.X2.vin1 a_40352_25076# X2.X1.X2.X2.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2252 vss a_8872_31700# a_8486_31700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2253 X1.X2.X1.X2.X2.X1.vout a_19722_7064# X1.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2254 X2.X2.X2.X1.X2.X1.X3.vin2 a_52792_12640# X2.X2.X2.X1.X2.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2255 a_2582_15634# a_2196_15634# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2256 X2.X2.X2.X1.X2.X1.X3.vin2 a_54606_13640# X2.X2.X2.X1.X2.X1.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2257 X1.X1.X1.X1.X2.X2.X3.vin1 a_4782_20446# X1.X1.X1.X1.X2.X2.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2258 X1.X1.X2.X2.X1.X1.X3.vin2 a_8872_20264# X1.X1.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2259 X1.X2.X2.X1.X2.X2.X3.vin2 a_25326_17452# X1.X2.X2.X1.X2.X2.X2.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2260 X1.X2.X2.X1.X1.X2.X2.vin1 a_25712_9828# X1.X2.X2.X1.X1.X2.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2261 X1.X2.X1.X1.X1.X1.X3.vin1 a_19422_31882# X1.X2.X1.X1.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2262 vss d0 a_40352_15546# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2263 X2.X1.X2.X1.X1.X2.X3.vin1 a_38152_8828# X2.X1.X2.X1.X1.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2264 X2.X2.X1.X2.X2.X1.X3.vin1 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2265 X1.X1.X2.X2.X3.vin1 a_8186_22210# X1.X1.X2.X2.X1.X1.vout vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2266 a_2582_8010# a_2196_8010# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2267 X2.X2.X1.X2.X2.X1.vout a_49002_7064# X2.X2.X1.X2.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2268 X1.X2.X1.X2.X2.X1.vout a_19036_9010# X1.X2.X1.X2.X2.X1.X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2269 a_48616_22312# d2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2270 X1.X2.X1.X3.vin2 a_19722_18540# X1.X2.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2271 X2.X1.X1.X1.X3.vin2 a_34362_26164# X2.X1.X1.X3.vin1 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2272 a_31862_25164# a_31476_25164# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2273 vss a_23512_20264# a_23126_20264# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2274 a_46502_32788# a_46116_32788# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2275 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2276 a_19722_14688# a_19336_14688# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2277 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin1 vss sky130_fd_pr__res_high_po_0p35 l=1.09
X2278 a_16836_19446# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2279 vdd a_54992_15546# a_54606_15546# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2280 a_46502_17540# a_46116_17540# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2281 vss d0 a_11072_32700# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2282 vss d3 a_37852_25982# vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2283 vdd a_25712_19358# a_25326_19358# vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2284 a_19422_5198# a_19036_5198# vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2285 X2.X2.X2.X2.X1.X1.X3.vin1 a_52792_20264# X2.X2.X2.X2.X1.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2286 X2.X1.X2.X3.vin1 a_37466_10734# X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2287 X2.X2.X2.X2.X1.X1.X3.vin2 a_54606_21264# X2.X2.X2.X2.X1.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2288 vout a_28096_892# X3.vin2 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2289 X2.X1.X2.X2.X2.X2.X3.vin1 a_38152_31700# X2.X1.X2.X2.X2.X2.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2290 X1.X2.X2.X2.X1.X2.X3.vin2 a_25326_25076# X1.X2.X2.X2.X2.vrefh vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2291 X1.X2.X2.X3.vin1 a_22826_10734# X1.X2.X2.X1.X3.vin2 vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2292 X2.X2.X1.X2.X3.vin2 a_48616_7064# X2.X2.X1.X2.X2.X1.vout vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2293 X2.X1.X2.X1.X2.X1.vout a_37766_12640# X2.X1.X2.X1.X2.X1.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2294 X1.X1.X2.X1.X1.X2.vout a_8486_8828# X1.X1.X2.X1.X1.X2.X3.vin1 vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
X2295 a_31476_23258# d0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 X1.X2.X1.X3.vin2 X1.X2.X2.X1.X3.vin2 7.46e-20
C1 X1.X1.X1.X1.X1.X2.vrefh vdd 0.43f
C2 X1.X2.X2.X3.vin1 a_22826_14586# 7.98e-19
C3 X2.X1.X1.X1.X2.vrefh d3 6.65e-20
C4 a_22826_6962# a_23212_6962# 0.419f
C5 a_48702_20446# X2.X2.X3.vin1 1.64e-19
C6 X2.X2.X1.X1.X2.X2.X3.vin2 a_49002_18540# 0.00846f
C7 d1 a_31862_6104# 3.41e-19
C8 a_4782_12822# d1 0.0749f
C9 X1.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin2 0.0128f
C10 X1.X2.X2.X2.X1.X2.X2.vin1 d1 1.03e-19
C11 a_5082_29936# X1.X1.X1.X1.X1.X1.X3.vin2 0.00815f
C12 a_5082_29936# vdd 0.477f
C13 X1.X1.X2.X2.X1.X2.vout X1.X1.X2.X2.X1.X1.vout 0.507f
C14 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.vout 0.326f
C15 d2 a_38152_8828# 0.00287f
C16 d3 X1.X1.X2.X3.vin2 0.511f
C17 a_39966_25076# d2 0.00792f
C18 X2.X1.X1.X2.vrefh vdd 0.414f
C19 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X1.vin2 0.216f
C20 X1.X1.X2.X1.X1.X1.X3.vin2 d0 4.34e-19
C21 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X2.X1.X1.vin1 0.668f
C22 d3 X2.X2.X1.X1.X2.X2.vout 8.47e-19
C23 X1.X1.X2.X2.X2.vrefh d3 6.65e-20
C24 X1.X2.X2.X2.X2.X2.X2.vin1 a_23512_31700# 5.34e-19
C25 X1.X1.X2.X1.X2.X2.X3.vin1 a_8872_16452# 0.199f
C26 X2.X2.X1.X2.X2.X1.vout a_48616_7064# 0.169f
C27 a_48702_9010# a_49002_7064# 4.19e-20
C28 X2.X2.X2.X1.X3.vin1 a_52492_10734# 0.169f
C29 a_25326_17452# X1.X2.X2.X1.X2.X2.X3.vin1 0.00207f
C30 X2.X2.X3.vin2 a_52406_8828# 2.33e-19
C31 X1.X1.X2.X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X3.vin1 0.00118f
C32 a_19336_10916# X1.X2.X1.X2.X2.X1.X3.vin1 0.00251f
C33 X2.X2.X1.X1.X1.X1.X2.vin1 X2.X2.X1.X1.X1.X1.X1.vin1 0.0689f
C34 X1.X1.X2.X2.X2.X1.X3.vin1 X1.X1.X2.X2.X2.X2.vrefh 0.00118f
C35 X2.X1.X2.X1.X2.vrefh a_40352_9828# 0.118f
C36 a_48316_31882# a_46502_32788# 1.06e-19
C37 X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X3.vin2 0.0533f
C38 X2.X2.X1.X2.X2.X1.vout vdd 0.775f
C39 a_52406_27888# a_52492_29834# 3.14e-19
C40 d2 a_10686_9828# 0.00792f
C41 X2.X2.X1.X2.X1.X2.X1.vin2 a_46502_11822# 8.88e-20
C42 X1.X2.X1.X2.vrefh vdd 0.414f
C43 d3 a_48702_12822# 0.00122f
C44 a_31862_32788# vdd 0.554f
C45 X1.X2.X1.X1.X3.vin2 d1 0.00807f
C46 X1.X2.X2.X2.X3.vin1 a_23212_25982# 0.17f
C47 X2.X2.X1.X1.X1.X2.vout X2.X2.X1.X1.X1.X1.vout 0.507f
C48 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin1 0.195f
C49 X1.X2.X2.X2.X2.X2.X2.vin1 d0 0.199f
C50 X1.X1.X2.X2.X1.X1.X3.vin2 a_11072_21264# 0.354f
C51 X1.X2.X1.X2.X3.vin2 d1 0.00807f
C52 a_25326_26982# d1 3.95e-19
C53 a_2582_21352# d1 3.41e-19
C54 a_54992_9828# vdd 1.05f
C55 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X2.vin1 0.564f
C56 X1.X1.X2.X2.X1.X2.X3.vin1 a_8872_24076# 0.199f
C57 X2.X2.X1.X2.X1.X2.X3.vin1 a_48316_12822# 0.199f
C58 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin2 7.84e-19
C59 X2.X2.X1.X1.X2.X1.X3.vin1 a_48316_24258# 0.199f
C60 a_16836_21352# d2 0.00274f
C61 a_46116_32788# d1 2.25e-20
C62 a_52406_8828# X2.X2.X2.X1.X1.X2.vout 0.418f
C63 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X3.vin1 0.206f
C64 d0 X1.X2.X1.X2.X2.X2.X1.vin2 0.276f
C65 X2.X1.X1.X2.X1.X1.X3.vin2 a_31862_15634# 0.567f
C66 X2.X1.X2.X1.X1.X2.X3.vin2 vdd 0.787f
C67 X1.X2.X2.X2.X2.X1.X1.vin1 a_25712_26982# 0.195f
C68 a_54606_32700# a_54992_32700# 0.419f
C69 d3 X2.X1.X1.X3.vin2 0.482f
C70 a_25326_25076# X1.X2.X2.X2.X1.X2.X3.vin1 0.00207f
C71 a_16836_25164# d0 0.518f
C72 d3 X2.X2.X1.X2.X1.X1.vout 0.00883f
C73 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X2.vin1 0.564f
C74 X2.X2.X2.X2.X2.X1.X3.vin1 d0 4.36e-19
C75 a_46502_32788# X2.X2.X1.X1.X1.X1.X1.vin1 0.42f
C76 a_46116_32788# X2.X2.X1.X1.X1.X1.X3.vin1 0.354f
C77 a_46502_19446# d1 0.00148f
C78 d2 X2.X1.X1.X2.X3.vin1 0.0014f
C79 X1.X1.X2.X2.X3.vin1 d4 3.38e-19
C80 X2.X1.X2.vrefh d5 0.00132f
C81 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X1.X2.vout 0.075f
C82 X2.X2.X1.X1.X2.X2.X1.vin1 vdd 0.592f
C83 X1.X2.X2.X1.X2.X2.X2.vin1 a_25712_17452# 0.197f
C84 d4 X1.X2.X2.X1.X2.X2.X2.vin1 8.68e-20
C85 X3.vin1 X3.vin2 0.514f
C86 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X3.vin2 8.93e-19
C87 a_10686_17452# d1 0.00148f
C88 X2.X2.X2.X1.X2.X1.vout a_52406_12640# 0.422f
C89 d3 X2.X1.X1.X1.X2.X1.vout 0.00226f
C90 X3.vin1 a_20672_892# 5.96e-19
C91 a_19336_18540# a_19422_16634# 3.21e-19
C92 a_19722_18540# a_19036_16634# 2.97e-19
C93 a_49002_10916# vdd 0.487f
C94 d3 X1.X1.X1.X2.X2.X1.vout 0.00146f
C95 a_31476_19446# d1 2.92e-22
C96 d3 X2.X2.X1.X1.X2.X1.X1.vin1 6.34e-20
C97 a_34062_28070# vdd 0.47f
C98 d2 X2.X1.X2.X1.X2.X1.X1.vin1 0.0105f
C99 a_38152_12640# a_37466_10734# 2.97e-19
C100 X1.X1.X1.X2.X1.X1.X3.vin1 d2 0.104f
C101 d2 a_23212_6962# 0.625f
C102 X1.X2.X2.X1.X1.X2.vrefh a_25712_6016# 0.118f
C103 a_46116_23258# d2 0.00464f
C104 a_8572_29834# X1.X1.X2.X2.X2.X1.X3.vin2 0.00546f
C105 X2.X2.X1.X1.X2.X1.vout d1 0.0238f
C106 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin2 0.12f
C107 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X3.vin1 2.33e-19
C108 X1.X1.X3.vin2 X1.X1.X2.X1.X2.X2.vout 3.38e-19
C109 a_8186_22210# X1.X1.X2.X2.X1.X1.vout 0.387f
C110 a_52492_10734# a_52406_8828# 3.3e-19
C111 X1.X1.X1.X2.X2.X2.X1.vin1 d1 0.0118f
C112 X1.X2.X2.X2.X1.X2.X2.vin1 a_25712_25076# 0.197f
C113 d0 X2.X1.X2.X2.X2.X2.X3.vin2 4.34e-19
C114 d2 X2.X2.X2.X1.X2.X2.X3.vin1 0.153f
C115 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin2 0.1f
C116 d2 a_19036_5198# 0.00393f
C117 a_25326_6016# X1.X2.X2.X1.X1.X1.X3.vin2 0.567f
C118 d0 a_40352_4110# 0.518f
C119 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X3.vin1 0.00118f
C120 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X3.vin2 8.93e-19
C121 a_17222_6104# d2 6.36e-19
C122 X2.X2.X2.X2.vrefh vdd 0.414f
C123 X2.X1.X1.X1.X1.X1.X1.vin2 a_31476_30882# 1.78e-19
C124 a_16836_19446# d1 2.92e-22
C125 d3 X2.X2.X1.X1.X1.X1.vout 0.0408f
C126 X1.X2.X1.X1.X2.X2.X1.vin2 a_17222_19446# 8.88e-20
C127 d0 X2.X1.X2.X1.X2.vrefh 0.848f
C128 d2 a_40352_15546# 0.00274f
C129 d3 X1.X2.X1.X2.X2.X1.X1.vin1 6.34e-20
C130 a_33976_18540# a_31862_17540# 5.36e-21
C131 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin1 0.52f
C132 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 0.234f
C133 X1.X2.X2.X2.X1.X2.X1.vin1 a_25712_21264# 1.64e-19
C134 d4 X2.X1.X3.vin1 0.287f
C135 X2.X2.X2.X1.X2.X1.X3.vin1 vdd 0.997f
C136 X2.X1.X1.X1.X2.X2.vout a_33676_20446# 0.36f
C137 a_34362_22312# a_34062_20446# 5.55e-20
C138 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.vrefh 2.33e-19
C139 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.vout 0.118f
C140 X1.X1.X2.X2.X2.X2.X3.vin1 a_8872_31700# 0.199f
C141 X1.X2.X2.X2.X2.X1.vout vdd 0.775f
C142 X2.X1.X2.X2.X1.X2.X3.vin1 d2 0.155f
C143 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin1 0.267f
C144 X1.X1.X2.X2.X1.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin2 0.0128f
C145 d0 a_31862_11822# 0.0489f
C146 X1.X1.X2.X1.X3.vin1 a_8486_8828# 9.54e-19
C147 a_17222_32788# d1 2.7e-19
C148 d2 X1.X1.X2.X1.X1.X2.X3.vin1 0.157f
C149 X1.X1.X2.X1.X2.X2.X1.vin2 a_10686_15546# 0.273f
C150 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 2.23e-19
C151 a_25712_23170# d2 0.00351f
C152 a_2196_19446# d1 2.92e-22
C153 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 1.22e-19
C154 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X3.vin1 2.33e-19
C155 X2.vrefh d2 0.0108f
C156 X2.X2.X3.vin1 a_52106_18358# 5.87e-20
C157 a_8486_24076# a_8572_22210# 3.38e-19
C158 X1.X1.X1.X1.X2.X2.X3.vin1 a_2582_19446# 0.00207f
C159 a_25326_32700# X1.X2.X2.X2.X2.X2.X1.vin2 8.88e-20
C160 X2.X2.X1.X2.X1.X2.X3.vin1 d1 0.146f
C161 X1.X2.X1.X1.X2.X1.X2.vin1 vdd 0.576f
C162 X1.X2.X1.X2.X2.X2.X2.vin1 a_16836_4198# 0.197f
C163 a_16836_6104# a_16836_4198# 0.00396f
C164 X1.X1.X3.vin1 X1.X1.X2.X1.X3.vin2 6.26e-19
C165 a_8872_27888# d1 0.521f
C166 a_22826_22210# a_23512_20264# 2.86e-19
C167 X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin1 4.41e-19
C168 X1.X1.X1.X1.X2.X1.X1.vin2 d1 4.01e-19
C169 X1.X2.X1.X2.X2.X2.X2.vin1 X1.X2.X2.vrefh 0.564f
C170 a_23126_5016# X1.X2.X2.X1.X1.X1.X3.vin1 0.428f
C171 a_23126_8828# a_23512_8828# 0.419f
C172 d2 X1.X2.X1.X2.X1.X1.vout 0.00169f
C173 X2.X2.X1.X1.X1.X2.X2.vin1 d1 1.03e-19
C174 a_52406_31700# X2.X2.X2.X2.X2.X2.X2.vin1 0.00351f
C175 a_37766_20264# a_37852_18358# 3.21e-19
C176 X2.X2.X2.X2.X2.X2.X3.vin1 a_54606_32700# 0.00207f
C177 d3 X1.X2.X2.X1.X3.vin2 0.387f
C178 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X1.vin2 0.1f
C179 d1 X3.vin1 0.0325f
C180 d2 X2.X2.X2.X2.X2.X2.X3.vin1 0.0571f
C181 a_19722_18540# vdd 0.478f
C182 X2.X2.X1.X1.X2.vrefh d2 0.158f
C183 d2 a_8486_27888# 0.00123f
C184 X1.X1.X1.X1.X2.X1.X1.vin1 d2 0.0105f
C185 a_31476_27070# X2.X1.X1.X1.X1.X2.X1.vin2 1.78e-19
C186 X2.X1.X1.X1.X1.X1.X3.vin2 a_31862_30882# 0.567f
C187 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X3.vin1 0.0131f
C188 X1.X2.X2.X1.X2.X2.X3.vin1 a_22826_14586# 0.00874f
C189 X1.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X3.vin1 0.0321f
C190 X1.X1.X2.X2.X1.X2.X1.vin2 a_10686_23170# 0.273f
C191 a_37466_10734# X2.X1.X2.X1.X3.vin1 0.385f
C192 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X1.vin2 0.216f
C193 d0 a_10686_11734# 0.0675f
C194 a_54606_25076# vdd 0.542f
C195 X2.X2.X2.X2.X1.X1.X3.vin2 d4 6.94e-19
C196 X2.X1.X1.X1.X1.X2.X3.vin2 a_31862_28976# 7.84e-19
C197 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X3.vin1 0.587f
C198 a_33676_28070# X2.X1.X1.X1.X1.X2.X3.vin1 0.199f
C199 X2.X2.X2.X1.X3.vin2 a_52492_14586# 0.363f
C200 d2 X1.X2.X1.X2.X2.X1.vout 0.0909f
C201 a_54992_7922# a_54992_6016# 0.00396f
C202 X1.X1.X2.X1.X1.X2.X1.vin2 a_10686_7922# 0.273f
C203 X2.X1.X1.X1.X2.X2.vout X2.X1.X1.X1.X2.X2.X3.vin1 0.335f
C204 a_33976_18540# a_33676_16634# 6.2e-19
C205 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X2.X3.vin1 0.0174f
C206 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.X3.vin1 1.22e-19
C207 d3 X1.X2.X2.X2.X1.X2.X3.vin1 2.1e-19
C208 X2.X1.X1.X2.X1.X2.vout d1 0.033f
C209 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin2 0.12f
C210 a_34362_26164# d4 6.91e-19
C211 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X3.vin2 0.449f
C212 a_8186_10734# a_8572_10734# 0.414f
C213 a_10686_23170# X1.X1.X2.X2.X1.X2.vrefh 8.22e-20
C214 a_22826_22210# X1.X2.X2.X2.X1.X1.X3.vin2 0.00815f
C215 d2 a_8572_10734# 0.0057f
C216 a_17222_27070# d2 0.00792f
C217 a_54992_19358# a_54992_17452# 0.00396f
C218 d0 a_43362_892# 1.37e-19
C219 X1.X2.X1.X1.X1.X2.X3.vin2 d1 0.171f
C220 X1.X1.X2.X2.X2.X1.vout a_8872_27888# 0.359f
C221 X2.X1.X3.vin1 a_37766_8828# 8.66e-20
C222 d0 X2.X1.X2.X1.X2.X1.X2.vin1 0.262f
C223 a_25326_9828# vdd 0.542f
C224 X1.X1.X3.vin1 X1.X1.X2.X1.X1.X2.vout 1.71e-19
C225 a_23212_18358# X1.X2.X2.X1.X2.X2.vout 7.93e-20
C226 a_34062_16634# X2.X1.X1.X2.X1.X1.X3.vin2 0.267f
C227 a_46502_9916# a_46502_8010# 0.00198f
C228 a_17222_6104# X1.X2.X1.X2.X2.X2.X1.vin2 0.273f
C229 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin1 0.52f
C230 X2.X2.X1.X1.X1.X2.X1.vin1 d0 0.267f
C231 d2 X1.X2.X1.X1.X1.X1.vout 0.0904f
C232 a_10686_25076# a_10686_23170# 0.00198f
C233 d3 X1.X1.X3.vin1 0.834f
C234 d3 a_23126_12640# 0.00195f
C235 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X3.vin2 0.0523f
C236 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 0.242f
C237 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X3.vin1 0.00118f
C238 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X3.vin2 0.17f
C239 a_31476_21352# vdd 1.05f
C240 X2.X2.X3.vin1 a_52106_10734# 3.93e-19
C241 a_2582_19446# a_4696_18540# 4.72e-20
C242 X1.X2.X2.X2.X2.X2.X2.vin1 X2.vrefh 0.597f
C243 X1.X2.X2.X2.X2.X2.X3.vin2 a_25712_32700# 0.354f
C244 d0 X2.X2.X1.X2.X1.X1.X1.vin2 0.276f
C245 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X3.vin2 0.552f
C246 X1.X3.vin1 a_13696_892# 0.195f
C247 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X3.vin2 0.161f
C248 a_46502_4198# vdd 0.541f
C249 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 5.19e-19
C250 a_19336_26164# vdd 1.05f
C251 d0 X2.X1.X1.X2.X1.X1.X3.vin1 4.36e-19
C252 X1.X2.X1.X2.X1.X2.X3.vin1 a_17222_11822# 0.00207f
C253 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X1.vin1 0.206f
C254 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X3.vin1 0.206f
C255 X2.X2.X2.X2.X2.X2.X3.vin2 vdd 0.738f
C256 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.vrefh 2.33e-19
C257 d3 X1.X1.X2.X1.X2.X1.X3.vin1 0.0195f
C258 a_8572_18358# a_8486_16452# 3.3e-19
C259 X2.X2.X2.X2.X1.X1.vout vdd 0.78f
C260 d1 X2.X1.X2.X1.X1.X2.vrefh 0.0738f
C261 a_46502_17540# X2.X2.X1.X2.X1.X1.X2.vin1 8.88e-20
C262 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X2.vrefh 0.267f
C263 X2.X2.X3.vin1 a_48702_5198# 2.12e-19
C264 X1.X1.X2.X2.X2.X2.X1.vin2 a_10686_30794# 0.273f
C265 X1.X2.X1.X2.X1.X1.X2.vin1 a_17222_15634# 0.402f
C266 X2.X2.X1.X1.X2.X1.X2.vin1 d2 0.0318f
C267 X1.X2.X1.X3.vin1 X1.X2.X3.vin2 7.53e-21
C268 a_4696_14688# X1.X1.X1.X2.X1.X2.vout 0.0929f
C269 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 0.581f
C270 a_10686_11734# a_10686_9828# 0.00198f
C271 X1.X2.X2.X3.vin1 X1.X2.X1.X2.X3.vin2 7.46e-20
C272 a_49002_29936# vdd 0.477f
C273 d3 X2.X2.X2.X3.vin2 0.481f
C274 X2.X1.X2.vrefh X3.vin2 3.04e-19
C275 a_52406_20264# X2.X2.X2.X2.X1.X1.X3.vin1 0.428f
C276 a_8186_14586# vdd 0.567f
C277 a_52492_6962# d2 0.625f
C278 X1.X1.X3.vin1 X1.X1.X2.vrefh 0.178f
C279 a_10686_25076# X1.X1.X2.X2.X1.X2.X2.vin1 0.402f
C280 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.vrefh 0.1f
C281 X2.X1.X1.X1.X1.X1.X1.vin2 a_33676_31882# 0.00113f
C282 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin1 0.195f
C283 d3 a_4782_16634# 4.67e-19
C284 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X3.vin2 0.161f
C285 a_38152_24076# a_37852_22210# 6.71e-19
C286 a_19722_18540# X1.X2.X1.X2.X1.X1.X3.vin1 0.00837f
C287 a_16836_23258# X1.X2.X1.X1.X2.X2.X1.vin1 1.64e-19
C288 a_17222_23258# a_17222_21352# 0.00198f
C289 a_37766_16452# a_37466_14586# 5.55e-20
C290 X1.X2.X1.X3.vin2 a_19722_14688# 0.00292f
C291 a_17222_4198# vdd 0.541f
C292 d4 X2.X1.X2.X1.X2.X2.X3.vin1 2.52e-19
C293 a_19722_7064# X1.X2.X1.X2.X2.X2.vout 0.263f
C294 X2.X2.X1.X1.X1.X2.X2.vin1 X2.X2.X1.X1.X1.X2.X3.vin2 0.234f
C295 a_48316_28070# a_48702_28070# 0.419f
C296 X2.X2.X2.X2.X1.X2.X3.vin1 d0 4.36e-19
C297 X1.X2.X1.X2.X1.X1.X3.vin2 d1 0.15f
C298 a_25712_17452# a_25712_15546# 0.00396f
C299 a_8872_12640# a_8572_10734# 6.2e-19
C300 X1.X1.X1.X1.X1.X1.X3.vin1 d1 0.0296f
C301 X2.X1.X2.X3.vin1 vdd 1.26f
C302 d0 X2.X1.X1.X2.X1.X2.X2.vin1 0.262f
C303 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.vrefh 2.33e-19
C304 d0 X2.X2.X2.X1.X1.X2.X1.vin2 0.276f
C305 d3 a_5082_26164# 0.284f
C306 a_40352_23170# d0 0.518f
C307 a_19336_14688# a_19036_12822# 6.71e-19
C308 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin2 7.84e-19
C309 d2 X2.X1.X1.X2.X2.X1.vout 0.0909f
C310 X1.X2.X3.vin2 d0 0.034f
C311 a_31862_13728# d1 3.41e-19
C312 X2.X1.X1.X2.X2.X2.X3.vin1 a_31862_4198# 0.00207f
C313 X1.X1.X2.X1.X2.X2.vout d1 0.033f
C314 X2.X1.X3.vin1 X2.X1.X1.X3.vin2 1.04f
C315 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin1 0.267f
C316 d2 a_46116_13728# 0.00351f
C317 a_38152_27888# a_37852_25982# 6.2e-19
C318 X2.X1.X1.X1.X2.X2.X2.vin1 X2.X1.X1.X2.vrefh 0.564f
C319 a_37766_20264# X2.X1.X2.X2.X1.X1.X3.vin1 0.428f
C320 X1.X2.X2.X1.X2.X1.X1.vin2 a_25712_11734# 0.12f
C321 a_25326_11734# X1.X2.X2.X1.X2.X1.X1.vin1 0.417f
C322 X2.X1.X2.X2.X2.X1.X2.vin1 d1 1.03e-19
C323 d3 X2.X1.X1.X1.X3.vin1 0.088f
C324 X1.X2.X1.X2.X2.X1.X3.vin2 d1 0.15f
C325 a_31476_23258# a_31862_23258# 0.419f
C326 d2 a_54606_28888# 0.00665f
C327 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X1.X2.X1.X2.X2.X1.vin1 0.668f
C328 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X1.vin1 5.19e-19
C329 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X1.vin2 0.668f
C330 X2.X2.X2.X2.X3.vin1 d4 8.41e-19
C331 a_34062_31882# X2.X1.X1.X1.X1.X1.X3.vin2 0.267f
C332 a_40352_17452# d1 2.92e-22
C333 a_4696_22312# a_4782_20446# 3.38e-19
C334 a_16836_15634# vdd 1.05f
C335 a_5082_22312# a_4396_20446# 3.31e-19
C336 a_52106_6962# a_52492_6962# 0.419f
C337 d2 X2.X1.X1.X2.X3.vin2 0.0501f
C338 X1.X2.X2.X2.X2.X1.X3.vin2 X1.X2.X2.X2.X2.X2.X1.vin1 5.19e-19
C339 a_8186_18358# a_8572_18358# 0.416f
C340 X1.X2.X2.X1.X2.X2.X3.vin2 d1 0.151f
C341 X2.X2.X2.X2.X1.X2.vrefh a_54606_21264# 0.3f
C342 X1.X2.X2.X1.X1.X1.X2.vin1 vdd 0.578f
C343 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X2.vrefh 0.076f
C344 d2 X2.X1.X2.X1.X2.X2.X2.vin1 0.0314f
C345 a_46502_8010# X2.X2.X1.X2.X2.X2.X1.vin1 8.22e-20
C346 X1.X2.X1.X1.X2.X1.X1.vin1 vdd 0.592f
C347 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X1.vin1 0.0689f
C348 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X1.vin1 0.0689f
C349 X1.X2.X1.X1.X1.X1.X3.vin2 d1 0.152f
C350 X2.X1.X2.X2.X1.X2.X3.vin2 a_39966_23170# 7.84e-19
C351 X2.X1.X2.X1.X2.X1.X3.vin2 a_39966_11734# 7.84e-19
C352 X2.X1.X1.X3.vin1 X2.X1.X2.X2.X3.vin2 7.46e-20
C353 d1 a_31476_4198# 2.81e-20
C354 X1.X1.X2.X2.X3.vin2 a_8486_27888# 0.00101f
C355 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X2.vin1 0.0689f
C356 a_46502_21352# a_48316_20446# 1.06e-19
C357 X2.X1.X2.X1.X2.X1.vout a_37852_14586# 0.169f
C358 X1.X1.X1.X1.X1.X2.X3.vin2 vdd 0.787f
C359 d1 X2.X1.X2.vrefh 0.258f
C360 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X1.vin2 0.668f
C361 d0 X1.X1.X1.X2.X1.X2.vrefh 0.844f
C362 d3 a_8872_24076# 0.00108f
C363 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.X1.vin1 0.206f
C364 X1.X2.X2.X2.X2.X1.X3.vin1 a_25326_26982# 0.52f
C365 X1.X1.X1.X2.X3.vin1 d1 0.00179f
C366 a_46502_19446# X2.X2.X1.X2.X1.X1.X1.vin1 8.22e-20
C367 X1.X2.X1.X1.X2.X2.X2.vin1 X1.X2.X1.X2.vrefh 0.564f
C368 X2.X1.X2.X2.X2.X1.X1.vin2 d0 0.276f
C369 X1.X2.X1.X2.X3.vin1 a_19336_10916# 0.17f
C370 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin2 7.84e-19
C371 a_23126_20264# X1.X2.X2.X2.X1.X1.X3.vin1 0.428f
C372 d0 X1.X2.X1.X2.X1.X2.X1.vin2 0.276f
C373 X1.X2.X1.X1.X1.X2.X2.vin1 d2 0.0329f
C374 X1.X2.X1.X1.X1.X1.X2.vin1 a_17222_30882# 0.402f
C375 X1.X1.X2.X2.X2.X2.vout d1 0.033f
C376 X1.X2.X2.X2.X1.X2.X1.vin2 X1.X2.X2.X2.X1.X2.X1.vin1 0.668f
C377 a_37466_25982# vdd 0.487f
C378 a_46502_9916# a_48316_9010# 1.06e-19
C379 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 5.19e-19
C380 a_8486_20264# a_8572_18358# 3.21e-19
C381 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X2.vin1 0.0689f
C382 d0 X1.X1.X1.X2.X1.X2.X3.vin1 4.36e-19
C383 a_31476_28976# d0 0.518f
C384 X2.X1.X2.X2.X1.X1.X3.vin2 a_37766_20264# 0.267f
C385 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X3.vin1 0.00117f
C386 a_2582_27070# X1.X1.X1.X1.X1.X2.X3.vin1 0.00207f
C387 d5 a_20286_892# 0.506f
C388 X1.X1.X1.X2.X1.X2.X3.vin2 a_2196_11822# 0.354f
C389 d2 a_19336_29936# 0.606f
C390 a_4782_12822# a_2582_11822# 4.77e-21
C391 d2 a_8486_31700# 0.00166f
C392 d3 X1.X2.X1.X1.X1.X1.X1.vin2 1.14e-19
C393 X1.X2.X1.X1.X2.X1.X1.vin2 a_17222_23258# 8.88e-20
C394 a_54606_17452# a_52406_16452# 4.77e-21
C395 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X3.vin1 0.0131f
C396 a_48702_12822# a_46502_11822# 4.77e-21
C397 X1.X2.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X2.X2.vrefh 0.117f
C398 X2.X2.X1.X2.X1.X2.X3.vin2 a_46116_11822# 0.354f
C399 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin2 0.12f
C400 a_16836_30882# vdd 1.05f
C401 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X3.vin2 0.161f
C402 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X2.X1.X1.X1.vin1 0.206f
C403 X2.X2.X2.X2.X1.X2.vout X2.X2.X2.X2.X1.X1.vout 0.507f
C404 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X2.vrefh 0.076f
C405 X1.X2.X2.X1.X2.X1.X3.vin2 a_23512_12640# 0.1f
C406 d1 a_2582_4198# 0.00148f
C407 a_33976_14688# vdd 1.05f
C408 X2.X1.X2.X1.X1.X2.X3.vin2 a_40352_9828# 0.354f
C409 a_17222_13728# a_19422_12822# 4.2e-20
C410 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X2.vin1 0.00117f
C411 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X3.vin1 0.206f
C412 X1.X2.X1.X1.X2.X2.vout vdd 0.865f
C413 a_33976_14688# a_34062_12822# 3.38e-19
C414 a_34362_14688# a_33676_12822# 3.31e-19
C415 X2.X1.X1.X3.vin1 a_34062_24258# 5.28e-19
C416 a_11072_26982# d0 0.518f
C417 X1.X2.X2.X2.X1.X2.vrefh d2 0.177f
C418 X2.X1.X1.X2.X2.X2.vout a_33676_5198# 0.36f
C419 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin2 7.84e-19
C420 a_34362_7064# a_34062_5198# 5.55e-20
C421 X1.X1.X1.X2.X2.X2.X3.vin1 a_4396_5198# 0.199f
C422 X1.X2.X2.X1.X1.X2.X1.vin2 a_25326_7922# 0.273f
C423 X1.X1.X3.vin2 a_5082_10916# 3.68e-19
C424 a_52106_10734# X2.X2.X2.X1.X1.X2.X3.vin2 0.00846f
C425 X1.X1.X1.X1.X1.X2.vrefh d0 0.844f
C426 a_8186_18358# d2 0.00146f
C427 X1.X2.X2.X2.X1.X1.X1.vin2 X1.X2.X2.X1.X2.X2.X3.vin2 3.94e-19
C428 X1.X2.X2.X2.X1.X1.X1.vin1 a_25326_17452# 8.22e-20
C429 X2.X1.X2.X1.X2.X1.X1.vin2 vdd 0.36f
C430 X1.X1.X2.X2.X2.X1.vout X1.X1.X2.X2.X2.X2.vout 0.514f
C431 a_2582_17540# vdd 0.553f
C432 a_10686_11734# a_8572_10734# 5.36e-21
C433 d3 X1.X2.X2.X2.X3.vin1 0.375f
C434 d1 X2.X1.X1.X2.X2.X1.X3.vin2 0.15f
C435 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X1.X3.vin2 3.94e-19
C436 a_46502_21352# X2.X2.X1.X1.X2.X2.X1.vin2 0.273f
C437 X2.X2.X2.X2.X2.X1.X3.vin1 a_54606_28888# 0.00207f
C438 d3 X1.X2.X2.X1.X3.vin1 0.0869f
C439 X2.X1.X1.X2.X1.X1.vout X2.X1.X1.X2.X3.vin1 0.131f
C440 a_8872_20264# d1 0.521f
C441 X1.X3.vin2 vdd 0.665f
C442 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X1.X2.X2.X2.X2.X1.vin1 0.668f
C443 X2.X1.X1.X2.vrefh d0 0.848f
C444 d5 a_49952_892# 0.0319f
C445 a_48702_16634# a_46502_15634# 4.77e-21
C446 a_10686_21264# X1.X1.X2.X2.X1.X1.X3.vin1 0.00207f
C447 X2.X2.X1.X1.X2.X1.vout X2.X2.X1.X1.X2.X1.X3.vin2 0.326f
C448 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X3.vin2 0.234f
C449 X1.X1.X2.X1.X2.X2.X1.vin2 d1 2.18e-19
C450 a_11072_6016# vdd 1.05f
C451 a_39966_15546# vdd 0.553f
C452 X1.X1.X3.vin1 a_5082_14688# 3.28e-19
C453 X2.X2.X1.X2.X2.X2.vrefh vdd 0.415f
C454 X1.X1.X1.X2.X2.X2.X3.vin1 a_4696_7064# 0.00329f
C455 d3 a_19722_14688# 0.0469f
C456 a_33976_26164# X2.X1.X1.X1.X3.vin2 0.0927f
C457 a_11072_13640# d1 2.92e-22
C458 a_31862_28976# X2.X1.X1.X1.X1.X2.vrefh 8.22e-20
C459 X1.X2.X1.X2.vrefh d0 0.848f
C460 X2.X1.X1.X3.vin1 d1 0.00955f
C461 a_37466_10734# d1 0.0318f
C462 a_11072_11734# vdd 1.05f
C463 a_31862_32788# d0 0.0394f
C464 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X2.vin1 0.0689f
C465 a_54606_17452# X2.X2.X2.X1.X2.X2.X3.vin2 0.567f
C466 a_31862_6104# a_33676_5198# 1.06e-19
C467 X1.X2.X1.X1.X1.X2.X1.vin2 d1 0.00406f
C468 X2.X1.X2.X2.X1.X2.X3.vin1 a_40352_23170# 0.354f
C469 a_31476_8010# vdd 1.05f
C470 X1.X1.X2.X1.X1.X2.X1.vin2 d1 0.00406f
C471 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X2.vrefh 0.0763f
C472 a_25326_23170# vdd 0.553f
C473 X2.X2.X2.X2.X1.X1.X3.vin2 X2.X2.X2.X2.X1.X1.X1.vin1 2.23e-19
C474 X1.X2.X1.X1.X2.X2.vrefh a_16836_23258# 0.118f
C475 X2.X2.X2.X2.X1.X1.X2.vin1 a_54992_19358# 1.78e-19
C476 X1.X1.X3.vin1 a_5646_892# 0.17f
C477 d2 X1.X1.X2.X1.X2.X1.X2.vin1 0.0318f
C478 d0 a_54992_9828# 0.515f
C479 a_52492_6962# a_52792_8828# 6.71e-19
C480 a_23212_14586# X1.X2.X2.X1.X2.X1.X3.vin2 0.00546f
C481 a_25326_26982# X1.X2.X2.X2.X2.X1.X3.vin2 7.84e-19
C482 d3 X2.X2.X3.vin1 0.834f
C483 d3 X2.X1.X1.X2.X2.vrefh 6.65e-20
C484 X1.X1.X1.X1.X1.X2.X3.vin1 d1 0.146f
C485 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.X1.X2.vin1 0.0689f
C486 a_33676_24258# a_31862_23258# 1.15e-20
C487 a_2196_6104# X1.X1.X1.X2.X2.X2.vrefh 1.64e-19
C488 X1.X1.X1.X2.X2.X2.X3.vin2 X1.X1.X2.vrefh 0.172f
C489 d0 X2.X1.X2.X1.X1.X2.X3.vin2 4.34e-19
C490 X2.X2.X2.X2.X1.X2.X1.vin1 a_54992_21264# 1.64e-19
C491 X1.X1.X2.X1.X2.X2.X3.vin2 a_10686_15546# 7.84e-19
C492 X1.X1.X1.X1.X2.X2.X3.vin2 a_2582_17540# 8.07e-19
C493 d2 X1.X2.X1.X1.X1.X2.X1.vin1 0.0114f
C494 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X1.vin1 0.0689f
C495 X1.X2.X2.X1.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin2 0.0128f
C496 a_48702_9010# X2.X2.X1.X2.X2.X1.X3.vin2 0.267f
C497 X1.X1.X1.X1.X1.X1.X3.vin1 a_4396_31882# 0.199f
C498 a_19036_16634# vdd 1.05f
C499 a_5082_10916# X1.X1.X1.X2.X3.vin2 0.263f
C500 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin1 0.267f
C501 X2.X1.X2.X2.X1.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin2 0.0128f
C502 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X2.vrefh 0.00118f
C503 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X1.vout 0.131f
C504 a_19036_20446# a_19336_18540# 6.48e-19
C505 a_52792_27888# vdd 1.05f
C506 a_2196_25164# vdd 1.05f
C507 d2 X1.X2.X1.X2.X1.X1.X1.vin2 0.231f
C508 d3 X1.X1.X2.X1.X2.vrefh 6.65e-20
C509 X1.X1.X2.X2.X2.X2.X1.vin2 d1 0.0985f
C510 X2.X2.X1.X1.X2.X2.X1.vin1 d0 0.267f
C511 a_48616_22312# a_49002_22312# 0.419f
C512 X1.X2.X1.X1.X1.X2.vrefh X1.X1.X2.X2.X2.X2.vrefh 0.117f
C513 X1.X1.X1.X2.X1.X1.vout a_4696_14688# 0.169f
C514 a_4782_16634# a_5082_14688# 4.19e-20
C515 a_39966_30794# vdd 0.553f
C516 d4 a_46502_32788# 8.99e-20
C517 a_54606_25076# X2.X2.X2.X2.X1.X2.X3.vin2 0.567f
C518 a_54606_9828# X2.X2.X2.X1.X1.X2.X3.vin1 0.00207f
C519 a_52406_20264# d1 0.0749f
C520 d2 a_37466_29834# 0.273f
C521 X1.X1.X1.X2.X1.X1.X3.vin2 vdd 0.905f
C522 d2 a_38152_5016# 0.00251f
C523 a_46502_15634# d1 0.00148f
C524 a_49002_26164# a_48702_24258# 5.25e-20
C525 X1.X2.X2.X1.X2.X1.vout X1.X2.X2.X1.X3.vin2 0.399f
C526 a_49002_14688# a_48702_12822# 5.55e-20
C527 a_48616_26164# X2.X2.X1.X1.X2.X1.vout 1.64e-19
C528 X2.X2.X1.X1.X2.X2.vrefh d1 0.0124f
C529 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.X1.vin1 0.206f
C530 d1 a_19722_7064# 0.0422f
C531 a_8186_22210# d4 1.54e-19
C532 X2.X2.X2.X1.X2.X2.X2.vin1 vdd 0.576f
C533 a_19036_9010# vdd 1.05f
C534 a_52106_14586# vdd 0.567f
C535 a_17222_17540# X1.X2.X1.X2.X1.X1.X1.vin2 0.273f
C536 a_37466_29834# a_37852_29834# 0.419f
C537 X2.X1.X1.X2.X2.X1.X2.vin1 a_31862_8010# 0.402f
C538 a_23126_27888# a_23212_29834# 3.14e-19
C539 a_31476_21352# X2.X1.X1.X1.X2.X2.X2.vin1 1.78e-19
C540 d4 X1.X1.X2.X1.X2.X2.X2.vin1 8.68e-20
C541 X1.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.vout 0.0866f
C542 X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.vout 4.93e-20
C543 X1.X1.X1.X1.X3.vin2 vdd 1.32f
C544 a_19722_26164# a_19036_24258# 2.97e-19
C545 a_37766_20264# d1 0.0749f
C546 a_25326_11734# d1 3.95e-19
C547 a_19336_26164# a_19422_24258# 3.21e-19
C548 a_52406_24076# a_52492_22210# 3.38e-19
C549 X2.X1.X2.X1.X1.X2.X3.vin2 a_38152_8828# 0.101f
C550 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X2.vrefh 0.076f
C551 X2.X2.X2.X1.X2.X1.X3.vin1 a_52792_12640# 0.199f
C552 X1.X1.X1.X2.vrefh a_2196_19446# 0.118f
C553 a_31476_23258# d1 2.92e-22
C554 a_52406_20264# a_54606_19358# 4.2e-20
C555 a_31476_19446# a_31476_17540# 0.00396f
C556 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 0.216f
C557 X2.X2.X2.X2.vrefh d0 0.844f
C558 X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X1.vin1 0.142f
C559 X1.X2.X1.X1.X2.vrefh vdd 0.426f
C560 X2.X2.X1.X2.X1.X1.vout a_49002_14688# 0.387f
C561 a_48702_16634# X2.X2.X1.X2.X3.vin1 1.52e-19
C562 a_40352_32700# vdd 1.05f
C563 a_31862_19446# d4 1.89e-19
C564 a_33976_18540# d2 0.0111f
C565 a_19036_31882# vdd 1.05f
C566 X1.X2.X1.X3.vin1 a_19722_18540# 0.389f
C567 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin2 0.12f
C568 X2.X2.X2.X2.X1.X2.X1.vin1 a_54992_23170# 0.195f
C569 a_39966_17452# X2.X1.X2.X1.X2.X2.X1.vin2 8.88e-20
C570 a_48702_31882# a_46502_30882# 4.77e-21
C571 d0 X2.X2.X2.X1.X2.X1.X3.vin1 4.36e-19
C572 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.vout 0.197f
C573 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 0.139f
C574 a_23126_20264# d1 0.0749f
C575 a_25326_21264# a_23126_20264# 4.77e-21
C576 d3 a_49002_26164# 0.284f
C577 a_25326_9828# X1.X2.X2.X1.X1.X2.X3.vin2 0.567f
C578 d3 X1.X2.X1.X2.X1.X2.X3.vin1 2.1e-19
C579 X2.X2.X2.X1.X2.X2.vrefh vdd 0.415f
C580 a_52406_20264# X2.X2.X3.vin2 7.93e-20
C581 a_48616_7064# vdd 1.05f
C582 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X1.vin2 0.076f
C583 X1.X2.X1.X2.X2.X1.X3.vin1 a_17222_8010# 0.00207f
C584 X2.X1.X2.X1.X2.X1.X3.vin2 a_40352_13640# 0.354f
C585 a_17222_19446# d4 1.89e-19
C586 X1.X1.X2.X2.X3.vin2 a_8486_31700# 9.7e-20
C587 X2.X1.X1.X1.X1.X1.X1.vin2 d2 1.68e-19
C588 a_33976_26164# a_31862_25164# 5.36e-21
C589 X1.X1.X1.X1.X1.X1.X3.vin2 vdd 0.939f
C590 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X1.X3.vin2 0.0943f
C591 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.X1.X1.vin2 3.94e-19
C592 a_46502_30882# d1 0.00148f
C593 a_28096_892# vdd 1.05f
C594 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X2.X1.X1.X2.vrefh 0.0128f
C595 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X2.vin1 0.0689f
C596 X1.X2.X2.X1.X2.X1.vout a_23126_12640# 0.422f
C597 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X3.vin1 0.206f
C598 a_4696_10916# X1.X1.X1.X2.X2.X1.vout 1.64e-19
C599 a_5082_10916# a_4782_9010# 5.25e-20
C600 a_2582_13728# a_4396_12822# 1.06e-19
C601 X2.X1.X3.vin1 X2.X1.X2.X1.X1.X1.vout 5.53e-20
C602 X1.X2.X1.X1.X2.X1.X2.vin1 d0 0.262f
C603 X2.X1.X1.X2.X2.X1.X1.vin1 d1 0.0118f
C604 a_20286_892# a_20672_892# 0.406f
C605 a_34062_12822# vdd 0.47f
C606 d1 X1.X2.X2.X1.X1.X2.X1.vin2 0.00406f
C607 X1.X1.X1.X1.X2.X1.X3.vin2 a_4696_22312# 0.00546f
C608 a_46502_30882# X2.X2.X1.X1.X1.X1.X3.vin1 0.00207f
C609 X2.X2.X2.X1.X1.X2.X1.vin1 vdd 0.592f
C610 d3 X2.X1.X2.X1.X2.X1.vout 0.00226f
C611 d2 a_46502_9916# 0.00328f
C612 X1.X1.X3.vin2 X1.X1.X2.X1.X2.X2.X3.vin2 0.0011f
C613 X2.X2.X1.X1.X1.X2.X3.vin1 X2.X2.X1.X1.X1.X2.X1.vin2 0.216f
C614 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X1.X2.X1.X2.X2.vrefh 0.1f
C615 a_33676_12822# X2.X1.X1.X2.X1.X2.X3.vin2 0.101f
C616 a_2582_19446# d4 1.89e-19
C617 X1.X2.X1.X1.X1.X1.X1.vin1 d4 0.00332f
C618 d3 a_34362_22312# 9.23e-19
C619 a_48316_16634# a_48702_16634# 0.419f
C620 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin1 0.195f
C621 X2.X1.X2.X2.X1.X1.X2.vin1 d1 1.03e-19
C622 a_54606_7922# a_54992_7922# 0.419f
C623 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X2.vrefh 0.00118f
C624 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X1.X3.vin1 0.581f
C625 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X2.vrefh 2.33e-19
C626 a_54606_21264# d2 0.0059f
C627 X1.X2.X1.X2.X1.X1.X3.vin1 a_19036_16634# 0.199f
C628 d2 a_2196_15634# 0.00414f
C629 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X2.vrefh 0.564f
C630 a_54606_25076# d0 0.0489f
C631 a_2582_9916# a_2582_8010# 0.00198f
C632 X1.X1.X1.X2.X1.X2.vout a_4782_12822# 0.418f
C633 X1.X2.X1.X2.X1.X1.X3.vin2 a_19336_14688# 0.00546f
C634 X1.X1.X1.X2.X2.X2.X1.vin2 a_2582_4198# 8.88e-20
C635 a_54992_21264# X2.X2.X2.X2.X1.X1.X1.vin2 1.78e-19
C636 a_8486_8828# a_8186_6962# 5.55e-20
C637 X2.X2.X1.X2.X3.vin1 d1 0.00179f
C638 X1.X2.X2.X2.X2.X1.X1.vin1 X2.X1.X1.X1.X2.vrefh 0.00437f
C639 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 5.19e-19
C640 a_23212_25982# d2 0.0057f
C641 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.X1.X3.vin1 0.206f
C642 a_5082_10916# d1 0.0316f
C643 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X2.X1.X2.X1.X1.X1.vin2 0.00232f
C644 a_19336_26164# X1.X2.X1.X3.vin1 0.356f
C645 a_46116_17540# a_46502_17540# 0.419f
C646 X2.X2.X2.vrefh a_54606_4110# 4.89e-19
C647 X2.X1.X2.X2.X2.X1.X3.vin1 d2 0.104f
C648 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.X3.vin1 0.587f
C649 a_48616_22312# d1 0.00613f
C650 X1.X1.X2.X1.X1.X1.X3.vin1 a_8872_5016# 0.199f
C651 X1.X2.vrefh vdd 0.419f
C652 a_33676_9010# vdd 1.05f
C653 d2 a_2196_8010# 0.00464f
C654 X1.X1.X1.X1.X2.X2.X3.vin2 vdd 0.761f
C655 a_16836_28976# a_16836_30882# 0.00396f
C656 d0 a_25326_9828# 0.0489f
C657 X1.X2.X1.X1.X2.X1.X3.vin1 a_19036_24258# 0.199f
C658 a_33676_24258# a_34062_24258# 0.419f
C659 a_46502_23258# a_46502_21352# 0.00198f
C660 a_10686_17452# a_8872_16452# 1.15e-20
C661 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X3.vin2 0.161f
C662 a_46116_23258# X2.X2.X1.X1.X2.X2.X1.vin1 1.64e-19
C663 a_37466_29834# a_38152_31700# 3.31e-19
C664 d2 a_2196_28976# 0.00351f
C665 X2.X1.X1.X1.X1.X2.vout X2.X1.X1.X1.X1.X2.X3.vin1 0.326f
C666 a_34362_26164# X2.X1.X1.X1.X3.vin1 0.385f
C667 X2.X2.X1.X2.X1.X2.X2.vin1 d1 1.03e-19
C668 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 0.242f
C669 a_39966_13640# a_37766_12640# 4.77e-21
C670 X2.X1.X2.X2.X2.X1.X1.vin1 vdd 0.592f
C671 a_39966_21264# a_39966_19358# 0.00198f
C672 d3 X1.X1.X1.X1.X2.X1.vout 0.00226f
C673 X2.X2.X2.X2.X1.X2.X1.vin1 d1 0.0118f
C674 X1.X2.X2.X1.X2.X1.X2.vin1 vdd 0.576f
C675 X2.X1.X2.X2.vrefh a_40352_17452# 0.118f
C676 X1.X2.X2.X2.X2.X2.X2.vin1 X2.X1.X1.X1.X1.X1.X1.vin2 0.00232f
C677 X1.X1.X2.X3.vin2 a_8186_22210# 0.00292f
C678 a_54992_17452# a_54992_15546# 0.00396f
C679 a_4396_9010# a_4782_9010# 0.419f
C680 d2 X2.X2.X1.X2.X2.vrefh 0.158f
C681 a_31476_21352# d0 0.518f
C682 a_46116_25164# a_46502_25164# 0.419f
C683 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X2.X1.X1.X2.X1.X1.vin2 0.00232f
C684 X2.X1.X1.X1.X1.X2.X1.vin1 vdd 0.592f
C685 X2.X1.X1.X2.X2.X2.vrefh X1.X2.X2.X1.X1.X2.vrefh 0.117f
C686 a_23212_25982# X1.X2.X2.X2.X1.X2.vout 7.93e-20
C687 d0 a_46502_4198# 0.049f
C688 a_37466_29834# X2.X1.X2.X2.X2.X2.X3.vin2 3.85e-19
C689 d1 a_20286_892# 4.67e-19
C690 a_33976_10916# vdd 1.05f
C691 X2.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X1.vin2 0.096f
C692 a_39966_9828# a_39966_7922# 0.00198f
C693 X2.X2.X3.vin2 X2.X2.X1.X2.X3.vin1 4.41e-19
C694 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 0.242f
C695 d0 X2.X2.X2.X2.X2.X2.X3.vin2 4.34e-19
C696 X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin2 6.26e-19
C697 d3 X2.X2.X2.X1.X1.X2.X3.vin2 0.0251f
C698 a_31476_15634# a_31476_13728# 0.00396f
C699 a_48316_16634# d1 0.521f
C700 X1.X2.X1.X2.X1.X2.X3.vin2 a_17222_9916# 8.07e-19
C701 a_52106_18358# d2 0.00146f
C702 X2.X1.X1.X2.X1.X1.X1.vin2 vdd 0.36f
C703 d2 X1.X1.X1.X1.X1.X2.vout 0.11f
C704 a_33676_12822# a_34362_10916# 3.08e-19
C705 a_34062_12822# a_33976_10916# 3.3e-19
C706 a_23212_29834# a_23126_31700# 3.38e-19
C707 X2.X2.X2.X2.X2.X1.X1.vin2 a_54992_26982# 0.12f
C708 X2.X1.X2.X2.X2.vrefh d3 6.65e-20
C709 a_54606_26982# X2.X2.X2.X2.X2.X1.X1.vin1 0.417f
C710 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X3.vin1 1.22e-19
C711 X2.X1.X2.X1.X2.X1.vout X2.X1.X2.X1.X2.X1.X3.vin1 0.118f
C712 X1.X2.X1.X2.X1.X1.X3.vin1 vdd 0.997f
C713 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X2.vin1 0.564f
C714 X1.X2.X1.X2.X1.X2.vout vdd 0.697f
C715 a_22826_29834# X1.X2.X2.X2.X3.vin2 0.422f
C716 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X3.vin1 0.00118f
C717 X1.X2.X1.X2.X1.X2.X3.vin2 d1 0.171f
C718 d2 a_17222_11822# 0.00792f
C719 a_33676_24258# d1 0.521f
C720 a_4782_5198# a_2582_4198# 4.77e-21
C721 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X1.vin2 0.076f
C722 X1.X1.X1.X2.X2.X2.X3.vin2 a_2196_4198# 0.354f
C723 a_8572_25982# a_8486_24076# 3.3e-19
C724 X1.X1.X2.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X1.vin2 8.93e-19
C725 X2.X1.X2.X1.X1.X1.X3.vin1 vdd 1.03f
C726 X2.X2.X2.X2.X2.X1.X3.vin2 X2.X2.X2.X2.X2.X2.X1.vin1 5.19e-19
C727 X1.X1.X2.X2.X1.X2.X3.vin1 d2 0.155f
C728 X1.X2.X1.X1.X2.X1.vout a_19722_22312# 0.383f
C729 X1.X1.X2.X1.X2.X1.X2.vin1 a_10686_11734# 8.88e-20
C730 a_31862_27070# d3 1.89e-19
C731 a_4396_9010# d1 0.521f
C732 d1 X2.X2.X1.X2.X2.X2.X1.vin2 0.0985f
C733 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X1.X2.X2.X2.X2.vrefh 0.1f
C734 a_46116_25164# d1 2.25e-20
C735 a_54992_25076# d2 0.00533f
C736 a_48316_31882# a_48702_31882# 0.419f
C737 d0 a_17222_4198# 0.049f
C738 d1 X2.X1.X1.X2.X2.X2.X3.vin1 0.149f
C739 X1.X2.X2.vrefh a_25326_4110# 4.89e-19
C740 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X1.vin1 5.19e-19
C741 a_16836_9916# a_17222_9916# 0.419f
C742 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X2.X1.X2.X2.X1.X1.vin2 0.00232f
C743 a_54606_26982# d1 3.95e-19
C744 d2 X2.X2.X1.X2.X2.X2.X1.vin1 9.24e-20
C745 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X3.vin2 0.449f
C746 X2.X2.X2.X2.X1.X2.vout vdd 0.697f
C747 d2 a_25326_15546# 0.00393f
C748 a_54606_6016# a_52406_5016# 4.77e-21
C749 X2.X1.X2.X2.X1.X2.X3.vin2 d2 0.121f
C750 X1.X1.X2.X1.X1.X1.vout vdd 0.78f
C751 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin2 0.12f
C752 d1 a_49952_892# 5.18e-19
C753 a_33976_10916# a_33676_9010# 6.2e-19
C754 a_19722_26164# X1.X2.X1.X1.X2.X1.X3.vin1 0.00837f
C755 a_39966_26982# a_40352_26982# 0.419f
C756 a_48316_31882# d1 0.511f
C757 a_25326_13640# X1.X2.X2.X1.X2.X1.X3.vin2 0.567f
C758 a_16836_9916# d1 2.25e-20
C759 a_19336_22312# a_19422_20446# 3.38e-19
C760 a_19722_22312# a_19036_20446# 3.31e-19
C761 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X3.vin1 0.587f
C762 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X3.vin1 0.0321f
C763 d2 a_25712_9828# 0.00533f
C764 d2 a_16836_8010# 0.00464f
C765 a_10686_28888# a_8872_27888# 1.15e-20
C766 X2.X1.X2.X2.X2.X1.X2.vin1 a_40352_28888# 0.197f
C767 a_48316_31882# X2.X2.X1.X1.X1.X1.X3.vin1 0.199f
C768 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X1.vin2 3.94e-19
C769 X1.X1.X2.X2.X2.vrefh a_10686_25076# 0.3f
C770 a_10686_26982# d3 0.00112f
C771 a_8186_10734# X1.X1.X2.X1.X1.X2.X3.vin2 0.00846f
C772 X2.X2.X1.X1.X2.X1.X1.vin2 a_46502_23258# 8.88e-20
C773 X1.X2.X1.X1.X2.X2.X1.vin2 d1 2.18e-19
C774 d2 X1.X1.X2.X1.X1.X2.X3.vin2 0.121f
C775 X1.X1.X1.X1.X1.X1.X2.vin1 d1 0.0144f
C776 X2.X1.X1.X1.X1.X1.X3.vin1 vdd 1.06f
C777 a_31862_28976# X2.X1.X1.X1.X1.X2.X3.vin1 0.52f
C778 a_2582_28976# X1.X1.X1.X1.X1.X2.X2.vin1 8.88e-20
C779 d0 a_16836_15634# 0.515f
C780 d2 a_52106_10734# 7.13e-19
C781 X1.X1.X1.X1.X2.X2.X3.vin1 d1 0.146f
C782 a_25712_26982# d1 2.25e-20
C783 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.vout 0.118f
C784 a_10686_15546# a_8572_14586# 2.68e-20
C785 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 0.587f
C786 X1.X2.X1.X1.X2.X2.X1.vin1 d2 0.0106f
C787 d1 a_52406_5016# 0.0752f
C788 a_25326_6016# a_25326_4110# 0.00198f
C789 X2.X2.X1.X1.X1.X1.X1.vin1 d1 1.51e-19
C790 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 0.242f
C791 d0 X1.X2.X2.X1.X1.X1.X2.vin1 0.262f
C792 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X1.X3.vin1 0.00789f
C793 a_46116_21352# a_46116_19446# 0.00396f
C794 X2.X2.X2.X2.X2.X2.X2.vin1 vrefl 0.597f
C795 X2.X2.X2.X2.X2.X2.X3.vin2 a_54992_32700# 0.354f
C796 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X3.vin1 0.587f
C797 X1.X2.X2.X2.X1.X1.X3.vin1 a_22826_18358# 0.00837f
C798 X1.X2.X2.X2.X2.X1.X1.vin2 X2.X1.X1.X1.X1.X2.X2.vin1 0.00232f
C799 X1.X2.X1.X1.X2.X1.X1.vin1 d0 0.267f
C800 a_48616_14688# X2.X2.X1.X2.X1.X2.vout 0.0929f
C801 d2 a_25326_30794# 6.36e-19
C802 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 0.0903f
C803 X2.X2.X3.vin2 a_49952_892# 0.239f
C804 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X2.vout 0.0898f
C805 X2.X2.X1.X2.X2.X2.X2.vin1 a_46502_4198# 0.402f
C806 d2 a_37852_14586# 0.526f
C807 X2.X2.X1.X1.X1.X1.X1.vin1 X2.X2.X1.X1.X1.X1.X3.vin1 0.206f
C808 X2.X2.X2.X2.X1.X1.X1.vin2 d1 1.49e-19
C809 d2 a_48702_5198# 0.00202f
C810 a_52406_5016# X2.X2.X2.X1.X1.X1.X3.vin1 0.428f
C811 X1.X1.X1.X1.X1.X2.X3.vin2 d0 4.34e-19
C812 X1.X1.X2.X2.X1.X1.vout d1 0.0238f
C813 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 0.139f
C814 a_23126_27888# a_25326_28888# 4.77e-21
C815 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.vrefh 2.33e-19
C816 X1.X1.X1.X1.X1.X2.vout a_4396_28070# 0.36f
C817 X2.X2.X1.X2.X3.vin2 a_49002_7064# 0.422f
C818 d6 a_43362_892# 0.0326f
C819 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.vout 0.2f
C820 X2.X2.X1.X1.X3.vin2 vdd 1.32f
C821 X1.X1.X2.X1.X2.X2.X3.vin2 d1 0.151f
C822 d3 a_48316_9010# 0.00178f
C823 X1.X2.X3.vin1 a_19422_16634# 2.92e-19
C824 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X1.X2.X1.X1.X1.X3.vin2 3.94e-19
C825 X2.X1.X2.X1.X1.X2.X1.vin1 a_39966_6016# 8.22e-20
C826 a_31476_25164# X2.X1.X1.X1.X2.X1.X2.vin1 1.78e-19
C827 X1.X1.X1.X2.X1.X2.X1.vin2 vdd 0.361f
C828 a_8186_29834# d1 0.0422f
C829 X2.X2.X2.X2.X1.X1.X1.vin2 a_54606_19358# 0.273f
C830 d2 a_34362_7064# 0.254f
C831 d1 X1.X2.X2.X1.X1.X1.X3.vin1 0.16f
C832 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X2.X3.vin1 1.22e-19
C833 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin2 7.84e-19
C834 X2.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.vrefh 0.117f
C835 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X1.vin2 0.668f
C836 a_16836_30882# d0 0.515f
C837 a_16836_28976# vdd 1.05f
C838 a_10686_23170# d1 3.41e-19
C839 X2.X2.X3.vin2 a_52406_5016# 2.33e-19
C840 a_8186_6962# a_8872_5016# 2.86e-19
C841 X2.X1.X1.X2.X2.X2.X2.vin1 a_31862_4198# 0.402f
C842 d3 a_39966_9828# 1.89e-19
C843 X1.X2.X3.vin1 a_19422_9010# 2.12e-19
C844 a_37466_22210# vdd 0.477f
C845 d2 X1.X2.X1.X2.X2.X2.X3.vin2 8.42e-19
C846 X1.X2.X1.X2.X2.X2.X3.vin1 d2 0.0577f
C847 d4 a_37852_18358# 0.63f
C848 a_33976_18540# X2.X1.X1.X2.X1.X1.X3.vin1 0.00232f
C849 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.X1.X1.X1.vin1 5.19e-19
C850 a_4696_18540# d1 0.00616f
C851 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X1.vin2 0.1f
C852 X1.X2.X1.X3.vin2 d2 4.4e-19
C853 a_2196_9916# X1.X1.X1.X2.X2.X1.X2.vin1 1.78e-19
C854 X2.X1.X1.X1.X2.X2.vout X2.X1.X1.X1.X2.X2.X3.vin2 0.08f
C855 X1.X1.X1.X2.X2.X2.vrefh a_2582_8010# 0.3f
C856 X2.X3.vin1 a_42976_892# 0.195f
C857 a_8872_8828# a_10686_7922# 1.06e-19
C858 d0 X2.X1.X2.X1.X2.X1.X1.vin2 0.276f
C859 a_38152_16452# a_37852_14586# 6.71e-19
C860 a_2582_17540# d0 0.0675f
C861 a_10686_15546# X1.X1.X2.X1.X2.X2.X1.vin1 0.417f
C862 d2 X1.X2.X1.X2.X1.X2.X2.vin1 0.0329f
C863 X1.X1.X2.X1.X2.X2.X1.vin2 a_11072_15546# 0.12f
C864 d3 a_37852_10734# 0.621f
C865 X2.X2.X1.X1.X2.X2.X2.vin1 vdd 0.576f
C866 X1.X2.X1.X1.X1.X1.X3.vin1 d1 0.0296f
C867 d2 a_39966_7922# 0.00479f
C868 a_52106_18358# a_52492_18358# 0.416f
C869 a_8186_29834# X1.X1.X2.X2.X2.X1.vout 0.383f
C870 a_52406_27888# a_52106_25982# 5.25e-20
C871 X2.X2.X1.X2.X1.X2.vrefh a_46116_15634# 0.118f
C872 X2.X1.X3.vin1 a_34062_5198# 2.12e-19
C873 X2.X1.X1.X1.X1.X2.X2.vin1 d3 8.68e-20
C874 d0 X1.X3.vin2 0.00479f
C875 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.X1.vin2 8.93e-19
C876 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.vrefh 0.161f
C877 X1.X2.X2.X2.X2.X2.X2.vin1 a_25326_30794# 8.88e-20
C878 a_19422_24258# vdd 0.561f
C879 a_19036_5198# a_17222_4198# 1.15e-20
C880 X1.X1.X2.X2.X1.X2.X2.vin1 d1 1.03e-19
C881 a_17222_6104# a_17222_4198# 0.00198f
C882 a_25712_26982# a_25712_25076# 0.00396f
C883 a_11072_15546# a_11072_13640# 0.00396f
C884 X1.X1.X2.X1.X2.X2.vout a_8872_16452# 0.36f
C885 a_11072_6016# d0 0.515f
C886 d2 a_4396_12822# 6.04e-19
C887 d0 a_39966_15546# 0.0675f
C888 a_25326_25076# d2 0.00792f
C889 a_48702_28070# d1 0.0749f
C890 a_46502_27070# d2 0.00792f
C891 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.X3.vin2 0.587f
C892 X1.X2.X2.X1.X2.X1.X1.vin2 X2.X1.X1.X2.X2.vrefh 0.0128f
C893 X2.X1.X1.X1.X2.X2.X2.vin1 vdd 0.576f
C894 d0 X2.X2.X1.X2.X2.X2.vrefh 0.848f
C895 a_8572_25982# X1.X1.X2.X2.X2.X1.X3.vin1 0.00251f
C896 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X2.X1.X2.X1.X2.X1.vin2 0.00232f
C897 a_16836_13728# a_17222_13728# 0.419f
C898 X1.X1.X2.X2.X1.X2.X1.vin2 a_11072_23170# 0.12f
C899 X1.X2.X3.vin2 d6 0.013f
C900 a_10686_23170# X1.X1.X2.X2.X1.X2.X1.vin1 0.417f
C901 X1.X1.X1.X2.X1.X1.X2.vin1 d1 1.03e-19
C902 d0 a_11072_11734# 0.518f
C903 X1.X1.X2.X2.X1.X1.X1.vin1 a_10686_17452# 8.22e-20
C904 X2.X2.X2.X2.X1.X2.X3.vin2 vdd 0.787f
C905 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X1.X2.X1.X2.X2.X3.vin2 3.94e-19
C906 a_25326_23170# d0 0.0675f
C907 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X1.X2.X3.vin1 0.587f
C908 d0 a_31476_8010# 0.515f
C909 a_10686_32700# X1.X1.X2.X2.X2.X2.X1.vin2 8.88e-20
C910 X1.X2.X1.X1.X2.X2.X2.vin1 vdd 0.576f
C911 X1.X1.X2.X2.X1.X2.vout a_8872_24076# 0.36f
C912 a_25326_28888# X1.X2.X2.X2.X2.X1.X2.vin1 0.402f
C913 a_10686_7922# X1.X1.X2.X1.X1.X2.X1.vin1 0.417f
C914 a_34362_18540# a_34062_16634# 5.25e-20
C915 a_33976_18540# X2.X1.X1.X2.X1.X1.vout 1.64e-19
C916 X1.X1.X2.X1.X1.X2.X1.vin2 a_11072_7922# 0.12f
C917 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X2.X3.vin1 0.00789f
C918 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X1.vin2 0.668f
C919 a_40352_9828# vdd 1.05f
C920 a_23512_16452# vdd 1.05f
C921 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X3.vin2 0.0523f
C922 d2 a_19722_10916# 7.13e-19
C923 a_17222_27070# a_19336_26164# 4.72e-20
C924 a_11072_23170# X1.X1.X2.X2.X1.X2.vrefh 1.64e-19
C925 a_31476_11822# a_31476_9916# 0.00396f
C926 a_8186_25982# X1.X1.X2.X2.X2.X1.X3.vin2 3.49e-19
C927 X1.X2.X2.X2.X2.X1.X1.vin2 d2 0.231f
C928 a_2196_21352# d2 0.00274f
C929 X2.X1.X1.X2.X2.vrefh a_31862_9916# 8.22e-20
C930 a_52106_22210# a_52492_22210# 0.419f
C931 X1.X2.X2.X1.X1.X2.X3.vin2 vdd 0.787f
C932 a_4696_18540# a_5082_18540# 0.413f
C933 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin2 0.12f
C934 X2.X2.X1.X2.X2.X2.vrefh a_46116_6104# 1.64e-19
C935 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X3.vin2 8.93e-19
C936 a_2196_25164# d0 0.518f
C937 X2.X2.X1.X2.X2.X1.X3.vin1 a_46502_8010# 0.00207f
C938 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X1.vin2 0.22f
C939 a_39966_30794# d0 0.0675f
C940 d3 a_8572_18358# 7.7e-20
C941 a_33976_29936# d1 0.00613f
C942 d2 X2.X2.X1.X1.X1.X2.vout 0.109f
C943 X1.X1.X2.X2.X1.X2.X3.vin2 a_10686_23170# 7.84e-19
C944 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X1.vin1 0.0689f
C945 a_52106_14586# a_52792_12640# 2.86e-19
C946 d0 X1.X1.X1.X2.X1.X1.X3.vin2 4.34e-19
C947 a_33976_14688# X2.X1.X1.X2.X3.vin1 0.363f
C948 a_46116_19446# d2 0.00441f
C949 X2.X1.X1.X1.X2.X2.X1.vin1 vdd 0.592f
C950 d2 X1.X1.X2.X1.X3.vin2 0.00194f
C951 X2.X2.X2.X1.X2.X1.X1.vin2 a_54606_11734# 0.273f
C952 X1.X1.X2.X1.X3.vin2 a_8186_10734# 0.241f
C953 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X2.vrefh 0.00118f
C954 d0 X2.X2.X2.X1.X2.X2.X2.vin1 0.262f
C955 X1.X1.X1.X1.X3.vin2 a_5082_22312# 0.423f
C956 X1.X3.vin1 X3.vin1 0.143f
C957 X2.X1.X2.X1.X2.X1.X3.vin1 a_37852_10734# 0.00251f
C958 X1.X1.X1.X2.X1.X1.X1.vin2 d2 0.231f
C959 X2.X2.X2.X1.X1.X1.X1.vin2 vdd 0.387f
C960 X1.X2.X1.X3.vin1 vdd 1.27f
C961 d3 X2.X1.X1.X1.X2.X1.X1.vin1 6.34e-20
C962 X2.X2.X2.X2.X1.X1.X3.vin1 d4 0.0194f
C963 X1.X2.X1.X1.X2.X2.vrefh d2 0.168f
C964 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin2 0.1f
C965 X2.X2.X3.vin1 a_49002_14688# 3.28e-19
C966 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.X2.vin1 0.00117f
C967 a_52106_10734# a_52792_8828# 3.08e-19
C968 d2 X2.X2.X2.X1.X2.X2.vout 0.00117f
C969 X1.X2.X2.X3.vin2 a_23212_18358# 0.0927f
C970 a_22826_18358# d1 0.0424f
C971 a_19422_16634# a_17222_15634# 4.77e-21
C972 a_46502_17540# a_48702_16634# 4.2e-20
C973 X1.X1.X2.X2.X2.X2.X1.vin2 a_11072_30794# 0.12f
C974 a_10686_30794# X1.X1.X2.X2.X2.X2.X1.vin1 0.417f
C975 d0 a_40352_32700# 0.515f
C976 X1.X2.X1.X1.X2.vrefh d0 0.848f
C977 a_25326_6016# a_25712_6016# 0.419f
C978 X1.X1.X1.X2.X3.vin2 a_4696_7064# 0.363f
C979 a_23512_31700# vdd 1.05f
C980 d2 X2.X2.X2.X1.X1.X2.vrefh 6.65e-20
C981 X2.X2.X1.X1.X2.X1.X3.vin2 a_48616_22312# 0.00546f
C982 a_10686_11734# X1.X1.X2.X1.X1.X2.X3.vin2 8.07e-19
C983 X2.X1.X2.X2.X3.vin1 a_37766_24076# 9.54e-19
C984 X2.X2.X1.X1.X1.X2.vrefh a_46116_30882# 0.118f
C985 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.vout 0.398f
C986 a_17222_25164# X1.X2.X1.X1.X2.X1.X1.vin2 0.273f
C987 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.vrefh 0.161f
C988 a_4696_18540# a_4396_16634# 6.2e-19
C989 a_2582_23258# d2 0.00665f
C990 X1.X1.X2.X1.X2.X2.X2.vin1 a_11072_17452# 0.197f
C991 X2.X1.X2.X2.X1.X1.X3.vin1 d4 0.0194f
C992 a_2582_6104# d2 6.36e-19
C993 a_52792_12640# vdd 1.05f
C994 a_5082_22312# vdd 0.567f
C995 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X3.vin2 0.234f
C996 X2.X1.X2.X2.X1.X2.vout d2 0.00124f
C997 a_2582_17540# X1.X1.X1.X2.X1.X1.X3.vin1 0.52f
C998 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X1.X2.X1.X2.X1.X1.vin1 0.668f
C999 d0 X2.X2.X2.X1.X2.X2.vrefh 0.844f
C1000 d3 X1.X1.X1.X2.X2.X1.X1.vin1 6.34e-20
C1001 X1.X1.X2.X2.X2.X2.vout a_8872_31700# 0.36f
C1002 a_54992_26982# a_54992_28888# 0.00396f
C1003 X1.X1.X1.X1.X1.X1.X3.vin2 d0 4.34e-19
C1004 d4 X1.X1.X3.vin2 0.288f
C1005 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 5.19e-19
C1006 d2 X1.X1.X2.X1.X1.X2.vout 0.106f
C1007 X1.X2.X2.X1.X1.X1.X1.vin2 vdd 0.387f
C1008 a_46116_28976# a_46116_30882# 0.00396f
C1009 X2.X1.X2.X1.X3.vin1 a_37766_8828# 9.54e-19
C1010 d0 vdd 70.3f
C1011 a_48702_28070# X2.X2.X1.X1.X1.X2.X3.vin2 0.277f
C1012 d0 a_28096_892# 2.73e-19
C1013 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin2 0.1f
C1014 X1.X1.X1.X2.X1.X2.vrefh a_2196_15634# 0.118f
C1015 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 0.0565f
C1016 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 0.216f
C1017 a_23126_8828# a_25326_7922# 4.2e-20
C1018 a_8872_24076# a_8186_22210# 3.31e-19
C1019 X1.X1.X1.X1.X2.X2.X1.vin2 a_2582_19446# 8.88e-20
C1020 a_52406_24076# a_52792_24076# 0.419f
C1021 X1.X2.X2.X2.X1.X1.X3.vin1 d4 0.0194f
C1022 d3 a_8186_10734# 0.284f
C1023 X2.X2.X1.X2.X1.X2.X1.vin2 d1 0.00406f
C1024 d3 d2 16.6f
C1025 a_19722_14688# a_19422_12822# 5.55e-20
C1026 d0 X2.X2.X2.X1.X1.X2.X1.vin1 0.267f
C1027 a_16836_32788# d2 3.9e-19
C1028 X2.X2.X1.X2.X1.X1.X2.vin1 X2.X2.X1.X2.X1.X2.vrefh 0.564f
C1029 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 0.581f
C1030 a_23126_5016# a_23512_5016# 0.419f
C1031 a_16836_19446# a_16836_17540# 0.00396f
C1032 a_48616_18540# a_48702_16634# 3.21e-19
C1033 a_37466_18358# X2.X1.X3.vin2 0.451f
C1034 a_49002_18540# a_48316_16634# 2.97e-19
C1035 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X2.X1.X1.X2.X2.vrefh 0.0128f
C1036 a_2582_15634# X1.X1.X1.X2.X1.X2.X1.vin1 8.22e-20
C1037 X2.X1.X1.X2.X1.X2.X3.vin1 d1 0.146f
C1038 a_17222_27070# X1.X2.X1.X1.X2.X1.X1.vin1 8.22e-20
C1039 d2 X2.X2.X2.X2.X2.X2.vout 0.106f
C1040 X2.X2.X1.X2.X1.X2.vout X2.X2.X1.X2.X1.X2.X3.vin1 0.326f
C1041 d2 X2.X2.X1.X2.X1.X2.X1.vin1 0.0114f
C1042 a_16836_6104# X1.X2.X1.X2.X2.X2.X2.vin1 1.78e-19
C1043 X1.X2.X1.X2.X2.vrefh vdd 0.426f
C1044 a_37766_27888# a_39966_26982# 4.2e-20
C1045 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X1.X1.vin2 0.216f
C1046 X1.X2.X2.X1.X2.X2.vout a_22826_14586# 0.263f
C1047 X1.X2.X2.X1.X2.X1.X1.vin1 a_25712_11734# 0.195f
C1048 a_39966_15546# a_40352_15546# 0.419f
C1049 d2 X2.X2.X2.X2.X2.X1.X3.vin2 0.177f
C1050 X1.X1.X1.X1.X2.X2.vrefh a_2196_23258# 0.118f
C1051 a_31862_28976# X2.X1.X1.X1.X1.X1.X3.vin2 8.07e-19
C1052 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.vout 0.075f
C1053 X2.X1.X2.X3.vin2 d2 4.4e-19
C1054 a_46502_17540# d1 3.95e-19
C1055 a_5082_22312# X1.X1.X1.X1.X2.X2.X3.vin2 3.85e-19
C1056 X1.X1.X1.X1.X2.X2.vout a_4782_20446# 0.418f
C1057 X2.X1.X2.X2.X1.X1.X3.vin2 d4 6.94e-19
C1058 a_46116_6104# vdd 1.05f
C1059 a_39966_25076# vdd 0.542f
C1060 a_4782_9010# a_4696_7064# 3.14e-19
C1061 a_4396_9010# a_5082_7064# 2.86e-19
C1062 d3 X1.X2.X2.X2.X1.X2.vout 0.0232f
C1063 d1 a_4396_5198# 0.522f
C1064 a_38152_8828# vdd 1.05f
C1065 X1.X2.X1.X1.X2.X1.X3.vin2 a_16836_23258# 0.354f
C1066 X1.X2.vrefh d0 0.0263f
C1067 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X3.vin2 0.161f
C1068 a_37852_25982# X2.X1.X2.X2.X3.vin2 0.0927f
C1069 a_52106_29834# d1 0.0422f
C1070 X1.X1.X1.X1.X2.X2.X3.vin2 d0 4.34e-19
C1071 a_8486_16452# a_8186_14586# 5.55e-20
C1072 a_23126_27888# d1 0.0749f
C1073 X2.X2.X3.vin1 a_49566_892# 0.17f
C1074 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin2 7.84e-19
C1075 X2.X2.X1.X1.X2.X2.X3.vin1 a_48316_20446# 0.199f
C1076 X2.X1.X2.X1.X1.X2.vrefh a_39966_6016# 0.3f
C1077 a_8572_14586# d1 0.00613f
C1078 X1.X2.X2.X2.X2.X1.X3.vin1 a_25712_26982# 0.354f
C1079 a_31862_32788# X2.X1.X1.X1.X1.X1.X1.vin2 0.273f
C1080 X2.X1.X2.X2.X2.X1.X1.vin1 d0 0.267f
C1081 a_10686_9828# vdd 0.542f
C1082 a_49002_22312# d4 1.99e-19
C1083 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 0.581f
C1084 d0 X1.X2.X2.X1.X2.X1.X2.vin1 0.262f
C1085 X2.X2.X1.X2.X1.X1.X3.vin2 a_46502_13728# 8.07e-19
C1086 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X3.vin2 0.552f
C1087 X1.X2.X2.X2.X1.X1.vout d2 0.00169f
C1088 a_19422_28070# d2 0.00202f
C1089 a_19422_31882# a_17222_30882# 4.77e-21
C1090 a_52106_25982# a_52406_24076# 4.41e-20
C1091 a_25326_23170# a_25712_23170# 0.419f
C1092 X2.X2.X1.X2.X2.X1.X3.vin1 a_48316_9010# 0.199f
C1093 a_10686_25076# a_8872_24076# 1.15e-20
C1094 X2.X1.X1.X1.X1.X2.X1.vin1 d0 0.267f
C1095 d5 d7 4.95e-19
C1096 d4 X2.X1.X2.X2.X3.vin2 0.0175f
C1097 a_48616_18540# d1 0.00616f
C1098 a_52792_16452# d1 0.521f
C1099 a_16836_21352# vdd 1.05f
C1100 d2 X1.X2.X1.X1.X3.vin1 0.0594f
C1101 a_39966_23170# a_39966_21264# 0.00198f
C1102 X1.X1.X2.X1.X2.vrefh a_11072_9828# 0.118f
C1103 a_2196_28976# X1.X1.X1.X1.X1.X2.vrefh 1.64e-19
C1104 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X3.vin1 0.00117f
C1105 d1 a_4696_7064# 0.00613f
C1106 d3 a_8872_12640# 0.00178f
C1107 X2.X1.X2.X2.X1.X1.X1.vin1 a_40352_17452# 1.64e-19
C1108 X2.X2.X2.X1.X2.X2.X3.vin2 a_52406_16452# 0.277f
C1109 X2.X1.X2.X3.vin1 X2.X1.X1.X2.X3.vin2 7.46e-20
C1110 d0 X2.X1.X1.X2.X1.X1.X1.vin2 0.276f
C1111 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X1.vin2 0.696f
C1112 a_54992_32700# vdd 1.05f
C1113 X1.X2.X1.X2.X1.X2.X1.vin2 a_17222_11822# 8.88e-20
C1114 X2.X2.X2.X1.X2.X2.X3.vin1 a_52106_14586# 0.00874f
C1115 X1.X2.X2.X1.X3.vin1 a_23126_5016# 1.52e-19
C1116 d1 X1.X1.X2.X1.X1.X1.X1.vin2 0.0985f
C1117 d2 X2.X1.X2.X1.X2.X1.X3.vin1 0.104f
C1118 a_37466_18358# X2.X1.X2.X1.X2.X2.X3.vin2 0.00846f
C1119 d0 X1.X2.X1.X2.X1.X1.X3.vin1 4.36e-19
C1120 X2.X1.X1.X2.X3.vin1 vdd 0.804f
C1121 X2.X2.X1.X2.X2.X2.X2.vin1 vdd 0.578f
C1122 a_4696_29936# a_2582_28976# 2.68e-20
C1123 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X3.vin2 8.93e-19
C1124 a_33976_29936# a_34362_29936# 0.419f
C1125 X1.X2.X1.X2.X1.X2.X3.vin1 a_19422_12822# 0.42f
C1126 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 2.23e-19
C1127 a_38152_24076# d1 0.521f
C1128 X2.X2.X2.X2.X2.X1.X3.vin1 d3 0.0195f
C1129 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X1.X2.X1.X2.X2.vrefh 0.1f
C1130 X1.X1.X1.X1.X1.X2.vrefh a_2196_30882# 0.118f
C1131 X1.X2.X2.X2.X1.X2.vout X1.X2.X2.X2.X1.X1.vout 0.507f
C1132 a_52406_20264# a_52792_20264# 0.419f
C1133 X2.X1.X1.X2.X3.vin1 a_34062_12822# 9.54e-19
C1134 a_34362_14688# X2.X1.X1.X2.X1.X2.X3.vin2 3.85e-19
C1135 d3 a_4396_28070# 0.00108f
C1136 d4 a_48702_16634# 0.00142f
C1137 a_19036_16634# X1.X2.X1.X2.X1.X1.vout 0.359f
C1138 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 0.587f
C1139 a_8872_8828# d1 0.521f
C1140 X2.X1.X1.X2.X2.X2.vout X2.X1.X1.X2.X2.X2.X3.vin2 0.08f
C1141 d0 X2.X1.X2.X1.X1.X1.X3.vin1 4.36e-19
C1142 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X1.vin2 0.076f
C1143 a_39966_23170# a_37852_22210# 2.68e-20
C1144 X2.X1.X2.X2.X2.X1.X1.vin1 a_39966_25076# 8.22e-20
C1145 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X1.X2.X3.vin2 3.94e-19
C1146 a_25326_7922# X1.X2.X2.X1.X1.X2.X1.vin1 0.417f
C1147 X1.X1.X2.X3.vin2 X1.X1.X3.vin2 0.171f
C1148 X1.X2.X2.X1.X1.X2.X1.vin2 a_25712_7922# 0.12f
C1149 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 2.23e-19
C1150 X2.X2.X1.X1.X1.X1.X2.vin1 X2.X2.X1.X1.X1.X2.vrefh 0.564f
C1151 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X3.vin1 0.199f
C1152 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 5.19e-19
C1153 X1.X1.X2.X1.X2.X2.vrefh a_11072_13640# 0.118f
C1154 a_4696_29936# a_2582_30882# 2.95e-20
C1155 a_2196_11822# d1 2.92e-22
C1156 X2.X1.X2.X1.X2.X1.X1.vin1 vdd 0.592f
C1157 a_46116_23258# vdd 1.05f
C1158 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin1 0.195f
C1159 X1.X1.X1.X2.X1.X1.X3.vin1 vdd 0.997f
C1160 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.vrefh 2.33e-19
C1161 a_23212_6962# vdd 1.05f
C1162 d4 X2.X1.X2.X1.X2.X2.vout 6.95e-19
C1163 a_34062_24258# d4 2.4e-19
C1164 a_52492_18358# X2.X2.X2.X1.X2.X2.vout 7.93e-20
C1165 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X1.X2.X2.X1.vin2 0.216f
C1166 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X1.X3.vin2 0.581f
C1167 a_39966_19358# a_37852_18358# 5.36e-21
C1168 a_23126_16452# d1 0.0749f
C1169 a_5082_29936# X1.X1.X1.X1.X1.X2.vout 0.254f
C1170 a_52792_31700# d1 0.515f
C1171 X2.X2.X2.X1.X2.X2.X3.vin1 vdd 0.962f
C1172 a_33676_24258# a_33976_22312# 6.1e-19
C1173 X1.X1.X1.X1.X1.X1.X1.vin2 d1 0.00147f
C1174 a_39966_30794# a_40352_30794# 0.419f
C1175 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X2.X1.vin2 0.1f
C1176 X1.X1.X2.X2.X1.X1.X3.vin2 X1.X1.X2.X2.X1.X1.X3.vin1 0.581f
C1177 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X2.vrefh 0.00118f
C1178 a_19036_5198# vdd 1.05f
C1179 a_17222_6104# vdd 0.553f
C1180 a_19036_24258# X1.X2.X1.X1.X2.X1.vout 0.359f
C1181 X1.X1.X2.X1.X2.X2.X1.vin1 d1 0.0118f
C1182 a_40352_15546# vdd 1.05f
C1183 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X2.vin1 0.564f
C1184 d1 X1.X2.X1.X2.X2.X2.vrefh 0.0124f
C1185 d3 X2.X1.X2.X2.X2.X2.X3.vin2 0.109f
C1186 X2.X1.X1.X2.X2.X2.X1.vin2 a_31862_4198# 8.88e-20
C1187 d3 X2.X1.X2.X1.X2.vrefh 6.65e-20
C1188 a_37766_20264# a_38152_20264# 0.419f
C1189 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.vout 0.335f
C1190 a_37852_25982# d1 0.0126f
C1191 X2.X1.X2.X2.X1.X2.X3.vin1 vdd 0.96f
C1192 X2.X1.X1.X1.X1.X2.X3.vin1 X2.X1.X1.X1.X1.X2.vrefh 2.33e-19
C1193 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X3.vin2 0.418f
C1194 a_17222_13728# d1 3.41e-19
C1195 a_8572_14586# a_8486_12640# 3.14e-19
C1196 a_23126_8828# d1 0.0749f
C1197 d2 a_31476_13728# 0.00351f
C1198 X2.X1.X1.X1.X1.X1.X3.vin1 d0 4.36e-19
C1199 a_19036_9010# X1.X2.X1.X2.X2.X1.vout 0.359f
C1200 a_22826_18358# X1.X2.X2.X3.vin1 0.374f
C1201 X1.X1.X2.X1.X1.X2.X3.vin1 vdd 0.96f
C1202 X1.X2.X1.X3.vin2 X1.X2.X3.vin2 3.82e-19
C1203 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin2 7.84e-19
C1204 X2.X1.X1.X2.X2.X2.X3.vin1 a_33676_5198# 0.199f
C1205 a_25712_23170# vdd 1.05f
C1206 X1.X2.X2.X2.X2.X1.X2.vin1 d1 1.03e-19
C1207 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.vrefh 0.00118f
C1208 a_33676_28070# a_33976_26164# 6.48e-19
C1209 X1.X1.X2.X1.X1.X2.X1.vin1 d1 0.0118f
C1210 a_40352_30794# a_40352_32700# 0.00396f
C1211 X2.vrefh vdd 0.419f
C1212 d3 a_31862_11822# 1.89e-19
C1213 d3 X1.X1.X2.X2.X3.vin2 0.417f
C1214 d2 a_39966_28888# 0.00665f
C1215 d3 a_52492_18358# 7.7e-20
C1216 a_25712_28888# X1.X2.X2.X2.X2.X2.X1.vin1 1.64e-19
C1217 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.vrefh 0.267f
C1218 d2 X2.X2.X2.X1.X3.vin2 0.00194f
C1219 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.X1.X1.X3.vin1 1.22e-19
C1220 a_25712_17452# d1 2.92e-22
C1221 d4 d1 0.151f
C1222 d4 X2.X1.X2.X2.X2.X2.vout 1.45e-19
C1223 a_54606_11734# d1 3.95e-19
C1224 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X1.X2.X2.X2.X2.vrefh 0.0128f
C1225 a_8186_25982# a_8572_25982# 0.414f
C1226 X1.X1.X2.X2.X3.vin1 d2 0.0014f
C1227 a_23212_22210# d1 0.00613f
C1228 X2.X1.X1.X2.X3.vin1 a_33976_10916# 0.17f
C1229 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.vout 0.118f
C1230 X1.X2.X1.X2.X1.X1.vout vdd 0.78f
C1231 a_23212_22210# a_25326_21264# 2.95e-20
C1232 a_23126_31700# d1 0.0489f
C1233 X2.X2.X2.X2.X2.X2.X3.vin1 vdd 0.993f
C1234 a_37852_29834# a_39966_28888# 2.95e-20
C1235 X1.X2.X1.X1.X2.X2.X3.vin2 a_19336_18540# 0.00504f
C1236 a_19422_20446# a_19722_18540# 4.41e-20
C1237 X1.X1.X3.vin2 X1.X1.X1.X2.X2.X1.vout 4.93e-20
C1238 X2.X2.X1.X1.X2.vrefh vdd 0.426f
C1239 X1.X1.X1.X2.X1.X1.vout X1.X1.X1.X2.X3.vin1 0.131f
C1240 d2 X1.X2.X2.X1.X2.X2.X2.vin1 0.0314f
C1241 X1.X1.X1.X1.X2.X1.X1.vin1 vdd 0.592f
C1242 a_8486_27888# vdd 0.561f
C1243 a_49002_22312# X2.X2.X1.X1.X2.X2.vout 0.263f
C1244 X1.X1.X2.X2.X2.X2.X1.vin1 d1 0.0118f
C1245 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X3.vin1 0.587f
C1246 a_23512_27888# a_25326_26982# 1.06e-19
C1247 a_40352_30794# vdd 1.05f
C1248 X1.X2.X1.X1.X2.vrefh a_17222_27070# 0.3f
C1249 d3 a_52792_8828# 0.00108f
C1250 a_23512_8828# a_22826_6962# 3.31e-19
C1251 a_23126_20264# a_23512_20264# 0.419f
C1252 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X3.vin2 0.17f
C1253 d1 X2.X1.X1.X2.X2.X2.X2.vin1 0.0144f
C1254 a_23212_25982# X1.X2.X2.X2.X2.X1.vout 1.64e-19
C1255 X1.X2.X1.X1.X1.X2.vout d1 0.033f
C1256 X2.X2.X2.X1.X2.X2.X1.vin2 d1 2.18e-19
C1257 X2.X1.X2.X1.X2.X2.X1.vin1 a_40352_13640# 1.64e-19
C1258 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.vout 0.038f
C1259 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 0.0565f
C1260 d0 X1.X1.X1.X2.X1.X2.X1.vin2 0.276f
C1261 a_54606_19358# d4 0.00112f
C1262 d3 a_10686_11734# 0.00112f
C1263 X1.X2.X1.X2.X2.X1.vout vdd 0.775f
C1264 d2 a_5082_14688# 0.0191f
C1265 a_2582_27070# X1.X1.X1.X1.X1.X2.X1.vin2 8.88e-20
C1266 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X1.X2.X2.X2.X2.vrefh 0.1f
C1267 X1.X2.X2.X1.X2.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin2 0.0128f
C1268 a_19036_31882# X1.X2.X1.X1.X1.X1.vout 0.359f
C1269 a_16836_28976# d0 0.518f
C1270 a_34062_9010# a_31862_8010# 4.77e-21
C1271 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X2.vin1 0.0689f
C1272 a_31862_21352# a_33676_20446# 1.06e-19
C1273 a_8572_10734# vdd 1.05f
C1274 a_25712_11734# d1 2.25e-20
C1275 X1.X2.X1.X3.vin1 a_19422_24258# 5.28e-19
C1276 a_17222_27070# vdd 0.542f
C1277 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.X1.X1.X1.vin1 0.206f
C1278 X2.X1.X2.X2.X2.vrefh a_40352_25076# 0.118f
C1279 d4 X2.X2.X3.vin2 0.297f
C1280 a_31862_19446# a_31862_17540# 0.00198f
C1281 a_31476_19446# X2.X1.X1.X2.X1.X1.X1.vin1 1.64e-19
C1282 X2.X1.X2.X2.X1.X1.X1.vin2 d4 3.99e-21
C1283 d4 X1.X1.X2.X2.X2.X1.vout 4.78e-20
C1284 X2.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X3.vin2 0.0533f
C1285 X2.X1.X3.vin1 d2 0.1f
C1286 a_23126_24076# d4 2.4e-19
C1287 X1.X2.X3.vin2 a_19722_10916# 3.68e-19
C1288 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X2.vin1 0.242f
C1289 a_48316_12822# a_48702_12822# 0.419f
C1290 X2.X2.X1.X2.X1.X2.X2.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 0.234f
C1291 X1.X2.X1.X1.X1.X1.vout vdd 0.781f
C1292 X2.X1.X2.X1.X2.X2.X2.vin1 a_39966_15546# 8.88e-20
C1293 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.X1.vin2 8.93e-19
C1294 a_23126_24076# a_23212_22210# 3.38e-19
C1295 a_54606_23170# X2.X2.X2.X2.X1.X2.vrefh 8.22e-20
C1296 a_4396_24258# d1 0.521f
C1297 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X1.vin2 0.668f
C1298 X1.X1.X3.vin1 d5 0.0576f
C1299 X2.X2.X2.X3.vin1 a_52406_12640# 5.28e-19
C1300 X1.X2.X2.X2.X1.X1.X3.vin2 a_23126_20264# 0.267f
C1301 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X3.vin1 0.00117f
C1302 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X2.vrefh 2.33e-19
C1303 a_54992_6016# a_54992_4110# 0.00396f
C1304 X1.X2.X2.X2.X1.X1.X1.vin2 d4 3.99e-21
C1305 X2.X2.X1.X1.X2.X2.X2.vin1 d0 0.262f
C1306 a_54606_9828# d1 0.00151f
C1307 a_33976_26164# X2.X1.X1.X1.X2.X1.X3.vin1 0.00251f
C1308 X2.X2.X2.X2.X2.X2.X1.vin2 d1 0.0985f
C1309 a_28096_892# vout 0.349f
C1310 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X2.X1.X1.X2.vrefh 0.00437f
C1311 d7 X3.vin2 4.93e-19
C1312 d4 a_5082_18540# 0.257f
C1313 d1 a_37766_8828# 0.0749f
C1314 vout vdd 0.362f
C1315 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.vout 0.399f
C1316 X1.X1.X1.X2.X1.X2.X3.vin1 a_4396_12822# 0.199f
C1317 a_52792_27888# a_54606_28888# 1.15e-20
C1318 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin2 7.84e-19
C1319 d1 X1.X2.X2.X1.X1.X2.X1.vin1 0.0118f
C1320 a_48702_28070# a_48616_26164# 3.3e-19
C1321 a_48316_28070# a_49002_26164# 3.08e-19
C1322 X2.X2.X1.X1.X2.X1.X2.vin1 vdd 0.576f
C1323 d2 X2.X2.X1.X2.X2.X1.X3.vin1 0.104f
C1324 X2.X1.X2.X2.X1.X1.X2.vin1 a_40352_21264# 0.197f
C1325 X2.X1.X2.X2.X1.X1.X3.vin1 a_39966_19358# 0.52f
C1326 X2.X2.X1.X1.X1.X2.X2.vin1 a_46502_28976# 8.88e-20
C1327 a_10686_21264# a_8872_20264# 1.15e-20
C1328 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X1.X2.X1.X2.X2.vrefh 0.267f
C1329 X1.X2.X1.X2.X1.X1.X1.vin2 a_16836_15634# 1.78e-19
C1330 X2.X1.X1.X1.X2.X2.X2.vin1 d0 0.262f
C1331 X1.X1.X2.X2.X1.X1.X1.vin2 d4 3.99e-21
C1332 a_48702_16634# X2.X2.X1.X2.X1.X1.vout 0.422f
C1333 a_2582_21352# X1.X1.X1.X1.X2.X2.X2.vin1 8.88e-20
C1334 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin1 0.52f
C1335 X2.X2.X2.X1.X1.X2.X1.vin2 X2.X2.X2.X1.X1.X2.vrefh 0.1f
C1336 X2.X2.X2.vrefh X2.X3.vin1 0.00136f
C1337 a_52492_6962# vdd 1.05f
C1338 X2.X2.X2.X2.X1.X1.X3.vin2 d2 0.169f
C1339 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.vout 0.118f
C1340 X2.X2.X2.X2.X1.X2.X3.vin2 d0 4.34e-19
C1341 d2 a_23512_8828# 0.00287f
C1342 X1.X1.X1.X2.X2.X1.X3.vin1 a_2582_8010# 0.00207f
C1343 X2.X1.X1.X1.X2.vrefh d1 0.00745f
C1344 X1.X2.X1.X2.X1.X1.vout X1.X2.X1.X2.X1.X2.vout 0.507f
C1345 a_52492_14586# d1 0.00613f
C1346 a_54606_17452# a_54992_17452# 0.419f
C1347 X1.X2.X1.X1.X2.X2.X2.vin1 d0 0.262f
C1348 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X1.vin2 0.076f
C1349 X1.X1.X2.X3.vin2 d1 0.0129f
C1350 X1.X2.X2.X1.X2.X1.X3.vin1 a_25326_11734# 0.52f
C1351 a_34362_26164# d2 7.13e-19
C1352 X2.X2.X2.vrefh a_54992_4110# 9.79e-19
C1353 a_46502_17540# X2.X2.X1.X2.X1.X1.X1.vin1 0.417f
C1354 a_46116_17540# X2.X2.X1.X2.X1.X1.X3.vin1 0.354f
C1355 X1.X1.X1.X1.X1.X2.X1.vin2 d1 0.00406f
C1356 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X1.vout 0.131f
C1357 d0 a_40352_9828# 0.515f
C1358 a_54606_11734# a_52492_10734# 5.36e-21
C1359 d3 X2.X2.X2.X2.X1.X2.X3.vin1 2.1e-19
C1360 X2.X2.X1.X1.X2.X2.vout d1 0.033f
C1361 d4 a_4396_16634# 0.00176f
C1362 X1.X1.X2.X2.X2.vrefh d1 0.00745f
C1363 X1.X1.X3.vin1 X1.X1.X3.vin2 3.25f
C1364 X2.X1.X1.X2.X2.X1.vout vdd 0.775f
C1365 X1.X1.X1.X3.vin2 X1.X1.X2.X3.vin1 1.22e-19
C1366 X1.X1.X1.X1.X1.X1.X1.vin2 a_4396_31882# 0.00113f
C1367 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.vrefh 0.161f
C1368 a_17222_28976# a_17222_30882# 0.00198f
C1369 d3 X2.X1.X1.X2.X1.X2.X2.vin1 8.68e-20
C1370 X1.X2.X1.X1.X1.X2.X1.vin1 a_16836_30882# 1.64e-19
C1371 a_25326_23170# X1.X2.X2.X2.X1.X2.vrefh 8.22e-20
C1372 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X1.X3.vin1 0.0425f
C1373 d0 X1.X2.X2.X1.X1.X2.X3.vin2 4.34e-19
C1374 X1.X2.X2.X2.X1.X1.X3.vin1 a_25326_19358# 0.52f
C1375 X1.X1.X1.X2.X2.X2.X2.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 0.234f
C1376 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.vout 0.118f
C1377 a_4396_5198# a_4782_5198# 0.419f
C1378 d3 X1.X2.X3.vin2 0.77f
C1379 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X2.vrefh 0.076f
C1380 X2.X2.X2.X1.X2.X1.X3.vin1 a_52106_10734# 0.00837f
C1381 a_34062_24258# X2.X1.X1.X1.X2.X1.vout 0.422f
C1382 X1.X1.X2.X1.X2.X2.X3.vin2 a_8872_16452# 0.101f
C1383 d2 X1.X1.X1.X1.X1.X2.X1.vin1 0.0114f
C1384 a_46116_13728# vdd 1.05f
C1385 a_23126_27888# a_22826_25982# 5.25e-20
C1386 d2 X1.X2.X2.X1.X2.X1.vout 0.00174f
C1387 d2 a_46502_11822# 0.00792f
C1388 a_48702_12822# d1 0.0749f
C1389 a_54606_25076# a_54992_25076# 0.419f
C1390 X2.X1.X2.X2.X1.X1.X3.vin2 a_39966_19358# 7.84e-19
C1391 X1.X2.X2.X3.vin1 a_23126_16452# 5.31e-19
C1392 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X3.vin1 0.00117f
C1393 X2.X1.X2.X1.X2.X1.X3.vin2 a_37766_12640# 0.267f
C1394 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X1.X2.X2.X1.X1.X1.vin1 0.0689f
C1395 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X1.vout 0.13f
C1396 a_54606_6016# X2.X2.X2.X1.X1.X1.X2.vin1 0.402f
C1397 X2.X1.X1.X1.X2.X2.X1.vin1 d0 0.267f
C1398 a_54606_28888# vdd 0.541f
C1399 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X1.X2.X1.X1.X2.vrefh 0.00437f
C1400 a_8486_16452# vdd 0.471f
C1401 a_4782_9010# X1.X1.X1.X2.X2.X1.vout 0.422f
C1402 a_46116_25164# X2.X2.X1.X1.X2.X1.X3.vin1 0.354f
C1403 d3 X2.X1.X1.X2.X1.X1.vout 0.00883f
C1404 a_52106_29834# X2.X2.X2.X2.X2.X1.vout 0.383f
C1405 a_46502_25164# X2.X2.X1.X1.X2.X1.X1.vin1 0.417f
C1406 X1.X2.X1.X1.X1.X2.X2.vin1 X1.X2.X1.X1.X2.vrefh 0.564f
C1407 a_23126_27888# X1.X2.X2.X2.X2.X1.X3.vin1 0.428f
C1408 d1 d7 2.34e-19
C1409 X2.X1.X1.X2.X3.vin2 vdd 1.29f
C1410 d0 X2.X2.X2.X1.X1.X1.X1.vin2 0.276f
C1411 a_31476_15634# X2.X1.X1.X2.X1.X2.X1.vin1 1.64e-19
C1412 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X1.vin1 0.0689f
C1413 X2.X1.X2.X1.X1.X2.X3.vin2 a_39966_7922# 7.84e-19
C1414 a_31862_15634# a_31862_13728# 0.00198f
C1415 X2.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X1.vin1 0.142f
C1416 d4 a_34362_29936# 0.00116f
C1417 X2.X1.X1.X3.vin2 d1 0.0129f
C1418 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X3.vin2 0.552f
C1419 d2 a_46116_15634# 0.00414f
C1420 X2.X2.X1.X2.X1.X1.vout d1 0.0238f
C1421 X2.X1.X1.X2.X1.X2.X3.vin2 a_34362_10916# 0.00846f
C1422 X2.X1.X2.X1.X2.X2.X2.vin1 vdd 0.576f
C1423 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X3.vin1 1.22e-19
C1424 d2 a_19336_7064# 0.608f
C1425 X1.X2.X2.X3.vin1 a_23126_8828# 1.64e-19
C1426 X1.X1.X2.X1.X3.vin1 a_8572_6962# 0.363f
C1427 X2.X2.X1.X2.vrefh a_46502_19446# 0.3f
C1428 a_52792_24076# a_52106_22210# 3.31e-19
C1429 X2.X2.X2.X2.X2.X1.X1.vin1 a_54992_26982# 0.195f
C1430 X1.X2.X2.X1.X1.X2.X1.vin2 X1.X2.X2.X1.X1.X2.vrefh 0.1f
C1431 a_4696_7064# a_4782_5198# 3.38e-19
C1432 a_4696_22312# X1.X1.X1.X1.X2.X2.vout 0.0929f
C1433 a_5082_7064# a_4396_5198# 3.31e-19
C1434 a_33676_9010# X2.X1.X1.X2.X2.X1.vout 0.359f
C1435 a_10686_6016# a_10686_7922# 0.00198f
C1436 a_19336_29936# a_19036_31882# 6.1e-19
C1437 X1.X1.X3.vin1 a_6032_892# 0.371f
C1438 X1.X1.X1.X1.X2.X2.X2.vin1 a_2196_19446# 0.197f
C1439 d2 X1.X2.X2.X1.X2.X1.X1.vin2 0.231f
C1440 X2.X1.X1.X1.X2.X1.vout d1 0.0238f
C1441 X2.X1.X2.X2.X2.X2.X2.vin1 a_38152_31700# 5.34e-19
C1442 X1.X2.X1.X1.X1.X2.X2.vin1 vdd 0.576f
C1443 X1.X1.X2.X1.X2.X1.X2.vin1 a_11072_11734# 1.78e-19
C1444 X1.X1.X2.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X1.vin1 2.23e-19
C1445 X1.X1.X1.X2.X2.X1.vout d1 0.0238f
C1446 X2.X1.X2.X2.X2.X1.X1.vin2 d3 3.99e-21
C1447 d4 X1.X2.X2.X3.vin1 0.0865f
C1448 d1 X2.X2.X2.X1.X1.X1.X2.vin1 0.0144f
C1449 a_52492_10734# a_54606_9828# 4.72e-20
C1450 X2.X2.X1.X1.X2.X1.X1.vin1 d1 0.0118f
C1451 a_25326_9828# a_25712_9828# 0.419f
C1452 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X2.vrefh 0.267f
C1453 X1.X2.X1.X2.X2.X1.X1.vin2 a_17222_8010# 8.88e-20
C1454 a_8186_29834# a_8872_31700# 3.31e-19
C1455 d2 X2.X1.X2.X1.X2.X2.X3.vin1 0.153f
C1456 X2.X1.X3.vin2 a_37766_5016# 2.33e-19
C1457 a_48702_31882# X2.X2.X1.X1.X1.X1.vout 0.422f
C1458 X1.X1.X3.vin1 X1.X1.X1.X2.X3.vin2 0.0816f
C1459 a_16836_21352# X1.X2.X1.X1.X2.X2.X2.vin1 1.78e-19
C1460 d0 X1.X2.X2.X1.X1.X1.X1.vin2 0.276f
C1461 a_19336_29936# vdd 1.05f
C1462 a_8486_31700# vdd 0.471f
C1463 d3 X1.X1.X1.X2.X1.X2.X3.vin1 2.1e-19
C1464 a_4696_26164# a_4396_24258# 6.2e-19
C1465 X1.X1.X1.X2.X2.X1.X3.vin2 a_2582_8010# 0.567f
C1466 X1.X2.X2.vrefh a_25712_4110# 9.79e-19
C1467 a_16836_9916# X1.X2.X1.X2.X2.X1.X3.vin1 0.354f
C1468 a_17222_9916# X1.X2.X1.X2.X2.X1.X1.vin1 0.417f
C1469 X2.X1.X2.X2.X1.X2.X3.vin1 a_37466_22210# 0.00874f
C1470 X2.X2.X2.X1.X1.X1.X3.vin2 a_52406_5016# 0.267f
C1471 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X1.vin2 0.668f
C1472 X2.X1.X1.X2.X1.X1.X3.vin2 a_34362_14688# 0.00815f
C1473 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X2.vrefh 0.00118f
C1474 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X3.vin1 0.00117f
C1475 a_22826_14586# a_23512_12640# 2.86e-19
C1476 d2 a_25712_15546# 0.00274f
C1477 a_54992_26982# d1 2.25e-20
C1478 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X3.vin2 0.237f
C1479 a_34362_10916# a_34062_9010# 5.25e-20
C1480 a_33976_10916# X2.X1.X1.X2.X2.X1.vout 1.64e-19
C1481 a_48616_18540# a_49002_18540# 0.413f
C1482 X2.X2.X1.X1.X1.X1.vout d1 0.0238f
C1483 a_46502_30882# X2.X2.X1.X1.X1.X1.X1.vin2 8.88e-20
C1484 d6 X1.X3.vin2 0.0894f
C1485 X1.X2.X1.X2.X2.X1.X1.vin1 d1 0.0118f
C1486 a_4696_7064# a_5082_7064# 0.419f
C1487 a_19722_22312# X1.X2.X1.X1.X2.X2.X3.vin2 3.85e-19
C1488 d3 X2.X2.X2.X2.X3.vin2 0.157f
C1489 X1.X2.X1.X1.X2.X2.vout a_19422_20446# 0.418f
C1490 X1.X2.X2.X2.X1.X2.vrefh vdd 0.414f
C1491 d2 a_31862_9916# 0.00328f
C1492 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X3.vin2 0.102f
C1493 d0 X1.X2.X1.X2.X2.vrefh 0.848f
C1494 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X2.vrefh 0.076f
C1495 X1.X1.X2.X2.X2.X1.X3.vin2 a_8872_27888# 0.1f
C1496 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X3.vin2 0.161f
C1497 X2.X2.X1.X1.X1.X1.vout X2.X2.X1.X1.X1.X1.X3.vin1 0.118f
C1498 a_8186_18358# vdd 0.476f
C1499 X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X2.vout 0.0866f
C1500 X1.X2.X2.X2.X1.X1.X2.vin1 d1 1.03e-19
C1501 X2.X1.X2.X2.X2.X1.X3.vin1 a_37466_25982# 0.00837f
C1502 a_25326_21264# X1.X2.X2.X2.X1.X1.X2.vin1 0.402f
C1503 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 0.242f
C1504 a_54606_13640# a_54606_11734# 0.00198f
C1505 X2.X2.X2.X2.X3.vin1 d2 0.0014f
C1506 X2.X1.X1.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X1.X2.vrefh 0.165f
C1507 X1.X2.X3.vin1 a_19422_5198# 2.12e-19
C1508 X1.X1.X2.X1.X1.X1.X1.vin2 a_10686_4110# 0.273f
C1509 a_2582_28976# a_4782_28070# 4.2e-20
C1510 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X2.X2.vin1 0.00117f
C1511 a_39966_21264# d2 0.0059f
C1512 a_8572_22210# a_8872_20264# 6.1e-19
C1513 a_22826_10734# a_23126_8828# 4.41e-20
C1514 a_33976_10916# X2.X1.X1.X2.X3.vin2 0.0927f
C1515 d0 a_46116_6104# 0.518f
C1516 a_37466_18358# a_37766_16452# 4.41e-20
C1517 a_19722_18540# X1.X2.X1.X3.vin2 0.233f
C1518 X2.X2.X2.X2.X3.vin2 X2.X2.X2.X2.X2.X1.X3.vin2 0.0533f
C1519 a_39966_25076# d0 0.0489f
C1520 a_37766_8828# a_37466_6962# 5.55e-20
C1521 X2.X1.X2.X1.X2.X1.X1.vin1 a_40352_9828# 1.64e-19
C1522 d2 X2.X1.X2.X2.X2.X2.X3.vin1 0.0571f
C1523 a_10686_26982# a_10686_25076# 0.00198f
C1524 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.vout 0.08f
C1525 a_38152_27888# d2 0.00251f
C1526 X1.X2.X2.X1.X1.X1.X3.vin2 a_25326_4110# 7.84e-19
C1527 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X1.vin1 0.0689f
C1528 a_46502_21352# a_46502_19446# 0.00198f
C1529 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.vout 0.398f
C1530 d2 a_49002_14688# 0.0191f
C1531 a_48702_5198# a_46502_4198# 4.77e-21
C1532 a_19336_14688# a_17222_13728# 2.68e-20
C1533 X2.X1.X2.X1.X2.X2.X3.vin1 a_38152_16452# 0.199f
C1534 X1.X2.X2.X1.X3.vin2 d1 0.00807f
C1535 a_8486_20264# vdd 0.561f
C1536 X2.X2.X1.X2.X2.X2.X3.vin2 a_46116_4198# 0.354f
C1537 a_22826_25982# d4 7.15e-19
C1538 X2.X2.X2.X2.X1.X1.X1.vin1 d1 0.011f
C1539 X1.X2.X2.X3.vin2 a_22826_22210# 0.00292f
C1540 a_2196_32788# vdd 1.05f
C1541 a_37852_29834# X2.X1.X2.X2.X2.X2.X3.vin1 0.00329f
C1542 X2.X2.X1.X2.X2.X2.X3.vin2 X2.X2.X2.vrefh 0.172f
C1543 X2.X1.X2.X1.X2.X2.vrefh a_40352_13640# 0.118f
C1544 d2 a_4696_10916# 0.0057f
C1545 d4 X2.X2.X1.X2.X1.X1.X1.vin1 6.34e-20
C1546 a_37852_22210# d2 0.526f
C1547 a_23126_27888# X1.X2.X2.X2.X2.X1.X3.vin2 0.267f
C1548 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X1.X2.vin1 0.00117f
C1549 a_38152_27888# a_37852_29834# 6.1e-19
C1550 X1.X2.X2.X1.X2.X2.X1.vin2 X2.X1.X1.X2.X1.X2.vrefh 0.0128f
C1551 X1.X1.X1.X1.X1.X2.vout X1.X1.X1.X1.X1.X2.X3.vin2 0.075f
C1552 d0 a_10686_9828# 0.0489f
C1553 X1.X1.X3.vin1 a_4782_9010# 2.12e-19
C1554 d3 X2.X2.X1.X2.X2.X1.vout 0.00146f
C1555 d4 X2.X2.X2.X2.X2.X1.vout 0.0233f
C1556 X1.X2.X2.X2.X2.X1.X3.vin1 d4 0.00851f
C1557 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X2.vin1 0.0689f
C1558 a_2196_11822# a_2582_11822# 0.419f
C1559 a_31862_25164# a_33676_24258# 1.06e-19
C1560 a_31476_13728# X2.X1.X1.X2.X1.X2.X2.vin1 1.78e-19
C1561 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X1.X3.vin2 5.19e-19
C1562 a_22826_14586# a_23212_14586# 0.419f
C1563 X1.X1.X2.X1.X2.X1.X2.vin1 vdd 0.576f
C1564 d3 a_31862_32788# 1.28e-19
C1565 a_39966_19358# d1 3.95e-19
C1566 a_16836_21352# d0 0.518f
C1567 a_54606_23170# d2 0.00479f
C1568 X2.X1.X2.X2.vrefh d4 6.65e-20
C1569 a_54606_19358# X2.X2.X2.X2.X1.X1.X1.vin1 0.417f
C1570 X2.X2.X3.vin1 d5 0.00767f
C1571 X1.X2.X2.X2.X1.X2.X3.vin1 d1 0.146f
C1572 X2.X2.X2.X2.X1.X1.X1.vin2 a_54992_19358# 0.12f
C1573 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 0.581f
C1574 d0 a_54992_32700# 0.515f
C1575 X1.X2.X1.X1.X1.X2.X1.vin1 vdd 0.592f
C1576 a_11072_23170# d1 2.25e-20
C1577 d3 X2.X1.X2.X1.X1.X2.X3.vin2 0.0251f
C1578 X2.X1.X1.X2.X2.X2.X3.vin2 a_31476_4198# 0.354f
C1579 a_34062_5198# a_31862_4198# 4.77e-21
C1580 X2.X1.X1.X1.X3.vin1 X2.X1.X2.X2.X3.vin2 0.0604f
C1581 X2.X2.X2.X1.X1.X1.vout X2.X2.X2.X1.X3.vin1 0.13f
C1582 d0 X2.X2.X1.X2.X2.X2.X2.vin1 0.262f
C1583 X1.X2.X1.X1.X2.X1.X3.vin2 d2 0.171f
C1584 X2.X1.X1.X2.X2.X2.X3.vin2 X2.X1.X2.vrefh 0.172f
C1585 X2.X2.X1.X2.X1.X1.X3.vin2 a_48616_14688# 0.00546f
C1586 a_39966_32700# X2.X1.X2.X2.X2.X2.X1.vin2 8.88e-20
C1587 X2.X1.X2.X1.X2.X1.vout a_38152_12640# 0.359f
C1588 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.X1.X1.vin1 5.19e-19
C1589 a_25326_21264# a_25326_19358# 0.00198f
C1590 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X1.vin2 3.94e-19
C1591 a_25326_19358# d1 3.95e-19
C1592 X2.X1.X3.vin2 X2.X1.X2.X1.X3.vin2 0.039f
C1593 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 0.242f
C1594 X1.X2.X1.X2.X1.X1.X1.vin2 vdd 0.36f
C1595 d2 X2.X2.X1.X2.X1.X1.X2.vin1 0.031f
C1596 X1.X2.X1.X2.X1.X1.X2.vin1 X1.X2.X1.X2.X1.X2.vrefh 0.564f
C1597 d4 a_49002_18540# 0.256f
C1598 a_23126_16452# X1.X2.X2.X1.X2.X2.X3.vin1 0.42f
C1599 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X2.X1.X2.X2.vrefh 0.0128f
C1600 X1.X1.X3.vin1 d1 0.046f
C1601 a_23126_12640# d1 0.0749f
C1602 a_2582_9916# a_4396_9010# 1.06e-19
C1603 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X2.vin1 0.0689f
C1604 a_37466_29834# vdd 0.477f
C1605 a_11072_13640# X1.X1.X2.X1.X2.X1.X1.vin2 1.78e-19
C1606 a_54992_28888# X2.X2.X2.X2.X2.X2.X1.vin1 1.64e-19
C1607 X1.X1.X2.X2.X1.X2.vout d2 0.00124f
C1608 a_38152_5016# vdd 1.05f
C1609 d2 X2.X2.X2.X1.X1.X2.X3.vin1 0.157f
C1610 X2.X3.vin1 X2.X3.vin2 0.514f
C1611 a_37466_25982# X2.X1.X2.X2.X1.X2.X3.vin2 0.00846f
C1612 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X1.vin1 5.19e-19
C1613 d0 X2.X1.X2.X1.X2.X1.X1.vin1 0.267f
C1614 X1.X1.X1.X2.X1.X1.X3.vin1 d0 4.36e-19
C1615 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X1.X2.X2.X2.X2.vrefh 0.0128f
C1616 a_46116_23258# d0 0.515f
C1617 d3 a_49002_10916# 0.29f
C1618 a_48702_20446# vdd 0.471f
C1619 X1.X1.X2.X1.X2.X2.X1.vin1 a_11072_15546# 0.195f
C1620 a_10686_19358# d1 3.95e-19
C1621 X2.X1.X1.X1.X2.X1.X2.vin1 d2 0.0318f
C1622 d2 a_40352_7922# 0.00351f
C1623 d1 X2.X1.X1.X2.X2.X2.X1.vin2 0.0985f
C1624 X1.X1.X2.X1.X2.X1.X3.vin1 d1 0.151f
C1625 a_52792_16452# a_54606_15546# 1.06e-19
C1626 X2.X1.X2.X2.X1.X1.X1.vin2 a_39966_19358# 0.273f
C1627 a_31476_25164# d1 2.25e-20
C1628 X1.X2.X2.X2.X2.X2.X2.vin1 a_25712_30794# 1.78e-19
C1629 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.X1.vin1 2.23e-19
C1630 a_34062_28070# d3 7.51e-19
C1631 d2 X1.X1.X1.X2.X2.X1.X2.vin1 0.0318f
C1632 d0 X2.X2.X2.X1.X2.X2.X3.vin1 4.36e-19
C1633 a_40352_25076# d2 0.00533f
C1634 a_22826_6962# a_23126_5016# 4.19e-20
C1635 a_23126_24076# X1.X2.X2.X2.X1.X2.X3.vin1 0.42f
C1636 X1.X2.X1.X2.X2.X2.X3.vin2 a_17222_4198# 0.567f
C1637 X1.X2.X1.X1.X2.X1.X2.vin1 X1.X2.X1.X1.X2.X2.vrefh 0.564f
C1638 X1.X2.X1.X2.X2.X2.X3.vin1 a_17222_4198# 0.00207f
C1639 a_25326_13640# a_25712_13640# 0.419f
C1640 d6 vdd 0.917f
C1641 d2 X1.X1.X1.X2.X1.X2.X3.vin2 0.121f
C1642 d2 X2.X1.X1.X2.X2.X2.X1.vin1 9.24e-20
C1643 X1.X1.X1.X2.X1.X1.X3.vin2 a_2196_15634# 0.354f
C1644 d6 a_28096_892# 0.00105f
C1645 a_17222_6104# d0 0.0675f
C1646 a_46116_6104# X2.X2.X1.X2.X2.X2.X2.vin1 1.78e-19
C1647 a_52492_14586# a_54606_13640# 2.95e-20
C1648 a_33976_18540# vdd 1.05f
C1649 d0 a_40352_15546# 0.518f
C1650 X1.X2.X2.X2.X1.X2.X3.vin2 d2 0.121f
C1651 X2.X2.X2.X2.X2.X1.X1.vin2 d2 0.231f
C1652 a_34062_20446# vdd 0.471f
C1653 X2.X2.X2.X3.vin2 d1 0.0129f
C1654 X1.X2.X2.X1.X2.X1.X1.vin1 X2.X1.X1.X2.X2.vrefh 0.00437f
C1655 a_16836_13728# X1.X2.X1.X2.X1.X2.X3.vin1 0.354f
C1656 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.vout 0.08f
C1657 a_17222_13728# X1.X2.X1.X2.X1.X2.X1.vin1 0.417f
C1658 X1.X1.X1.X2.vrefh d4 6.65e-20
C1659 X2.X1.X2.X2.X2.X1.X1.vin2 a_39966_28888# 8.88e-20
C1660 X2.X1.X2.X2.X1.X2.X3.vin1 d0 4.36e-19
C1661 X1.X1.X2.X2.X1.X2.X1.vin1 a_11072_23170# 0.195f
C1662 d4 X1.X2.X2.X1.X2.X2.X3.vin1 2.52e-19
C1663 a_2196_9916# d1 2.25e-20
C1664 a_48316_31882# X2.X2.X1.X1.X1.X1.X1.vin2 0.00113f
C1665 a_10686_32700# d4 8.99e-20
C1666 a_23126_8828# X1.X2.X2.X1.X1.X2.X3.vin1 0.42f
C1667 d2 X2.X2.X1.X1.X1.X1.X2.vin1 6e-20
C1668 a_52492_29834# a_52406_31700# 3.38e-19
C1669 d3 X2.X2.X2.X1.X2.X1.X3.vin1 0.0195f
C1670 X1.X1.X3.vin2 X1.X1.X1.X2.X2.X2.vout 1.5e-19
C1671 a_4782_16634# d1 0.0749f
C1672 d2 a_11072_9828# 0.00533f
C1673 d0 X1.X1.X2.X1.X1.X2.X3.vin1 4.36e-19
C1674 X2.X1.X2.X2.X2.X2.X3.vin1 a_38152_31700# 0.199f
C1675 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 5.19e-19
C1676 X2.X1.X1.X1.X1.X1.X1.vin2 vdd 0.399f
C1677 a_25712_23170# d0 0.518f
C1678 a_31862_28976# X2.X1.X1.X1.X1.X2.X1.vin2 0.273f
C1679 d3 X1.X2.X2.X2.X2.X1.vout 0.0015f
C1680 a_19422_20446# vdd 0.471f
C1681 X2.vrefh d0 0.0263f
C1682 X1.X1.X2.X2.X2.X2.X2.vin1 a_10686_30794# 8.88e-20
C1683 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.X1.vin2 8.93e-19
C1684 X1.X2.X2.X2.X2.X2.X1.vin2 X2.X1.X1.X1.X1.X2.vrefh 0.0128f
C1685 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X2.vrefh 2.33e-19
C1686 X1.X1.X1.X1.X2.X2.X1.vin2 d1 2.18e-19
C1687 X2.X1.X1.X1.X2.X2.vrefh a_31476_23258# 0.118f
C1688 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X3.vin2 8.93e-19
C1689 X1.X1.X1.X1.X2.X1.X3.vin2 a_2196_23258# 0.354f
C1690 X1.X2.X2.X2.X2.X1.X2.vin1 X1.X2.X2.X2.X2.X1.X3.vin2 0.234f
C1691 X2.X1.X3.vin1 X2.X1.X1.X2.X1.X1.vout 2.91e-19
C1692 X1.X2.X2.X2.X1.X1.X1.vin2 a_25326_19358# 0.273f
C1693 X1.X1.X2.X1.X1.X2.X1.vin1 a_11072_7922# 0.195f
C1694 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X3.vin1 0.00118f
C1695 a_5082_26164# d1 0.0318f
C1696 a_52106_6962# X2.X2.X2.X1.X1.X2.X3.vin1 0.00874f
C1697 a_46502_9916# vdd 0.553f
C1698 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X2.vout 0.2f
C1699 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.vout 0.075f
C1700 a_8872_16452# a_8572_14586# 6.71e-19
C1701 a_23512_20264# a_22826_18358# 2.97e-19
C1702 a_31476_11822# X2.X1.X1.X2.X2.X1.X1.vin1 1.64e-19
C1703 X1.X1.X1.X1.X2.X2.X1.vin1 d2 0.0106f
C1704 a_31862_11822# a_31862_9916# 0.00198f
C1705 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.X3.vin2 0.587f
C1706 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X2.X3.vin1 0.0131f
C1707 X2.X2.X2.X2.X2.X2.X3.vin1 d0 4.36e-19
C1708 X1.X2.X2.X2.X2.X1.X1.vin1 d2 0.0105f
C1709 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 1.22e-19
C1710 d2 a_46502_32788# 1.95e-19
C1711 X2.X2.X1.X1.X2.vrefh d0 0.848f
C1712 X2.X2.X1.X1.X1.X1.X1.vin1 X2.X2.X1.X1.X1.X1.X1.vin2 0.696f
C1713 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X3.vin1 2.33e-19
C1714 d4 X1.X2.X2.X2.X2.X1.X3.vin2 0.0533f
C1715 a_5082_18540# X1.X1.X3.vin1 0.47f
C1716 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin1 0.267f
C1717 X1.X1.X1.X1.X2.X1.X1.vin1 d0 0.267f
C1718 a_52406_5016# a_52792_5016# 0.419f
C1719 a_35312_892# vdd 0.475f
C1720 a_19722_22312# X1.X2.X1.X1.X2.X2.X3.vin1 0.00874f
C1721 a_40352_30794# d0 0.518f
C1722 a_33976_26164# X2.X1.X1.X1.X1.X2.vout 7.93e-20
C1723 a_54606_21264# vdd 0.541f
C1724 X2.X2.X2.X3.vin2 X2.X2.X3.vin2 0.171f
C1725 a_52492_25982# a_52792_24076# 6.48e-19
C1726 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X1.X3.vin2 1.22e-19
C1727 d3 a_19722_18540# 0.0469f
C1728 a_2196_15634# vdd 1.05f
C1729 X2.X1.X1.X1.X3.vin1 d1 0.00179f
C1730 a_5082_14688# X1.X1.X1.X2.X1.X2.X3.vin1 0.00874f
C1731 a_11072_17452# d1 2.92e-22
C1732 a_39966_25076# X2.X1.X2.X2.X1.X2.X3.vin1 0.00207f
C1733 d1 X2.X1.X2.X1.X1.X1.vout 0.0239f
C1734 X1.X2.X1.X1.X1.X2.X2.vin1 a_16836_28976# 1.78e-19
C1735 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.X1.vin2 0.216f
C1736 X1.X1.X3.vin1 a_8486_12640# 8.66e-20
C1737 d4 X1.X2.X2.X2.X2.X2.X3.vin1 0.00851f
C1738 X2.X2.X2.X1.X2.X1.X1.vin2 a_54992_11734# 0.12f
C1739 a_54606_11734# X2.X2.X2.X1.X2.X1.X1.vin1 0.417f
C1740 a_8186_22210# d2 0.0191f
C1741 a_23126_31700# X1.X2.X2.X2.X2.X2.X3.vin1 0.42f
C1742 X1.X2.X1.X1.X1.X1.X2.vin1 X1.X2.X1.X1.X1.X2.vrefh 0.564f
C1743 d3 a_54606_25076# 1.89e-19
C1744 a_4782_31882# d1 0.0394f
C1745 X2.X2.X1.X2.X1.X1.X1.vin2 a_46116_15634# 1.78e-19
C1746 a_23212_25982# vdd 1.05f
C1747 X1.X1.X2.X1.X2.X2.X2.vin1 d2 0.0314f
C1748 a_49002_29936# X2.X2.X1.X1.X1.X2.vout 0.254f
C1749 X2.X2.X2.X1.X1.X1.X1.vin1 vdd 0.592f
C1750 X2.X1.X2.X2.X2.X1.X3.vin1 vdd 0.997f
C1751 d1 a_23512_5016# 0.522f
C1752 X1.X1.X2.X2.X1.X1.X1.vin2 a_10686_19358# 0.273f
C1753 X1.X1.X1.X2.X1.X2.X2.vin1 X1.X1.X1.X2.X2.vrefh 0.564f
C1754 a_2196_8010# vdd 1.05f
C1755 a_8486_12640# X1.X1.X2.X1.X2.X1.X3.vin1 0.428f
C1756 a_31862_19446# d2 0.00583f
C1757 a_17222_27070# d0 0.0489f
C1758 X1.X2.X2.X2.X1.X1.X3.vin2 a_22826_18358# 3.49e-19
C1759 a_10686_6016# d1 0.00148f
C1760 a_8186_14586# X1.X1.X2.X1.X3.vin2 0.423f
C1761 X1.X1.X2.X2.X2.X2.X1.vin1 a_11072_30794# 0.195f
C1762 X2.X2.X1.X2.X1.X1.X3.vin1 a_48702_16634# 0.428f
C1763 d2 a_23126_5016# 0.00123f
C1764 X2.X1.X2.X1.X1.X1.X3.vin1 a_38152_5016# 0.199f
C1765 a_2196_28976# vdd 1.05f
C1766 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X2.vout 0.0866f
C1767 X1.X2.X2.X1.X1.X1.X3.vin2 a_25712_6016# 0.354f
C1768 X2.X1.X2.X1.X3.vin2 a_37766_12640# 0.00101f
C1769 a_10686_23170# a_10686_21264# 0.00198f
C1770 a_52792_31700# a_54606_30794# 1.06e-19
C1771 a_8872_24076# d1 0.521f
C1772 a_10686_9828# X1.X1.X2.X1.X1.X2.X3.vin1 0.00207f
C1773 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X1.vin2 0.216f
C1774 d3 a_25326_9828# 1.89e-19
C1775 a_5082_18540# a_4782_16634# 5.25e-20
C1776 X1.X1.X2.X2.X1.X2.X1.vin2 d2 0.226f
C1777 a_4696_18540# X1.X1.X1.X2.X1.X1.vout 1.64e-19
C1778 a_39966_15546# a_37852_14586# 2.68e-20
C1779 X1.X1.X1.X1.X2.X2.vrefh a_2582_21352# 8.22e-20
C1780 X1.X1.X1.X2.X2.X2.X3.vin1 d2 0.0577f
C1781 X2.X2.X1.X2.X2.vrefh vdd 0.426f
C1782 X1.X1.X1.X1.X1.X1.X3.vin2 a_2196_30882# 0.354f
C1783 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X1.X1.vin2 0.216f
C1784 d2 X1.X2.X2.X1.X2.X2.vrefh 0.168f
C1785 X1.X2.X1.X1.X2.X1.X3.vin2 a_19336_22312# 0.00546f
C1786 a_52406_27888# a_54606_26982# 4.2e-20
C1787 a_17222_19446# d2 0.00583f
C1788 a_39966_11734# a_40352_11734# 0.419f
C1789 X2.X2.X2.X1.X2.X2.X1.vin2 a_54606_15546# 0.273f
C1790 a_2196_30882# vdd 1.05f
C1791 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X3.vin2 0.418f
C1792 X1.X2.X3.vin2 X1.X2.X2.X1.X2.X1.vout 3.2e-19
C1793 X1.X2.X2.X2.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin2 0.0128f
C1794 X2.X2.X1.X1.X1.X2.X1.vin1 a_46116_30882# 1.64e-19
C1795 a_2196_13728# a_2196_11822# 0.00396f
C1796 a_46502_28976# a_46502_30882# 0.00198f
C1797 X1.X2.X2.X1.X1.X1.X1.vin1 vdd 0.592f
C1798 X1.X2.X1.X1.X1.X1.X1.vin2 d1 0.00147f
C1799 X1.X1.X1.X3.vin1 a_4696_18540# 0.17f
C1800 a_4782_24258# d4 2.4e-19
C1801 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X2.vin1 0.564f
C1802 a_52106_18358# vdd 0.476f
C1803 X1.X1.X1.X1.X1.X2.vout vdd 0.696f
C1804 a_25712_32700# X1.X2.X2.X2.X2.X2.X1.vin2 1.78e-19
C1805 a_52106_25982# a_52492_25982# 0.414f
C1806 X1.X1.X2.X2.X1.X2.vrefh d2 0.177f
C1807 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.X1.vin1 0.206f
C1808 d3 a_19336_26164# 0.621f
C1809 X2.X2.X1.X1.X2.X1.X2.vin1 d0 0.262f
C1810 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 0.0565f
C1811 X2.X2.X2.X1.X2.X1.X2.vin1 d1 1.03e-19
C1812 a_2582_19446# d2 0.00583f
C1813 X1.X2.X1.X1.X1.X1.X1.vin1 d2 0.00798f
C1814 d3 X2.X2.X2.X2.X1.X1.vout 0.00883f
C1815 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.X1.X1.X1.vin1 5.19e-19
C1816 a_17222_19446# a_17222_17540# 0.00198f
C1817 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X2.X1.X1.X2.X2.vrefh 0.00437f
C1818 X2.X2.X3.vin1 a_48702_16634# 2.92e-19
C1819 X1.X2.X1.X2.X2.X1.X2.vin1 a_17222_8010# 0.402f
C1820 X2.X2.X1.X2.X2.X1.X3.vin2 a_49002_7064# 0.00815f
C1821 X2.X2.X2.X2.X2.X2.vout X2.X2.X2.X2.X2.X2.X3.vin2 0.08f
C1822 a_17222_11822# vdd 0.542f
C1823 X2.X2.X2.X1.X2.X1.X1.vin1 a_54606_9828# 8.22e-20
C1824 X2.X2.X2.X1.X2.X1.X1.vin2 X2.X2.X2.X1.X1.X2.X3.vin2 3.94e-19
C1825 a_8572_25982# a_8872_27888# 6.2e-19
C1826 a_17222_6104# a_19036_5198# 1.06e-19
C1827 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X2.vin1 0.0689f
C1828 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin1 0.195f
C1829 d3 a_49002_29936# 0.00177f
C1830 a_10686_25076# d2 0.00792f
C1831 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X1.X1.vin1 0.206f
C1832 X1.X2.X2.X1.X2.X1.X1.vin2 X2.X1.X1.X2.X1.X2.X2.vin1 0.00232f
C1833 X1.X1.X2.X2.X1.X2.X3.vin1 vdd 0.96f
C1834 a_4396_16634# a_4782_16634# 0.419f
C1835 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.vout 0.0857f
C1836 a_48316_28070# d2 0.00393f
C1837 d3 a_8186_14586# 9.23e-19
C1838 a_8572_10734# a_10686_9828# 4.72e-20
C1839 a_54992_25076# vdd 1.05f
C1840 X2.X1.X1.X1.X1.X2.X3.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 1.22e-19
C1841 a_31862_8010# a_33976_7064# 2.95e-20
C1842 d2 X1.X2.X2.X2.X2.X2.vrefh 0.168f
C1843 X1.X2.X2.X2.X3.vin1 d1 0.00179f
C1844 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X1.X2.X1.vin2 8.93e-19
C1845 X1.X2.X2.X1.X3.vin1 d1 0.00179f
C1846 X2.X2.X1.X2.X1.X1.X3.vin1 d1 0.146f
C1847 X2.X2.X1.X2.X2.X2.X1.vin1 vdd 0.592f
C1848 a_25326_15546# vdd 0.553f
C1849 X2.X1.X2.X2.X1.X2.X3.vin2 vdd 0.787f
C1850 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 2.23e-19
C1851 d1 X1.X1.X1.X2.X2.X2.X3.vin2 0.214f
C1852 d4 a_8872_16452# 0.00119f
C1853 X1.X1.X1.X2.X2.X1.vout a_5082_7064# 0.383f
C1854 X1.X2.X2.X3.vin1 a_23126_12640# 5.28e-19
C1855 X2.X2.X2.X1.X1.X2.X3.vin1 a_52792_8828# 0.199f
C1856 d3 X2.X1.X2.X3.vin1 0.676f
C1857 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin1 0.195f
C1858 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 5.19e-19
C1859 a_4396_24258# a_4782_24258# 0.419f
C1860 d1 a_39966_4110# 0.00107f
C1861 a_25712_9828# vdd 1.05f
C1862 d0 a_46116_13728# 0.518f
C1863 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 0.587f
C1864 X2.X2.X1.X2.X2.X1.X1.vin2 a_46502_8010# 8.88e-20
C1865 a_16836_8010# vdd 1.05f
C1866 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X3.vin2 0.165f
C1867 X2.X2.X1.X1.X3.vin2 a_48702_20446# 9.7e-20
C1868 a_19722_14688# d1 0.0422f
C1869 X1.X2.X2.X1.X3.vin2 a_22826_10734# 0.241f
C1870 X1.X2.X1.X1.X3.vin2 a_19722_22312# 0.423f
C1871 a_4696_26164# a_5082_26164# 0.414f
C1872 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.X1.vin2 0.23f
C1873 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X3.vin1 1.22e-19
C1874 a_19422_28070# a_19336_26164# 3.3e-19
C1875 a_19036_28070# a_19722_26164# 3.08e-19
C1876 X1.X1.X2.X1.X1.X2.X3.vin2 vdd 0.787f
C1877 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X3.vin1 0.0174f
C1878 a_54606_28888# d0 0.0489f
C1879 X2.X2.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X3.vin1 0.0321f
C1880 X1.X2.X2.vrefh X3.vin1 0.0274f
C1881 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.vout 0.118f
C1882 a_52106_10734# vdd 0.489f
C1883 X1.X1.X1.X3.vin2 a_4782_12822# 6.03e-19
C1884 a_10686_28888# X1.X1.X2.X2.X2.X2.X1.vin1 8.22e-20
C1885 X1.X1.X2.X2.X1.X2.X3.vin2 a_8872_24076# 0.101f
C1886 a_54606_15546# a_52492_14586# 2.68e-20
C1887 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X2.vrefh 0.076f
C1888 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X2.X1.vin2 3.94e-19
C1889 d2 a_23212_29834# 0.627f
C1890 X1.X2.X1.X1.X2.X2.X1.vin1 vdd 0.592f
C1891 X2.X2.X3.vin1 d1 0.0901f
C1892 X2.X1.X1.X2.X2.vrefh d1 0.00745f
C1893 X2.X2.X1.X2.X1.X2.vrefh d1 0.0071f
C1894 a_19336_26164# X1.X2.X1.X1.X3.vin1 0.169f
C1895 X2.X1.X2.X3.vin2 X2.X1.X2.X3.vin1 0.559f
C1896 a_38152_12640# a_37852_10734# 6.2e-19
C1897 a_39966_23170# X2.X1.X2.X2.X1.X1.X3.vin2 8.07e-19
C1898 X1.X2.X2.X2.vrefh d1 0.00964f
C1899 d1 X1.X1.X1.X2.X2.X2.vout 0.0331f
C1900 a_31476_8010# a_31476_6104# 0.00396f
C1901 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 0.242f
C1902 a_48616_7064# a_48702_5198# 3.38e-19
C1903 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.vrefh 0.267f
C1904 X1.X2.X2.X2.X3.vin1 a_23126_24076# 9.54e-19
C1905 a_49002_7064# a_48316_5198# 3.31e-19
C1906 a_25326_25076# a_25326_23170# 0.00198f
C1907 d0 X2.X1.X2.X1.X2.X2.X2.vin1 0.262f
C1908 a_52792_20264# d4 0.00161f
C1909 a_54606_9828# X2.X2.X2.X1.X1.X2.X2.vin1 0.402f
C1910 a_25326_30794# vdd 0.553f
C1911 X2.X1.X1.X2.X2.X1.X2.vin1 X2.X1.X1.X2.X2.X2.vrefh 0.564f
C1912 a_37766_8828# X2.X1.X2.X1.X1.X2.X3.vin1 0.42f
C1913 a_37852_14586# vdd 1.05f
C1914 X1.X2.X2.X2.X1.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin1 0.00437f
C1915 X2.X2.X2.X2.X2.X2.X1.vin2 a_54606_30794# 0.273f
C1916 X1.X1.X2.X2.X1.X1.vout a_8572_22210# 0.169f
C1917 d1 X1.X1.X2.X1.X1.X1.X1.vin1 0.013f
C1918 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X2.vin1 0.242f
C1919 a_48702_5198# vdd 0.47f
C1920 d3 X1.X2.X1.X1.X2.X1.X1.vin1 6.34e-20
C1921 a_4696_29936# X1.X1.X1.X1.X1.X2.X3.vin1 0.00329f
C1922 X1.X1.X2.X1.X2.vrefh d1 0.00745f
C1923 a_34362_29936# X2.X1.X1.X1.X3.vin1 0.434f
C1924 a_31476_15634# d1 2.92e-22
C1925 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X2.vrefh 0.267f
C1926 X1.X2.X1.X1.X1.X2.X2.vin1 d0 0.262f
C1927 X2.X1.X3.vin2 a_34362_14688# 2.04e-19
C1928 X1.X1.X2.X2.vrefh d1 0.00964f
C1929 d3 X1.X1.X1.X1.X1.X2.X3.vin2 0.0251f
C1930 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X3.vin1 0.00118f
C1931 X1.X2.X2.X1.X2.X2.X1.vin2 X1.X2.X2.X1.X2.X1.X3.vin2 3.94e-19
C1932 X1.X2.X2.X1.X2.X2.X1.vin1 a_25326_13640# 8.22e-20
C1933 a_31476_9916# X2.X1.X1.X2.X2.X1.X2.vin1 1.78e-19
C1934 a_39966_19358# X2.X1.X2.X2.vrefh 8.22e-20
C1935 X1.X2.X2.X1.X1.X2.X1.vin1 a_25712_7922# 0.195f
C1936 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 5.19e-19
C1937 a_38152_20264# d4 0.00161f
C1938 X1.X1.X2.X2.X1.X2.X2.vin1 a_11072_25076# 0.197f
C1939 a_37466_6962# X2.X1.X2.X1.X1.X1.vout 0.386f
C1940 a_23126_12640# a_22826_10734# 5.25e-20
C1941 a_2582_17540# X1.X1.X1.X2.X1.X1.X1.vin2 0.273f
C1942 d3 a_37466_25982# 0.292f
C1943 X1.X1.X3.vin1 a_4782_5198# 2.12e-19
C1944 a_16836_23258# d1 2.92e-22
C1945 a_34362_7064# vdd 0.477f
C1946 X2.X1.X2.X1.X2.X2.vout X2.X1.X2.X1.X2.X1.vout 0.514f
C1947 a_2582_25164# X1.X1.X1.X1.X2.X1.X3.vin1 0.52f
C1948 a_10686_23170# a_8572_22210# 2.68e-20
C1949 X2.X2.X2.X2.X1.X2.X3.vin1 a_54606_23170# 0.52f
C1950 a_49002_10916# X2.X2.X1.X2.X2.X1.X3.vin1 0.00837f
C1951 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X2.vrefh 0.00118f
C1952 a_4396_31882# a_4782_31882# 0.419f
C1953 X2.X2.X3.vin1 X2.X2.X3.vin2 3.25f
C1954 X2.X2.X1.X3.vin2 X2.X2.X2.X3.vin1 1.22e-19
C1955 a_23512_20264# d4 0.00161f
C1956 a_34062_24258# a_34362_22312# 4.19e-20
C1957 X1.X1.X2.X2.X2.X2.X2.vin1 d1 7.58e-19
C1958 X2.X1.X1.X1.X2.X1.vout a_33976_22312# 0.169f
C1959 X2.X2.X1.X1.X1.X2.vrefh d1 0.0738f
C1960 X2.X2.X1.X1.X2.X1.X2.vin1 a_46116_23258# 0.197f
C1961 a_8186_6962# a_8572_6962# 0.419f
C1962 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X1.vout 0.038f
C1963 a_23212_22210# a_23512_20264# 6.1e-19
C1964 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X2.X1.vin1 0.267f
C1965 X1.X2.X1.X2.X2.X2.X3.vin1 vdd 0.993f
C1966 X1.X2.X1.X2.X2.X2.X3.vin2 vdd 0.725f
C1967 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X3.vin2 8.93e-19
C1968 a_16836_32788# a_16836_30882# 0.00396f
C1969 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X1.X3.vin1 0.0131f
C1970 X1.X2.X2.X2.X1.X2.vrefh d0 0.848f
C1971 d3 a_33976_14688# 7.7e-20
C1972 X2.X1.X1.X2.X1.X2.X1.vin2 d1 0.00406f
C1973 X1.X2.X1.X3.vin2 vdd 0.716f
C1974 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X1.X3.vin1 0.00118f
C1975 a_37466_25982# X2.X1.X2.X3.vin2 0.452f
C1976 a_49002_26164# d1 0.0318f
C1977 d3 X1.X2.X1.X1.X2.X2.vout 8.47e-19
C1978 a_31476_30882# d1 2.92e-22
C1979 X1.X2.X1.X2.X1.X2.X3.vin1 d1 0.146f
C1980 X2.X2.X3.vin1 X2.X2.X2.X1.X1.X2.vout 1.71e-19
C1981 X2.X1.X1.X1.X2.vrefh a_31476_27070# 0.118f
C1982 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X3.vin2 1.42e-20
C1983 a_46116_28976# d1 2.25e-20
C1984 X1.X2.X2.X2.X1.X1.X1.vin2 X1.X2.X2.X2.vrefh 0.1f
C1985 d2 X2.X1.X1.X2.X1.X2.X1.vin1 0.0114f
C1986 X1.X2.X1.X1.X1.X2.X3.vin2 a_17222_25164# 8.07e-19
C1987 X2.X1.X2.X1.X3.vin1 a_37852_10734# 0.169f
C1988 d2 a_54992_28888# 0.00464f
C1989 X1.X2.X1.X2.X1.X2.X2.vin1 vdd 0.576f
C1990 a_39966_7922# vdd 0.553f
C1991 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 0.587f
C1992 X1.X1.X3.vin1 a_5082_7064# 9.8e-19
C1993 X2.X1.X1.X1.X1.X2.X3.vin2 a_33976_26164# 0.00535f
C1994 a_34062_28070# a_34362_26164# 4.41e-20
C1995 a_52406_8828# a_54606_7922# 4.2e-20
C1996 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X3.vin2 0.552f
C1997 d3 X2.X1.X2.X1.X2.X1.X1.vin2 3.99e-21
C1998 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 0.216f
C1999 d2 X2.X1.X2.X2.X2.X1.X3.vin2 0.177f
C2000 a_2196_19446# a_2196_17540# 0.00396f
C2001 a_19722_10916# a_19036_9010# 2.97e-19
C2002 a_19336_10916# a_19422_9010# 3.21e-19
C2003 a_31862_17540# d1 3.95e-19
C2004 X2.X1.X1.X1.X3.vin2 d4 0.0401f
C2005 a_34062_9010# a_33976_7064# 3.14e-19
C2006 a_33676_9010# a_34362_7064# 2.86e-19
C2007 X2.X1.X2.X1.X2.X1.vout d1 0.0238f
C2008 a_31476_6104# vdd 1.05f
C2009 X1.X2.X2.X2.X1.X1.X3.vin2 d4 6.94e-19
C2010 a_4396_12822# vdd 1.05f
C2011 X2.X2.X2.X2.X1.X2.vrefh a_54992_21264# 0.118f
C2012 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X3.vin2 0.552f
C2013 a_40352_25076# a_40352_23170# 0.00396f
C2014 a_40352_13640# a_40352_11734# 0.00396f
C2015 X1.X1.X2.X2.X2.X2.X3.vin2 a_8186_29834# 3.85e-19
C2016 a_54992_11734# d1 2.25e-20
C2017 a_25326_25076# vdd 0.542f
C2018 d2 a_46116_17540# 0.00256f
C2019 a_34362_22312# d1 0.0422f
C2020 a_46502_27070# vdd 0.542f
C2021 a_23212_22210# X1.X2.X2.X2.X1.X1.X3.vin2 0.00546f
C2022 a_2196_32788# d0 0.511f
C2023 a_37852_29834# X2.X1.X2.X2.X2.X1.X3.vin2 0.00546f
C2024 X1.X1.X2.X1.X2.X1.vout X1.X1.X2.X1.X2.X1.X3.vin2 0.326f
C2025 X2.X2.X1.X1.X2.X2.vrefh a_46502_21352# 8.22e-20
C2026 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X3.vin2 8.93e-19
C2027 d1 a_34062_5198# 0.0751f
C2028 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X1.X2.X2.vrefh 0.1f
C2029 X2.X1.X2.vrefh X2.X2.X2.vrefh 0.0959f
C2030 X2.X2.X2.X1.X2.X2.X1.vin1 d1 0.0118f
C2031 X2.X2.X2.X3.vin1 X2.X2.X1.X2.X3.vin2 7.46e-20
C2032 a_14082_892# X1.X3.vin2 0.255f
C2033 d0 X1.X1.X2.X1.X2.X1.X2.vin1 0.262f
C2034 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X1.X2.X2.X2.X2.vrefh 0.267f
C2035 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.vrefh 0.1f
C2036 X1.X2.X1.X1.X1.X2.X1.vin1 d0 0.267f
C2037 a_19722_10916# vdd 0.487f
C2038 a_31862_21352# X2.X1.X1.X1.X2.X2.X3.vin2 7.84e-19
C2039 X2.X1.X1.X1.X2.X2.X3.vin1 a_33676_20446# 0.199f
C2040 X1.X2.X2.X2.X2.X1.X1.vin2 vdd 0.36f
C2041 a_2196_21352# vdd 1.05f
C2042 X2.X2.X2.X1.X2.X2.vout a_52106_14586# 0.263f
C2043 a_39966_23170# d1 3.41e-19
C2044 d1 a_46502_8010# 0.00148f
C2045 a_37852_18358# d2 0.0113f
C2046 d2 a_38152_12640# 3.82e-19
C2047 d0 X1.X2.X1.X2.X1.X1.X1.vin2 0.276f
C2048 X2.X1.X2.X2.X1.X1.X1.vin1 d4 6.34e-20
C2049 a_48702_12822# X2.X2.X1.X2.X1.X2.X3.vin2 0.277f
C2050 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X3.vin1 0.199f
C2051 X2.X2.X1.X1.X1.X2.vout vdd 0.696f
C2052 X1.X1.X1.X1.X2.X1.vout d1 0.0238f
C2053 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.X1.vin1 2.23e-19
C2054 X2.X1.X2.X1.X2.X2.X2.vin1 a_40352_15546# 1.78e-19
C2055 a_52792_27888# d3 0.00178f
C2056 a_54992_23170# X2.X2.X2.X2.X1.X2.vrefh 1.64e-19
C2057 a_46116_19446# vdd 1.05f
C2058 a_54606_13640# X2.X2.X2.X1.X2.X1.X2.vin1 0.402f
C2059 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X3.vin2 8.93e-19
C2060 X1.X1.X2.X1.X3.vin2 vdd 1.32f
C2061 X1.X2.X2.vrefh X2.X1.X2.vrefh 0.0959f
C2062 a_33676_16634# d1 0.521f
C2063 X1.X2.X2.X2.X1.X1.X1.vin1 a_25712_17452# 1.64e-19
C2064 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X1.X3.vin1 0.0425f
C2065 X1.X1.X1.X2.X1.X1.X1.vin2 vdd 0.36f
C2066 X1.X2.X2.X2.X1.X1.X1.vin1 d4 6.34e-20
C2067 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X3.vin1 0.0131f
C2068 a_37766_16452# X2.X1.X2.X1.X3.vin2 9.7e-20
C2069 X2.X2.X2.X1.X1.X2.X3.vin2 d1 0.171f
C2070 X1.X2.X1.X3.vin1 a_19422_20446# 5.31e-19
C2071 X1.X2.X3.vin1 a_22826_14586# 2.24e-19
C2072 X2.X2.X1.X1.X2.X2.vrefh X2.X1.X2.X2.X1.X2.vrefh 0.117f
C2073 a_46116_27070# X2.X2.X1.X1.X1.X2.X1.vin2 1.78e-19
C2074 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X2.vout 0.197f
C2075 X2.X2.X2.X2.X2.X2.X1.vin1 d1 0.0118f
C2076 d3 a_19036_9010# 0.00178f
C2077 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 0.587f
C2078 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 0.216f
C2079 a_25326_9828# a_23512_8828# 1.15e-20
C2080 X1.X2.X1.X1.X2.X2.vrefh vdd 0.415f
C2081 a_37766_12640# a_39966_11734# 4.2e-20
C2082 a_52792_27888# X2.X2.X2.X2.X2.X1.X3.vin2 0.1f
C2083 d3 a_52106_14586# 9.23e-19
C2084 X2.X2.X2.X1.X2.X2.vout vdd 0.865f
C2085 X2.X2.X1.X1.X1.X2.X3.vin2 a_49002_26164# 0.00846f
C2086 X2.X1.X2.X2.X2.vrefh d1 0.00745f
C2087 a_48702_28070# X2.X2.X1.X3.vin1 1.64e-19
C2088 a_48702_24258# vdd 0.561f
C2089 X2.X2.X2.X1.X1.X2.vrefh vdd 0.43f
C2090 d0 d6 4.97e-19
C2091 X1.X1.X2.X2.X1.X1.X3.vin2 a_8872_20264# 0.1f
C2092 X2.X2.X1.X1.X1.X2.X2.vin1 X2.X2.X1.X1.X1.X2.X3.vin1 0.00117f
C2093 d3 X1.X1.X1.X1.X3.vin2 0.387f
C2094 X2.X1.X2.X2.X1.X1.X3.vin1 a_40352_19358# 0.354f
C2095 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X2.vrefh 0.076f
C2096 a_48702_28070# a_46502_28976# 4.2e-20
C2097 X2.X1.X2.X2.X1.X2.X3.vin2 a_37466_22210# 3.85e-19
C2098 d3 a_40352_32700# 2.56e-19
C2099 X1.X1.X2.X2.X1.X1.X1.vin1 d4 6.34e-20
C2100 X1.X2.X1.X1.X2.vrefh d3 6.65e-20
C2101 a_2582_23258# vdd 0.541f
C2102 a_2582_6104# vdd 0.553f
C2103 a_2582_21352# a_4782_20446# 4.2e-20
C2104 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X1.X2.X2.X2.vin1 0.00117f
C2105 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X2.vrefh 0.267f
C2106 X2.X1.X3.vin1 X2.X1.X2.X3.vin1 3.45e-19
C2107 X1.X2.X3.vin2 a_23126_5016# 2.33e-19
C2108 X2.X2.X1.X2.X3.vin2 X2.X2.X2.X1.X3.vin1 0.0604f
C2109 a_31862_27070# d1 0.00151f
C2110 X2.X1.X2.X2.X1.X2.vout vdd 0.697f
C2111 a_17222_32788# X1.X2.X1.X1.X1.X1.X2.vin1 8.88e-20
C2112 d2 a_10686_15546# 0.00393f
C2113 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X2.vrefh 0.1f
C2114 X2.X2.X2.X2.X1.X1.vout X2.X2.X2.X2.X1.X1.X3.vin2 0.342f
C2115 X2.X1.X1.X1.X1.X1.X1.vin2 d0 0.201f
C2116 a_37852_18358# a_38152_16452# 6.48e-19
C2117 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 0.242f
C2118 a_10686_6016# a_10686_4110# 0.00198f
C2119 X1.X1.X2.X1.X1.X2.vout vdd 0.696f
C2120 a_2582_13728# d1 3.41e-19
C2121 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X2.vrefh 0.076f
C2122 X2.X2.X2.X1.X2.X2.X3.vin2 a_54992_17452# 0.354f
C2123 a_52406_27888# a_52106_29834# 4.19e-20
C2124 a_33676_31882# d1 0.511f
C2125 a_48616_22312# a_46502_21352# 2.68e-20
C2126 a_22826_25982# X1.X2.X2.X2.X3.vin1 0.372f
C2127 X2.X2.X2.X1.X1.X1.X1.vin2 X2.X2.X2.X1.X1.X1.X1.vin1 0.668f
C2128 X1.X2.X1.X1.X3.vin2 X1.X2.X2.X3.vin2 7.46e-20
C2129 X2.X2.X1.X2.X3.vin1 a_48616_10916# 0.17f
C2130 X1.X2.X2.X1.X2.X1.X3.vin1 a_25712_11734# 0.354f
C2131 d2 a_16836_13728# 0.00351f
C2132 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X3.vin2 0.0523f
C2133 d2 X2.X1.X2.X1.X3.vin1 0.0619f
C2134 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X3.vin1 0.206f
C2135 X1.X1.X2.X2.X2.X1.X2.vin1 d1 1.03e-19
C2136 a_22826_10734# X1.X2.X2.X1.X3.vin1 0.385f
C2137 X1.X1.X3.vin2 a_8572_18358# 0.355f
C2138 d0 a_46502_9916# 0.0675f
C2139 d3 vdd 16.1f
C2140 d4 X1.X1.X1.X2.X1.X1.vout 0.00145f
C2141 a_25712_26982# a_25712_28888# 0.00396f
C2142 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.X1.X1.X1.vin2 3.94e-19
C2143 a_16836_32788# vdd 1.05f
C2144 a_11072_17452# a_11072_15546# 0.00396f
C2145 d2 a_25326_28888# 0.00665f
C2146 d2 a_10686_7922# 0.00479f
C2147 d3 a_34062_12822# 0.00122f
C2148 a_25712_23170# X1.X2.X2.X2.X1.X2.vrefh 1.64e-19
C2149 X1.X2.X2.X2.X1.X1.X3.vin1 a_25712_19358# 0.354f
C2150 X2.X2.X2.X2.X2.X2.vout vdd 0.698f
C2151 a_33976_29936# a_31862_30882# 2.95e-20
C2152 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X2.vin1 0.564f
C2153 a_4782_5198# X1.X1.X1.X2.X2.X2.X3.vin2 0.277f
C2154 X2.X2.X1.X2.X1.X2.X1.vin1 vdd 0.592f
C2155 X1.X1.X2.X3.vin1 a_8486_8828# 1.64e-19
C2156 d0 a_35312_892# 3.19e-19
C2157 a_54606_21264# d0 0.0489f
C2158 d0 a_2196_15634# 0.515f
C2159 a_10686_26982# d1 3.95e-19
C2160 d4 X2.X2.X1.X1.X1.X1.X1.vin2 8.21e-20
C2161 X2.X2.X2.X2.X1.X2.X3.vin2 a_54992_25076# 0.354f
C2162 d2 X2.X2.X2.X1.X2.X1.X1.vin2 0.231f
C2163 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.vout 0.075f
C2164 X1.X1.X1.X3.vin1 d4 1f
C2165 X2.X2.X2.X2.X1.X2.vrefh d1 0.0071f
C2166 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X2.vin1 0.564f
C2167 X2.X2.X2.X2.X2.X1.X3.vin2 vdd 0.903f
C2168 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X3.vin2 0.234f
C2169 a_14082_892# vdd 0.473f
C2170 X1.X2.X1.X1.X1.X2.X2.vin1 a_17222_27070# 0.402f
C2171 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X3.vin1 0.206f
C2172 X2.X1.X2.X3.vin2 vdd 0.716f
C2173 d2 a_10686_30794# 6.36e-19
C2174 X2.X1.X2.X1.X1.X1.X1.vin2 a_39966_4110# 0.273f
C2175 X2.X2.X2.X2.X1.X1.X3.vin1 d2 0.104f
C2176 X2.X1.X2.X2.X2.X1.X3.vin1 d0 4.36e-19
C2177 d0 X2.X2.X2.X1.X1.X1.X1.vin1 0.269f
C2178 a_52106_22210# a_52406_20264# 4.19e-20
C2179 a_49002_18540# X2.X2.X1.X2.X1.X1.X3.vin1 0.00837f
C2180 X1.X1.X2.vrefh vdd 0.704f
C2181 d0 a_2196_8010# 0.515f
C2182 a_19336_14688# a_19722_14688# 0.419f
C2183 X1.X2.X1.X2.X1.X2.vrefh a_17222_15634# 0.3f
C2184 a_23512_16452# a_25326_15546# 1.06e-19
C2185 X2.X1.X3.vin2 a_34362_10916# 3.68e-19
C2186 d2 X1.X2.X1.X2.X2.X2.vout 0.11f
C2187 a_8186_29834# X1.X1.X2.X2.X2.X1.X3.vin2 0.00815f
C2188 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X2.vrefh 0.267f
C2189 d3 X1.X2.vrefh 0.00665f
C2190 a_54606_26982# X2.X2.X2.X2.X2.vrefh 8.22e-20
C2191 a_2196_28976# d0 0.518f
C2192 d3 a_33676_9010# 0.00178f
C2193 d4 X1.X1.X1.X1.X1.X1.vout 0.0336f
C2194 X1.X1.X1.X2.X2.X2.vout a_4782_5198# 0.418f
C2195 a_5082_7064# X1.X1.X1.X2.X2.X2.X3.vin2 3.85e-19
C2196 X1.X1.X2.X1.X1.X1.X3.vin2 a_10686_7922# 8.07e-19
C2197 a_19722_29936# a_19422_31882# 4.19e-20
C2198 a_19336_29936# X1.X2.X1.X1.X1.X1.vout 0.169f
C2199 a_4396_20446# a_2582_19446# 1.15e-20
C2200 X2.X1.X2.X2.X1.X1.X3.vin1 d2 0.104f
C2201 X2.X1.X1.X2.X1.X2.vout a_33676_12822# 0.36f
C2202 a_40352_17452# X2.X1.X2.X1.X2.X2.X1.vin2 1.78e-19
C2203 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X1.vout 0.399f
C2204 a_19422_28070# vdd 0.47f
C2205 X1.X2.X2.X2.X1.X1.vout vdd 0.78f
C2206 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 0.0903f
C2207 d2 X1.X2.X2.X1.X2.X1.X1.vin1 0.0105f
C2208 a_23512_24076# a_22826_22210# 3.31e-19
C2209 d1 a_48316_9010# 0.521f
C2210 d0 X2.X2.X1.X2.X2.vrefh 0.848f
C2211 a_31862_23258# d2 0.00665f
C2212 X1.X2.X1.X2.X1.X1.X2.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 0.234f
C2213 X2.X1.X2.X2.X2.X1.X1.vin1 d3 6.34e-20
C2214 a_2196_30882# d0 0.515f
C2215 a_52492_10734# X2.X2.X2.X1.X1.X2.X3.vin2 0.00535f
C2216 X1.X2.X2.X1.X1.X2.X3.vin2 a_25712_9828# 0.354f
C2217 X1.X1.X3.vin2 d2 0.1f
C2218 X1.X1.X3.vin2 a_8186_10734# 6.66e-19
C2219 X1.X2.X2.X1.X1.X1.X1.vin2 X1.X2.X2.X1.X1.X1.X1.vin1 0.668f
C2220 a_31476_27070# a_31476_25164# 0.00396f
C2221 X1.X2.X1.X1.X3.vin1 vdd 0.805f
C2222 a_17222_21352# a_19036_20446# 1.06e-19
C2223 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X2.vin1 0.0689f
C2224 X1.X1.X1.X1.X2.X1.X2.vin1 d2 0.0318f
C2225 d0 X1.X2.X2.X1.X1.X1.X1.vin1 0.269f
C2226 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X3.vin1 0.206f
C2227 a_5082_26164# a_4782_24258# 5.25e-20
C2228 a_4696_26164# X1.X1.X1.X1.X2.X1.vout 1.64e-19
C2229 a_16836_19446# X1.X2.X1.X2.X1.X1.X1.vin1 1.64e-19
C2230 X2.X1.X1.X1.X2.vrefh a_31862_25164# 8.22e-20
C2231 X1.X2.X2.X2.X1.X1.X3.vin1 d2 0.104f
C2232 d3 a_33976_10916# 0.621f
C2233 a_39966_9828# d1 0.00151f
C2234 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.vout 0.399f
C2235 X2.X2.X1.X2.X1.X1.X3.vin2 a_46502_15634# 0.567f
C2236 a_49002_18540# X2.X2.X3.vin1 0.47f
C2237 X2.X1.X2.X1.X2.X1.X3.vin1 vdd 0.997f
C2238 d2 X2.X2.X1.X2.X2.X1.X1.vin2 0.231f
C2239 a_38152_20264# a_39966_19358# 1.06e-19
C2240 a_5082_7064# X1.X1.X1.X2.X2.X2.vout 0.263f
C2241 X2.X1.X1.X2.vrefh a_31862_19446# 0.3f
C2242 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin1 0.449f
C2243 X1.X2.X1.X1.X2.X1.X2.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 0.234f
C2244 X1.X1.X3.vin1 X1.X1.X1.X2.X1.X2.vout 3.08e-19
C2245 a_25326_32700# d4 8.99e-20
C2246 d0 a_17222_11822# 0.0489f
C2247 a_39966_28888# a_39966_30794# 0.00198f
C2248 a_25326_32700# a_23126_31700# 4.77e-21
C2249 d2 X2.X1.X1.X2.X2.X1.X3.vin1 0.104f
C2250 a_31862_21352# X2.X1.X1.X1.X2.X2.X1.vin2 0.273f
C2251 d2 a_25326_7922# 0.00479f
C2252 a_46116_21352# d1 2.25e-20
C2253 X1.X1.X2.X2.X1.X2.X3.vin1 d0 4.36e-19
C2254 d3 X1.X2.X1.X2.X1.X2.vout 0.0232f
C2255 a_37766_20264# a_37466_18358# 5.25e-20
C2256 a_54992_21264# d2 0.00414f
C2257 a_54606_25076# a_54606_23170# 0.00198f
C2258 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X1.vin1 0.0689f
C2259 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 0.242f
C2260 X2.X2.X2.X1.X2.X1.X3.vin2 a_54606_11734# 7.84e-19
C2261 a_48616_29936# a_46502_30882# 2.95e-20
C2262 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X3.vin2 0.234f
C2263 a_37852_10734# d1 0.0126f
C2264 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 2.23e-19
C2265 X1.X1.X1.X2.X2.X1.X1.vin2 a_2582_8010# 8.88e-20
C2266 a_10686_4110# X1.X1.X2.X1.X1.X1.X1.vin1 0.417f
C2267 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X1.vout 0.131f
C2268 a_54992_25076# d0 0.515f
C2269 X1.X1.X1.X1.X1.X2.X3.vin1 a_4782_28070# 0.42f
C2270 X1.X1.X2.X1.X1.X1.X1.vin2 a_11072_4110# 0.12f
C2271 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.X3.vin1 0.0174f
C2272 X1.X2.X1.X2.X2.X1.X2.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 0.234f
C2273 a_52406_27888# d4 2.4e-19
C2274 X2.X1.X2.X2.X1.X1.X3.vin2 d2 0.169f
C2275 a_5082_10916# X1.X1.X1.X2.X2.X1.X3.vin1 0.00837f
C2276 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X3.vin1 0.0131f
C2277 X1.X1.X2.X1.X1.X2.vout X1.X1.X2.X1.X1.X1.vout 0.507f
C2278 X2.X1.X1.X1.X1.X2.X2.vin1 d1 1.03e-19
C2279 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X3.vin2 0.0523f
C2280 d0 X2.X2.X1.X2.X2.X2.X1.vin1 0.267f
C2281 d0 a_25326_15546# 0.0675f
C2282 X2.X1.X2.X2.X1.X2.X3.vin2 d0 4.34e-19
C2283 X1.X2.X1.X2.X2.vrefh a_17222_11822# 0.3f
C2284 a_23512_12640# a_25326_11734# 1.06e-19
C2285 a_10686_26982# X1.X1.X2.X2.X1.X2.X3.vin2 8.07e-19
C2286 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin2 0.12f
C2287 a_52106_14586# X2.X2.X2.X1.X3.vin2 0.423f
C2288 X2.X1.X1.X1.X2.X1.X3.vin2 a_31476_23258# 0.354f
C2289 d3 X2.X2.X2.X2.X1.X2.vout 0.0232f
C2290 X2.X2.X1.X1.X2.X2.X3.vin1 a_46502_19446# 0.00207f
C2291 X2.X2.X2.X1.X2.X2.X1.vin1 a_54606_13640# 8.22e-20
C2292 X2.X2.X2.X1.X2.X2.X1.vin2 X2.X2.X2.X1.X2.X1.X3.vin2 3.94e-19
C2293 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X3.vin2 2.23e-19
C2294 a_19336_14688# X1.X2.X1.X2.X1.X2.X3.vin1 0.00329f
C2295 a_39966_17452# X2.X1.X2.X1.X2.X2.X3.vin2 0.567f
C2296 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X3.vin1 0.00118f
C2297 X1.X2.X1.X2.vrefh a_17222_19446# 0.3f
C2298 a_23512_20264# a_25326_19358# 1.06e-19
C2299 d0 a_25712_9828# 0.515f
C2300 X2.X2.X2.X2.X2.X2.vrefh d2 0.168f
C2301 a_52792_12640# a_52106_10734# 2.97e-19
C2302 d0 a_16836_8010# 0.515f
C2303 X1.X1.X1.X1.X1.X1.X1.vin1 vdd 0.596f
C2304 X1.X1.X1.X3.vin1 X1.X1.X2.X3.vin2 1.22e-19
C2305 d2 X1.X1.X1.X2.X3.vin2 0.0501f
C2306 a_49002_22312# d2 0.0191f
C2307 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X3.vin1 0.0131f
C2308 X1.X2.X2.X1.X2.X2.X1.vin1 X2.X1.X1.X2.X1.X2.vrefh 0.00437f
C2309 a_23512_31700# a_25326_30794# 1.06e-19
C2310 X1.X1.X1.X2.X1.X1.X3.vin2 a_5082_14688# 0.00815f
C2311 X1.X2.X1.X1.X1.X2.vrefh a_17222_30882# 0.3f
C2312 d0 X1.X1.X2.X1.X1.X2.X3.vin2 4.34e-19
C2313 X2.X2.X1.X2.X2.X1.X3.vin2 a_46502_6104# 8.07e-19
C2314 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X2.vrefh 0.00118f
C2315 a_31476_13728# vdd 1.05f
C2316 a_33976_29936# a_34062_31882# 3.14e-19
C2317 X2.vrefh X2.X1.X1.X1.X1.X1.X1.vin2 0.109f
C2318 a_34362_29936# a_33676_31882# 2.86e-19
C2319 d2 X2.X1.X2.X2.X3.vin2 0.0685f
C2320 X2.X2.X1.X3.vin1 a_48616_18540# 0.17f
C2321 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X2.vin1 0.0689f
C2322 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin2 0.12f
C2323 a_31862_13728# a_33676_12822# 1.06e-19
C2324 X2.X2.X1.X2.X1.X2.vout a_48702_12822# 0.418f
C2325 X2.X1.X1.X1.X2.X1.X3.vin1 a_33676_24258# 0.199f
C2326 X2.X2.X1.X1.X3.vin2 a_48702_24258# 0.00101f
C2327 a_49002_26164# X2.X2.X1.X1.X2.X1.X3.vin2 3.49e-19
C2328 a_2582_27070# d2 0.00792f
C2329 a_39966_28888# vdd 0.541f
C2330 a_40352_19358# d1 2.25e-20
C2331 a_23126_27888# a_23512_27888# 0.419f
C2332 d1 a_22826_6962# 0.0422f
C2333 X1.X2.X1.X1.X2.X2.X1.vin1 d0 0.267f
C2334 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin1 0.195f
C2335 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X1.X3.vin2 1.22e-19
C2336 d2 a_48316_12822# 6.04e-19
C2337 a_54992_23170# d2 0.00351f
C2338 X2.X2.X2.X2.X1.X1.X1.vin1 a_54992_19358# 0.195f
C2339 X1.X2.X1.X1.X1.X1.X2.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 0.234f
C2340 a_39966_25076# X2.X1.X2.X2.X1.X2.X3.vin2 0.567f
C2341 X2.X2.X2.X1.X3.vin2 vdd 1.32f
C2342 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X3.vin1 0.00118f
C2343 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X1.vin2 3.94e-19
C2344 X2.X1.X2.X2.X3.vin2 a_37852_29834# 0.363f
C2345 a_25326_30794# d0 0.0675f
C2346 X1.X1.X2.X2.X3.vin1 vdd 0.804f
C2347 a_8186_18358# a_8486_16452# 4.41e-20
C2348 X2.X1.X2.X2.X2.X2.X2.vin1 a_39966_30794# 8.88e-20
C2349 X2.X2.X1.X2.X1.X1.vout X2.X2.X1.X2.X1.X2.vout 0.507f
C2350 X1.X2.X2.X1.X2.X2.X2.vin1 vdd 0.576f
C2351 X1.X2.X2.X2.X1.X1.X3.vin2 a_25326_19358# 7.84e-19
C2352 a_25712_19358# d1 2.25e-20
C2353 X1.X2.X2.X2.X1.X1.X2.vin1 X1.X2.X2.X2.X1.X1.X1.vin1 0.0689f
C2354 a_8572_18358# d1 0.00638f
C2355 X2.X1.X2.X1.X2.X1.X1.vin1 X2.X2.X1.X2.X2.vrefh 0.00437f
C2356 X1.X2.X1.X3.vin1 X1.X2.X1.X3.vin2 0.552f
C2357 X2.X2.X1.X1.X2.X2.X2.vin1 a_46116_19446# 0.197f
C2358 X2.X2.X1.X1.X1.X1.X3.vin2 a_46502_30882# 0.567f
C2359 X1.X1.X1.X2.X2.X1.X3.vin1 a_4396_9010# 0.199f
C2360 a_10686_32700# X1.X1.X2.X2.X2.X2.X2.vin1 0.402f
C2361 X1.X2.X3.vin1 X1.X2.X1.X2.X3.vin2 0.0816f
C2362 d3 X2.X2.X1.X1.X3.vin2 0.433f
C2363 X2.X2.X1.X2.X2.X2.vout d2 0.11f
C2364 X2.X2.X2.X2.X1.X1.X3.vin1 a_52492_18358# 0.00255f
C2365 X1.X1.X1.X1.X2.X1.X3.vin2 a_2582_21352# 8.07e-19
C2366 a_31476_17540# a_31476_15634# 0.00396f
C2367 a_5082_14688# vdd 0.477f
C2368 d2 X2.X1.X2.X1.X2.X2.vout 0.00117f
C2369 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X2.X1.X2.X1.X1.X2.vin1 0.00232f
C2370 a_8572_29834# X1.X1.X2.X2.X2.X2.X3.vin1 0.00329f
C2371 d1 X2.X1.X2.X1.X1.X1.X2.vin1 0.0144f
C2372 a_11072_19358# d1 2.25e-20
C2373 X2.X1.X1.X1.X2.X1.X1.vin1 d1 0.0118f
C2374 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin2 0.12f
C2375 X2.X1.X2.X2.X1.X2.vout a_37466_22210# 0.254f
C2376 X2.X2.X1.X2.X2.X2.X1.vin2 a_46116_4198# 1.78e-19
C2377 a_39966_19358# X2.X1.X2.X2.X1.X1.X1.vin1 0.417f
C2378 X2.X1.X2.X2.X1.X1.X1.vin2 a_40352_19358# 0.12f
C2379 X1.X2.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X3.vin1 0.0321f
C2380 X2.X1.X2.X2.X2.X2.X2.vin1 a_40352_32700# 0.197f
C2381 d2 a_54606_6016# 4.64e-19
C2382 a_39966_32700# X2.X2.vrefh 0.3f
C2383 d2 a_4782_9010# 7.51e-19
C2384 a_5082_10916# X1.X1.X1.X2.X2.X1.X3.vin2 3.49e-19
C2385 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X2.vrefh 0.076f
C2386 a_46502_25164# d2 0.00328f
C2387 X2.X2.X2.X3.vin1 a_52406_16452# 5.31e-19
C2388 a_10686_9828# X1.X1.X2.X1.X1.X2.X3.vin2 0.567f
C2389 X1.X2.X2.X1.X1.X1.vout X1.X2.X2.X1.X1.X1.X3.vin1 0.118f
C2390 X1.X2.X2.vrefh a_20286_892# 7.23e-19
C2391 X1.X2.X1.X2.X2.X2.X3.vin1 d0 4.36e-19
C2392 d0 X1.X2.X1.X2.X2.X2.X3.vin2 4.34e-19
C2393 X1.X2.X2.X1.X2.X1.X3.vin2 a_25712_13640# 0.354f
C2394 a_46502_6104# a_48316_5198# 1.06e-19
C2395 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X2.vin1 0.0689f
C2396 d5 a_43362_892# 4.95e-19
C2397 a_52492_14586# X2.X2.X2.X1.X2.X1.X3.vin2 0.00546f
C2398 X2.X1.X3.vin1 vdd 0.854f
C2399 X2.X2.X2.X2.X2.X1.X1.vin1 d2 0.0105f
C2400 a_48616_26164# a_49002_26164# 0.414f
C2401 a_5646_892# vdd 1.05f
C2402 X2.X1.X2.X1.X2.X1.X3.vin2 a_37466_10734# 3.49e-19
C2403 d3 a_37466_22210# 0.0474f
C2404 a_48316_16634# X2.X2.X1.X2.X1.X1.X3.vin2 0.1f
C2405 X2.X2.X2.vrefh a_49952_892# 7.3e-19
C2406 a_2196_4198# vdd 1.05f
C2407 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X3.vin1 0.206f
C2408 X2.X1.X3.vin1 a_34062_12822# 2.12e-19
C2409 a_39966_26982# X2.X1.X2.X2.X2.X1.X2.vin1 8.88e-20
C2410 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X2.X1.X3.vin2 8.93e-19
C2411 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X2.X1.X1.X2.X1.X2.vin1 0.00232f
C2412 X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin2 0.0128f
C2413 X1.X1.X2.X2.X2.X2.X3.vin2 d4 1.57e-19
C2414 X1.X1.X1.X2.X2.X1.X1.vin1 d1 0.0118f
C2415 X1.X1.X2.X2.X2.vrefh a_11072_25076# 0.118f
C2416 d2 a_48702_31882# 9.83e-19
C2417 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X2.vrefh 0.00118f
C2418 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 2.23e-19
C2419 d2 a_17222_9916# 0.00328f
C2420 a_38152_27888# a_37466_25982# 2.97e-19
C2421 d0 X1.X2.X1.X2.X1.X2.X2.vin1 0.262f
C2422 X2.X1.X2.X2.X2.X2.X2.vin1 vdd 0.578f
C2423 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X2.vin1 0.242f
C2424 X2.X1.X1.X1.X1.X2.X3.vin1 X2.X1.X1.X1.X1.X2.X1.vin2 0.216f
C2425 d0 a_39966_7922# 0.0675f
C2426 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.X1.vin1 2.23e-19
C2427 X1.X2.X2.X2.X2.X2.X1.vin1 X2.X1.X1.X1.X1.X2.vrefh 0.00437f
C2428 X1.X1.X2.X2.X2.X2.X2.vin1 a_11072_30794# 1.78e-19
C2429 a_8486_8828# a_8572_6962# 3.38e-19
C2430 X1.X1.X2.X2.X1.X1.X2.vin1 d1 1.03e-19
C2431 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin1 0.195f
C2432 X1.X1.X3.vin1 X1.X3.vin1 0.273f
C2433 a_48616_29936# a_48316_31882# 6.1e-19
C2434 X2.X2.X1.X3.vin1 d4 0.509f
C2435 a_54606_32700# d1 0.00148f
C2436 a_25326_21264# d2 0.0059f
C2437 a_25326_19358# X1.X2.X2.X2.X1.X1.X1.vin1 0.417f
C2438 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X2.X1.X2.X2.X1.X2.vin1 0.00232f
C2439 d2 X2.X1.X2.X2.X2.X2.vout 0.102f
C2440 X1.X2.X2.X2.X1.X1.X1.vin2 a_25712_19358# 0.12f
C2441 d2 d1 29.2f
C2442 a_8186_10734# d1 0.0318f
C2443 X2.X1.X2.X1.X2.X2.X3.vin1 a_39966_15546# 0.52f
C2444 X2.X1.X2.X3.vin2 a_37466_22210# 0.00292f
C2445 a_19722_26164# X1.X2.X1.X1.X3.vin2 0.241f
C2446 d0 a_31476_6104# 0.518f
C2447 X2.X2.X1.X2.X2.X1.X3.vin1 vdd 0.997f
C2448 a_25326_25076# d0 0.0489f
C2449 a_46502_27070# d0 0.0489f
C2450 a_2582_27070# a_4396_28070# 1.15e-20
C2451 d3 a_19422_24258# 0.00195f
C2452 a_23126_12640# X1.X2.X2.X1.X2.X1.X3.vin1 0.428f
C2453 X2.X1.X2.X1.X2.X2.vout a_38152_16452# 0.36f
C2454 X2.X1.X1.X2.X1.X1.X2.vin1 a_31476_15634# 0.197f
C2455 X1.X2.X1.X2.X1.X2.X2.vin1 X1.X2.X1.X2.X2.vrefh 0.564f
C2456 d2 X2.X2.X1.X1.X1.X1.X3.vin1 0.00317f
C2457 a_33676_24258# X2.X1.X1.X1.X2.X1.X3.vin2 0.1f
C2458 a_37852_29834# d1 0.00613f
C2459 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 2.23e-19
C2460 a_37852_29834# X2.X1.X2.X2.X2.X2.vout 0.0929f
C2461 d2 X2.X2.X2.X1.X1.X1.X3.vin1 3e-19
C2462 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X3.vin1 0.546f
C2463 a_37466_14586# X2.X1.X2.X1.X2.X1.vout 0.383f
C2464 X1.X2.X2.X1.X2.X2.X2.vin1 X2.X1.X1.X2.X1.X1.X1.vin2 0.00232f
C2465 X2.X2.X2.X2.X1.X1.X3.vin2 vdd 0.905f
C2466 a_31476_17540# a_31862_17540# 0.419f
C2467 d4 X2.X1.X1.X2.X1.X1.X1.vin1 6.34e-20
C2468 a_23512_8828# vdd 1.05f
C2469 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X3.vin1 0.587f
C2470 X2.X1.X3.vin2 a_34926_892# 0.0927f
C2471 a_17222_17540# d1 3.95e-19
C2472 X1.X1.X2.X2.X1.X1.vout X1.X1.X2.X2.X1.X1.X3.vin2 0.342f
C2473 a_54606_19358# d2 0.00309f
C2474 a_19036_28070# a_17222_28976# 1.06e-19
C2475 X1.X2.X1.X1.X1.X2.X2.vin1 X1.X2.X1.X1.X1.X2.X1.vin1 0.0689f
C2476 X2.X2.X2.X1.X2.X1.X1.vin1 a_54992_11734# 0.195f
C2477 a_4396_9010# X1.X1.X1.X2.X2.X1.X3.vin2 0.1f
C2478 a_33676_28070# a_33976_29936# 6.71e-19
C2479 X2.X1.X2.X1.X1.X2.X1.vin1 a_40352_6016# 1.64e-19
C2480 X2.X1.X1.X1.X2.X2.vout d4 9.49e-19
C2481 X2.X2.X1.X2.vrefh a_46502_17540# 8.22e-20
C2482 d3 X2.X2.X2.X2.X1.X2.X3.vin2 0.0247f
C2483 a_38152_8828# a_39966_7922# 1.06e-19
C2484 a_34362_26164# vdd 0.489f
C2485 a_33976_22312# a_34362_22312# 0.419f
C2486 a_4696_22312# a_2582_21352# 2.68e-20
C2487 X2.X1.X1.X2.X2.X2.vrefh a_31862_8010# 0.3f
C2488 X1.X2.X2.X2.X1.X2.vout d1 0.033f
C2489 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 0.139f
C2490 a_8486_20264# a_8186_18358# 5.25e-20
C2491 a_19036_9010# a_19336_7064# 6.1e-19
C2492 X1.X2.X2.X1.X1.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin2 0.0128f
C2493 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X3.vin2 8.93e-19
C2494 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.vout 0.038f
C2495 a_10686_19358# X1.X1.X2.X2.X1.X1.X1.vin1 0.417f
C2496 X1.X1.X2.X2.X1.X1.X1.vin2 a_11072_19358# 0.12f
C2497 d2 X1.X1.X2.X2.X2.X1.vout 0.115f
C2498 a_2196_21352# d0 0.518f
C2499 X2.X2.X3.vin2 d2 0.1f
C2500 X1.X2.X2.X2.X2.X1.X1.vin2 d0 0.276f
C2501 X2.X1.X2.X2.X1.X1.X1.vin2 d2 0.231f
C2502 X1.X1.X2.X1.X1.X1.X3.vin2 d1 0.154f
C2503 X1.X2.X3.vin2 d5 0.0348f
C2504 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X2.X1.X1.X1.X1.X2.vin1 0.00232f
C2505 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X1.X3.vin2 5.19e-19
C2506 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X1.vin2 0.076f
C2507 X1.X2.X2.X2.X1.X2.X2.vin1 X2.X1.X1.X1.X2.X1.X1.vin2 0.00232f
C2508 a_31476_25164# a_31862_25164# 0.419f
C2509 X1.X1.X1.X1.X1.X2.X1.vin1 vdd 0.592f
C2510 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.X3.vin1 0.587f
C2511 a_10686_23170# X1.X1.X2.X2.X1.X1.X3.vin2 8.07e-19
C2512 X2.X1.X1.X2.X2.X1.X2.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 0.234f
C2513 X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.vout 2.91e-19
C2514 a_52106_6962# d1 0.0422f
C2515 d3 X1.X2.X2.X1.X1.X2.X3.vin2 0.0251f
C2516 a_23126_16452# X1.X2.X2.X1.X2.X2.vout 0.418f
C2517 X1.X2.X2.X1.X2.X1.vout vdd 0.805f
C2518 a_46502_11822# vdd 0.542f
C2519 X1.X1.X2.X2.X1.X2.X1.vin1 d2 0.0114f
C2520 a_38152_16452# d1 0.521f
C2521 a_52406_24076# d4 2.4e-19
C2522 X1.X2.X2.X2.X2.X1.vout a_23212_29834# 0.169f
C2523 X2.X1.X1.X2.X2.X2.X2.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 0.234f
C2524 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X3.vin1 2.33e-19
C2525 a_46116_19446# d0 0.515f
C2526 a_33676_5198# a_34062_5198# 0.419f
C2527 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X1.X1.vin1 0.206f
C2528 X1.X1.X3.vin2 a_8486_5016# 2.33e-19
C2529 d2 X2.X2.X2.X1.X1.X2.vout 0.106f
C2530 X1.X2.X2.X2.X1.X1.X1.vin2 d2 0.231f
C2531 X2.X2.X2.X1.X1.X1.vout a_52406_5016# 0.422f
C2532 a_54606_15546# X2.X2.X2.X1.X2.X2.X1.vin1 0.417f
C2533 X2.X2.X2.X1.X2.X2.X1.vin2 a_54992_15546# 0.12f
C2534 X1.X1.X1.X2.X1.X1.X1.vin2 d0 0.276f
C2535 a_5082_18540# d2 0.00132f
C2536 X1.X2.X2.X2.X2.X2.X2.vin1 d1 7.58e-19
C2537 a_48316_31882# X2.X2.X1.X1.X1.X1.X3.vin2 0.1f
C2538 a_2582_13728# a_2582_11822# 0.00198f
C2539 X1.X1.X1.X3.vin1 X1.X1.X3.vin1 0.188f
C2540 a_8872_12640# d1 0.521f
C2541 X1.X1.X1.X3.vin2 a_5082_10916# 0.452f
C2542 X1.X2.X1.X1.X2.X2.vrefh d0 0.848f
C2543 a_46116_15634# vdd 1.05f
C2544 a_31862_17540# X2.X1.X1.X2.X1.X1.X2.vin1 8.88e-20
C2545 a_19336_7064# vdd 1.05f
C2546 d4 a_34062_16634# 0.00142f
C2547 d3 X1.X2.X1.X3.vin1 0.702f
C2548 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 0.242f
C2549 d1 X1.X2.X1.X2.X2.X2.X1.vin2 0.0985f
C2550 a_10686_21264# a_10686_19358# 0.00198f
C2551 d0 X2.X2.X2.X1.X1.X2.vrefh 0.844f
C2552 a_23126_24076# X1.X2.X2.X2.X1.X2.vout 0.418f
C2553 a_16836_25164# d1 2.25e-20
C2554 X1.X1.X2.X2.X1.X1.X1.vin2 d2 0.231f
C2555 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X1.X3.vin1 0.0321f
C2556 a_8486_12640# a_8186_10734# 5.25e-20
C2557 X2.X2.X2.X2.X2.X1.X3.vin1 d1 0.151f
C2558 a_19422_9010# a_17222_8010# 4.77e-21
C2559 a_25712_25076# d2 0.00533f
C2560 X1.X2.X3.vin2 X1.X2.X1.X2.X2.X2.vout 1.5e-19
C2561 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 5.19e-19
C2562 a_4396_28070# d1 0.521f
C2563 a_2582_23258# d0 0.0489f
C2564 a_2196_9916# a_2582_9916# 0.419f
C2565 a_2582_6104# d0 0.0675f
C2566 X1.X2.X2.X1.X2.X1.X1.vin2 vdd 0.36f
C2567 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin2 7.84e-19
C2568 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin2 0.12f
C2569 a_19036_5198# X1.X2.X1.X2.X2.X2.X3.vin2 0.101f
C2570 X1.X2.X1.X2.X2.X2.X3.vin1 a_19036_5198# 0.199f
C2571 X2.X1.X2.X2.X2.X2.X3.vin1 a_39966_30794# 0.52f
C2572 X2.X2.X3.vin2 a_52106_6962# 0.00111f
C2573 X1.X1.X2.X2.X1.X2.X3.vin2 d2 0.121f
C2574 a_17222_6104# X1.X2.X1.X2.X2.X2.X3.vin1 0.52f
C2575 d4 X1.X2.X2.X1.X2.X2.vout 6.95e-19
C2576 d2 X1.X1.X1.X1.X2.vrefh 0.158f
C2577 a_23126_8828# X1.X2.X2.X1.X1.X2.vout 0.418f
C2578 a_4782_16634# X1.X1.X1.X2.X1.X1.vout 0.422f
C2579 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X1.X1.vin1 2.23e-19
C2580 a_49002_7064# X2.X2.X1.X2.X2.X2.X3.vin1 0.00874f
C2581 X2.X2.X1.X1.X1.X2.X3.vin2 d2 0.122f
C2582 a_10686_13640# X1.X1.X2.X1.X2.X1.X3.vin2 0.567f
C2583 X2.X1.X2.X2.X2.X2.vout a_38152_31700# 0.36f
C2584 X2.X1.X2.X2.X1.X2.X1.vin2 a_39966_23170# 0.273f
C2585 d3 a_52792_12640# 0.00178f
C2586 a_8572_10734# X1.X1.X2.X1.X1.X2.X3.vin2 0.00535f
C2587 X2.X1.X2.X1.X2.X2.X3.vin1 vdd 0.962f
C2588 X2.X1.X1.X1.X1.X1.X2.vin1 a_31476_30882# 0.197f
C2589 X1.X1.X1.X1.X2.X2.X2.vin1 d4 8.68e-20
C2590 d3 a_5082_22312# 9.23e-19
C2591 a_46116_8010# a_46502_8010# 0.419f
C2592 a_38152_31700# d1 0.515f
C2593 X1.X1.X2.X2.X1.X1.X1.vin1 a_11072_17452# 1.64e-19
C2594 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.vout 0.2f
C2595 a_25712_15546# vdd 1.05f
C2596 d2 a_52492_10734# 0.0057f
C2597 a_11072_32700# X1.X1.X2.X2.X2.X2.X1.vin2 1.78e-19
C2598 X1.X2.X2.X2.X2.X1.X2.vin1 a_25712_28888# 0.197f
C2599 d3 d0 7.67e-19
C2600 d2 a_4396_16634# 3.82e-19
C2601 a_48702_28070# a_48616_29936# 3.38e-19
C2602 a_48316_28070# a_49002_29936# 3.31e-19
C2603 a_52106_6962# X2.X2.X2.X1.X1.X2.vout 0.254f
C2604 a_16836_32788# d0 0.511f
C2605 a_22826_14586# X1.X2.X2.X1.X2.X1.X3.vin2 0.00815f
C2606 X1.X1.X2.X2.X2.X2.X2.vin1 a_8872_31700# 5.34e-19
C2607 a_17222_28976# X1.X2.X1.X1.X1.X2.X3.vin1 0.52f
C2608 X2.X1.X2.X2.X2.X2.vout X2.X1.X2.X2.X2.X2.X3.vin2 0.08f
C2609 a_46116_30882# vdd 1.05f
C2610 d1 a_40352_4110# 5.03e-20
C2611 X2.X1.X2.X2.X2.X2.X3.vin2 d1 0.0135f
C2612 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin2 0.1f
C2613 d4 a_34062_31882# 2.4e-19
C2614 a_4782_24258# X1.X1.X1.X1.X2.X1.vout 0.422f
C2615 a_31862_9916# vdd 0.553f
C2616 X3.vin2 a_43362_892# 0.472f
C2617 d0 X2.X2.X1.X2.X1.X2.X1.vin1 0.267f
C2618 a_25326_6016# X1.X2.X2.X1.X1.X1.X3.vin1 0.00207f
C2619 X2.X1.X2.X1.X2.vrefh d1 0.00745f
C2620 a_4696_26164# d2 0.0057f
C2621 a_19336_22312# d1 0.00613f
C2622 a_19422_28070# X1.X2.X1.X3.vin1 1.64e-19
C2623 X1.X2.X1.X1.X1.X2.X3.vin2 a_19722_26164# 0.00846f
C2624 a_5082_26164# X1.X1.X1.X3.vin1 0.509f
C2625 X2.X2.X2.X2.X3.vin1 vdd 0.804f
C2626 a_11072_25076# a_11072_23170# 0.00396f
C2627 d3 X1.X2.X1.X2.X2.vrefh 6.65e-20
C2628 X2.X2.X2.X2.X2.X1.X3.vin2 d0 4.34e-19
C2629 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X1.vin2 0.076f
C2630 d0 a_14082_892# 1.37e-19
C2631 d4 X1.X2.X2.X2.X2.X2.vout 0.0955f
C2632 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X1.vout 0.0524f
C2633 X1.X2.X3.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 8.36e-19
C2634 a_39966_21264# vdd 0.541f
C2635 a_23126_31700# X1.X2.X2.X2.X2.X2.vout 0.418f
C2636 X1.X1.X2.X2.X3.vin2 d1 0.00807f
C2637 a_31862_11822# d1 0.00151f
C2638 a_52492_18358# d1 0.00638f
C2639 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X2.X1.vin1 5.19e-19
C2640 d2 a_34362_29936# 0.254f
C2641 X2.X1.X2.X2.X2.X2.X3.vin1 vdd 0.993f
C2642 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X3.vin1 0.199f
C2643 a_38152_27888# vdd 1.05f
C2644 X1.X2.X1.X1.X2.X2.vrefh a_16836_21352# 1.64e-19
C2645 d2 a_37466_6962# 0.272f
C2646 a_31862_8010# a_31862_6104# 0.00198f
C2647 d0 X1.X1.X2.vrefh 4.73f
C2648 a_31476_8010# X2.X1.X1.X2.X2.X2.X1.vin1 1.64e-19
C2649 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 0.242f
C2650 a_49002_7064# X2.X2.X1.X2.X2.X2.X3.vin2 3.85e-19
C2651 a_25326_13640# a_25326_11734# 0.00198f
C2652 X1.X2.X2.X2.X1.X2.X3.vin2 a_25326_23170# 7.84e-19
C2653 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 0.234f
C2654 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X1.vin1 0.0689f
C2655 d3 a_39966_25076# 1.89e-19
C2656 X2.X2.X1.X2.vrefh d4 6.65e-20
C2657 d3 a_38152_8828# 0.00108f
C2658 a_54606_30794# X2.X2.X2.X2.X2.X2.X1.vin1 0.417f
C2659 a_8572_6962# a_8872_5016# 6.1e-19
C2660 a_8486_12640# a_8872_12640# 0.419f
C2661 a_25712_30794# vdd 1.05f
C2662 X2.X2.X2.X2.X2.X2.X1.vin2 a_54992_30794# 0.12f
C2663 d2 a_4396_31882# 0.00167f
C2664 a_49002_14688# vdd 0.477f
C2665 a_23126_27888# a_22826_29834# 4.19e-20
C2666 a_4696_10916# vdd 1.05f
C2667 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.X3.vin1 0.0174f
C2668 a_25326_11734# a_23212_10734# 5.36e-21
C2669 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 0.049f
C2670 a_11072_11734# a_11072_9828# 0.00396f
C2671 a_37852_22210# vdd 1.05f
C2672 d1 a_52792_8828# 0.521f
C2673 a_54606_19358# a_52492_18358# 5.36e-21
C2674 X1.X2.X2.X3.vin1 d2 6.42e-19
C2675 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X2.vin1 0.0689f
C2676 a_49002_26164# X2.X2.X1.X1.X2.X1.X3.vin1 0.00837f
C2677 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 5.19e-19
C2678 X1.X1.X1.X2.X2.X2.X1.vin2 d2 7.2e-20
C2679 a_31862_9916# a_33676_9010# 1.06e-19
C2680 X2.X2.X1.X1.X2.vrefh a_46502_27070# 0.3f
C2681 a_40352_19358# X2.X1.X2.X2.vrefh 1.64e-19
C2682 X1.X2.X2.X1.X1.X2.X1.vin2 X2.X1.X1.X2.X2.X1.X2.vin1 0.00232f
C2683 d3 a_10686_9828# 1.89e-19
C2684 X2.X3.vin2 a_49952_892# 0.684f
C2685 a_23212_18358# a_25326_17452# 4.72e-20
C2686 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X1.vin2 0.216f
C2687 a_54606_26982# a_52492_25982# 5.36e-21
C2688 a_10686_11734# d1 3.95e-19
C2689 a_48316_20446# X2.X2.X1.X1.X2.X2.X3.vin2 0.101f
C2690 X1.X2.X2.X3.vin2 a_23126_20264# 5.21e-19
C2691 a_39966_17452# a_37766_16452# 4.77e-21
C2692 a_54606_23170# vdd 0.553f
C2693 X2.X2.X2.X2.X1.X2.X3.vin1 a_54992_23170# 0.354f
C2694 X2.X2.X3.vin2 a_52492_18358# 0.355f
C2695 X1.X1.X2.X2.X2.X1.vout X1.X1.X2.X2.X3.vin2 0.399f
C2696 a_4782_31882# X1.X1.X1.X1.X1.X1.vout 0.422f
C2697 a_52406_27888# X2.X2.X2.X3.vin2 7.93e-20
C2698 a_48316_24258# a_46502_23258# 1.15e-20
C2699 X2.X1.X1.X1.X2.X1.vout X2.X1.X1.X1.X2.X2.vout 0.514f
C2700 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 0.0565f
C2701 d0 X2.X1.X2.X1.X2.X1.X3.vin1 4.36e-19
C2702 X1.X2.X1.X1.X2.X1.X3.vin2 vdd 0.903f
C2703 a_31476_32788# d4 1.8e-19
C2704 d1 a_43362_892# 2.34e-19
C2705 a_33976_10916# a_31862_9916# 5.36e-21
C2706 X2.X2.X1.X2.X1.X1.X2.vin1 vdd 0.576f
C2707 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.vout 0.335f
C2708 a_17222_32788# a_17222_30882# 0.00198f
C2709 X2.X1.X2.X1.X2.X1.X2.vin1 d1 1.03e-19
C2710 d3 X2.X1.X1.X2.X3.vin1 0.375f
C2711 a_16836_9916# X1.X2.X1.X2.X2.X1.X2.vin1 1.78e-19
C2712 X1.X2.X3.vin2 a_20672_892# 0.239f
C2713 a_31476_27070# a_31862_27070# 0.419f
C2714 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 0.242f
C2715 d2 a_54606_13640# 0.00665f
C2716 a_39966_6016# a_39966_4110# 0.00198f
C2717 X1.X1.X2.X2.X1.X2.vout vdd 0.697f
C2718 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X1.X2.X1.X1.X2.vrefh 0.1f
C2719 X2.X2.X1.X1.X1.X2.X1.vin1 d1 0.0118f
C2720 X2.X2.X2.X1.X1.X2.X3.vin1 vdd 0.96f
C2721 X1.X2.X2.X2.X1.X1.X1.vin1 X1.X2.X2.X2.vrefh 0.267f
C2722 a_34062_20446# a_33976_18540# 3.3e-19
C2723 a_33676_20446# a_34362_18540# 3.08e-19
C2724 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.X1.X3.vin1 1.22e-19
C2725 a_33676_20446# X2.X1.X1.X1.X2.X2.X3.vin2 0.101f
C2726 a_10686_6016# X1.X1.X2.X1.X1.X1.X2.vin1 0.402f
C2727 a_19422_12822# vdd 0.47f
C2728 X2.X1.X1.X1.X2.X1.X2.vin1 vdd 0.576f
C2729 a_4696_26164# a_4396_28070# 6.48e-19
C2730 a_40352_7922# vdd 1.05f
C2731 X2.X1.X1.X1.X1.X2.X1.vin2 X2.X1.X1.X1.X1.X1.X3.vin2 3.94e-19
C2732 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.X1.vin1 0.206f
C2733 X2.X2.X1.X2.X1.X1.X1.vin2 d1 1.49e-19
C2734 a_2196_13728# a_2582_13728# 0.419f
C2735 d3 X2.X1.X2.X1.X2.X1.X1.vin1 6.34e-20
C2736 a_40352_25076# vdd 1.05f
C2737 X1.X1.X1.X2.X2.X1.X2.vin1 vdd 0.576f
C2738 X1.X2.X1.X2.X3.vin2 a_19422_9010# 0.00101f
C2739 X2.X1.X1.X3.vin2 a_34062_16634# 5.21e-19
C2740 a_34362_18540# X2.X1.X1.X2.X1.X1.X3.vin2 3.49e-19
C2741 a_2196_19446# X1.X1.X1.X2.X1.X1.X1.vin1 1.64e-19
C2742 a_2582_19446# a_2582_17540# 0.00198f
C2743 d1 a_8486_5016# 0.0752f
C2744 X2.X1.X1.X2.X1.X1.X3.vin1 d1 0.146f
C2745 X2.X2.X1.X2.X2.X1.X2.vin1 a_46502_8010# 0.402f
C2746 X2.X2.X2.X1.X1.X2.vout a_52792_8828# 0.36f
C2747 X2.X1.X1.X2.X2.X1.vout a_34362_7064# 0.383f
C2748 a_2196_32788# a_2196_30882# 0.00396f
C2749 X2.X1.X2.X1.X3.vin2 a_37466_10734# 0.241f
C2750 a_22826_25982# d2 7.13e-19
C2751 X2.X1.X1.X2.X2.X2.X1.vin1 vdd 0.592f
C2752 X1.X1.X1.X2.X1.X2.X3.vin2 vdd 0.787f
C2753 d2 X2.X2.X1.X2.X1.X1.X1.vin1 0.0116f
C2754 X1.X2.X2.X2.X1.X2.X3.vin2 vdd 0.787f
C2755 d2 a_22826_10734# 7.13e-19
C2756 X2.X2.X2.X2.X2.X1.X1.vin2 vdd 0.36f
C2757 X2.X1.X1.X1.X3.vin2 a_34362_22312# 0.423f
C2758 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.vout 0.326f
C2759 a_49566_892# vdd 1.05f
C2760 X1.X1.X2.X1.X2.X2.vout X1.X1.X2.X1.X2.X1.vout 0.514f
C2761 d2 a_4782_5198# 0.00202f
C2762 X1.X1.X1.X1.X1.X1.X1.vin1 d0 0.0488f
C2763 a_4696_18540# X1.X1.X1.X3.vin2 0.0927f
C2764 a_10686_28888# X1.X1.X2.X2.X2.X1.X2.vin1 0.402f
C2765 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X3.vin2 8.93e-19
C2766 X2.X1.X2.X1.X1.X2.vrefh a_40352_6016# 0.118f
C2767 a_17222_28976# X1.X2.X1.X1.X1.X2.vrefh 8.22e-20
C2768 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X1.vin2 3.94e-19
C2769 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.vout 0.326f
C2770 X2.X2.X1.X1.X1.X1.X2.vin1 vdd 0.578f
C2771 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X3.vin1 2.33e-19
C2772 a_37766_27888# X2.X1.X2.X2.X2.X1.vout 0.422f
C2773 d2 X2.X2.X2.X2.X2.X1.vout 0.115f
C2774 d0 a_31476_13728# 0.518f
C2775 a_11072_9828# vdd 1.05f
C2776 X1.X2.X2.X2.X2.X1.X3.vin1 d2 0.104f
C2777 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X2.vout 0.398f
C2778 a_34362_14688# X2.X1.X1.X2.X1.X2.vout 0.254f
C2779 d3 X2.X1.X2.X2.X1.X2.X3.vin1 2.1e-19
C2780 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X1.X2.X2.vrefh 0.267f
C2781 d6 a_35312_892# 0.00114f
C2782 a_2196_17540# X1.X1.X1.X2.X1.X1.X2.vin1 1.78e-19
C2783 X1.X1.X2.X1.X3.vin2 a_8572_10734# 0.0927f
C2784 d2 a_19336_14688# 0.526f
C2785 X1.X2.X2.X1.X1.X2.X3.vin1 a_22826_6962# 0.00874f
C2786 a_19036_20446# X1.X2.X1.X1.X2.X2.X3.vin2 0.101f
C2787 a_39966_28888# d0 0.0489f
C2788 X2.X1.X2.X2.vrefh d2 0.173f
C2789 d3 X1.X1.X2.X1.X1.X2.X3.vin1 2.1e-19
C2790 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.X1.X2.vin1 0.242f
C2791 X2.X1.X1.X2.X3.vin2 a_34362_7064# 0.422f
C2792 a_10686_26982# a_10686_28888# 0.00198f
C2793 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.vrefh 0.267f
C2794 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 0.216f
C2795 a_8486_12640# a_10686_11734# 4.2e-20
C2796 X2.X2.X2.X2.X1.X2.X3.vin1 d1 0.146f
C2797 d3 X2.vrefh 0.00665f
C2798 a_52406_12640# a_54606_11734# 4.2e-20
C2799 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X2.X1.X1.vin2 0.216f
C2800 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 0.587f
C2801 X2.X1.X1.X2.X1.X2.X2.vin1 d1 1.03e-19
C2802 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X3.vin1 0.449f
C2803 X1.X1.X1.X1.X2.X2.X1.vin1 vdd 0.592f
C2804 X2.X2.X3.vin1 X2.X2.X1.X2.X1.X2.vout 3.08e-19
C2805 X1.X2.X2.X2.X2.X1.X1.vin1 vdd 0.592f
C2806 d4 a_22826_29834# 0.00116f
C2807 X2.X1.X1.X2.X1.X2.vrefh a_31862_13728# 8.22e-20
C2808 d1 X2.X2.X2.X1.X1.X2.X1.vin2 0.00406f
C2809 a_40352_23170# d1 2.25e-20
C2810 a_37766_8828# X2.X1.X2.X1.X1.X2.vout 0.418f
C2811 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.vrefh 2.33e-19
C2812 a_49002_18540# d2 0.00132f
C2813 X1.X2.X3.vin2 d1 0.0804f
C2814 a_46502_32788# vdd 0.554f
C2815 X1.X2.X1.X2.X1.X1.X3.vin2 a_17222_15634# 0.567f
C2816 d0 X1.X2.X2.X1.X2.X2.X2.vin1 0.262f
C2817 a_22826_29834# a_23126_31700# 5.55e-20
C2818 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin1 0.195f
C2819 a_52492_10734# a_52792_8828# 6.48e-19
C2820 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin2 7.84e-19
C2821 d2 a_5082_7064# 0.254f
C2822 X1.X1.X2.X2.X2.X1.X1.vin2 a_10686_26982# 0.273f
C2823 X2.X2.X1.X1.X2.X1.X3.vin2 d2 0.171f
C2824 a_39966_9828# X2.X1.X2.X1.X1.X2.X3.vin1 0.00207f
C2825 d3 X1.X2.X1.X2.X1.X1.vout 0.00883f
C2826 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X3.vin1 0.0131f
C2827 X2.X2.X1.X1.X2.vrefh d3 6.65e-20
C2828 d3 X1.X1.X1.X1.X2.X1.X1.vin1 6.34e-20
C2829 d3 a_8486_27888# 0.00195f
C2830 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 0.234f
C2831 a_2582_11822# X1.X1.X1.X2.X2.X1.X1.vin1 8.22e-20
C2832 X2.X1.X1.X2.X1.X1.vout d1 0.0238f
C2833 X2.X1.X2.X2.X2.X1.X1.vin1 a_40352_25076# 1.64e-19
C2834 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.vout 0.335f
C2835 a_8186_22210# vdd 0.477f
C2836 a_8186_25982# a_8486_24076# 4.41e-20
C2837 X1.X1.X2.X1.X2.X2.X2.vin1 vdd 0.576f
C2838 d4 a_19336_18540# 0.63f
C2839 a_8572_10734# X1.X1.X2.X1.X1.X2.vout 7.93e-20
C2840 a_34926_892# X2.X3.vin1 0.354f
C2841 a_2582_25164# X1.X1.X1.X1.X2.X1.X1.vin2 0.273f
C2842 d3 X1.X2.X1.X2.X2.X1.vout 0.00146f
C2843 X2.X2.X2.X2.X2.X1.X3.vin2 X2.X2.X2.X2.X2.X2.X3.vin1 1.22e-19
C2844 X2.X1.X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X2.X1.X1.vin1 0.206f
C2845 X1.X2.X2.X1.X1.X2.X3.vin2 a_23512_8828# 0.101f
C2846 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X2.vrefh 0.076f
C2847 a_31862_19446# vdd 0.541f
C2848 d2 a_2582_11822# 0.00792f
C2849 a_8872_24076# a_8572_22210# 6.71e-19
C2850 a_23126_5016# vdd 0.562f
C2851 X2.X2.X1.X3.vin1 X2.X2.X2.X3.vin2 1.22e-19
C2852 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X1.X2.X1.vin1 2.23e-19
C2853 X1.X2.X1.X2.X1.X2.vout a_19422_12822# 0.418f
C2854 d3 a_8572_10734# 0.621f
C2855 a_48702_28070# X2.X2.X1.X1.X1.X2.X3.vin1 0.42f
C2856 a_17222_27070# d3 1.89e-19
C2857 X2.X1.X3.vin1 d0 0.04f
C2858 a_4396_20446# d1 0.521f
C2859 d0 a_5646_892# 2.73e-19
C2860 a_25326_17452# X1.X2.X2.X1.X2.X2.X1.vin2 8.88e-20
C2861 d2 X1.X2.X2.X1.X2.X2.X3.vin1 0.153f
C2862 X1.X1.X2.X2.X1.X2.X1.vin2 vdd 0.361f
C2863 X2.X1.X2.X3.vin1 a_37852_18358# 0.17f
C2864 X1.X1.X1.X2.vrefh d2 0.173f
C2865 d0 a_2196_4198# 0.515f
C2866 X2.X2.X1.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X1.X1.vin2 0.076f
C2867 X1.X1.X1.X1.X2.X2.X3.vin1 a_4782_20446# 0.42f
C2868 a_52792_31700# X2.X2.X2.X2.X2.X2.X2.vin1 5.34e-19
C2869 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 2.23e-19
C2870 a_10686_32700# d2 1.95e-19
C2871 X1.X1.X1.X2.X2.X2.X3.vin1 vdd 0.993f
C2872 X1.X1.X1.X2.X1.X2.vrefh d1 0.0071f
C2873 X1.X2.X2.X1.X2.X2.vrefh vdd 0.415f
C2874 X1.X1.X2.X1.X1.X1.X1.vin2 X1.X2.X2.vrefh 0.0128f
C2875 X1.X2.X3.vin1 a_19722_7064# 9.8e-19
C2876 d2 a_11072_15546# 0.00274f
C2877 X2.X1.X2.X2.X2.X1.X1.vin2 d1 4.01e-19
C2878 d3 X1.X2.X1.X1.X1.X1.vout 0.0408f
C2879 X1.X2.X1.X2.X1.X2.X1.vin2 d1 0.00406f
C2880 a_37466_25982# X2.X1.X2.X2.X2.X1.X3.vin2 3.49e-19
C2881 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.X2.vin1 0.00117f
C2882 a_17222_32788# a_19422_31882# 4.2e-20
C2883 X1.X2.X2.X1.X2.X2.vout X1.X2.X2.X1.X3.vin2 0.0866f
C2884 a_17222_19446# vdd 0.541f
C2885 a_46116_11822# a_46116_9916# 0.00396f
C2886 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X1.vin1 0.0689f
C2887 X2.X2.X1.X2.X2.vrefh a_46502_9916# 8.22e-20
C2888 X2.X1.X2.X2.X2.X2.X2.vin1 d0 0.199f
C2889 X1.X1.X2.X1.X1.X1.X3.vin2 a_10686_4110# 7.84e-19
C2890 X1.X1.X1.X2.X1.X2.X3.vin1 d1 0.146f
C2891 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X3.vin2 8.93e-19
C2892 X2.X1.X1.X1.X1.X2.X2.vin1 a_31476_27070# 0.197f
C2893 a_48616_22312# X2.X2.X1.X1.X2.X2.X3.vin1 0.00329f
C2894 X2.X1.X1.X1.X1.X1.vout d1 0.0238f
C2895 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X1.vout 0.118f
C2896 a_48616_26164# d2 0.0057f
C2897 a_31476_28976# d1 2.25e-20
C2898 d2 a_40352_28888# 0.00464f
C2899 d2 X1.X2.X1.X2.X1.X2.X1.vin1 0.0114f
C2900 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X3.vin2 0.552f
C2901 a_54606_4110# a_54992_4110# 0.419f
C2902 d2 X1.X2.X2.X1.X1.X2.X3.vin1 0.157f
C2903 X1.X1.X1.X2.X2.X1.X3.vin2 a_4696_7064# 0.00546f
C2904 X1.X1.X2.X2.X1.X2.vrefh vdd 0.414f
C2905 X1.X2.X1.X1.X1.X1.X1.vin1 vdd 0.596f
C2906 d0 X2.X2.X1.X2.X2.X1.X3.vin1 4.36e-19
C2907 a_2582_19446# vdd 0.541f
C2908 d2 X1.X2.X2.X2.X2.X1.X3.vin2 0.177f
C2909 d2 a_11072_7922# 0.00351f
C2910 X2.X2.X1.X2.X2.X2.vout X2.X2.X1.X2.X2.X1.vout 0.514f
C2911 X2.X2.X2.X2.X3.vin2 d1 0.00807f
C2912 a_8486_16452# X1.X1.X2.X1.X3.vin2 9.7e-20
C2913 X1.X1.X2.X2.X1.X1.X3.vin2 d4 6.94e-19
C2914 a_10686_25076# vdd 0.542f
C2915 d2 a_31476_17540# 0.00256f
C2916 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X2.vrefh 0.564f
C2917 d2 a_37466_14586# 0.0191f
C2918 X2.X2.X2.X2.X1.X1.X3.vin2 d0 4.34e-19
C2919 a_11072_26982# d1 2.25e-20
C2920 d2 X2.X2.X2.X1.X2.X1.X1.vin1 0.0105f
C2921 a_48316_28070# vdd 1.05f
C2922 a_48702_12822# a_48616_10916# 3.3e-19
C2923 a_48316_12822# a_49002_10916# 3.08e-19
C2924 a_33976_22312# d2 0.526f
C2925 d2 X1.X2.X2.X2.X2.X2.X3.vin1 0.0571f
C2926 a_52106_22210# d4 2.94e-19
C2927 X1.X1.X1.X1.X1.X2.vrefh d1 0.0738f
C2928 X2.X2.X2.X3.vin2 a_52406_24076# 6.03e-19
C2929 X1.X2.X1.X1.X1.X1.X3.vin2 a_17222_30882# 0.567f
C2930 a_52492_14586# a_52406_12640# 3.14e-19
C2931 a_37466_22210# a_37852_22210# 0.419f
C2932 X3.vin1 a_28482_892# 0.426f
C2933 a_19422_28070# a_17222_27070# 4.77e-21
C2934 X1.X2.X1.X1.X1.X2.X3.vin2 a_16836_27070# 0.354f
C2935 X1.X2.X2.X2.X2.X2.vrefh vdd 0.415f
C2936 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 2.23e-19
C2937 X1.X2.X2.X1.X2.X1.X1.vin1 a_25326_9828# 8.22e-20
C2938 X1.X2.X2.X1.X2.X1.X1.vin2 X1.X2.X2.X1.X1.X2.X3.vin2 3.94e-19
C2939 a_39966_4110# X2.X1.X2.X1.X1.X1.X1.vin1 0.417f
C2940 X2.X1.X2.X1.X1.X1.X1.vin2 a_40352_4110# 0.12f
C2941 d2 a_33676_5198# 0.00393f
C2942 X2.X2.X2.X2.X1.X1.vout X2.X2.X2.X2.X1.X1.X3.vin1 0.118f
C2943 a_5082_29936# d1 0.0422f
C2944 a_4782_20446# a_4696_18540# 3.3e-19
C2945 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X3.vin1 0.199f
C2946 a_19722_14688# X1.X2.X1.X2.X3.vin1 0.436f
C2947 a_2196_28976# a_2196_30882# 0.00396f
C2948 a_4396_20446# a_5082_18540# 3.08e-19
C2949 d2 a_54606_15546# 0.00393f
C2950 X2.X1.X1.X2.vrefh d1 0.00964f
C2951 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X2.vin1 0.564f
C2952 a_8572_18358# a_8872_16452# 6.48e-19
C2953 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin2 1.42e-20
C2954 d3 X2.X1.X1.X2.X2.X1.vout 0.00146f
C2955 X1.X1.X1.X1.X1.X2.X1.vin1 d0 0.267f
C2956 a_54992_26982# X2.X2.X2.X2.X2.vrefh 1.64e-19
C2957 X1.X2.vrefh X1.X2.X1.X1.X1.X1.X1.vin1 0.108f
C2958 X2.X1.X3.vin2 X2.X1.X2.X1.X2.X2.X3.vin2 0.0011f
C2959 a_33976_29936# X2.X1.X1.X1.X1.X2.vout 0.0929f
C2960 X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 0.0565f
C2961 X1.X1.X1.X1.X2.X2.X3.vin2 a_2582_19446# 0.567f
C2962 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.vout 0.13f
C2963 d0 a_46502_11822# 0.0489f
C2964 X2.X1.X1.X2.X1.X2.vout X2.X1.X1.X2.X1.X2.X3.vin2 0.075f
C2965 d4 X2.X2.X1.X2.X1.X1.X3.vin2 4.77e-19
C2966 d2 a_46116_8010# 0.00464f
C2967 d1 X2.X2.X1.X2.X2.X1.vout 0.0238f
C2968 X2.X1.X2.X2.X1.X2.X1.vin2 d2 0.226f
C2969 d4 a_37466_18358# 0.281f
C2970 X2.X1.X3.vin1 X2.X1.X1.X2.X3.vin1 7.18e-19
C2971 a_19422_16634# X1.X2.X1.X2.X1.X1.X3.vin2 0.267f
C2972 X1.X2.X1.X2.vrefh d1 0.00964f
C2973 a_31862_32788# d1 2.7e-19
C2974 d3 a_8486_16452# 4.67e-19
C2975 a_23212_29834# vdd 1.05f
C2976 a_31476_27070# X2.X1.X1.X1.X2.X1.X1.vin1 1.64e-19
C2977 X1.X2.X1.X1.X2.X2.X3.vin1 a_19036_20446# 0.199f
C2978 a_16836_15634# a_16836_13728# 0.00396f
C2979 a_31862_27070# a_31862_25164# 0.00198f
C2980 a_25326_4110# a_25712_4110# 0.419f
C2981 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin2 7.84e-19
C2982 a_25326_9828# a_25326_7922# 0.00198f
C2983 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X1.vin2 0.242f
C2984 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin1 0.195f
C2985 a_54992_9828# d1 2.92e-22
C2986 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 1.22e-19
C2987 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X1.vout 0.038f
C2988 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X3.vin1 2.33e-19
C2989 a_38152_16452# a_37466_14586# 3.31e-19
C2990 d0 a_46116_15634# 0.515f
C2991 d2 X2.X1.X1.X2.X1.X1.X2.vin1 0.031f
C2992 d3 X2.X1.X1.X2.X3.vin2 0.156f
C2993 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X3.vin2 8.93e-19
C2994 X2.X1.X1.X2.X2.vrefh a_31476_11822# 0.118f
C2995 X2.X1.X2.X1.X1.X2.X3.vin2 d1 0.171f
C2996 X2.X2.X2.X2.X2.X2.X1.vin2 X2.X2.X2.X2.X2.X2.X2.vin1 0.242f
C2997 a_54606_30794# a_54606_32700# 0.00198f
C2998 X1.X1.X3.vin2 a_8186_14586# 3.67e-19
C2999 d2 X2.X2.X2.X1.X1.X2.X2.vin1 0.0329f
C3000 X2.X2.X1.X1.X1.X2.X2.vin1 X2.X2.X1.X1.X1.X2.X1.vin2 0.242f
C3001 d2 X2.X1.X2.X1.X1.X2.X3.vin1 0.157f
C3002 d2 a_54606_30794# 6.36e-19
C3003 a_54606_28888# X2.X2.X2.X2.X2.X1.X3.vin2 0.567f
C3004 X2.X1.X3.vin2 a_37766_12640# 2.33e-19
C3005 X1.X2.X2.X2.X2.X2.X3.vin2 d4 0.0535f
C3006 a_19422_24258# X1.X2.X1.X1.X2.X1.X3.vin2 0.267f
C3007 d0 X1.X2.X2.X1.X2.X1.X1.vin2 0.276f
C3008 X2.X1.X2.X2.X2.X1.X3.vin2 a_39966_30794# 8.07e-19
C3009 X1.X2.X2.X2.X2.X2.X3.vin2 a_23126_31700# 0.277f
C3010 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X2.vin1 0.242f
C3011 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X1.X2.X2.X1.vin2 0.216f
C3012 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X3.vin1 0.00117f
C3013 X2.X2.X1.X1.X2.X2.X1.vin1 d1 0.0118f
C3014 d2 a_25712_7922# 0.00351f
C3015 a_8186_25982# X1.X1.X2.X2.X2.X1.X3.vin1 0.00837f
C3016 X1.X2.X1.X1.X1.X2.X2.vin1 d3 8.68e-20
C3017 X1.X2.X3.vin1 a_20286_892# 0.17f
C3018 X2.X1.X1.X1.X1.X2.X1.vin1 X1.X2.X2.X2.X2.X2.vrefh 0.00437f
C3019 d0 X2.X1.X2.X1.X2.X2.X3.vin1 4.36e-19
C3020 X2.X2.X2.X2.X1.X2.X3.vin2 a_54606_23170# 7.84e-19
C3021 a_23126_16452# a_23212_14586# 3.38e-19
C3022 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X1.vin1 0.0689f
C3023 X2.X2.X3.vin2 X2.X2.X1.X2.X2.X1.vout 4.93e-20
C3024 X1.X1.X2.X1.X1.X1.X1.vin1 a_11072_4110# 0.195f
C3025 a_49002_10916# d1 0.0316f
C3026 a_19422_9010# X1.X2.X1.X2.X2.X1.X3.vin2 0.267f
C3027 X1.X2.X2.X2.X1.X1.X1.vin2 X2.X1.X1.X2.vrefh 0.0128f
C3028 X1.X2.X2.X3.vin1 X1.X2.X3.vin2 1.16f
C3029 d2 a_8872_16452# 6.04e-19
C3030 d4 a_4782_28070# 2.4e-19
C3031 d0 a_25712_15546# 0.518f
C3032 a_31476_27070# d2 0.00533f
C3033 a_34062_28070# d1 0.0749f
C3034 a_31476_15634# a_31862_15634# 0.419f
C3035 d3 a_8486_31700# 4.75e-19
C3036 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X1.vin2 0.668f
C3037 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X1.X3.vin2 0.0943f
C3038 a_46116_30882# d0 0.515f
C3039 d2 a_2196_13728# 0.00351f
C3040 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 5.19e-19
C3041 X1.X1.X2.X3.vin2 a_8572_25982# 0.355f
C3042 d2 X2.X1.X1.X1.X1.X1.X2.vin1 6e-20
C3043 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X3.vin1 0.0174f
C3044 X2.X2.X2.X2.vrefh d1 0.00964f
C3045 d0 a_31862_9916# 0.0675f
C3046 a_8572_29834# a_8872_27888# 6.1e-19
C3047 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X1.X2.X1.X2.vrefh 0.1f
C3048 d2 a_10686_28888# 0.00665f
C3049 X2.X1.X1.X2.X1.X2.X1.vin2 a_31476_11822# 1.78e-19
C3050 X2.X1.X1.X1.X2.X1.X1.vin2 a_31476_23258# 1.78e-19
C3051 a_23512_8828# a_23212_6962# 6.71e-19
C3052 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.X3.vin1 1.22e-19
C3053 X2.X2.X2.X1.X2.X1.X3.vin1 d1 0.151f
C3054 a_40352_21264# a_40352_19358# 0.00396f
C3055 X2.X1.X1.X2.X1.X2.X1.vin1 vdd 0.592f
C3056 X2.X2.X2.X1.X1.X1.X2.vin1 a_54992_6016# 0.197f
C3057 X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin2 0.0128f
C3058 a_54992_28888# vdd 1.05f
C3059 a_33976_29936# a_31862_28976# 2.68e-20
C3060 X1.X2.X2.X2.X2.X1.vout d1 0.0238f
C3061 a_34362_29936# X2.X1.X1.X1.X1.X1.vout 0.386f
C3062 d3 a_8186_18358# 0.0469f
C3063 a_39966_21264# d0 0.0489f
C3064 X2.X1.X1.X1.X3.vin1 a_34062_31882# 1.52e-19
C3065 X2.X2.X1.X3.vin1 X2.X2.X3.vin1 0.188f
C3066 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X1.vin2 0.668f
C3067 X2.X1.X1.X2.X1.X2.X3.vin1 a_33676_12822# 0.199f
C3068 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X2.X1.X2.vrefh 0.0128f
C3069 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin2 7.84e-19
C3070 X2.X2.X3.vin2 a_49002_10916# 3.68e-19
C3071 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.vout 0.118f
C3072 d2 X1.X1.X1.X2.X1.X2.vout 0.00124f
C3073 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin1 0.52f
C3074 X1.X1.X2.X2.X2.X1.X1.vin2 d2 0.231f
C3075 X2.X1.X2.X2.X2.X1.X3.vin2 vdd 0.903f
C3076 X2.X1.X2.X2.X2.X2.X3.vin1 d0 4.36e-19
C3077 X1.X2.X2.X1.X2.X2.X1.vin2 X1.X2.X2.X1.X2.X2.X1.vin1 0.668f
C3078 a_19722_22312# d4 1.99e-19
C3079 d2 X2.X2.X1.X2.X1.X2.X3.vin2 0.121f
C3080 a_16836_23258# a_17222_23258# 0.419f
C3081 a_52792_20264# d2 3.82e-19
C3082 a_54606_19358# X2.X2.X2.X2.vrefh 8.22e-20
C3083 a_40352_9828# a_40352_7922# 0.00396f
C3084 X2.X2.X2.X2.X2.X1.X1.vin1 a_54606_25076# 8.22e-20
C3085 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X1.X2.X3.vin2 3.94e-19
C3086 a_19422_31882# X1.X2.X1.X1.X1.X1.X3.vin2 0.267f
C3087 d2 a_8872_31700# 0.00293f
C3088 X2.X1.X1.X2.X2.X1.X3.vin2 a_31862_8010# 0.567f
C3089 d5 X1.X3.vin2 0.0478f
C3090 a_25712_30794# d0 0.518f
C3091 X2.X1.X2.X2.X3.vin1 a_37766_20264# 1.52e-19
C3092 a_54606_17452# a_52792_16452# 1.15e-20
C3093 a_46116_17540# vdd 1.05f
C3094 X1.X2.X1.X1.X2.X1.X2.vin1 d1 1.03e-19
C3095 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 0.0903f
C3096 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X1.vout 0.399f
C3097 X1.X1.X1.X2.X2.X2.X2.vin1 vdd 0.578f
C3098 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X3.vin1 0.0131f
C3099 X2.X1.X2.X2.X2.X2.X2.vin1 a_40352_30794# 1.78e-19
C3100 X1.X2.X2.X3.vin2 a_22826_18358# 0.263f
C3101 X1.X2.X2.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin1 0.00437f
C3102 d3 a_8486_20264# 4.67e-19
C3103 a_19722_18540# d1 0.0424f
C3104 X1.X2.X3.vin2 a_22826_10734# 6.66e-19
C3105 a_19036_28070# a_19722_29936# 3.31e-19
C3106 a_19422_28070# a_19336_29936# 3.38e-19
C3107 a_48316_20446# a_46502_19446# 1.15e-20
C3108 a_38152_20264# d2 3.82e-19
C3109 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X3.vin2 0.237f
C3110 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.vout 0.118f
C3111 a_31862_4198# vdd 0.541f
C3112 a_8486_5016# a_10686_4110# 4.2e-20
C3113 X1.X1.X2.X1.X1.X1.X3.vin1 X1.X1.X2.X1.X1.X1.X1.vin2 0.22f
C3114 X1.X2.X2.X1.X1.X2.X1.vin2 X1.X2.X2.X1.X1.X1.X3.vin2 3.94e-19
C3115 X1.X2.X2.X1.X1.X2.X1.vin1 a_25326_6016# 8.22e-20
C3116 a_54606_25076# d1 0.00151f
C3117 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X3.vin1 1.22e-19
C3118 a_31862_17540# a_31862_15634# 0.00198f
C3119 a_19336_29936# X1.X2.X1.X1.X3.vin1 0.363f
C3120 a_54606_23170# d0 0.0675f
C3121 d2 X2.X2.X1.X2.X2.X1.X2.vin1 0.0318f
C3122 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X1.vin2 0.668f
C3123 X2.X1.X2.X2.X1.X1.X1.vin1 a_40352_19358# 0.195f
C3124 d2 X2.X2.X2.X1.X1.X1.X3.vin2 0.0682f
C3125 a_23512_20264# d2 3.82e-19
C3126 a_46502_28976# X2.X2.X1.X1.X1.X2.vrefh 8.22e-20
C3127 X2.X2.X1.X1.X2.X1.X3.vin1 d2 0.104f
C3128 d4 X1.X1.X1.X3.vin2 0.134f
C3129 X1.X2.X1.X1.X2.X1.X3.vin2 d0 4.34e-19
C3130 a_23212_25982# a_25326_25076# 4.72e-20
C3131 a_4696_29936# a_4782_31882# 3.14e-19
C3132 a_5082_29936# a_4396_31882# 2.86e-19
C3133 a_38152_12640# vdd 1.05f
C3134 a_46502_6104# X2.X2.X1.X2.X2.X2.X3.vin2 7.84e-19
C3135 X1.X2.X2.vrefh d7 3.76e-19
C3136 a_37852_18358# vdd 1.05f
C3137 X2.X2.X1.X2.X2.X2.X3.vin1 a_48316_5198# 0.199f
C3138 d2 X1.X1.X2.X1.X2.X2.vrefh 0.168f
C3139 d0 X2.X2.X1.X2.X1.X1.X2.vin1 0.262f
C3140 a_19336_7064# a_19036_5198# 6.71e-19
C3141 a_25326_9828# d1 0.00151f
C3142 a_49002_26164# X2.X2.X1.X3.vin1 0.509f
C3143 a_17222_6104# a_19336_7064# 2.68e-20
C3144 a_31476_30882# a_31862_30882# 0.419f
C3145 X2.X2.X1.X2.X1.X1.vout X2.X2.X1.X2.X1.X1.X3.vin2 0.342f
C3146 a_40352_26982# X2.X1.X2.X2.X2.X1.X2.vin1 1.78e-19
C3147 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.X1.X3.vin2 2.23e-19
C3148 d2 X2.X1.X1.X2.X2.X1.X1.vin2 0.231f
C3149 X2.X1.X1.X1.X2.X2.X2.vin1 a_31862_19446# 0.402f
C3150 a_34362_18540# X2.X1.X3.vin2 6.58e-20
C3151 X1.X2.X1.X2.X2.X1.X2.vin1 X1.X2.X1.X2.X2.X2.vrefh 0.564f
C3152 a_46116_28976# a_46502_28976# 0.419f
C3153 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X2.X1.X1.X1.X2.X1.vin2 0.00232f
C3154 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 1.22e-19
C3155 d0 X2.X2.X2.X1.X1.X2.X3.vin1 4.36e-19
C3156 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X3.vin1 0.00118f
C3157 d3 a_37466_29834# 0.00329f
C3158 d2 X1.X2.X1.X2.X2.X1.X3.vin1 0.104f
C3159 X1.X2.X2.X2.X1.X1.X2.vin1 a_25712_21264# 0.197f
C3160 a_31476_21352# d1 2.25e-20
C3161 X2.X1.X1.X1.X2.X1.X2.vin1 d0 0.262f
C3162 d0 a_40352_7922# 0.518f
C3163 a_40352_21264# d2 0.00414f
C3164 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.vout 0.398f
C3165 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X2.vout 0.2f
C3166 a_17222_21352# X1.X2.X1.X1.X2.X2.X3.vin1 0.52f
C3167 a_40352_25076# d0 0.515f
C3168 d0 X1.X1.X1.X2.X2.X1.X2.vin1 0.262f
C3169 d1 a_46502_4198# 0.0015f
C3170 X2.X1.X2.X1.X1.X2.vout X2.X1.X2.X1.X1.X1.vout 0.507f
C3171 d3 a_48702_20446# 4.67e-19
C3172 X2.X1.X1.X1.X3.vin2 d2 0.00194f
C3173 a_48616_29936# X2.X2.X1.X1.X1.X1.vout 0.169f
C3174 a_19336_26164# d1 0.0126f
C3175 a_49002_29936# a_48702_31882# 4.19e-20
C3176 X1.X2.X2.X2.X1.X1.X1.vin1 a_25712_19358# 0.195f
C3177 a_25712_6016# a_25712_4110# 0.00396f
C3178 X1.X2.X2.X2.X1.X1.X3.vin2 d2 0.169f
C3179 X2.X2.X2.X2.X2.X2.X3.vin2 d1 0.0135f
C3180 d0 X2.X1.X1.X2.X2.X2.X1.vin1 0.267f
C3181 X2.X2.X1.X1.X2.X2.X1.vin2 a_46502_19446# 8.88e-20
C3182 X2.X1.X2.X1.X2.X2.X3.vin1 a_40352_15546# 0.354f
C3183 X2.X1.X2.X1.X1.X2.X3.vin2 a_37466_6962# 3.85e-19
C3184 X2.X2.X2.X2.X1.X1.vout d1 0.0238f
C3185 d0 X1.X1.X1.X2.X1.X2.X3.vin2 4.34e-19
C3186 X1.X2.X2.X2.X1.X2.X3.vin2 d0 4.34e-19
C3187 a_2582_27070# X1.X1.X1.X1.X1.X2.X3.vin2 0.567f
C3188 X2.X2.X2.X2.X2.X1.X1.vin2 d0 0.276f
C3189 X1.X2.X1.X2.X1.X2.X2.vin1 a_17222_11822# 0.402f
C3190 a_39966_17452# a_40352_17452# 0.419f
C3191 a_33676_16634# a_31862_15634# 1.15e-20
C3192 d0 a_49566_892# 2.73e-19
C3193 X1.X2.X2.X2.X2.X2.X1.vin2 X1.X2.X2.X2.X2.X2.X1.vin1 0.668f
C3194 a_16836_27070# X1.X2.X1.X1.X1.X2.X1.vin2 1.78e-19
C3195 a_37466_25982# X2.X1.X2.X2.X3.vin2 0.263f
C3196 d4 a_54606_17452# 1.89e-19
C3197 X2.X1.X1.X1.X2.X1.vout X2.X1.X1.X1.X2.X1.X3.vin2 0.326f
C3198 a_23126_27888# X1.X2.X2.X3.vin2 7.93e-20
C3199 d3 a_33976_18540# 7.7e-20
C3200 X2.X2.X2.X1.X2.X1.X3.vin1 a_52492_10734# 0.00251f
C3201 X1.X1.X1.X2.X1.X1.X1.vin2 a_2196_15634# 1.78e-19
C3202 a_52106_6962# X2.X2.X2.X1.X1.X1.X3.vin2 0.00815f
C3203 a_49002_29936# d1 0.0422f
C3204 d2 X1.X1.X2.X2.X2.X2.vrefh 0.168f
C3205 a_31476_17540# X2.X1.X1.X2.X1.X1.X3.vin1 0.354f
C3206 d3 a_34062_20446# 4.67e-19
C3207 a_31862_17540# X2.X1.X1.X2.X1.X1.X1.vin1 0.417f
C3208 X1.X2.X1.X1.X2.X2.X2.vin1 a_17222_19446# 0.402f
C3209 a_10686_15546# vdd 0.553f
C3210 X2.X2.X1.X1.X1.X1.X2.vin1 d0 0.262f
C3211 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.vout 0.0215f
C3212 d0 a_11072_9828# 0.515f
C3213 a_8186_14586# d1 0.0422f
C3214 a_48316_5198# X2.X2.X1.X2.X2.X2.X3.vin2 0.101f
C3215 X2.X1.X3.vin2 X2.X3.vin1 0.238f
C3216 X1.X2.X1.X1.X1.X2.X3.vin2 a_17222_28976# 7.84e-19
C3217 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X2.vrefh 0.076f
C3218 a_19036_28070# X1.X2.X1.X1.X1.X2.X3.vin1 0.199f
C3219 a_54992_19358# d2 0.00256f
C3220 a_54606_11734# X2.X2.X2.X1.X2.vrefh 8.22e-20
C3221 X1.X2.X1.X2.X2.X2.X1.vin1 a_17222_8010# 8.22e-20
C3222 X1.X1.X1.X2.X2.X1.vout X1.X1.X1.X2.X2.X1.X3.vin2 0.326f
C3223 a_34062_28070# a_34362_29936# 5.55e-20
C3224 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X3.vin1 2.33e-19
C3225 X2.X2.X2.X2.X2.X1.vout X2.X2.X2.X2.X3.vin2 0.399f
C3226 a_16836_13728# vdd 1.05f
C3227 a_34362_22312# X2.X1.X1.X1.X2.X2.vout 0.263f
C3228 a_4696_22312# X1.X1.X1.X1.X2.X2.X3.vin1 0.00329f
C3229 d3 X2.X1.X1.X1.X1.X1.X1.vin2 1.14e-19
C3230 d1 a_17222_4198# 0.0015f
C3231 a_54606_17452# X2.X2.X2.X1.X2.X2.X1.vin2 8.88e-20
C3232 X2.X1.X2.X1.X3.vin1 vdd 0.805f
C3233 d5 vdd 13.3f
C3234 d5 a_28096_892# 9.9e-19
C3235 d3 a_19422_20446# 4.67e-19
C3236 a_19722_29936# X1.X2.X1.X1.X1.X2.X3.vin1 0.00874f
C3237 d6 a_14082_892# 0.0338f
C3238 a_19422_9010# a_19722_7064# 4.19e-20
C3239 X1.X2.X1.X2.X2.X1.vout a_19336_7064# 0.169f
C3240 a_39966_25076# a_40352_25076# 0.419f
C3241 d4 X2.X1.X1.X1.X1.X2.vout 0.0921f
C3242 X1.X1.X2.X2.X1.X1.X1.vin1 a_11072_19358# 0.195f
C3243 a_25326_28888# vdd 0.541f
C3244 a_39966_6016# X2.X1.X2.X1.X1.X1.X2.vin1 0.402f
C3245 X1.X2.X2.X2.X2.X1.X1.vin1 d0 0.267f
C3246 X2.X1.X2.X3.vin1 d1 0.00955f
C3247 a_10686_7922# vdd 0.553f
C3248 X1.X1.X1.X1.X2.X2.X1.vin1 d0 0.267f
C3249 a_2196_25164# X1.X1.X1.X1.X2.X1.X2.vin1 1.78e-19
C3250 X2.X1.X2.X2.X1.X1.X1.vin1 d2 0.0116f
C3251 a_31862_25164# X2.X1.X1.X1.X2.X1.X1.vin1 0.417f
C3252 a_31476_25164# X2.X1.X1.X1.X2.X1.X3.vin1 0.354f
C3253 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X3.vin1 0.00836f
C3254 X2.X1.X3.vin1 X2.X1.X1.X2.X3.vin2 0.0816f
C3255 a_52792_24076# a_52492_22210# 6.71e-19
C3256 d3 a_46502_9916# 0.00112f
C3257 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X1.vin2 0.076f
C3258 d0 a_46502_32788# 0.0394f
C3259 X1.X1.X2.vrefh d6 4.63e-19
C3260 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X3.vin1 0.00789f
C3261 a_34062_9010# X2.X1.X1.X2.X2.X1.X3.vin2 0.267f
C3262 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 0.0903f
C3263 X2.X2.X2.X1.X2.X1.X1.vin2 vdd 0.36f
C3264 a_34062_5198# X2.X1.X1.X2.X2.X2.X3.vin2 0.277f
C3265 X1.X2.X2.X2.X1.X1.X1.vin1 d2 0.0116f
C3266 a_10686_30794# vdd 0.553f
C3267 a_52792_20264# a_52492_18358# 6.2e-19
C3268 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin1 0.195f
C3269 X2.X2.X2.X1.X2.X2.X1.vin1 a_54992_15546# 0.195f
C3270 a_33976_7064# X2.X1.X1.X2.X2.X2.vout 0.0929f
C3271 X1.X1.X2.X1.X2.X2.X2.vin1 d0 0.262f
C3272 X2.X2.X2.X2.X1.X1.X3.vin1 vdd 0.997f
C3273 X1.X1.X1.X2.X1.X2.X3.vin1 a_2582_11822# 0.00207f
C3274 d2 X1.X2.X2.X1.X2.X1.X3.vin1 0.104f
C3275 X1.X1.X3.vin1 X1.X1.X2.X1.X3.vin1 0.00304f
C3276 X2.X2.X1.X1.X1.X1.vout X2.X2.X1.X1.X1.X1.X3.vin2 0.342f
C3277 a_8572_29834# X1.X1.X2.X2.X2.X2.vout 0.0929f
C3278 a_16836_15634# d1 2.92e-22
C3279 d3 a_23212_25982# 0.621f
C3280 X2.X1.X2.X2.X1.X2.X3.vin1 a_37852_22210# 0.00329f
C3281 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X2.vin1 0.00117f
C3282 X2.X1.X2.X2.X2.X1.X3.vin1 d3 0.0332f
C3283 a_31862_17540# a_34062_16634# 4.2e-20
C3284 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X2.vrefh 0.564f
C3285 X1.X1.X2.X2.X1.X1.X3.vin2 a_10686_19358# 7.84e-19
C3286 X1.X2.X1.X2.X2.X2.vout vdd 0.698f
C3287 a_31862_19446# d0 0.0489f
C3288 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X1.vin1 0.0689f
C3289 d2 X1.X2.X2.X1.X1.X2.vrefh 6.65e-20
C3290 d1 X1.X2.X2.X1.X1.X1.X2.vin1 0.0144f
C3291 X1.X2.X2.X1.X1.X1.vout a_23512_5016# 0.359f
C3292 a_34362_10916# X2.X1.X1.X2.X2.X1.X3.vin2 3.49e-19
C3293 a_10686_9828# a_11072_9828# 0.419f
C3294 X1.X2.X1.X1.X2.X1.X1.vin1 d1 0.0118f
C3295 d2 a_39966_6016# 4.64e-19
C3296 X1.X1.X2.X2.X1.X1.X1.vin1 d2 0.0116f
C3297 a_48616_18540# X2.X2.X1.X3.vin2 0.0927f
C3298 a_31862_25164# d2 0.00328f
C3299 X1.X3.vin2 a_20672_892# 0.684f
C3300 X1.X1.X2.X2.X1.X2.X1.vin2 d0 0.276f
C3301 X2.X2.X2.X1.X2.vrefh a_54606_9828# 0.3f
C3302 a_39966_26982# a_37852_25982# 5.36e-21
C3303 X2.X1.X2.X2.X1.X1.X3.vin1 vdd 0.997f
C3304 a_2582_9916# X1.X1.X1.X2.X2.X1.X1.vin1 0.417f
C3305 X1.X1.X1.X1.X1.X2.X3.vin2 d1 0.171f
C3306 a_2196_9916# X1.X1.X1.X2.X2.X1.X3.vin1 0.354f
C3307 X1.X2.X2.X1.X2.X1.X1.vin1 vdd 0.592f
C3308 X1.X1.X1.X2.X2.X2.X3.vin1 d0 4.36e-19
C3309 a_31862_23258# vdd 0.541f
C3310 X2.X1.X2.X2.X2.X2.X3.vin1 a_40352_30794# 0.354f
C3311 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X1.vin2 0.668f
C3312 X2.X1.X2.X2.X2.X1.X1.vin2 a_40352_28888# 1.78e-19
C3313 X1.X1.X2.X2.X3.vin1 a_8486_20264# 1.52e-19
C3314 d0 X1.X2.X2.X1.X2.X2.vrefh 0.848f
C3315 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 0.587f
C3316 a_11072_32700# d4 1.8e-19
C3317 a_17222_19446# d0 0.0489f
C3318 X1.X1.X3.vin2 vdd 0.834f
C3319 d3 X2.X2.X1.X2.X2.vrefh 6.65e-20
C3320 X2.X1.X2.X2.X1.X2.X1.vin2 a_40352_23170# 0.12f
C3321 a_37466_25982# d1 0.0316f
C3322 a_39966_23170# X2.X1.X2.X2.X1.X2.X1.vin1 0.417f
C3323 a_4782_20446# d4 9.67e-19
C3324 a_33676_31882# a_31862_30882# 1.15e-20
C3325 X1.X1.X1.X1.X2.X1.X2.vin1 vdd 0.576f
C3326 X2.X2.X2.X3.vin2 a_52106_22210# 0.00292f
C3327 X2.X2.X3.vin1 a_48702_9010# 2.12e-19
C3328 a_8186_14586# a_8486_12640# 4.19e-20
C3329 a_23212_10734# a_23126_8828# 3.3e-19
C3330 X2.X1.X2.X1.X1.X1.vout X2.X1.X2.X1.X1.X1.X3.vin2 0.342f
C3331 X1.X2.X2.X2.X1.X1.X3.vin1 vdd 0.997f
C3332 d2 a_2582_9916# 0.00328f
C3333 X2.X1.X3.vin2 a_37766_16452# 3.98e-19
C3334 a_8872_8828# a_8186_6962# 3.31e-19
C3335 d2 X1.X1.X1.X2.X1.X1.vout 0.00169f
C3336 X1.X2.X3.vin1 a_22826_18358# 5.87e-20
C3337 a_37766_8828# a_37852_6962# 3.38e-19
C3338 a_54606_13640# X2.X2.X2.X1.X2.X1.X3.vin1 0.00207f
C3339 X2.X2.X1.X1.X1.X2.X3.vin2 a_49002_29936# 3.85e-19
C3340 X1.X1.X2.X2.X1.X2.vrefh d0 0.848f
C3341 a_48702_28070# X2.X2.X1.X1.X3.vin1 9.54e-19
C3342 X1.X2.X1.X1.X1.X1.X1.vin1 d0 0.0488f
C3343 a_33976_7064# a_31862_6104# 2.68e-20
C3344 a_10686_21264# X1.X1.X2.X2.X1.X1.X2.vin1 0.402f
C3345 a_16836_30882# d1 2.92e-22
C3346 X2.X2.X1.X2.X2.X1.X1.vin2 vdd 0.36f
C3347 d3 X1.X1.X1.X1.X1.X2.vout 6.83e-19
C3348 d3 a_52106_18358# 0.0469f
C3349 a_2582_19446# d0 0.0489f
C3350 a_10686_21264# d2 0.0059f
C3351 a_33976_14688# d1 0.00613f
C3352 d2 X2.X2.X1.X2.X1.X2.vout 0.00124f
C3353 X1.X2.X2.X3.vin2 d4 1.03f
C3354 a_23126_12640# a_23512_12640# 0.419f
C3355 X2.X1.X1.X2.X2.X1.X3.vin1 vdd 0.997f
C3356 d2 a_52792_5016# 0.00251f
C3357 X1.X2.X2.X1.X1.X1.X3.vin2 X1.X2.X2.X1.X1.X1.X3.vin1 0.581f
C3358 a_10686_25076# d0 0.0489f
C3359 d2 X2.X2.X1.X1.X1.X1.X1.vin2 1.68e-19
C3360 a_46116_15634# a_46116_13728# 0.00396f
C3361 X1.X2.X1.X1.X2.X2.vout d1 0.033f
C3362 a_25326_7922# vdd 0.553f
C3363 X1.X1.X1.X3.vin1 d2 6.42e-19
C3364 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X1.vin2 0.242f
C3365 a_54606_9828# a_54606_7922# 0.00198f
C3366 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X1.vin1 5.19e-19
C3367 d3 a_17222_11822# 1.89e-19
C3368 a_54992_21264# vdd 1.05f
C3369 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 0.049f
C3370 d3 X1.X1.X2.X2.X1.X2.X3.vin1 2.1e-19
C3371 a_17222_28976# X1.X2.X1.X1.X1.X1.X3.vin2 8.07e-19
C3372 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.vout 0.075f
C3373 a_33676_16634# a_34062_16634# 0.419f
C3374 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X1.X2.X1.X1.X2.X1.vin1 0.668f
C3375 X2.X1.X2.X2.X1.X1.X3.vin2 vdd 0.905f
C3376 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X1.vin1 5.19e-19
C3377 X1.X2.X2.X2.X2.X2.vrefh d0 0.848f
C3378 X2.X1.X2.X1.X2.X1.X1.vin2 d1 4.01e-19
C3379 d4 X1.X2.X1.X2.X1.X1.X1.vin1 6.34e-20
C3380 X1.X2.X2.X1.X3.vin2 a_23212_14586# 0.363f
C3381 a_2582_17540# d1 3.95e-19
C3382 a_6032_892# vdd 0.475f
C3383 X1.X1.X2.X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X1.vin2 0.076f
C3384 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin1 0.267f
C3385 a_16836_17540# d2 0.00256f
C3386 d3 X2.X1.X2.X2.X1.X2.X3.vin2 0.0247f
C3387 d1 X1.X3.vin2 0.00146f
C3388 X1.X2.X2.X1.X2.X1.X3.vin2 a_25326_11734# 7.84e-19
C3389 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X1.vin1 0.0689f
C3390 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X1.vout 0.13f
C3391 d2 X1.X1.X1.X1.X1.X1.vout 0.0903f
C3392 a_23212_29834# a_23512_31700# 6.71e-19
C3393 X2.X2.X2.X2.X2.X2.X1.vin1 a_54992_30794# 0.195f
C3394 X2.X2.X2.X2.X2.X2.vrefh vdd 0.415f
C3395 X1.X1.X1.X2.X3.vin2 vdd 1.29f
C3396 a_11072_6016# d1 2.92e-22
C3397 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X1.vout 0.118f
C3398 a_39966_15546# d1 3.41e-19
C3399 X2.X1.X1.X2.X1.X1.X3.vin2 a_31862_13728# 8.07e-19
C3400 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.vout 0.075f
C3401 X1.X2.X1.X2.X3.vin2 a_19422_5198# 9.7e-20
C3402 a_49002_22312# vdd 0.567f
C3403 d1 X2.X2.X1.X2.X2.X2.vrefh 0.0124f
C3404 d4 X1.X1.X1.X1.X3.vin1 0.0378f
C3405 d4 X2.X2.X1.X3.vin2 0.12f
C3406 a_16836_17540# a_17222_17540# 0.419f
C3407 X2.X1.X1.X2.vrefh a_31476_17540# 1.64e-19
C3408 X2.X1.X1.X2.X2.X1.X3.vin1 a_33676_9010# 0.199f
C3409 X1.X1.X2.X1.X1.X1.X2.vin1 d2 6e-20
C3410 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X1.vin2 0.1f
C3411 X1.X2.X1.X3.vin2 a_19722_10916# 0.452f
C3412 a_31476_32788# a_31476_30882# 0.00396f
C3413 X2.X1.X2.X2.X3.vin2 vdd 1.29f
C3414 a_8572_25982# a_8872_24076# 6.48e-19
C3415 a_23212_18358# X1.X2.X2.X1.X2.X2.X3.vin2 0.00517f
C3416 d3 X1.X1.X2.X1.X1.X2.X3.vin2 0.0251f
C3417 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X3.vin2 0.102f
C3418 a_11072_11734# d1 2.25e-20
C3419 a_25326_23170# d1 3.41e-19
C3420 a_48316_12822# vdd 1.05f
C3421 X2.X2.X3.vin1 a_52406_12640# 8.66e-20
C3422 a_52106_6962# a_52792_5016# 2.86e-19
C3423 a_25326_23170# a_25326_21264# 0.00198f
C3424 a_2582_27070# vdd 0.542f
C3425 X2.X1.X2.X1.X2.X2.X3.vin2 a_37766_16452# 0.277f
C3426 a_54992_23170# vdd 1.05f
C3427 d1 a_31476_8010# 2.92e-22
C3428 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X3.vin1 0.00117f
C3429 X1.X1.X1.X1.X1.X2.X3.vin2 X1.X1.X1.X1.X2.vrefh 0.161f
C3430 d3 a_52106_10734# 0.284f
C3431 a_19036_12822# a_19336_10916# 6.48e-19
C3432 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X2.vin1 0.564f
C3433 a_28096_892# X3.vin2 0.0927f
C3434 X1.X2.X1.X2.X2.X2.vrefh X1.X1.X2.X1.X1.X2.vrefh 0.117f
C3435 X3.vin2 vdd 0.614f
C3436 a_23212_14586# a_23126_12640# 3.14e-19
C3437 X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.vout 1.5e-19
C3438 a_20672_892# vdd 0.477f
C3439 a_23212_6962# a_23126_5016# 3.14e-19
C3440 X2.X1.X1.X1.X1.X1.X1.vin1 d4 0.00332f
C3441 a_25326_32700# d2 1.95e-19
C3442 a_19036_16634# d1 0.521f
C3443 X1.X2.X1.X1.X1.X1.X3.vin1 a_17222_30882# 0.00207f
C3444 a_33976_10916# X2.X1.X1.X2.X2.X1.X3.vin1 0.00251f
C3445 a_48702_16634# vdd 0.561f
C3446 a_52792_27888# d1 0.521f
C3447 X2.X2.X1.X2.X2.X2.vout a_48616_7064# 0.0929f
C3448 X2.X2.X2.X1.X2.X1.X1.vin1 a_54992_9828# 1.64e-19
C3449 a_2196_25164# d1 2.25e-20
C3450 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X2.vin1 0.0689f
C3451 d2 X2.X2.X2.X1.X2.X1.X3.vin2 0.171f
C3452 X2.X1.X2.X1.X1.X1.X3.vin2 a_39966_4110# 7.84e-19
C3453 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X1.vin1 0.0689f
C3454 a_17222_9916# a_19036_9010# 1.06e-19
C3455 a_11072_25076# d2 0.00533f
C3456 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X1.X2.X1.X1.X2.vrefh 0.267f
C3457 a_39966_30794# d1 3.41e-19
C3458 a_48616_14688# a_46502_13728# 2.68e-20
C3459 X1.X1.X1.X2.X1.X2.vrefh a_2196_13728# 1.64e-19
C3460 a_34062_20446# X2.X1.X3.vin1 1.64e-19
C3461 a_52406_27888# d2 0.00123f
C3462 X2.X2.X1.X2.X2.X2.vout vdd 0.698f
C3463 X1.X1.X1.X2.X1.X1.X3.vin2 d1 0.15f
C3464 X2.X1.X1.X1.X2.X2.X3.vin2 a_34362_18540# 0.00846f
C3465 a_33976_18540# X2.X1.X3.vin1 0.354f
C3466 a_31476_27070# a_31476_28976# 0.00396f
C3467 X2.X1.X2.X1.X2.X2.vout vdd 0.865f
C3468 a_10686_13640# a_11072_13640# 0.419f
C3469 d2 X1.X1.X1.X1.X1.X2.X2.vin1 0.0329f
C3470 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.vout 0.033f
C3471 a_5082_26164# a_4782_28070# 4.41e-20
C3472 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X3.vin2 0.234f
C3473 a_34062_24258# vdd 0.561f
C3474 a_4696_26164# X1.X1.X1.X1.X1.X2.X3.vin2 0.00535f
C3475 X2.X1.X2.X2.X2.X1.X3.vin1 a_39966_28888# 0.00207f
C3476 a_19036_9010# d1 0.521f
C3477 X2.X2.X2.X1.X2.X2.X2.vin1 d1 1.03e-19
C3478 a_4782_9010# vdd 0.561f
C3479 a_2582_13728# X1.X1.X1.X2.X1.X2.X1.vin1 0.417f
C3480 a_2196_13728# X1.X1.X1.X2.X1.X2.X3.vin1 0.354f
C3481 a_54606_6016# vdd 0.541f
C3482 X2.X2.X1.X1.X2.X2.X3.vin1 d4 2.08e-19
C3483 a_46502_25164# vdd 0.553f
C3484 a_52106_14586# d1 0.0422f
C3485 a_25326_26982# X1.X2.X2.X2.X2.vrefh 8.22e-20
C3486 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X1.vin2 0.216f
C3487 a_33676_31882# a_34062_31882# 0.419f
C3488 a_23126_24076# a_25326_23170# 4.2e-20
C3489 a_48702_9010# a_46502_8010# 4.77e-21
C3490 X2.X1.X2.vrefh a_34926_892# 7.23e-19
C3491 X1.X1.X1.X1.X3.vin2 d1 0.00807f
C3492 a_2582_32788# a_2582_30882# 0.00198f
C3493 a_52492_6962# X2.X2.X2.X1.X1.X2.X3.vin1 0.00329f
C3494 X2.X2.X2.X1.X1.X2.X1.vin1 a_54606_6016# 8.22e-20
C3495 X2.X2.X2.X1.X1.X2.X1.vin2 X2.X2.X2.X1.X1.X1.X3.vin2 3.94e-19
C3496 a_17222_28976# X1.X2.X1.X1.X1.X2.X1.vin2 0.273f
C3497 a_40352_32700# d1 2.92e-22
C3498 a_19336_10916# X1.X2.X1.X2.X3.vin2 0.0927f
C3499 X2.X2.X2.X2.X2.X1.X1.vin1 vdd 0.592f
C3500 X1.X2.X1.X1.X2.vrefh d1 0.00745f
C3501 a_2582_15634# a_4696_14688# 2.95e-20
C3502 X1.X1.X3.vin1 X1.X1.X1.X3.vin2 1.04f
C3503 X2.X1.X1.X1.X1.X2.X3.vin2 d4 0.0533f
C3504 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X3.vin2 0.234f
C3505 a_25326_6016# a_23512_5016# 1.15e-20
C3506 X1.X2.X1.X1.X1.X2.X3.vin1 X1.X2.X1.X1.X1.X2.vrefh 2.33e-19
C3507 a_19036_31882# d1 0.511f
C3508 a_48702_31882# vdd 0.565f
C3509 X2.X2.X2.X2.X1.X1.X1.vin1 a_54606_17452# 8.22e-20
C3510 X2.X2.X2.X2.X1.X1.X1.vin2 X2.X2.X2.X1.X2.X2.X3.vin2 3.94e-19
C3511 a_17222_9916# vdd 0.553f
C3512 X2.X2.vrefh X2.X2.X1.X1.X1.X1.X1.vin1 0.108f
C3513 d0 X2.X1.X1.X2.X1.X2.X1.vin1 0.267f
C3514 d3 X1.X2.X1.X3.vin2 0.483f
C3515 a_54992_28888# d0 0.515f
C3516 X1.X1.X1.X2.X1.X2.vout X1.X1.X1.X2.X1.X2.X3.vin1 0.326f
C3517 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X2.X1.X2.X2.X2.X1.vin2 0.00232f
C3518 X2.X2.X2.X1.X2.X2.vrefh d1 0.0124f
C3519 d2 X1.X2.X1.X2.X3.vin1 0.0014f
C3520 d1 a_48616_7064# 0.00613f
C3521 a_2582_17540# a_4396_16634# 1.06e-19
C3522 X1.X2.X3.vin1 a_23126_16452# 8.66e-20
C3523 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X2.vin1 0.0689f
C3524 X2.X1.X3.vin1 a_35312_892# 0.371f
C3525 a_11072_28888# X1.X1.X2.X2.X2.X2.X1.vin1 1.64e-19
C3526 a_8572_22210# d2 0.526f
C3527 X2.X1.X2.X2.X2.X1.X3.vin2 d0 4.34e-19
C3528 d3 X1.X2.X1.X2.X1.X2.X2.vin1 8.68e-20
C3529 X1.X2.X2.X2.X2.X1.vout X1.X2.X2.X2.X2.X1.X3.vin2 0.326f
C3530 X1.X1.X1.X1.X1.X1.X3.vin2 d1 0.152f
C3531 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.X1.X2.vin1 0.0689f
C3532 a_10686_26982# X1.X1.X2.X2.X2.X1.X3.vin2 7.84e-19
C3533 a_25326_21264# vdd 0.541f
C3534 X2.X1.X2.X2.X2.X2.vout vdd 0.698f
C3535 X1.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin2 0.0128f
C3536 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X2.X1.X1.vin1 0.206f
C3537 d1 vdd 65f
C3538 a_40352_23170# a_40352_21264# 0.00396f
C3539 d1 a_28096_892# 4.67e-19
C3540 a_25326_32700# X1.X2.X2.X2.X2.X2.X2.vin1 0.402f
C3541 d0 a_46116_17540# 0.518f
C3542 X2.X2.X3.vin2 a_52106_14586# 3.67e-19
C3543 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X2.X1.X1.vin1 0.206f
C3544 X2.X2.X2.X1.X1.X2.X2.vin1 a_54992_9828# 0.197f
C3545 a_34062_12822# d1 0.0749f
C3546 d2 a_31476_11822# 0.00533f
C3547 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X3.vin1 2.33e-19
C3548 d3 a_4396_12822# 0.00108f
C3549 d0 X1.X1.X1.X2.X2.X2.X2.vin1 0.262f
C3550 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 0.581f
C3551 X1.X1.X1.X3.vin1 X1.X1.X2.X2.X3.vin2 7.46e-20
C3552 d1 X2.X2.X2.X1.X1.X2.X1.vin1 0.0118f
C3553 X1.X1.X2.X1.X2.X1.vout a_8572_14586# 0.169f
C3554 X2.X2.X3.vin1 X2.X2.X2.vrefh 0.178f
C3555 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin1 0.52f
C3556 X2.X2.X1.X1.X1.X1.X3.vin1 vdd 1.06f
C3557 d3 a_25326_25076# 1.89e-19
C3558 X2.X2.X2.X1.X1.X1.X3.vin1 vdd 1.03f
C3559 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.X3.vin1 0.587f
C3560 a_46502_27070# d3 1.89e-19
C3561 X1.X1.X2.X2.X2.X1.X1.vin2 a_11072_26982# 0.12f
C3562 a_10686_26982# X1.X1.X2.X2.X2.X1.X1.vin1 0.417f
C3563 X1.X2.X3.vin1 a_23126_8828# 8.66e-20
C3564 d0 a_31862_4198# 0.049f
C3565 X1.X1.X1.X3.vin2 a_4782_16634# 5.21e-19
C3566 a_5082_18540# X1.X1.X1.X2.X1.X1.X3.vin2 3.49e-19
C3567 X1.X2.X2.X1.X2.X2.X1.vin1 a_25712_13640# 1.64e-19
C3568 a_54606_19358# vdd 0.553f
C3569 d2 a_31862_15634# 0.0059f
C3570 X2.X1.X2.X2.X1.X1.vout a_37766_20264# 0.422f
C3571 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X3.vin1 0.0174f
C3572 X2.X1.X1.X1.X2.X2.vrefh d2 0.168f
C3573 X2.X2.X1.X3.vin2 a_48702_12822# 6.03e-19
C3574 X1.X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin2 0.0128f
C3575 d4 X1.X2.X3.vin1 0.286f
C3576 X2.X2.X1.X1.X1.X2.X2.vin1 a_46116_27070# 0.197f
C3577 X1.X1.X2.X2.X2.X1.X3.vin1 a_8872_27888# 0.199f
C3578 a_2196_25164# X1.X1.X1.X1.X2.vrefh 1.64e-19
C3579 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X1.vin2 0.216f
C3580 a_31862_32788# X2.X1.X1.X1.X1.X1.X2.vin1 8.88e-20
C3581 X2.X2.X2.X2.X2.X1.X1.vin2 a_54606_28888# 8.88e-20
C3582 d2 X1.X1.X1.X2.X2.X2.vrefh 0.168f
C3583 a_52406_27888# X2.X2.X2.X2.X2.X1.X3.vin1 0.428f
C3584 a_54606_21264# X2.X2.X2.X2.X1.X1.X3.vin2 0.567f
C3585 X1.X1.X2.X2.X2.X1.vout vdd 0.775f
C3586 d2 X1.X1.X2.X1.X2.X1.X1.vin2 0.231f
C3587 X2.X2.X2.X3.vin2 a_52492_25982# 0.355f
C3588 X2.X2.X3.vin2 vdd 0.76f
C3589 X2.X1.X2.X2.X1.X1.X1.vin2 vdd 0.36f
C3590 X1.X2.vrefh d1 7.29e-21
C3591 a_17222_23258# d2 0.00665f
C3592 d1 a_33676_9010# 0.521f
C3593 a_23126_24076# vdd 0.47f
C3594 d3 a_19722_10916# 0.29f
C3595 X1.X1.X1.X1.X2.X2.X3.vin2 d1 0.151f
C3596 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X1.vin2 8.93e-19
C3597 X1.X2.X2.X2.X2.X1.X1.vin2 d3 3.99e-21
C3598 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.vrefh 0.161f
C3599 a_25326_9828# X1.X2.X2.X1.X1.X2.X3.vin1 0.00207f
C3600 X1.X2.X2.X1.X2.X2.X2.vin1 a_25326_15546# 8.88e-20
C3601 X2.X2.X3.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 8.36e-19
C3602 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X1.vout 0.0524f
C3603 a_39966_23170# X2.X1.X2.X2.X1.X2.vrefh 8.22e-20
C3604 X1.X1.X2.X2.X1.X2.X1.vin1 vdd 0.592f
C3605 a_48316_24258# X2.X2.X1.X1.X2.X1.vout 0.359f
C3606 X1.X1.X2.X2.X2.X2.X3.vin2 d2 0.00427f
C3607 X1.X1.X2.X1.X1.X1.X1.vin1 X1.X2.X2.vrefh 0.00437f
C3608 d3 X2.X2.X1.X1.X1.X2.vout 0.125f
C3609 X2.X1.X2.X2.X2.X1.X1.vin1 d1 0.0118f
C3610 a_4396_16634# X1.X1.X1.X2.X1.X1.X3.vin2 0.1f
C3611 X1.X2.X2.X1.X2.X1.X2.vin1 d1 1.03e-19
C3612 a_46502_11822# a_46502_9916# 0.00198f
C3613 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X2.X3.vin1 0.0131f
C3614 X1.X2.X2.X2.X1.X1.X1.vin2 vdd 0.36f
C3615 X2.X2.X2.X1.X1.X2.vout vdd 0.696f
C3616 X1.X2.X1.X1.X1.X1.X3.vin1 a_19422_31882# 0.428f
C3617 a_46116_11822# X2.X2.X1.X2.X2.X1.X1.vin1 1.64e-19
C3618 d3 X1.X1.X2.X1.X3.vin2 0.387f
C3619 X2.X2.X3.vin1 X2.X2.X2.X1.X1.X1.vout 5.53e-20
C3620 d2 a_39966_13640# 0.00665f
C3621 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X3.vin1 2.33e-19
C3622 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.X1.X1.vin2 3.94e-19
C3623 a_33676_28070# a_31862_27070# 1.15e-20
C3624 a_5082_18540# vdd 0.478f
C3625 X2.X2.X2.X1.X3.vin2 a_52106_10734# 0.241f
C3626 X2.X2.X1.X3.vin1 d2 6.42e-19
C3627 X2.X2.X1.X1.X2.X2.vout X2.X2.X1.X1.X2.X2.X3.vin1 0.335f
C3628 X2.X1.X1.X1.X1.X2.X1.vin1 d1 0.0118f
C3629 d2 a_31862_30882# 4.64e-19
C3630 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.vrefh 0.161f
C3631 a_33976_10916# d1 0.0126f
C3632 X2.X2.X1.X1.X3.vin2 a_49002_22312# 0.423f
C3633 d2 a_46502_28976# 0.00479f
C3634 a_34362_14688# X2.X1.X1.X2.X1.X2.X3.vin1 0.00874f
C3635 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin1 0.195f
C3636 a_37466_22210# X2.X1.X2.X2.X1.X1.X3.vin2 0.00815f
C3637 X2.X1.X1.X2.X1.X1.X1.vin2 d1 1.49e-19
C3638 X1.X1.X2.X2.X1.X1.X1.vin2 vdd 0.36f
C3639 a_8486_12640# vdd 0.561f
C3640 a_23126_20264# a_23212_18358# 3.21e-19
C3641 a_25712_25076# vdd 1.05f
C3642 d3 X2.X2.X2.X1.X2.X2.vout 8.47e-19
C3643 a_4396_24258# X1.X1.X1.X1.X2.X1.X3.vin2 0.1f
C3644 X1.X2.X1.X2.X1.X1.X3.vin1 d1 0.146f
C3645 d3 a_48702_24258# 0.00195f
C3646 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X1.X2.X1.X1.X2.vrefh 0.1f
C3647 d2 X2.X1.X1.X2.X1.X1.X1.vin1 0.0116f
C3648 X1.X2.X1.X2.X1.X2.vout d1 0.033f
C3649 X1.X1.X2.X2.X1.X2.X3.vin2 vdd 0.787f
C3650 X1.X1.X1.X1.X2.vrefh vdd 0.426f
C3651 a_48316_9010# a_48702_9010# 0.419f
C3652 X1.X2.X2.X1.X3.vin2 a_23212_10734# 0.0927f
C3653 d0 a_10686_15546# 0.0675f
C3654 a_19722_26164# d4 3.47e-19
C3655 a_37466_29834# X2.X1.X2.X2.X2.X2.X3.vin1 0.00874f
C3656 a_4696_26164# X1.X1.X1.X1.X3.vin2 0.0927f
C3657 X2.X2.X2.X2.X1.X1.X3.vin2 a_52106_18358# 3.49e-19
C3658 X2.X2.X1.X1.X1.X2.X3.vin2 vdd 0.787f
C3659 a_38152_27888# a_37466_29834# 2.86e-19
C3660 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin2 0.1f
C3661 X2.X2.X1.X2.X1.X2.X3.vin2 a_49002_10916# 0.00846f
C3662 a_10686_17452# X1.X1.X2.X1.X2.X2.X3.vin1 0.00207f
C3663 X2.X1.X1.X1.X2.X2.vout d2 0.00117f
C3664 d1 X2.X1.X2.X1.X1.X1.X3.vin1 0.16f
C3665 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin1 0.195f
C3666 a_23512_27888# d2 0.00251f
C3667 d3 X2.X1.X2.X2.X1.X2.vout 0.0232f
C3668 d0 a_16836_13728# 0.518f
C3669 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 5.19e-19
C3670 a_52492_10734# vdd 1.05f
C3671 X1.X2.X2.X1.X1.X2.vout a_22826_6962# 0.254f
C3672 X1.X1.X1.X1.X2.X1.X1.vin2 a_2196_23258# 1.78e-19
C3673 X2.X1.X2.X1.X1.X1.X1.vin1 a_40352_4110# 0.195f
C3674 d0 d5 0.533f
C3675 a_4396_16634# vdd 1.05f
C3676 d3 X1.X1.X2.X1.X1.X2.vout 6.06e-19
C3677 d4 X2.X2.X1.X1.X3.vin1 0.00246f
C3678 d2 X2.X1.X1.X2.X2.X2.X3.vin2 8.42e-19
C3679 X2.X2.X2.X2.X1.X2.vout d1 0.033f
C3680 X1.X1.X1.X2.X2.vrefh a_2196_11822# 0.118f
C3681 a_2582_28976# a_2582_30882# 0.00198f
C3682 a_4782_20446# X1.X1.X3.vin1 1.64e-19
C3683 X1.X1.X1.X1.X2.X2.X3.vin2 a_5082_18540# 0.00846f
C3684 d2 a_54992_15546# 0.00274f
C3685 X1.X1.X1.X1.X1.X2.X1.vin1 a_2196_30882# 1.64e-19
C3686 d1 X1.X1.X2.X1.X1.X1.vout 0.0239f
C3687 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X3.vin1 0.0131f
C3688 a_25326_28888# d0 0.0489f
C3689 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X3.vin2 8.93e-19
C3690 X2.X2.X1.X2.X2.vrefh a_46502_11822# 0.3f
C3691 d0 a_10686_7922# 0.0675f
C3692 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 5.19e-19
C3693 X2.X1.X2.X2.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin2 0.0128f
C3694 a_48616_22312# a_48316_20446# 6.71e-19
C3695 d3 a_16836_32788# 2.56e-19
C3696 a_31862_23258# X2.X1.X1.X1.X2.X2.X1.vin1 8.22e-20
C3697 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X2.vout 0.398f
C3698 a_4696_26164# vdd 1.05f
C3699 d3 X2.X2.X2.X2.X2.X2.vout 1.05e-19
C3700 a_25326_13640# a_23126_12640# 4.77e-21
C3701 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.vout 0.197f
C3702 d0 X2.X2.X2.X1.X2.X1.X1.vin2 0.276f
C3703 X2.X1.X2.X2.X1.X2.X1.vin1 d2 0.0114f
C3704 X2.X1.X2.X3.vin1 a_37466_14586# 7.98e-19
C3705 X2.X1.X1.X3.vin2 X2.X1.X2.X1.X3.vin2 7.46e-20
C3706 a_39966_9828# X2.X1.X2.X1.X1.X2.X2.vin1 0.402f
C3707 a_48616_10916# a_48316_9010# 6.2e-19
C3708 a_10686_6016# X1.X1.X2.X1.X1.X1.X3.vin1 0.00207f
C3709 X2.X2.X2.X1.X2.X1.X2.vin1 a_54992_13640# 0.197f
C3710 a_10686_30794# d0 0.0675f
C3711 X2.X1.X2.X1.X1.X1.vout a_37852_6962# 0.169f
C3712 a_39966_32700# a_37766_31700# 4.77e-21
C3713 d3 X2.X2.X2.X2.X2.X1.X3.vin2 7.71e-19
C3714 X2.X1.X1.X1.X1.X1.X3.vin1 d1 0.0296f
C3715 a_23126_12640# a_23212_10734# 3.21e-19
C3716 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X2.vrefh 0.165f
C3717 X1.X2.X2.X1.X1.X2.X3.vin2 a_25326_7922# 7.84e-19
C3718 a_34362_29936# vdd 0.477f
C3719 a_16836_15634# X1.X2.X1.X2.X1.X2.X1.vin1 1.64e-19
C3720 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X1.vin1 0.0689f
C3721 a_17222_15634# a_17222_13728# 0.00198f
C3722 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 0.587f
C3723 X2.X2.X2.X2.X1.X1.X3.vin1 d0 4.36e-19
C3724 d3 X2.X1.X2.X3.vin2 0.511f
C3725 a_46502_13728# X2.X2.X1.X2.X1.X2.X3.vin1 0.52f
C3726 a_37466_6962# vdd 0.477f
C3727 a_31476_11822# a_31862_11822# 0.419f
C3728 a_8186_29834# a_8572_29834# 0.419f
C3729 a_37852_10734# X2.X1.X2.X1.X1.X2.vout 7.93e-20
C3730 a_4396_31882# X1.X1.X1.X1.X1.X1.X3.vin2 0.1f
C3731 a_4396_31882# vdd 1.05f
C3732 X2.X1.X1.X1.X2.X1.X3.vin2 a_34362_22312# 0.00815f
C3733 X2.X1.X2.X2.X1.X1.X2.vin1 X2.X2.X1.X1.X2.X2.X1.vin2 0.00232f
C3734 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X2.X2.vin1 0.0689f
C3735 X2.X1.X3.vin1 a_34362_7064# 9.8e-19
C3736 a_46116_21352# a_46502_21352# 0.419f
C3737 a_54606_30794# X2.X2.X2.X2.X2.X2.X3.vin2 7.84e-19
C3738 a_52406_16452# a_52792_16452# 0.419f
C3739 X2.X1.X2.X2.X1.X1.X3.vin1 d0 4.36e-19
C3740 d0 X1.X2.X2.X1.X2.X1.X1.vin1 0.267f
C3741 a_13696_892# X3.vin1 0.369f
C3742 d2 X1.X2.X2.X1.X2.X2.vout 0.00117f
C3743 a_31862_23258# d0 0.0489f
C3744 a_4396_24258# a_4696_22312# 6.1e-19
C3745 X1.X2.X2.X3.vin1 vdd 1.26f
C3746 X1.X1.X1.X2.X2.X2.X1.vin2 vdd 0.387f
C3747 X2.X1.X2.X2.X3.vin1 a_37852_25982# 0.17f
C3748 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X2.X1.X2.X1.X2.vrefh 0.0128f
C3749 X2.X2.X1.X1.X3.vin2 d1 0.00807f
C3750 a_17222_23258# a_19336_22312# 2.95e-20
C3751 X1.X1.X3.vin2 d0 0.0368f
C3752 a_19422_28070# d3 0.00107f
C3753 d3 X1.X2.X2.X2.X1.X1.vout 0.00883f
C3754 X1.X1.X1.X1.X2.X2.X2.vin1 d2 0.0314f
C3755 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X2.vin1 0.242f
C3756 a_10686_9828# a_10686_7922# 0.00198f
C3757 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 0.242f
C3758 X1.X1.X1.X1.X2.X1.X2.vin1 d0 0.262f
C3759 X1.X1.X2.X1.X1.X1.X1.vin2 X1.X2.X1.X2.X2.X2.X2.vin1 0.00232f
C3760 X1.X2.X2.X2.X1.X1.X1.vin1 X2.X1.X1.X2.vrefh 0.00437f
C3761 a_52106_29834# a_52406_31700# 5.55e-20
C3762 X1.X1.X1.X2.X1.X2.X1.vin2 d1 0.00406f
C3763 X1.X2.X2.X2.X1.X1.X3.vin1 d0 4.36e-19
C3764 X1.X1.X3.vin1 a_8186_6962# 6.45e-19
C3765 a_52792_27888# X2.X2.X2.X2.X2.X1.vout 0.359f
C3766 a_19036_16634# a_19336_14688# 6.1e-19
C3767 X2.X1.X2.X2.X2.X1.X3.vin1 a_38152_27888# 0.199f
C3768 a_4696_14688# a_4782_12822# 3.38e-19
C3769 d2 X1.X2.X2.X1.X1.X2.vout 0.106f
C3770 a_5082_14688# a_4396_12822# 3.31e-19
C3771 d3 X1.X2.X1.X1.X3.vin1 0.153f
C3772 a_8186_22210# a_8486_20264# 4.19e-20
C3773 d0 X2.X2.X1.X2.X2.X1.X1.vin2 0.276f
C3774 a_16836_28976# d1 2.25e-20
C3775 X2.X1.X1.X2.X2.X1.X3.vin2 a_33976_7064# 0.00546f
C3776 X1.X1.X1.X2.vrefh a_2582_17540# 8.22e-20
C3777 d2 X1.X1.X1.X2.X1.X2.X1.vin1 0.0114f
C3778 d2 a_34062_31882# 7.66e-19
C3779 X2.X2.X2.X1.X2.X2.vrefh a_54606_13640# 0.3f
C3780 X2.X1.X2.X2.X3.vin1 d4 3.38e-19
C3781 d2 a_25712_28888# 0.00464f
C3782 d3 X2.X1.X2.X1.X2.X1.X3.vin1 0.0195f
C3783 a_37466_22210# d1 0.0422f
C3784 d0 X2.X1.X1.X2.X2.X1.X3.vin1 4.36e-19
C3785 a_37766_24076# a_38152_24076# 0.419f
C3786 a_8872_16452# a_8186_14586# 3.31e-19
C3787 d0 a_25326_7922# 0.0675f
C3788 a_54606_13640# vdd 0.541f
C3789 d2 X1.X1.X2.X2.X2.X1.X3.vin2 0.177f
C3790 a_54606_23170# a_54606_21264# 0.00198f
C3791 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X2.vrefh 0.267f
C3792 X2.X2.X3.vin1 X2.X3.vin2 0.12f
C3793 a_54992_21264# d0 0.515f
C3794 a_8486_8828# a_8872_8828# 0.419f
C3795 d2 X1.X2.X2.X2.X2.X2.vout 0.106f
C3796 a_33976_29936# X2.X1.X1.X1.X1.X2.X3.vin1 0.00329f
C3797 X2.X1.X2.X2.X1.X1.X3.vin2 d0 4.34e-19
C3798 a_52106_25982# a_52792_24076# 3.08e-19
C3799 X2.X2.X1.X1.X2.X2.X2.vin1 d1 1.03e-19
C3800 a_10686_26982# a_8572_25982# 5.36e-21
C3801 d0 a_6032_892# 3.19e-19
C3802 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 0.587f
C3803 X1.X1.X2.X2.X1.X1.X1.vin1 X1.X2.X1.X2.vrefh 0.00437f
C3804 X1.X1.X2.X1.X2.X1.X1.vin2 a_10686_11734# 0.273f
C3805 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin1 0.199f
C3806 X1.X1.X2.X2.X2.X1.X1.vin1 d2 0.0105f
C3807 a_25326_15546# a_25712_15546# 0.419f
C3808 a_16836_6104# X1.X2.X1.X2.X2.X2.vrefh 1.64e-19
C3809 a_54992_19358# X2.X2.X2.X2.vrefh 1.64e-19
C3810 X2.X2.X1.X2.vrefh d2 0.173f
C3811 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 5.19e-19
C3812 X2.X2.X2.X2.X1.X1.vout a_52792_20264# 0.359f
C3813 a_22826_25982# vdd 0.487f
C3814 a_19036_28070# X1.X2.X1.X1.X1.X2.X3.vin2 0.101f
C3815 X2.X2.X2.X1.X2.X2.X3.vin2 a_52792_16452# 0.101f
C3816 X2.X2.X1.X2.X1.X1.X1.vin1 vdd 0.592f
C3817 a_22826_10734# vdd 0.489f
C3818 a_19422_24258# d1 0.0749f
C3819 X2.X2.X2.X1.X2.X2.vout X2.X2.X2.X1.X3.vin2 0.0866f
C3820 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X2.X1.X2.X1.X1.X1.vin2 0.00232f
C3821 X2.X2.X2.X2.X2.X2.vrefh d0 0.844f
C3822 a_4782_5198# vdd 0.47f
C3823 d4 X1.X1.X1.X2.X1.X1.X1.vin1 6.34e-20
C3824 X2.X1.X1.X1.X2.X2.X2.vin1 d1 1.03e-19
C3825 d2 a_4696_29936# 0.606f
C3826 a_11072_6016# a_11072_7922# 0.00396f
C3827 a_5082_26164# X1.X1.X1.X1.X3.vin1 0.385f
C3828 X2.X2.X1.X1.X2.X2.X3.vin2 a_46502_19446# 0.567f
C3829 X1.X2.X1.X1.X1.X2.X3.vin2 a_19722_29936# 3.85e-19
C3830 a_37852_25982# a_37766_24076# 3.3e-19
C3831 a_19422_28070# X1.X2.X1.X1.X3.vin1 9.54e-19
C3832 X2.X2.X2.X2.X2.X1.vout vdd 0.775f
C3833 X1.X1.X2.X1.X1.X1.X3.vin1 X1.X1.X2.X1.X1.X1.X1.vin1 0.206f
C3834 X1.X2.X2.X2.X2.X1.X3.vin1 vdd 0.997f
C3835 X2.X1.X2.X1.X1.X1.X1.vin2 vdd 0.387f
C3836 X2.X1.X2.X1.X1.X1.vout a_37766_5016# 0.422f
C3837 X1.X2.X2.X1.X1.X2.X1.vin1 X1.X2.X2.X1.X1.X1.X3.vin2 5.19e-19
C3838 d4 a_52406_16452# 8.66e-19
C3839 a_19336_14688# vdd 1.05f
C3840 X2.X1.X1.X2.X1.X1.X3.vin1 a_31862_15634# 0.00207f
C3841 X2.X1.X2.X2.vrefh vdd 0.414f
C3842 X2.X2.X2.X2.X1.X2.X3.vin2 d1 0.171f
C3843 a_52406_31700# a_52792_31700# 0.419f
C3844 a_2582_27070# d0 0.0489f
C3845 a_42976_892# a_43362_892# 0.419f
C3846 a_54992_23170# d0 0.518f
C3847 X2.X1.X3.vin2 X2.X1.X2.vrefh 0.15f
C3848 X1.X2.X1.X1.X2.X2.X2.vin1 d1 1.03e-19
C3849 a_54606_6016# X2.X2.X2.X1.X1.X1.X1.vin2 8.88e-20
C3850 X2.X1.X2.X1.X2.X2.X3.vin1 a_37852_14586# 0.00329f
C3851 X1.X1.X2.X1.X1.X2.X3.vin1 a_10686_7922# 0.52f
C3852 d2 a_48702_9010# 7.51e-19
C3853 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin2 0.1f
C3854 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X2.X1.X1.X2.X2.X2.vin1 0.00232f
C3855 X1.X2.X3.vin2 X1.X2.X1.X2.X3.vin1 4.41e-19
C3856 X1.X2.X3.vin1 X1.X2.X2.X1.X3.vin2 6.26e-19
C3857 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X2.X1.X1.X1.X2.vrefh 0.0128f
C3858 X2.X2.X1.X1.X2.X2.vrefh a_46502_23258# 0.3f
C3859 X2.X2.X1.X1.X1.X2.X3.vin1 X2.X2.X1.X1.X1.X2.vrefh 2.33e-19
C3860 d0 X3.vin2 1.31e-19
C3861 a_22826_6962# X1.X2.X2.X1.X1.X1.vout 0.386f
C3862 a_39966_13640# X2.X1.X2.X1.X2.X1.X2.vin1 0.402f
C3863 a_31476_32788# d2 3.9e-19
C3864 X1.X1.X1.X2.X2.X1.X2.vin1 a_2196_8010# 0.197f
C3865 a_23212_25982# X1.X2.X2.X2.X1.X2.X3.vin2 0.00535f
C3866 a_40352_9828# d1 2.92e-22
C3867 a_23512_16452# d1 0.521f
C3868 a_5082_29936# X1.X1.X1.X1.X1.X1.vout 0.386f
C3869 d3 X2.X2.X2.X1.X3.vin2 0.387f
C3870 X1.X1.X1.X1.X3.vin1 a_4782_31882# 1.52e-19
C3871 d0 a_20672_892# 3.19e-19
C3872 X2.X2.X1.X1.X2.X1.X3.vin2 vdd 0.903f
C3873 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 0.587f
C3874 a_49002_18540# vdd 0.478f
C3875 a_5082_7064# vdd 0.477f
C3876 X2.X1.X1.X2.X1.X2.X2.vin1 a_31476_11822# 0.197f
C3877 d3 X1.X1.X2.X2.X3.vin1 0.376f
C3878 X1.X2.X1.X2.X2.X2.vout a_19036_5198# 0.36f
C3879 d2 X2.X1.X2.X1.X1.X2.vout 0.106f
C3880 a_19722_7064# a_19422_5198# 5.55e-20
C3881 a_54606_28888# a_54992_28888# 0.419f
C3882 X1.X2.X2.X1.X1.X2.X3.vin2 d1 0.171f
C3883 X2.X2.X2.X2.X2.vrefh d2 0.158f
C3884 a_25712_32700# d4 1.8e-19
C3885 X1.X2.X1.X2.X2.X2.X3.vin1 a_19336_7064# 0.00329f
C3886 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.vout 0.335f
C3887 d2 X2.X1.X2.X1.X1.X2.X2.vin1 0.0329f
C3888 a_31862_19446# a_33976_18540# 4.72e-20
C3889 a_34062_20446# a_31862_19446# 4.77e-21
C3890 a_10686_4110# vdd 0.553f
C3891 X2.X1.X1.X1.X2.X2.X3.vin2 a_31476_19446# 0.354f
C3892 X1.X2.X1.X2.vrefh a_16836_17540# 1.64e-19
C3893 a_46502_28976# X2.X2.X1.X1.X1.X2.X1.vin1 0.417f
C3894 a_46116_28976# X2.X2.X1.X1.X1.X2.X3.vin1 0.354f
C3895 a_8186_25982# a_8872_27888# 2.97e-19
C3896 X2.X1.X1.X1.X2.X2.X1.vin1 d1 0.0118f
C3897 a_54992_13640# a_54992_11734# 0.00396f
C3898 X2.X2.X2.X3.vin1 a_52406_8828# 1.64e-19
C3899 d4 a_19422_16634# 0.00142f
C3900 a_46502_21352# d2 0.00393f
C3901 d4 a_52406_31700# 2.4e-19
C3902 X2.X1.X2.X1.X2.X1.vout X2.X1.X2.X1.X2.X1.X3.vin2 0.326f
C3903 d3 a_5082_14688# 0.0469f
C3904 a_52406_27888# X2.X2.X2.X2.X3.vin2 0.00101f
C3905 d0 a_54606_6016# 0.0489f
C3906 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X1.vout 0.13f
C3907 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X3.vin2 0.449f
C3908 X2.X2.X1.X2.X2.X2.vrefh a_46116_8010# 0.118f
C3909 a_46502_25164# d0 0.0675f
C3910 d1 X2.X2.X2.X1.X1.X1.X1.vin2 0.0985f
C3911 X1.X2.X2.X2.X1.X1.X1.vin2 X2.X1.X1.X1.X2.X2.X2.vin1 0.00232f
C3912 a_11072_26982# a_11072_25076# 0.00396f
C3913 X1.X2.X1.X3.vin1 d1 0.00955f
C3914 a_2582_11822# vdd 0.542f
C3915 d2 a_48616_10916# 0.0057f
C3916 X1.X2.X2.X1.X3.vin1 a_23212_10734# 0.169f
C3917 X2.X2.X2.X1.X2.X2.X1.vin1 a_54992_13640# 1.64e-19
C3918 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.vout 0.326f
C3919 X1.X2.X1.X2.X1.X2.X3.vin2 a_16836_11822# 0.354f
C3920 X1.X2.X3.vin1 a_23126_12640# 8.66e-20
C3921 a_19422_12822# a_17222_11822# 4.77e-21
C3922 X2.X2.X2.X2.X2.X1.X1.vin1 d0 0.267f
C3923 a_52406_5016# a_54606_4110# 4.2e-20
C3924 X2.X1.X2.X1.X2.X2.X3.vin2 a_40352_17452# 0.354f
C3925 a_33676_28070# d2 0.00393f
C3926 X2.X2.X2.X1.X1.X1.X3.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 0.22f
C3927 X1.X1.X1.X2.vrefh vdd 0.414f
C3928 X1.X2.X2.X1.X2.X2.X3.vin1 vdd 0.962f
C3929 a_23512_31700# d1 0.515f
C3930 a_25326_30794# a_25712_30794# 0.419f
C3931 d4 X2.X2.X2.X1.X2.X2.X3.vin2 0.0264f
C3932 X2.X1.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin2 0.0128f
C3933 a_25326_7922# a_23212_6962# 2.68e-20
C3934 a_10686_32700# vdd 0.541f
C3935 d3 X2.X1.X3.vin1 0.834f
C3936 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.X3.vin1 0.00836f
C3937 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X3.vin1 0.206f
C3938 a_11072_15546# vdd 1.05f
C3939 X1.X2.X1.X1.X2.X2.X3.vin2 a_16836_19446# 0.354f
C3940 d0 a_17222_9916# 0.0675f
C3941 a_19422_20446# a_17222_19446# 4.77e-21
C3942 a_52792_12640# d1 0.521f
C3943 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.X1.vin2 3.94e-19
C3944 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X1.X2.X3.vin1 0.587f
C3945 a_5082_22312# d1 0.0422f
C3946 a_4696_29936# a_4396_28070# 6.71e-19
C3947 d4 X2.X2.vrefh 0.00449f
C3948 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X3.vin1 0.0565f
C3949 a_54992_11734# X2.X2.X2.X1.X2.vrefh 1.64e-19
C3950 a_48616_26164# vdd 1.05f
C3951 X1.X2.X1.X2.X1.X2.X1.vin1 vdd 0.592f
C3952 X1.X1.X1.X1.X2.X2.vout X1.X1.X1.X1.X2.X2.X3.vin1 0.335f
C3953 d1 X1.X2.X2.X1.X1.X1.X1.vin2 0.0985f
C3954 X1.X2.X2.X1.X1.X2.X3.vin1 vdd 0.96f
C3955 X2.X2.X2.X1.X2.X2.X2.vin1 a_54606_15546# 8.88e-20
C3956 a_46502_6104# X2.X2.X1.X2.X2.X2.X1.vin2 0.273f
C3957 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X1.vin2 8.93e-19
C3958 a_40352_28888# vdd 1.05f
C3959 a_25326_21264# d0 0.0489f
C3960 X1.X2.X1.X2.X2.X1.vout X1.X2.X1.X2.X2.X2.vout 0.514f
C3961 d0 d1 11.2f
C3962 a_10686_6016# X1.X1.X2.X1.X1.X2.vrefh 0.3f
C3963 X2.X1.X2.X2.X1.X2.X3.vin2 a_40352_25076# 0.354f
C3964 a_52492_22210# a_52406_20264# 3.14e-19
C3965 d2 a_22826_29834# 0.273f
C3966 a_16836_11822# a_16836_9916# 0.00396f
C3967 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X2.X1.X1.X2.X2.X2.vin1 0.00232f
C3968 X1.X2.X2.X2.X2.X1.X3.vin2 vdd 0.903f
C3969 a_19336_14688# X1.X2.X1.X2.X1.X2.vout 0.0929f
C3970 X2.X1.X1.X3.vin1 X2.X1.X3.vin2 7.53e-21
C3971 a_11072_7922# vdd 1.05f
C3972 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X3.vin2 0.234f
C3973 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X1.vin1 5.19e-19
C3974 X2.X1.X2.X2.X1.X2.vrefh d2 0.177f
C3975 X2.X1.X3.vin2 a_37466_10734# 6.66e-19
C3976 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X1.X3.vin1 0.0425f
C3977 X1.X2.X1.X2.X2.vrefh a_17222_9916# 8.22e-20
C3978 d2 X1.X2.X2.X1.X1.X1.vout 0.115f
C3979 X2.X1.X2.X1.X1.X1.X3.vin1 X2.X1.X2.X1.X1.X1.X1.vin2 0.22f
C3980 a_52406_16452# a_52492_14586# 3.38e-19
C3981 d3 X2.X2.X1.X2.X2.X1.X3.vin1 0.0195f
C3982 a_37766_5016# a_39966_4110# 4.2e-20
C3983 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X3.vin1 0.206f
C3984 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X2.vin1 0.0689f
C3985 X2.X1.X1.X2.X2.X2.vrefh a_31862_6104# 8.22e-20
C3986 X1.X1.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X1.X3.vin2 0.0533f
C3987 a_2582_25164# a_4396_24258# 1.06e-19
C3988 d0 X2.X2.X1.X1.X1.X1.X3.vin1 4.36e-19
C3989 a_46502_23258# a_48616_22312# 2.95e-20
C3990 d0 X2.X2.X2.X1.X1.X1.X3.vin1 4.36e-19
C3991 a_25712_21264# a_25712_19358# 0.00396f
C3992 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X2.vout 0.2f
C3993 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X1.X3.vin2 1.22e-19
C3994 a_37466_14586# vdd 0.567f
C3995 a_31476_17540# vdd 1.05f
C3996 X2.X2.X2.X1.X3.vin1 a_52406_8828# 9.54e-19
C3997 a_19722_29936# X1.X2.X1.X1.X1.X1.X3.vin2 0.00815f
C3998 X1.X1.X2.vrefh a_5646_892# 7.23e-19
C3999 X2.X2.X2.X1.X2.X1.X1.vin1 vdd 0.592f
C4000 X1.X2.X1.X2.X2.vrefh d1 0.00745f
C4001 a_10686_32700# X1.X2.vrefh 0.3f
C4002 X1.X1.X2.X2.X2.X2.X2.vin1 a_11072_32700# 0.197f
C4003 X1.X2.X2.X2.X2.X2.X3.vin1 vdd 0.993f
C4004 a_33976_22312# vdd 1.05f
C4005 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.vrefh 0.161f
C4006 a_23512_24076# a_23212_22210# 6.71e-19
C4007 a_54606_19358# d0 0.0675f
C4008 X1.X1.X2.vrefh a_2196_4198# 0.119f
C4009 X1.X1.X1.X2.X2.X2.X1.vin1 a_2582_8010# 8.22e-20
C4010 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.vrefh 2.33e-19
C4011 X2.X1.X1.X3.vin2 a_34362_14688# 0.00292f
C4012 a_54606_15546# X2.X2.X2.X1.X2.X2.vrefh 8.22e-20
C4013 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin1 0.52f
C4014 d3 a_23512_8828# 0.00108f
C4015 a_11072_30794# vdd 1.05f
C4016 a_19336_18540# d2 0.0111f
C4017 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X1.vin2 3.94e-19
C4018 a_33676_5198# vdd 1.05f
C4019 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.vout 0.335f
C4020 a_5082_26164# X1.X1.X1.X1.X2.X1.X3.vin2 3.49e-19
C4021 X1.X1.X1.X1.X3.vin2 a_4782_24258# 0.00101f
C4022 d1 a_46116_6104# 2.25e-20
C4023 d3 a_34362_26164# 0.284f
C4024 a_54606_15546# vdd 0.553f
C4025 a_39966_25076# d1 0.00151f
C4026 d1 a_38152_8828# 0.521f
C4027 X2.X1.X1.X2.X1.X1.X3.vin1 a_34062_16634# 0.428f
C4028 X2.X2.X3.vin2 d0 0.034f
C4029 X2.X1.X2.X2.X1.X1.X1.vin2 d0 0.276f
C4030 X2.X2.X1.X1.X2.X1.X1.vin2 d2 0.231f
C4031 X1.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin1 0.00437f
C4032 X1.X2.X2.X1.X1.X1.X3.vin1 a_25326_4110# 0.52f
C4033 X2.X2.X3.vin1 X2.X2.X1.X3.vin2 1.04f
C4034 X1.X1.X2.X1.X1.X2.X3.vin2 a_11072_9828# 0.354f
C4035 d2 X2.X1.X2.X1.X1.X1.X3.vin2 0.0682f
C4036 a_8486_16452# a_10686_15546# 4.2e-20
C4037 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 0.216f
C4038 a_19336_18540# a_17222_17540# 5.36e-21
C4039 X2.X1.X1.X1.X2.X1.X3.vin1 d2 0.104f
C4040 X1.X1.X2.X2.X1.X2.X3.vin1 a_8186_22210# 0.00874f
C4041 a_52406_24076# X2.X2.X2.X2.X1.X2.X3.vin1 0.42f
C4042 X1.X1.X2.X2.X1.X2.X1.vin1 d0 0.267f
C4043 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X3.vin1 0.206f
C4044 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X3.vin2 0.161f
C4045 X1.X1.X1.X1.X2.X2.vout a_4696_18540# 7.93e-20
C4046 X2.X1.X2.X2.X1.X2.X1.vin2 vdd 0.361f
C4047 a_46116_8010# vdd 1.05f
C4048 a_4396_12822# a_4696_10916# 6.48e-19
C4049 d3 X1.X2.X2.X1.X2.X1.vout 0.00226f
C4050 a_10686_9828# d1 0.00151f
C4051 d3 a_46502_11822# 1.89e-19
C4052 X1.X2.X2.X2.X1.X1.X1.vin2 d0 0.276f
C4053 a_37766_20264# X2.X1.X3.vin2 7.93e-20
C4054 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X2.X3.vin1 2.33e-19
C4055 d2 X1.X2.X1.X2.X2.X1.X1.vin2 0.231f
C4056 X2.X1.X2.X2.X1.X2.X1.vin1 a_40352_23170# 0.195f
C4057 X1.X1.X2.X1.X2.X1.vout X1.X1.X2.X1.X2.X1.X3.vin1 0.118f
C4058 a_4782_24258# vdd 0.561f
C4059 a_22826_18358# a_23212_18358# 0.416f
C4060 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X2.vin1 0.564f
C4061 d2 X1.X1.X1.X2.X2.X1.X3.vin1 0.104f
C4062 a_17222_21352# X1.X2.X1.X1.X2.X2.X1.vin2 0.273f
C4063 a_16836_21352# d1 2.25e-20
C4064 X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X3.vin1 0.0604f
C4065 X2.X1.X1.X2.X1.X1.X2.vin1 vdd 0.576f
C4066 a_8486_24076# a_10686_23170# 4.2e-20
C4067 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X3.vin1 1.42e-20
C4068 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X1.vin2 0.216f
C4069 X2.X2.X2.X1.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X3.vin1 0.581f
C4070 a_54992_32700# d1 2.92e-22
C4071 a_25712_21264# d2 0.00414f
C4072 X2.X2.X1.X3.vin1 X2.X2.X2.X2.X3.vin2 7.46e-20
C4073 X2.X2.X2.X1.X2.X1.vout a_52492_14586# 0.169f
C4074 X1.X1.X2.X2.X1.X1.X1.vin2 d0 0.276f
C4075 a_33976_7064# X2.X1.X1.X2.X2.X2.X3.vin1 0.00329f
C4076 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X3.vin2 0.234f
C4077 X2.X2.X2.X1.X1.X2.X2.vin1 vdd 0.576f
C4078 a_25712_25076# d0 0.515f
C4079 a_54606_30794# vdd 0.553f
C4080 X1.X2.X1.X3.vin2 a_19422_12822# 6.03e-19
C4081 a_2582_27070# X1.X1.X1.X1.X2.X1.X1.vin1 8.22e-20
C4082 X1.X1.X2.X2.X1.X1.X3.vin2 d2 0.169f
C4083 X2.X1.X2.X1.X1.X2.X3.vin1 vdd 0.96f
C4084 X2.X2.X1.X2.X2.X1.X2.vin1 X2.X2.X1.X2.X2.X2.vrefh 0.564f
C4085 d1 X2.X2.X1.X2.X2.X2.X2.vin1 0.0144f
C4086 X2.X1.X1.X2.X3.vin1 d1 0.00179f
C4087 a_8572_25982# d2 0.0057f
C4088 a_54606_32700# X2.X2.X2.X2.X2.X2.X2.vin1 0.402f
C4089 d4 X2.X1.X1.X1.X1.X2.X3.vin1 0.00851f
C4090 X1.X1.X2.X2.X1.X2.X3.vin2 d0 4.34e-19
C4091 d2 X1.X1.X2.X1.X3.vin1 0.0619f
C4092 X1.X1.X1.X1.X2.vrefh d0 0.844f
C4093 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X1.vin1 0.0689f
C4094 X2.X2.X2.X1.X1.X2.X3.vin2 a_54606_7922# 7.84e-19
C4095 a_46502_15634# a_46502_13728# 0.00198f
C4096 a_46116_15634# X2.X2.X1.X2.X1.X2.X1.vin1 1.64e-19
C4097 a_8186_10734# X1.X1.X2.X1.X3.vin1 0.385f
C4098 a_52106_22210# d2 0.0191f
C4099 a_52792_12640# a_52492_10734# 6.2e-19
C4100 a_25712_7922# vdd 1.05f
C4101 a_8572_14586# a_10686_13640# 2.95e-20
C4102 a_25326_15546# X1.X2.X2.X1.X2.X2.vrefh 8.22e-20
C4103 d3 X1.X2.X2.X1.X2.X1.X1.vin2 3.99e-21
C4104 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin2 0.12f
C4105 a_37466_29834# X2.X1.X2.X2.X2.X1.X3.vin2 0.00815f
C4106 X2.X2.X1.X1.X1.X2.X3.vin2 d0 4.34e-19
C4107 d4 a_39966_17452# 1.89e-19
C4108 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.vrefh 2.33e-19
C4109 a_34062_16634# X2.X1.X1.X2.X1.X1.vout 0.422f
C4110 X1.X2.X1.X1.X1.X2.X3.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 1.22e-19
C4111 X1.X2.X3.vin2 X1.X2.X2.X1.X2.X2.vout 3.38e-19
C4112 a_39966_7922# a_40352_7922# 0.419f
C4113 a_25326_17452# X1.X2.X2.X1.X2.X2.X3.vin2 0.567f
C4114 a_33976_29936# X2.X1.X1.X1.X1.X1.X3.vin2 0.00546f
C4115 a_8872_16452# vdd 1.05f
C4116 d2 a_48616_29936# 0.606f
C4117 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 2.23e-19
C4118 X1.X1.X1.X2.X1.X1.X3.vin1 d1 0.146f
C4119 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X1.X3.vin2 0.0533f
C4120 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin2 0.1f
C4121 X2.X1.X2.X1.X2.X1.X1.vin1 d1 0.0118f
C4122 a_31476_27070# vdd 1.05f
C4123 X2.X1.X1.X1.X2.X2.X1.vin2 a_31476_19446# 1.78e-19
C4124 a_46116_23258# d1 2.92e-22
C4125 d1 a_23212_6962# 0.00613f
C4126 X2.X2.X3.vin1 X2.X2.X1.X2.X3.vin2 0.0816f
C4127 a_10686_25076# X1.X1.X2.X2.X1.X2.X3.vin1 0.00207f
C4128 a_2196_13728# vdd 1.05f
C4129 X2.X2.X2.X1.X2.X2.X3.vin1 d1 0.146f
C4130 X2.X1.X1.X1.X1.X1.X2.vin1 vdd 0.578f
C4131 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X2.X1.X1.X2.vrefh 0.0128f
C4132 a_37766_12640# a_37466_10734# 5.25e-20
C4133 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X2.vin1 0.564f
C4134 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.vout 0.0898f
C4135 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin2 0.12f
C4136 X2.X1.X1.X2.X2.X1.X1.vin2 a_31476_8010# 1.78e-19
C4137 a_17222_6104# d1 3.41e-19
C4138 d1 a_19036_5198# 0.522f
C4139 a_46116_27070# a_46116_25164# 0.00396f
C4140 a_31476_6104# X2.X1.X1.X2.X2.X2.X1.vin1 0.195f
C4141 a_40352_15546# d1 2.25e-20
C4142 a_4396_12822# X1.X1.X1.X2.X1.X2.X3.vin2 0.101f
C4143 a_10686_28888# vdd 0.541f
C4144 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X3.vin1 1.22e-19
C4145 X2.X2.X1.X1.X2.vrefh a_46502_25164# 8.22e-20
C4146 X1.X1.X3.vin2 a_8486_16452# 3.98e-19
C4147 a_11072_23170# a_11072_21264# 0.00396f
C4148 d2 X2.X2.X1.X2.X1.X1.X3.vin2 0.169f
C4149 d3 a_31862_9916# 0.00112f
C4150 a_25326_25076# X1.X2.X2.X2.X1.X2.X3.vin2 0.567f
C4151 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.vrefh 0.161f
C4152 a_37466_18358# d2 0.00146f
C4153 a_4696_14688# X1.X1.X1.X2.X3.vin1 0.363f
C4154 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.vout 0.118f
C4155 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin1 0.267f
C4156 a_31862_32788# a_31862_30882# 0.00198f
C4157 X2.X1.X2.X2.X1.X2.X3.vin1 d1 0.146f
C4158 X1.X1.X2.X2.X1.X1.X3.vin1 a_8872_20264# 0.199f
C4159 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 2.23e-19
C4160 X1.X2.X3.vin1 X1.X2.X2.X1.X3.vin1 0.00304f
C4161 a_48316_24258# a_48616_22312# 6.1e-19
C4162 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 0.22f
C4163 a_8486_31700# a_10686_30794# 4.2e-20
C4164 d3 X2.X2.X2.X2.X3.vin1 0.375f
C4165 X1.X1.X1.X1.X2.X2.vrefh d2 0.168f
C4166 X1.X1.X2.X1.X1.X2.X3.vin1 d1 0.146f
C4167 X1.X1.X1.X2.X2.vrefh a_2196_9916# 1.64e-19
C4168 X1.X1.X2.X2.X2.X1.X1.vin2 vdd 0.36f
C4169 X1.X1.X1.X2.X1.X2.vout vdd 0.697f
C4170 a_25326_23170# X1.X2.X2.X2.X1.X1.X3.vin2 8.07e-19
C4171 X2.X2.X2.X1.X1.X1.vout d2 0.115f
C4172 X2.X2.X1.X2.X1.X2.X3.vin2 vdd 0.787f
C4173 a_25712_23170# d1 2.25e-20
C4174 X1.X1.X1.X2.X1.X2.X1.vin2 a_2582_11822# 8.88e-20
C4175 d2 a_23512_12640# 3.82e-19
C4176 a_52792_20264# vdd 1.05f
C4177 a_19422_12822# a_19722_10916# 4.41e-20
C4178 X1.X2.X1.X2.X1.X2.X3.vin2 a_19336_10916# 0.00535f
C4179 X2.vrefh d1 7.29e-21
C4180 X2.X1.X1.X1.X2.X1.X3.vin2 d2 0.171f
C4181 a_8872_31700# vdd 1.05f
C4182 X2.X1.X2.X2.X1.X2.vout a_37852_22210# 0.0929f
C4183 d3 X2.X1.X2.X2.X2.X2.X3.vin1 0.0137f
C4184 X1.X1.X2.X2.X1.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin1 0.00437f
C4185 a_48316_20446# a_48616_18540# 6.48e-19
C4186 d2 X1.X1.X1.X2.X2.X1.X3.vin2 0.175f
C4187 a_39966_26982# X2.X1.X2.X2.X2.vrefh 8.22e-20
C4188 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X2.vin1 0.242f
C4189 vout X3.vin2 0.0726f
C4190 a_38152_27888# d3 0.00178f
C4191 X1.X2.X3.vin1 a_19722_14688# 3.28e-19
C4192 d7 a_28482_892# 0.00777f
C4193 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.vrefh 0.161f
C4194 X1.X2.X2.X2.X2.X2.X3.vin2 d2 0.00427f
C4195 X1.X2.X1.X2.X1.X1.vout d1 0.0238f
C4196 d3 a_49002_14688# 0.0469f
C4197 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X3.vin1 0.0321f
C4198 X2.X2.X2.X2.X2.X2.X3.vin1 d1 0.147f
C4199 a_38152_20264# vdd 1.05f
C4200 X2.X2.X1.X1.X2.vrefh d1 0.00745f
C4201 X1.X1.X2.X1.X2.X2.X1.vin1 a_10686_13640# 8.22e-20
C4202 d3 a_4696_10916# 0.621f
C4203 a_48616_26164# X2.X2.X1.X1.X3.vin2 0.0927f
C4204 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X1.X2.X1.X2.X1.X3.vin2 3.94e-19
C4205 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin2 0.12f
C4206 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X1.X2.X3.vin2 3.94e-19
C4207 a_22826_22210# a_23126_20264# 4.19e-20
C4208 d3 a_37852_22210# 7.7e-20
C4209 X1.X2.X2.X2.X2.X1.X1.vin1 a_25326_25076# 8.22e-20
C4210 X1.X1.X1.X1.X2.X1.X1.vin1 d1 0.0118f
C4211 a_8486_27888# d1 0.0749f
C4212 X1.X1.X1.X2.X2.X2.X1.vin2 d0 0.276f
C4213 X1.X2.X1.X2.X2.X1.X3.vin1 a_19036_9010# 0.199f
C4214 d2 a_25326_6016# 4.64e-19
C4215 X1.X3.vin1 X1.X3.vin2 0.514f
C4216 a_17222_25164# d2 0.00328f
C4217 a_40352_30794# d1 2.25e-20
C4218 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X3.vin2 0.102f
C4219 a_22826_10734# X1.X2.X2.X1.X1.X2.X3.vin2 0.00846f
C4220 a_48616_14688# X2.X2.X1.X2.X1.X2.X3.vin1 0.00329f
C4221 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X1.vin1 0.267f
C4222 d2 X2.X2.X1.X1.X1.X1.X3.vin2 0.0661f
C4223 a_5082_18540# X1.X1.X1.X2.X1.X1.X3.vin1 0.00837f
C4224 X1.X1.X2.X1.X2.X1.X3.vin2 a_11072_13640# 0.354f
C4225 d2 a_4782_28070# 0.00202f
C4226 a_31862_27070# a_31862_28976# 0.00198f
C4227 X1.X2.X1.X2.X2.X1.vout d1 0.0238f
C4228 X2.X2.X1.X2.X2.X1.X2.vin1 vdd 0.576f
C4229 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X1.X3.vin2 0.581f
C4230 a_16836_17540# a_16836_15634# 0.00396f
C4231 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X3.vin1 0.00118f
C4232 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X3.vin1 0.206f
C4233 a_23512_20264# vdd 1.05f
C4234 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.vrefh 2.33e-19
C4235 X2.X2.X2.X1.X1.X1.X3.vin2 vdd 0.937f
C4236 a_25326_30794# X1.X2.X2.X2.X2.X2.vrefh 8.22e-20
C4237 a_37466_18358# a_38152_16452# 3.08e-19
C4238 X2.X2.X2.X2.X2.X2.vrefh a_54606_28888# 0.3f
C4239 a_25712_26982# X1.X2.X2.X2.X2.vrefh 1.64e-19
C4240 a_38152_8828# a_37466_6962# 3.31e-19
C4241 X2.X2.X1.X1.X2.X1.X3.vin1 vdd 0.997f
C4242 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X1.vin1 0.206f
C4243 a_34062_31882# X2.X1.X1.X1.X1.X1.vout 0.422f
C4244 a_54606_13640# a_52792_12640# 1.15e-20
C4245 X2.X1.X2.vrefh X2.X3.vin1 0.0451f
C4246 X1.X1.X1.X1.X1.X1.X3.vin1 a_2582_30882# 0.00207f
C4247 a_8572_10734# d1 0.0126f
C4248 a_52106_6962# X2.X2.X2.X1.X1.X1.vout 0.386f
C4249 X1.X1.X2.X1.X2.X2.vrefh vdd 0.415f
C4250 a_46502_25164# X2.X2.X1.X1.X2.X1.X2.vin1 8.88e-20
C4251 a_17222_27070# d1 0.00151f
C4252 X1.X2.X1.X1.X1.X2.X3.vin1 X1.X2.X1.X1.X1.X2.X1.vin2 0.216f
C4253 X2.X2.X2.X1.X1.X2.X1.vin1 X2.X2.X2.X1.X1.X1.X3.vin2 5.19e-19
C4254 X1.X2.X1.X1.X2.X1.X2.vin1 a_17222_23258# 0.402f
C4255 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X3.vin1 0.00118f
C4256 a_8186_18358# X1.X1.X3.vin2 0.451f
C4257 d3 X1.X2.X1.X1.X2.X1.X3.vin2 2.81e-19
C4258 a_46502_13728# X2.X2.X1.X2.X1.X2.X2.vin1 8.88e-20
C4259 X1.X2.X1.X2.X2.X2.X1.vin2 a_16836_4198# 1.78e-19
C4260 X2.X1.X1.X2.X2.X1.X1.vin2 vdd 0.36f
C4261 a_2196_21352# X1.X1.X1.X1.X2.X2.X1.vin1 0.195f
C4262 d0 a_54606_13640# 0.0489f
C4263 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X3.vin1 0.00118f
C4264 X1.X2.X2.X1.X1.X1.X3.vin2 a_23512_5016# 0.1f
C4265 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X2.X1.X1.vin1 0.668f
C4266 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X2.vrefh 0.076f
C4267 X1.X2.X1.X1.X1.X1.vout d1 0.0238f
C4268 a_52492_6962# a_54606_6016# 2.95e-20
C4269 X1.X1.X2.X2.X2.X1.vout a_8486_27888# 0.422f
C4270 X2.X1.X2.X1.X2.X1.vout X2.X1.X2.X1.X3.vin2 0.399f
C4271 X2.X1.X1.X3.vin2 a_34062_9010# 7.93e-20
C4272 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 5.19e-19
C4273 X1.X2.X1.X2.X2.X1.X3.vin1 vdd 0.997f
C4274 X1.X1.X3.vin1 a_8486_8828# 8.66e-20
C4275 d2 a_23212_14586# 0.526f
C4276 d3 X1.X1.X2.X2.X1.X2.vout 0.0232f
C4277 a_23212_18358# a_23126_16452# 3.3e-19
C4278 d3 X2.X2.X2.X1.X1.X2.X3.vin1 2.1e-19
C4279 a_40352_21264# vdd 1.05f
C4280 X1.X1.X1.X2.X1.X1.X3.vin1 a_4396_16634# 0.199f
C4281 a_19722_22312# d2 0.0191f
C4282 X2.X1.X2.X2.X1.X1.vout d4 0.00132f
C4283 X1.X2.X2.X1.X2.X2.X3.vin2 a_22826_14586# 3.85e-19
C4284 a_52106_29834# a_52492_29834# 0.419f
C4285 d3 a_19422_12822# 0.00122f
C4286 X1.X2.X1.X1.X1.X1.X3.vin2 X1.X2.X1.X1.X1.X2.vrefh 0.165f
C4287 a_23212_29834# a_25326_30794# 2.68e-20
C4288 X1.X2.X2.X2.X1.X1.X3.vin2 vdd 0.905f
C4289 a_8486_20264# X1.X1.X3.vin2 7.93e-20
C4290 X2.X1.X1.X1.X3.vin2 vdd 1.32f
C4291 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X3.vin2 0.237f
C4292 a_25712_25076# a_25712_23170# 0.00396f
C4293 d0 X2.X2.X1.X2.X1.X1.X1.vin1 0.267f
C4294 a_8572_25982# X1.X1.X2.X2.X3.vin2 0.0927f
C4295 d5 d6 0.00219f
C4296 a_2196_17540# d2 0.00256f
C4297 X2.X2.X1.X1.X2.X1.X2.vin1 d1 1.03e-19
C4298 d3 X1.X1.X1.X2.X1.X2.X3.vin2 0.0247f
C4299 X2.X1.X1.X3.vin1 a_34362_18540# 0.389f
C4300 a_23512_27888# X1.X2.X2.X2.X2.X1.vout 0.359f
C4301 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 0.139f
C4302 a_48316_20446# d4 0.00107f
C4303 X2.X1.X1.X3.vin2 a_34362_10916# 0.452f
C4304 d3 X1.X2.X2.X2.X1.X2.X3.vin2 0.0247f
C4305 X1.X1.X2.X2.X2.X2.vrefh vdd 0.415f
C4306 X2.X2.X2.X2.X2.X1.X1.vin2 d3 3.99e-21
C4307 X1.X1.X2.X2.X2.X1.X1.vin1 a_11072_26982# 0.195f
C4308 X2.X1.X1.X1.X2.X2.vrefh a_31476_21352# 1.64e-19
C4309 a_52492_6962# d1 0.00613f
C4310 X1.X2.X2.X1.X2.X2.X3.vin1 a_23512_16452# 0.199f
C4311 X1.X2.X2.X2.X2.X1.X3.vin1 d0 4.36e-19
C4312 d0 X2.X1.X2.X1.X1.X1.X1.vin2 0.276f
C4313 a_54992_19358# vdd 1.05f
C4314 a_2582_23258# X1.X1.X1.X1.X2.X2.X1.vin1 8.22e-20
C4315 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X2.X1.X2.X1.X2.vrefh 0.0128f
C4316 X2.X1.X2.X2.vrefh d0 0.848f
C4317 a_16836_25164# a_17222_25164# 0.419f
C4318 d2 X2.X1.X2.X1.X2.X2.X1.vin2 0.231f
C4319 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X2.X1.X1.X2.X1.X1.vin2 0.00232f
C4320 d4 a_23212_18358# 0.63f
C4321 a_33676_20446# d4 0.00107f
C4322 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.X2.vin1 0.00117f
C4323 a_48316_28070# a_46502_27070# 1.15e-20
C4324 X1.X1.X1.X3.vin2 d2 4.4e-19
C4325 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.vrefh 0.267f
C4326 a_31862_32788# a_34062_31882# 4.2e-20
C4327 a_54606_26982# X2.X2.X2.X2.X2.X1.X2.vin1 8.88e-20
C4328 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X2.X1.X3.vin2 8.93e-19
C4329 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.vrefh 0.161f
C4330 X1.X1.X1.X1.X1.X2.X2.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 0.234f
C4331 X2.X1.X2.X2.X1.X1.X1.vin1 vdd 0.592f
C4332 d2 X1.X1.X2.X1.X2.X1.X1.vin1 0.0105f
C4333 a_4396_28070# a_4782_28070# 0.419f
C4334 X1.X2.X2.X2.X1.X2.X1.vin2 d2 0.226f
C4335 d1 X2.X1.X1.X2.X2.X1.vout 0.0238f
C4336 X2.X2.X1.X1.X2.X1.X3.vin2 d0 4.34e-19
C4337 X1.X2.X2.X2.X1.X2.X3.vin1 a_23512_24076# 0.199f
C4338 d4 X2.X1.X1.X2.X1.X1.X3.vin2 4.77e-19
C4339 X1.X2.X2.X1.X2.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X1.vin1 2.23e-19
C4340 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X3.vin1 0.587f
C4341 X1.X2.X1.X1.X1.X1.X1.vin2 a_17222_30882# 8.88e-20
C4342 X1.X2.X2.X2.X2.X1.X1.vin1 d3 6.34e-20
C4343 a_4696_29936# a_5082_29936# 0.419f
C4344 X1.X2.X2.X1.X2.X2.X2.vin1 a_25712_15546# 1.78e-19
C4345 a_8486_12640# a_8572_10734# 3.21e-19
C4346 a_40352_23170# X2.X1.X2.X2.X1.X2.vrefh 1.64e-19
C4347 a_19036_20446# d4 0.00107f
C4348 X1.X2.X1.X2.X2.X1.X3.vin2 a_17222_8010# 0.567f
C4349 X1.X3.vin1 vdd 1.78f
C4350 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X2.X1.X1.X2.X2.vrefh 0.0128f
C4351 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X1.vout 0.033f
C4352 a_46116_13728# d1 2.25e-20
C4353 d5 a_35312_892# 0.04f
C4354 d3 a_46502_32788# 1.28e-19
C4355 d0 a_10686_4110# 0.0675f
C4356 d2 a_54992_13640# 0.00464f
C4357 X1.X1.X1.X2.X1.X1.vout X1.X1.X1.X2.X1.X1.X3.vin2 0.342f
C4358 X1.X2.X2.X2.X1.X1.X1.vin1 vdd 0.592f
C4359 d2 X1.X2.X1.X2.X1.X1.X2.vin1 0.031f
C4360 X2.X2.X2.vrefh a_43362_892# 2.22e-19
C4361 X1.X1.X1.X1.X1.X2.X1.vin2 a_2196_27070# 1.78e-19
C4362 a_54606_28888# d1 0.00148f
C4363 a_8486_16452# d1 0.0749f
C4364 a_52492_29834# a_52792_31700# 6.71e-19
C4365 d2 X2.X1.X2.X1.X2.X1.X3.vin2 0.171f
C4366 X1.X2.X2.X1.X2.X1.X3.vin1 vdd 0.997f
C4367 X1.X1.X2.X1.X1.X1.X2.vin1 a_11072_6016# 0.197f
C4368 a_52492_25982# d2 0.0057f
C4369 d3 a_8186_22210# 0.0474f
C4370 a_37766_27888# a_37852_25982# 3.21e-19
C4371 a_33976_26164# X2.X1.X1.X3.vin1 0.356f
C4372 X2.X1.X1.X1.X1.X2.X3.vin2 a_31862_27070# 0.567f
C4373 a_38152_27888# a_39966_28888# 1.15e-20
C4374 d2 X2.X1.X2.X2.X2.X2.X1.vin2 7.2e-20
C4375 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin2 0.12f
C4376 X2.X1.X1.X2.X3.vin2 d1 0.00807f
C4377 d0 a_2582_11822# 0.0489f
C4378 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X2.X2.vrefh 0.076f
C4379 d2 X2.X2.X1.X1.X1.X2.X3.vin1 0.158f
C4380 a_2582_6104# X1.X1.X1.X2.X2.X2.X3.vin1 0.52f
C4381 a_54606_25076# a_52406_24076# 4.77e-21
C4382 X1.X2.X1.X1.X2.X2.vrefh X1.X1.X2.X2.X1.X2.vrefh 0.117f
C4383 X2.X1.X1.X1.X1.X2.X2.vin1 a_31862_28976# 8.88e-20
C4384 X1.X2.X2.X1.X1.X2.vrefh vdd 0.43f
C4385 a_48316_28070# X2.X2.X1.X1.X1.X2.vout 0.36f
C4386 X2.X1.X1.X2.X1.X2.vrefh a_31476_15634# 0.118f
C4387 X1.X2.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X3.vin2 0.0533f
C4388 X1.X1.X2.X2.X1.X1.X1.vin1 vdd 0.592f
C4389 X2.X1.X2.X1.X2.X2.X2.vin1 d1 1.03e-19
C4390 a_39966_6016# vdd 0.541f
C4391 a_17222_17540# X1.X2.X1.X2.X1.X1.X2.vin1 8.88e-20
C4392 a_52492_6962# X2.X2.X2.X1.X1.X2.vout 0.0929f
C4393 d2 X1.X2.X1.X2.X2.X1.X2.vin1 0.0318f
C4394 X2.X1.X1.X1.X2.X2.X3.vin1 d4 2.08e-19
C4395 a_49002_26164# X2.X2.X1.X1.X3.vin1 0.385f
C4396 X1.X1.X1.X2.vrefh d0 0.844f
C4397 d2 a_54606_17452# 0.00583f
C4398 a_31862_25164# vdd 0.553f
C4399 d0 X1.X2.X2.X1.X2.X2.X3.vin1 4.36e-19
C4400 a_10686_32700# d0 0.0489f
C4401 X1.X1.X1.X1.X2.X1.vout X1.X1.X1.X1.X2.X1.X3.vin2 0.326f
C4402 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X1.X2.X1.X1.X2.vrefh 0.267f
C4403 X1.X1.X2.X1.X3.vin1 a_8486_5016# 1.52e-19
C4404 d2 X1.X1.X2.X1.X1.X1.X3.vin1 3e-19
C4405 d4 X2.X1.X1.X1.X1.X1.X3.vin2 0.0533f
C4406 a_54606_21264# X2.X2.X2.X2.X1.X1.X3.vin1 0.00207f
C4407 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X2.vrefh 0.1f
C4408 a_48702_9010# X2.X2.X1.X2.X2.X1.vout 0.422f
C4409 X1.X1.X2.X2.X2.X1.X2.vin1 a_11072_28888# 0.197f
C4410 X1.X2.X1.X1.X1.X2.X2.vin1 d1 1.03e-19
C4411 d0 a_11072_15546# 0.518f
C4412 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X3.vin2 0.418f
C4413 d2 X2.X2.X2.X1.X2.vrefh 0.158f
C4414 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.X3.vin1 0.587f
C4415 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin1 0.52f
C4416 a_31476_32788# a_31862_32788# 0.419f
C4417 d2 X1.X2.X1.X1.X1.X1.X2.vin1 6e-20
C4418 d0 X1.X2.X1.X2.X1.X2.X1.vin1 0.267f
C4419 a_2582_9916# vdd 0.553f
C4420 a_19336_29936# d1 0.00613f
C4421 d0 X1.X2.X2.X1.X1.X2.X3.vin1 4.36e-19
C4422 X1.X2.X2.X2.X2.X2.X3.vin1 a_23512_31700# 0.199f
C4423 X2.X1.X2.X1.X1.X1.X1.vin2 X2.X2.X1.X2.X2.X2.X2.vin1 0.00232f
C4424 a_40352_28888# d0 0.515f
C4425 X1.X1.X1.X2.X1.X1.vout vdd 0.78f
C4426 a_8486_31700# d1 0.0489f
C4427 d2 X2.X1.X1.X1.X1.X2.vout 0.11f
C4428 X1.X2.X2.X2.X2.X1.X3.vin2 d0 4.34e-19
C4429 d2 a_37852_6962# 0.625f
C4430 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X2.X1.X1.X1.X2.vrefh 0.0128f
C4431 d0 a_11072_7922# 0.518f
C4432 X1.X1.X1.X1.X2.X2.vout d4 9.49e-19
C4433 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin2 0.1f
C4434 a_10686_21264# vdd 0.541f
C4435 d3 X1.X2.X1.X1.X1.X1.X1.vin1 0.00492f
C4436 a_39966_19358# a_39966_17452# 0.00198f
C4437 a_19336_22312# a_19722_22312# 0.419f
C4438 X2.X2.X1.X2.X1.X2.vout vdd 0.697f
C4439 X2.X2.X1.X1.X2.X2.vout a_48316_20446# 0.36f
C4440 a_49002_22312# a_48702_20446# 5.55e-20
C4441 a_16836_32788# X1.X2.X1.X1.X1.X1.X1.vin1 0.195f
C4442 X2.X2.X1.X1.X1.X1.X1.vin2 vdd 0.399f
C4443 X1.X2.X2.X2.X2.X1.vout X1.X2.X2.X2.X2.X2.vout 0.514f
C4444 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X1.X3.vin2 8.93e-19
C4445 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.vrefh 0.161f
C4446 a_37466_29834# X2.X1.X2.X2.X3.vin2 0.422f
C4447 a_23126_27888# X1.X2.X2.X2.X3.vin2 0.00101f
C4448 d0 a_31476_17540# 0.518f
C4449 a_46502_9916# X2.X2.X1.X2.X2.X1.X1.vin2 0.273f
C4450 a_52792_5016# vdd 1.05f
C4451 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X3.vin1 0.00117f
C4452 X1.X2.X2.X1.X2.X1.X3.vin2 a_23126_12640# 0.267f
C4453 X1.X1.X1.X3.vin1 vdd 1.27f
C4454 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.vout 0.075f
C4455 a_37852_14586# a_38152_12640# 6.1e-19
C4456 X1.X2.X2.X2.X1.X2.vrefh d1 0.0071f
C4457 d0 X2.X2.X2.X1.X2.X1.X1.vin1 0.267f
C4458 X1.X2.X2.X2.X1.X2.vrefh a_25326_21264# 0.3f
C4459 X2.X2.X2.X2.X1.X2.X3.vin1 a_52106_22210# 0.00874f
C4460 d2 a_33676_12822# 6.04e-19
C4461 X1.X2.X2.X2.X2.X2.X3.vin1 d0 4.36e-19
C4462 d3 a_10686_25076# 1.89e-19
C4463 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X3.vin2 0.234f
C4464 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X1.X3.vin1 0.0321f
C4465 d2 a_54606_7922# 0.00479f
C4466 a_8186_18358# d1 0.0424f
C4467 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X2.vrefh 0.00118f
C4468 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X3.vin1 0.581f
C4469 a_48616_10916# X2.X2.X1.X2.X2.X1.vout 1.64e-19
C4470 a_49002_10916# a_48702_9010# 5.25e-20
C4471 a_11072_30794# d0 0.518f
C4472 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X3.vin1 0.00117f
C4473 a_48316_28070# d3 0.00108f
C4474 a_37466_22210# a_38152_20264# 2.86e-19
C4475 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X2.vout 0.398f
C4476 a_16836_17540# vdd 1.05f
C4477 X2.X2.X2.X2.X1.X1.X3.vin1 a_52106_18358# 0.00837f
C4478 a_31862_15634# a_33976_14688# 2.95e-20
C4479 d0 a_54606_15546# 0.0675f
C4480 X1.X1.X1.X1.X1.X1.vout X1.X1.X1.X1.X1.X1.X3.vin2 0.342f
C4481 a_8186_29834# X1.X1.X2.X2.X2.X2.X3.vin1 0.00874f
C4482 a_52406_27888# a_52792_27888# 0.419f
C4483 X2.X2.X2.X2.X2.X1.X3.vin1 a_52492_25982# 0.00251f
C4484 a_54606_21264# a_54992_21264# 0.419f
C4485 X1.X1.X1.X1.X1.X1.vout vdd 0.781f
C4486 X2.X2.X1.X1.X2.X1.X3.vin2 a_46116_23258# 0.354f
C4487 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X1.X3.vin2 5.19e-19
C4488 a_8486_20264# d1 0.0749f
C4489 a_46502_21352# X2.X2.X1.X1.X2.X2.X1.vin1 0.417f
C4490 a_46116_21352# X2.X2.X1.X1.X2.X2.X3.vin1 0.354f
C4491 d6 X3.vin2 3.1f
C4492 a_25712_17452# X1.X2.X2.X1.X2.X2.X1.vin2 1.78e-19
C4493 a_2196_32788# d1 2.25e-20
C4494 a_2582_32788# X1.X1.X1.X1.X1.X1.X2.vin1 8.88e-20
C4495 X2.X2.X3.vin1 a_52406_16452# 8.66e-20
C4496 X2.X1.X2.X2.X1.X2.X1.vin2 d0 0.276f
C4497 d6 a_20672_892# 0.00114f
C4498 X1.X1.X1.X1.X2.X1.vout a_4696_22312# 0.169f
C4499 a_25326_11734# X1.X2.X2.X1.X2.vrefh 8.22e-20
C4500 a_52106_14586# X2.X2.X2.X1.X2.X1.X3.vin2 0.00815f
C4501 a_4782_24258# a_5082_22312# 4.19e-20
C4502 X1.X1.X2.X1.X1.X1.X2.vin1 vdd 0.578f
C4503 d0 a_46116_8010# 0.515f
C4504 a_11072_32700# d2 3.9e-19
C4505 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 0.139f
C4506 X2.X1.X1.X1.X1.X2.vrefh a_31476_30882# 0.118f
C4507 d2 X2.X1.X1.X2.X2.X1.X2.vin1 0.0318f
C4508 X2.X1.X2.X1.X2.X2.X1.vin1 X2.X2.X1.X2.X1.X2.vrefh 0.00437f
C4509 X1.X2.X3.vin2 X1.X2.X2.vrefh 0.15f
C4510 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 0.139f
C4511 X1.X2.X1.X1.X1.X1.X1.vin2 a_19422_31882# 0.00743f
C4512 X1.X1.X2.X1.X1.X2.X3.vin2 a_10686_7922# 7.84e-19
C4513 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X1.vin1 0.0689f
C4514 a_11072_6016# a_11072_4110# 0.00396f
C4515 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin2 0.1f
C4516 a_48616_10916# a_49002_10916# 0.414f
C4517 X1.X1.X2.X1.X2.X1.X2.vin1 d1 1.03e-19
C4518 a_39966_6016# X2.X1.X2.X1.X1.X1.X3.vin1 0.00207f
C4519 d0 X2.X1.X1.X2.X1.X1.X2.vin1 0.262f
C4520 a_5082_14688# X1.X1.X1.X2.X1.X2.X3.vin2 3.85e-19
C4521 a_19422_16634# a_19722_14688# 4.19e-20
C4522 d2 a_25326_13640# 0.00665f
C4523 a_39966_26982# d2 0.00328f
C4524 X1.X2.X1.X2.X1.X1.vout a_19336_14688# 0.169f
C4525 X1.X1.X1.X2.X3.vin1 a_4782_12822# 9.54e-19
C4526 X1.X1.X2.X2.X1.X1.vout X1.X1.X2.X2.X1.X1.X3.vin1 0.118f
C4527 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X3.vin2 0.0533f
C4528 X1.X2.X1.X1.X1.X2.X1.vin1 d1 0.0118f
C4529 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X1.vin2 0.076f
C4530 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X1.X3.vin2 0.0943f
C4531 d0 X2.X2.X2.X1.X1.X2.X2.vin1 0.262f
C4532 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X1.X2.X2.X2.X2.X3.vin2 8.93e-19
C4533 X2.X1.X1.X1.X1.X2.X2.vin1 X2.X1.X1.X1.X1.X2.X3.vin2 0.234f
C4534 a_33676_28070# a_34062_28070# 0.419f
C4535 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X3.vin2 0.161f
C4536 a_54606_30794# d0 0.0675f
C4537 a_25326_32700# vdd 0.541f
C4538 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X3.vin1 2.33e-19
C4539 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X1.X2.X2.X3.vin2 1.22e-19
C4540 X2.X1.X2.X1.X3.vin2 a_37852_10734# 0.0927f
C4541 d0 X2.X1.X2.X1.X1.X2.X3.vin1 4.36e-19
C4542 X1.X2.X2.X3.vin2 d2 4.4e-19
C4543 d2 a_31862_28976# 0.00479f
C4544 a_25326_28888# a_25326_30794# 0.00198f
C4545 d2 a_23212_10734# 0.0057f
C4546 X1.X2.X1.X2.X1.X1.X1.vin2 d1 1.49e-19
C4547 X2.X2.X2.X1.X2.X1.X3.vin2 vdd 0.903f
C4548 d0 a_25712_7922# 0.518f
C4549 a_54606_23170# X2.X2.X2.X2.X1.X1.X3.vin2 8.07e-19
C4550 X1.X2.X2.X1.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin1 0.00437f
C4551 a_39966_25076# X2.X1.X2.X2.X1.X2.X1.vin2 8.88e-20
C4552 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X1.vin2 0.076f
C4553 a_39966_13640# X2.X1.X2.X1.X2.X1.X1.vin2 8.88e-20
C4554 a_46116_8010# a_46116_6104# 0.00396f
C4555 a_11072_25076# vdd 1.05f
C4556 X3.vin2 a_35312_892# 5.64e-19
C4557 a_37466_29834# d1 0.0422f
C4558 a_37466_29834# X2.X1.X2.X2.X2.X2.vout 0.263f
C4559 X2.X1.X2.X2.X1.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin1 0.00437f
C4560 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X3.vin2 0.0321f
C4561 a_52406_27888# vdd 0.561f
C4562 d2 X1.X2.X1.X2.X1.X1.X1.vin1 0.0116f
C4563 d1 a_38152_5016# 0.522f
C4564 X1.X1.X1.X1.X1.X2.X2.vin1 vdd 0.576f
C4565 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X2.X3.vin1 0.0174f
C4566 a_46116_19446# a_46116_17540# 0.00396f
C4567 X1.X1.X2.X1.X2.X1.X1.vin2 a_11072_11734# 0.12f
C4568 a_10686_11734# X1.X1.X2.X1.X2.X1.X1.vin1 0.417f
C4569 a_31476_27070# d0 0.515f
C4570 X1.X2.X2.X1.X2.X1.X1.vin1 a_25712_9828# 1.64e-19
C4571 X1.X2.X2.X1.X1.X2.X3.vin1 a_23212_6962# 0.00329f
C4572 a_48702_20446# d1 0.0749f
C4573 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.vrefh 0.267f
C4574 X1.X1.X2.X2.X3.vin1 a_8186_22210# 0.436f
C4575 a_39966_15546# a_39966_13640# 0.00198f
C4576 d2 a_37766_5016# 0.00123f
C4577 X2.X2.X2.X2.X2.vrefh a_54606_25076# 0.3f
C4578 d0 a_2196_13728# 0.518f
C4579 a_52492_18358# a_54606_17452# 4.72e-20
C4580 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X2.vout 0.197f
C4581 X2.X1.X1.X1.X1.X1.X2.vin1 d0 0.262f
C4582 X1.X1.X1.X2.X1.X2.X2.vin1 a_2196_11822# 0.197f
C4583 a_46502_15634# a_48616_14688# 2.95e-20
C4584 d4 X1.X2.X2.X2.X3.vin2 0.0939f
C4585 a_16836_17540# X1.X2.X1.X2.X1.X1.X3.vin1 0.354f
C4586 X2.X1.X2.X1.X1.X2.X3.vin1 a_38152_8828# 0.199f
C4587 d1 d6 4.67e-19
C4588 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.X3.vin2 0.0523f
C4589 a_17222_17540# X1.X2.X1.X2.X1.X1.X1.vin1 0.417f
C4590 a_10686_28888# d0 0.0489f
C4591 a_33976_18540# d1 0.00616f
C4592 X1.X2.X2.X2.X3.vin2 a_23126_31700# 9.7e-20
C4593 X2.X2.X1.X3.vin2 d2 4.4e-19
C4594 X2.X2.X1.X2.X1.X2.X2.vin1 a_46116_11822# 0.197f
C4595 a_34062_20446# d1 0.0749f
C4596 d2 X1.X1.X1.X1.X3.vin1 0.0594f
C4597 X2.X1.X1.X2.X2.X1.X3.vin2 a_31862_6104# 8.07e-19
C4598 a_52406_12640# X2.X2.X2.X1.X2.X1.X3.vin1 0.428f
C4599 d2 a_8186_6962# 0.272f
C4600 X1.X2.X2.X1.X1.X2.X1.vin2 X2.X1.X1.X2.X2.X2.vrefh 0.0128f
C4601 X2.X1.X2.X1.X1.X1.X1.vin1 vdd 0.592f
C4602 a_10686_6016# a_8872_5016# 1.15e-20
C4603 a_16836_13728# X1.X2.X1.X2.X1.X2.X2.vin1 1.78e-19
C4604 X1.X2.X1.X2.X3.vin1 vdd 0.804f
C4605 a_8572_22210# vdd 1.05f
C4606 a_33976_26164# a_33676_24258# 6.2e-19
C4607 a_22826_29834# X1.X2.X2.X2.X2.X1.vout 0.383f
C4608 X1.X1.X2.X2.X2.X1.X1.vin2 d0 0.276f
C4609 a_31476_9916# X2.X1.X1.X2.X2.X1.X1.vin1 0.195f
C4610 X2.X1.X1.X1.X1.X1.X1.vin2 d1 0.00147f
C4611 d0 X2.X2.X1.X2.X1.X2.X3.vin2 4.34e-19
C4612 a_2582_6104# X1.X1.X1.X2.X2.X2.X2.vin1 8.88e-20
C4613 X1.X1.X2.X3.vin2 a_8486_24076# 6.03e-19
C4614 a_43362_892# X2.X3.vin2 0.255f
C4615 a_46502_13728# X2.X2.X1.X2.X1.X2.X1.vin2 0.273f
C4616 a_19422_20446# d1 0.0749f
C4617 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X3.vin2 8.93e-19
C4618 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X2.X1.X1.X1.X2.vrefh 0.00437f
C4619 X1.X1.X2.X1.X1.X2.X3.vin1 a_11072_7922# 0.354f
C4620 X2.X2.X2.X1.X1.X1.X3.vin2 X2.X2.X2.X1.X1.X1.X1.vin2 8.93e-19
C4621 X2.X2.X2.X1.X1.X1.X2.vin1 a_54606_4110# 8.88e-20
C4622 X2.X2.X3.vin1 a_49002_7064# 9.8e-19
C4623 d3 X2.X1.X2.X2.X2.X1.X3.vin2 0.0952f
C4624 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 0.234f
C4625 a_10686_13640# X1.X1.X2.X1.X2.X1.X3.vin1 0.00207f
C4626 X2.X1.X1.X1.X1.X1.X1.vin1 d2 0.00798f
C4627 a_31476_11822# vdd 1.05f
C4628 a_4396_9010# a_2582_8010# 1.15e-20
C4629 a_46502_9916# d1 3.95e-19
C4630 X2.X2.X2.X1.X2.X2.X3.vin1 a_54606_15546# 0.52f
C4631 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.X1.X1.vin1 5.19e-19
C4632 a_33676_16634# a_34362_14688# 2.86e-19
C4633 a_33676_12822# a_31862_11822# 1.15e-20
C4634 a_34062_16634# a_33976_14688# 3.14e-19
C4635 X2.X2.X2.X2.X2.X2.X1.vin2 vrefl 0.0763f
C4636 X2.X2.X1.X2.X1.X1.X2.vin1 a_46116_15634# 0.197f
C4637 X1.X2.X1.X2.X2.X2.vout X1.X2.X1.X2.X2.X2.X3.vin2 0.08f
C4638 X2.X2.X2.X2.X2.X1.X3.vin2 a_54992_28888# 0.354f
C4639 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.vout 0.335f
C4640 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.vrefh 0.161f
C4641 d1 a_35312_892# 5.18e-19
C4642 X2.vrefh X1.X2.X2.X2.X2.X2.X3.vin1 0.00118f
C4643 a_40352_28888# a_40352_30794# 0.00396f
C4644 a_54606_21264# d1 0.00148f
C4645 X2.X2.X1.X1.X2.X1.X2.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 0.234f
C4646 a_11072_4110# vdd 1.05f
C4647 X1.X1.X2.X1.X1.X1.X3.vin2 a_8186_6962# 0.00815f
C4648 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X2.X3.vin1 0.206f
C4649 a_2196_15634# d1 2.92e-22
C4650 X1.X2.X3.vin1 a_22826_6962# 6.45e-19
C4651 a_31862_15634# vdd 0.541f
C4652 X2.X1.X1.X1.X2.X2.vrefh vdd 0.415f
C4653 a_54992_25076# a_54992_23170# 0.00396f
C4654 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin2 7.84e-19
C4655 d2 X1.X1.X2.X1.X1.X2.vrefh 6.65e-20
C4656 X1.X1.X1.X2.X2.X2.vrefh vdd 0.415f
C4657 X2.X2.X1.X1.X2.X2.X3.vin1 d2 0.153f
C4658 d0 X2.X2.X1.X2.X2.X1.X2.vin1 0.262f
C4659 a_23212_25982# d1 0.0126f
C4660 d0 X2.X2.X2.X1.X1.X1.X3.vin2 4.34e-19
C4661 X2.X1.X2.X2.X2.X1.X3.vin1 d1 0.151f
C4662 X2.X2.X1.X1.X2.X1.X3.vin1 d0 4.36e-19
C4663 a_52792_8828# a_54606_7922# 1.06e-19
C4664 a_25326_19358# a_23212_18358# 5.36e-21
C4665 d1 X2.X2.X2.X1.X1.X1.X1.vin1 0.0118f
C4666 X1.X1.X2.X1.X2.X1.X1.vin2 vdd 0.36f
C4667 d2 X2.X2.X1.X2.X3.vin2 0.0501f
C4668 a_17222_23258# vdd 0.541f
C4669 a_2196_8010# d1 2.92e-22
C4670 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 0.216f
C4671 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X1.vin2 0.242f
C4672 a_37766_24076# a_39966_23170# 4.2e-20
C4673 d0 X1.X1.X2.X1.X2.X2.vrefh 0.848f
C4674 a_19336_18540# a_19722_18540# 0.413f
C4675 a_37852_22210# a_39966_21264# 2.95e-20
C4676 a_54606_21264# a_54606_19358# 0.00198f
C4677 X2.X2.X2.X1.X1.X1.X3.vin1 X2.X2.X2.X1.X1.X1.X1.vin1 0.206f
C4678 d3 a_37852_18358# 7.7e-20
C4679 d3 a_38152_12640# 0.00178f
C4680 a_2196_28976# d1 2.25e-20
C4681 X2.X1.X1.X1.X1.X2.X3.vin2 d2 0.122f
C4682 X1.X2.X2.X2.X2.X1.X1.vin2 a_25326_28888# 8.88e-20
C4683 d0 X2.X1.X1.X2.X2.X1.X1.vin2 0.276f
C4684 X1.X1.X1.X2.X2.X2.X2.vin1 X1.X1.X2.vrefh 0.564f
C4685 X1.X1.X2.X1.X2.X2.X3.vin1 a_8572_14586# 0.00329f
C4686 a_8486_5016# X1.X1.X2.X1.X1.X1.X3.vin1 0.428f
C4687 X1.X1.X2.X2.X2.X2.X3.vin2 vdd 0.738f
C4688 a_48616_14688# X2.X2.X1.X2.X3.vin1 0.363f
C4689 a_10686_17452# X1.X1.X2.X1.X2.X2.X1.vin2 8.88e-20
C4690 d2 a_11072_28888# 0.00464f
C4691 d2 X2.X1.X2.X1.X3.vin2 0.00194f
C4692 d0 X1.X2.X1.X2.X2.X1.X3.vin1 4.36e-19
C4693 a_42976_892# vdd 1.05f
C4694 X2.X2.X1.X2.X2.vrefh d1 0.00745f
C4695 a_39966_13640# vdd 0.541f
C4696 a_5082_29936# a_4782_28070# 5.55e-20
C4697 a_40352_21264# d0 0.515f
C4698 a_2196_30882# d1 2.92e-22
C4699 a_2582_30882# X1.X1.X1.X1.X1.X1.X2.vin1 0.402f
C4700 X2.X2.X1.X3.vin1 vdd 1.27f
C4701 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X3.vin2 8.93e-19
C4702 a_31862_30882# vdd 0.541f
C4703 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X2.vin1 0.564f
C4704 d1 X1.X2.X2.X1.X1.X1.X1.vin1 0.013f
C4705 X2.X2.X2.X1.X2.X2.X2.vin1 a_54992_15546# 1.78e-19
C4706 a_46502_28976# vdd 0.553f
C4707 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X1.vin1 2.23e-19
C4708 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.vrefh 0.165f
C4709 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X1.vin2 0.22f
C4710 X1.X2.X2.X2.X1.X1.X3.vin2 d0 4.34e-19
C4711 X2.X1.X2.X3.vin2 a_37852_18358# 0.0927f
C4712 a_17222_11822# a_17222_9916# 0.00198f
C4713 X1.X1.X1.X1.X1.X2.vout d1 0.033f
C4714 a_52106_18358# d1 0.0424f
C4715 a_16836_11822# X1.X2.X1.X2.X2.X1.X1.vin1 1.64e-19
C4716 X2.X2.X2.X2.X2.X1.X1.vin1 a_54992_25076# 1.64e-19
C4717 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X3.vin1 2.33e-19
C4718 a_23212_25982# a_23126_24076# 3.3e-19
C4719 X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.vout 0.398f
C4720 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 1.22e-19
C4721 X2.X1.X2.X1.X1.X1.X3.vin1 X2.X1.X2.X1.X1.X1.X1.vin1 0.206f
C4722 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X3.vin1 2.33e-19
C4723 X1.X1.X1.X1.X2.X1.X3.vin1 a_4396_24258# 0.199f
C4724 X1.X2.X1.X2.X3.vin2 a_19722_7064# 0.422f
C4725 X1.X1.X2.X2.X2.X2.vrefh d0 0.848f
C4726 X2.X1.X1.X2.X1.X1.X1.vin1 vdd 0.592f
C4727 a_17222_11822# d1 0.00151f
C4728 a_19036_24258# d2 3.82e-19
C4729 X2.X2.X2.X2.X2.X2.X3.vin1 a_54606_30794# 0.52f
C4730 X1.X1.X2.X2.X1.X2.X3.vin1 d1 0.146f
C4731 a_54992_19358# d0 0.518f
C4732 X1.X1.X2.X2.X2.X2.X3.vin2 X1.X2.vrefh 0.183f
C4733 a_23512_27888# vdd 1.05f
C4734 X2.X1.X1.X1.X2.X2.vout vdd 0.865f
C4735 a_48316_16634# a_48616_14688# 6.1e-19
C4736 X1.X2.X2.X1.X1.X2.X1.vin1 a_25712_6016# 1.64e-19
C4737 d4 X2.X1.X3.vin2 0.288f
C4738 a_37466_6962# a_38152_5016# 2.86e-19
C4739 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X3.vin1 0.0131f
C4740 a_54992_25076# d1 2.92e-22
C4741 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X1.vin2 0.076f
C4742 a_54992_15546# X2.X2.X2.X1.X2.X2.vrefh 1.64e-19
C4743 X2.X2.X1.X1.X1.X1.X2.vin1 a_46116_30882# 0.197f
C4744 X2.X1.X1.X2.X1.X1.X1.vin2 a_31862_15634# 8.88e-20
C4745 X1.X2.X3.vin1 d2 0.1f
C4746 X2.X2.X2.X2.X1.X2.X1.vin2 X2.X2.X2.X2.X1.X2.X1.vin1 0.668f
C4747 X1.X1.X2.X1.X1.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin2 0.0128f
C4748 d1 X2.X2.X1.X2.X2.X2.X1.vin1 0.0118f
C4749 X2.X1.X1.X2.X2.X2.X3.vin2 vdd 0.725f
C4750 a_25326_15546# d1 3.41e-19
C4751 X1.X1.X1.X1.X2.X1.X3.vin2 d2 0.171f
C4752 X2.X1.X2.X1.X2.X2.vout a_37852_14586# 0.0929f
C4753 X2.X1.X2.X2.X1.X2.X3.vin2 d1 0.171f
C4754 X2.X2.X1.X2.X2.X2.vout a_48702_5198# 0.418f
C4755 a_54992_15546# vdd 1.05f
C4756 X2.X1.X2.X2.X1.X1.X1.vin1 d0 0.267f
C4757 d3 X2.X1.X2.X1.X3.vin1 0.0869f
C4758 X2.X2.X1.X1.X1.X2.X1.vin2 X2.X2.X1.X1.X1.X2.vrefh 0.1f
C4759 a_52106_18358# X2.X2.X3.vin2 0.451f
C4760 X2.X2.X2.X2.X1.X2.X2.vin1 d2 0.0329f
C4761 X2.X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X2.X2.vrefh 0.117f
C4762 X1.X1.X1.X1.X3.vin1 X1.X1.X2.X2.X3.vin2 0.0604f
C4763 X1.X2.X2.X1.X1.X1.X3.vin1 a_25712_4110# 0.354f
C4764 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X3.vin2 8.93e-19
C4765 a_52406_24076# vdd 0.47f
C4766 a_31476_13728# X2.X1.X1.X2.X1.X2.X1.vin1 0.195f
C4767 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X2.X2.X1.vin1 0.206f
C4768 X1.X1.X3.vin2 X1.X1.X2.X1.X3.vin2 0.039f
C4769 X2.X1.X2.X1.X2.X1.X3.vin1 a_38152_12640# 0.199f
C4770 a_25712_9828# d1 2.92e-22
C4771 d0 X1.X3.vin1 0.0254f
C4772 d1 a_16836_8010# 2.92e-22
C4773 X2.X1.X2.X2.X1.X2.X1.vin1 vdd 0.592f
C4774 X1.X1.X1.X2.X1.X2.X3.vin2 a_4696_10916# 0.00535f
C4775 a_4782_12822# a_5082_10916# 4.41e-20
C4776 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X2.vrefh 0.00118f
C4777 X1.X1.X1.X2.X1.X1.X2.vin1 a_2582_15634# 0.402f
C4778 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin2 0.12f
C4779 X1.X2.X2.X2.X1.X1.X1.vin1 d0 0.267f
C4780 d3 X2.X2.X2.X1.X2.X1.X1.vin2 3.99e-21
C4781 X1.X1.X2.X1.X1.X2.X3.vin2 d1 0.171f
C4782 X1.X1.X2.X2.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin2 0.0128f
C4783 d2 X1.X2.X2.X1.X1.X2.X2.vin1 0.0329f
C4784 d5 a_14082_892# 4.95e-19
C4785 X2.X1.X1.X1.X1.X2.X1.vin1 a_31862_30882# 8.22e-20
C4786 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X2.X1.X1.X2.X1.X2.vin1 0.00232f
C4787 d0 X1.X2.X2.X1.X2.X1.X3.vin1 4.36e-19
C4788 X2.X2.X2.X1.X1.X2.X1.vin2 a_54606_7922# 0.273f
C4789 a_39966_28888# X2.X1.X2.X2.X2.X1.X3.vin2 0.567f
C4790 X2.X1.X1.X1.X2.vrefh X1.X2.X2.X2.X2.vrefh 0.117f
C4791 a_10686_28888# a_8486_27888# 4.77e-21
C4792 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X1.vin1 5.19e-19
C4793 a_52106_10734# d1 0.0318f
C4794 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X2.X1.X3.vin1 2.33e-19
C4795 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X1.X2.X2.X1.vin2 0.216f
C4796 X1.X2.X1.X1.X2.X2.X1.vin1 d1 0.0118f
C4797 a_34062_16634# vdd 0.561f
C4798 a_52492_25982# X2.X2.X2.X2.X3.vin2 0.0927f
C4799 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X1.vin2 0.076f
C4800 d0 X1.X2.X2.X1.X1.X2.vrefh 0.848f
C4801 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X1.vin2 0.076f
C4802 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X1.vin1 0.206f
C4803 X1.X1.X2.vrefh d5 0.00132f
C4804 a_31862_21352# d2 0.00393f
C4805 X1.X1.X2.X2.X1.X1.X1.vin1 d0 0.267f
C4806 X2.X2.X2.X1.X3.vin1 a_52406_5016# 1.52e-19
C4807 X2.X1.X1.X2.X2.X2.vout X2.X1.X1.X2.X2.X2.X3.vin1 0.335f
C4808 d4 X1.X1.X2.X1.X2.X2.X3.vin1 2.52e-19
C4809 a_25326_30794# d1 3.41e-19
C4810 d0 a_39966_6016# 0.0489f
C4811 X1.X1.X1.X1.X2.X1.X2.vin1 a_2582_23258# 0.402f
C4812 a_39966_11734# a_39966_9828# 0.00198f
C4813 a_54992_30794# vdd 1.05f
C4814 a_46116_4198# a_46502_4198# 0.419f
C4815 a_37852_14586# d1 0.00613f
C4816 a_31862_25164# d0 0.0675f
C4817 d1 a_48702_5198# 0.0751f
C4818 X2.X2.X2.vrefh a_46502_4198# 0.301f
C4819 a_22826_6962# X1.X2.X2.X1.X1.X1.X3.vin2 0.00815f
C4820 a_10686_32700# a_8486_31700# 4.77e-21
C4821 X1.X2.X2.X1.X2.X2.vout vdd 0.865f
C4822 a_19722_26164# d2 7.13e-19
C4823 X2.X2.X2.X2.X2.X2.X2.vin1 X2.X2.X2.X2.X2.X2.X3.vin2 0.237f
C4824 X2.X1.X3.vin2 a_37766_8828# 2.33e-19
C4825 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.vout 0.0898f
C4826 a_19036_12822# X1.X2.X1.X2.X1.X2.X3.vin2 0.101f
C4827 a_25712_15546# X1.X2.X2.X1.X2.X2.vrefh 1.64e-19
C4828 a_8572_14586# X1.X1.X2.X1.X2.X1.X3.vin2 0.00546f
C4829 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X1.vin2 0.668f
C4830 X1.X1.X1.X1.X2.X2.X2.vin1 vdd 0.576f
C4831 d3 X1.X2.X2.X1.X2.X1.X1.vin1 6.34e-20
C4832 d4 X2.X1.X2.X1.X2.X2.X3.vin2 0.0264f
C4833 a_52106_22210# X2.X2.X2.X2.X1.X1.vout 0.387f
C4834 a_17222_25164# X1.X2.X1.X1.X2.X1.X2.vin1 8.88e-20
C4835 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X1.X2.X1.vin2 8.93e-19
C4836 d3 X1.X1.X3.vin2 0.77f
C4837 X2.X1.X1.X1.X1.X2.vout X2.X1.X1.X1.X1.X1.vout 0.507f
C4838 d0 a_2582_9916# 0.0675f
C4839 d2 X2.X2.X1.X1.X3.vin1 0.0594f
C4840 a_39966_11734# a_37852_10734# 5.36e-21
C4841 X2.X2.X3.vin2 a_52106_10734# 6.66e-19
C4842 d1 a_34362_7064# 0.0422f
C4843 X1.X2.X2.X1.X1.X2.vout vdd 0.696f
C4844 d2 X1.X1.X2.X1.X2.X1.vout 0.00174f
C4845 a_54992_17452# X2.X2.X2.X1.X2.X2.X1.vin2 1.78e-19
C4846 X2.X2.X1.X1.X2.X2.X3.vin2 a_46502_17540# 8.07e-19
C4847 a_4696_22312# d2 0.526f
C4848 a_22826_22210# d4 2.94e-19
C4849 X1.X1.X1.X3.vin1 a_5082_22312# 7.98e-19
C4850 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X3.vin1 0.587f
C4851 a_25712_28888# vdd 1.05f
C4852 a_22826_22210# a_23212_22210# 0.419f
C4853 X1.X1.X1.X2.X1.X2.X1.vin1 vdd 0.592f
C4854 X2.X1.X2.X1.X1.X1.X2.vin1 a_40352_6016# 0.197f
C4855 a_34062_31882# vdd 0.565f
C4856 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X2.X1.X1.X2.vrefh 0.00437f
C4857 a_10686_21264# d0 0.0489f
C4858 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X1.X3.vin1 0.0425f
C4859 a_48616_29936# a_49002_29936# 0.419f
C4860 d1 X1.X2.X1.X2.X2.X2.X3.vin2 0.214f
C4861 X2.X1.X2.vrefh a_31476_4198# 0.119f
C4862 d0 X2.X2.X1.X1.X1.X1.X1.vin2 0.201f
C4863 X2.X1.X1.X1.X2.X1.X1.vin1 X2.X1.X1.X1.X2.X1.X1.vin2 0.668f
C4864 X1.X2.X1.X2.X2.X2.X3.vin1 d1 0.149f
C4865 d3 X2.X2.X1.X2.X2.X1.X1.vin2 3.99e-21
C4866 a_46116_27070# X2.X2.X1.X1.X2.X1.X1.vin1 1.64e-19
C4867 X1.X1.X2.X2.X2.X1.X3.vin2 vdd 0.903f
C4868 a_46502_27070# a_46502_25164# 0.00198f
C4869 a_31862_6104# X2.X1.X1.X2.X2.X2.X3.vin1 0.52f
C4870 d4 a_19722_29936# 5.68e-19
C4871 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X3.vin1 2.33e-19
C4872 a_8186_6962# a_8486_5016# 4.19e-20
C4873 X1.X2.X2.X3.vin2 X1.X2.X3.vin2 0.171f
C4874 d3 X2.X1.X1.X2.X2.X1.X3.vin1 0.0195f
C4875 X1.X2.X1.X3.vin2 d1 0.0129f
C4876 a_4696_26164# X1.X1.X1.X1.X1.X2.vout 7.93e-20
C4877 a_19036_28070# X1.X2.X1.X1.X1.X2.vout 0.36f
C4878 X1.X2.X2.X2.X2.X2.vout vdd 0.698f
C4879 X2.X2.X1.X1.X1.X2.vrefh X2.X1.X2.X2.X2.X2.vrefh 0.117f
C4880 X2.X1.X1.X1.X1.X1.X3.vin1 a_31862_30882# 0.00207f
C4881 a_48702_24258# a_49002_22312# 4.19e-20
C4882 X2.X2.X1.X1.X2.X1.vout a_48616_22312# 0.169f
C4883 X1.X1.X2.X2.X2.X2.X3.vin1 X1.X1.X2.X2.X2.X2.X1.vin1 0.206f
C4884 X1.X1.X3.vin2 X1.X1.X2.vrefh 0.15f
C4885 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X1.vin1 0.267f
C4886 X1.X1.X2.X2.X2.X1.X1.vin1 vdd 0.592f
C4887 a_2582_32788# X1.X1.X1.X1.X1.X1.X1.vin2 0.273f
C4888 X1.X2.X1.X2.X1.X2.X2.vin1 d1 1.03e-19
C4889 a_4396_20446# a_4782_20446# 0.419f
C4890 X1.X1.X1.X2.X2.X2.X2.vin1 a_2196_4198# 0.197f
C4891 X1.X1.X1.X1.X2.X2.X2.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 0.234f
C4892 d1 a_39966_7922# 3.41e-19
C4893 a_16836_17540# d0 0.518f
C4894 d2 X2.X1.X1.X2.X1.X2.vrefh 0.177f
C4895 a_54606_28888# a_54606_30794# 0.00198f
C4896 a_19722_29936# X1.X2.X1.X1.X1.X2.vout 0.254f
C4897 a_19036_24258# a_19336_22312# 6.1e-19
C4898 X2.X2.X1.X2.vrefh vdd 0.414f
C4899 X2.X2.X1.X1.X2.X2.X3.vin2 a_48616_18540# 0.00504f
C4900 a_40352_26982# X2.X1.X2.X2.X2.vrefh 1.64e-19
C4901 d4 X1.X1.X2.X3.vin1 0.0865f
C4902 a_16836_4198# a_17222_4198# 0.419f
C4903 a_48702_20446# a_49002_18540# 4.41e-20
C4904 d1 a_31476_6104# 2.25e-20
C4905 a_11072_21264# a_11072_19358# 0.00396f
C4906 a_23512_5016# a_25326_4110# 1.06e-19
C4907 a_4396_12822# d1 0.521f
C4908 X1.X2.X1.X1.X2.X2.vout a_19336_18540# 7.93e-20
C4909 a_4696_29936# X1.X1.X1.X1.X1.X1.X3.vin2 0.00546f
C4910 a_25326_25076# d1 0.00151f
C4911 X1.X2.X2.vrefh a_17222_4198# 0.301f
C4912 a_4696_29936# vdd 1.05f
C4913 a_46502_27070# d1 0.00151f
C4914 d2 X1.X1.X1.X2.X2.vrefh 0.158f
C4915 X1.X1.X2.X2.X1.X2.vout a_8186_22210# 0.254f
C4916 d2 a_17222_15634# 0.0059f
C4917 a_52406_24076# X2.X2.X2.X2.X1.X2.vout 0.418f
C4918 X2.X1.X1.X1.X2.X1.X1.vin2 d2 0.231f
C4919 X1.X1.X1.X2.X2.X1.X1.vin1 X1.X1.X1.X2.X2.X1.X1.vin2 0.668f
C4920 d3 X1.X1.X1.X2.X3.vin2 0.156f
C4921 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X3.vin2 0.418f
C4922 X2.X2.X2.X1.X2.vrefh a_54992_9828# 0.118f
C4923 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 5.19e-19
C4924 X1.X2.X2.X2.X1.X1.vout X1.X2.X2.X2.X1.X1.X3.vin1 0.118f
C4925 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 5.19e-19
C4926 X1.X1.X2.X1.X1.X1.X2.vin1 d0 0.262f
C4927 d3 a_49002_22312# 9.23e-19
C4928 a_8486_16452# a_8872_16452# 0.419f
C4929 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.vout 0.118f
C4930 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X1.X3.vin2 0.0943f
C4931 d2 X1.X2.X2.X1.X1.X1.X3.vin2 0.0682f
C4932 X2.X1.X2.X2.X2.X1.X1.vin2 a_39966_26982# 0.273f
C4933 a_19336_26164# a_17222_25164# 5.36e-21
C4934 a_25326_32700# a_23512_31700# 1.15e-20
C4935 X2.X1.X1.X3.vin2 X2.X1.X3.vin2 3.82e-19
C4936 a_37466_18358# X2.X1.X2.X3.vin1 0.374f
C4937 a_48316_9010# a_49002_7064# 2.86e-19
C4938 X1.X2.X1.X1.X2.X1.X3.vin1 d2 0.104f
C4939 a_48702_9010# a_48616_7064# 3.14e-19
C4940 X2.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X3.vin1 0.0174f
C4941 a_52106_10734# a_52492_10734# 0.414f
C4942 a_25326_17452# a_23126_16452# 4.77e-21
C4943 X1.X1.X2.X2.X1.X1.X3.vin1 d4 0.0194f
C4944 d3 X2.X1.X2.X2.X3.vin2 0.417f
C4945 a_31862_27070# X2.X1.X1.X1.X1.X2.X3.vin1 0.00207f
C4946 a_48702_9010# vdd 0.561f
C4947 a_17222_17540# a_17222_15634# 0.00198f
C4948 X1.X1.X2.X1.X2.X1.vout a_8872_12640# 0.359f
C4949 X2.X2.X1.X1.X1.X1.X2.vin1 a_46502_32788# 8.88e-20
C4950 d2 X1.X1.X1.X2.X2.X1.X1.vin2 0.231f
C4951 X2.X2.X1.X2.X1.X2.X1.vin2 a_46116_11822# 1.78e-19
C4952 d3 a_48316_12822# 0.00108f
C4953 a_25712_30794# X1.X2.X2.X2.X2.X2.vrefh 1.64e-19
C4954 a_2582_27070# d3 1.89e-19
C4955 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X1.X3.vin2 0.161f
C4956 X1.X1.X2.vrefh a_6032_892# 7.3e-19
C4957 a_49002_29936# X2.X2.X1.X1.X1.X1.X3.vin2 0.00815f
C4958 X1.X2.X2.X2.X2.X1.X2.vin1 X2.X1.X1.X1.X1.X2.X1.vin2 0.00232f
C4959 a_31476_32788# vdd 1.05f
C4960 a_31476_28976# a_31862_28976# 0.419f
C4961 a_22826_25982# a_23212_25982# 0.414f
C4962 X2.X2.X2.X1.X2.X1.X3.vin2 a_52792_12640# 0.1f
C4963 d2 X2.X1.X1.X1.X1.X2.vrefh 6.65e-20
C4964 X2.X1.X2.X2.X3.vin1 d2 0.0014f
C4965 a_25326_32700# d0 0.0489f
C4966 a_19722_10916# d1 0.0316f
C4967 a_2196_21352# d1 2.25e-20
C4968 X1.X2.X2.X2.X2.X1.X1.vin2 d1 4.01e-19
C4969 X1.X1.X2.X2.X1.X1.X2.vin1 a_11072_21264# 0.197f
C4970 X2.X1.X2.X1.X1.X2.vout vdd 0.696f
C4971 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X2.vin1 0.00117f
C4972 a_46502_25164# a_48702_24258# 4.2e-20
C4973 X2.X2.X2.X2.X2.vrefh vdd 0.426f
C4974 a_8486_24076# a_8872_24076# 0.419f
C4975 a_19422_24258# a_17222_23258# 4.77e-21
C4976 a_46502_13728# a_48702_12822# 4.2e-20
C4977 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X2.vin1 0.00117f
C4978 X2.X2.X2.X1.X1.X2.vrefh a_54606_6016# 0.3f
C4979 a_11072_21264# d2 0.00414f
C4980 X2.X1.X1.X2.X1.X1.X3.vin2 a_31476_15634# 0.354f
C4981 X2.X1.X2.X1.X1.X2.X2.vin1 vdd 0.576f
C4982 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin1 0.52f
C4983 d0 X2.X2.X2.X1.X2.X1.X3.vin2 4.34e-19
C4984 a_52492_6962# X2.X2.X2.X1.X1.X1.X3.vin2 0.00546f
C4985 a_37852_25982# X2.X1.X2.X2.X2.X1.vout 1.64e-19
C4986 a_25326_25076# a_23126_24076# 4.77e-21
C4987 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X3.vin2 0.17f
C4988 X2.X2.X1.X1.X1.X2.vout d1 0.033f
C4989 a_25326_26982# a_25712_26982# 0.419f
C4990 d3 a_48702_16634# 4.67e-19
C4991 a_11072_25076# d0 0.515f
C4992 X2.X2.X2.X2.vrefh a_54606_17452# 0.3f
C4993 d2 a_17222_30882# 4.64e-19
C4994 X1.X2.X2.X2.X2.X1.X3.vin1 a_23212_25982# 0.00251f
C4995 a_46116_19446# d1 2.92e-22
C4996 X1.X1.X2.X1.X3.vin2 d1 0.00807f
C4997 a_46116_32788# X2.X2.X1.X1.X1.X1.X1.vin1 0.195f
C4998 a_8186_25982# d4 3.58e-19
C4999 X1.X2.X1.X1.X1.X2.X1.vin2 X1.X2.X1.X1.X1.X1.X3.vin2 3.94e-19
C5000 X1.X1.X1.X1.X1.X2.X2.vin1 d0 0.262f
C5001 d2 a_34362_14688# 0.0191f
C5002 a_46502_21352# vdd 0.553f
C5003 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.vout 0.118f
C5004 a_25326_17452# a_25712_17452# 0.419f
C5005 a_34062_28070# X2.X1.X1.X1.X1.X2.vout 0.418f
C5006 d4 a_25326_17452# 1.89e-19
C5007 X1.X1.X1.X2.X1.X1.X1.vin2 d1 1.49e-19
C5008 d3 X2.X1.X2.X1.X2.X2.vout 8.47e-19
C5009 a_52106_14586# a_52406_12640# 4.19e-20
C5010 X1.X1.X1.X1.X1.X1.X1.vin2 vrefh 0.0964f
C5011 X3.vin1 a_20286_892# 5.17e-19
C5012 d3 a_34062_24258# 0.00195f
C5013 a_19336_18540# a_19036_16634# 6.2e-19
C5014 X1.X2.X1.X1.X2.X2.vrefh d1 0.0124f
C5015 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X3.vin1 0.00118f
C5016 a_48616_10916# vdd 1.05f
C5017 X1.X2.X1.X2.X2.X1.X3.vin2 a_19722_7064# 0.00815f
C5018 d3 a_4782_9010# 0.00148f
C5019 X1.X2.X1.X1.X1.X2.vout X1.X2.X1.X1.X1.X2.X3.vin1 0.326f
C5020 a_25712_13640# a_25712_11734# 0.00396f
C5021 d4 X2.X1.X2.X2.X2.X1.vout 4.78e-20
C5022 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X2.vrefh 2.33e-19
C5023 d3 a_46502_25164# 0.00112f
C5024 X2.X2.X2.X1.X2.X2.vout d1 0.033f
C5025 X1.X1.X1.X2.X1.X1.X1.vin1 d2 0.0116f
C5026 a_46116_17540# a_46116_15634# 0.00396f
C5027 a_33676_28070# vdd 1.05f
C5028 d2 a_39966_11734# 0.00328f
C5029 d1 X2.X2.X2.X1.X1.X2.vrefh 0.0738f
C5030 a_48702_24258# d1 0.0749f
C5031 X2.X1.X3.vin1 d5 0.0551f
C5032 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X2.X1.X1.X1.X2.X2.vin1 0.00232f
C5033 d5 a_5646_892# 0.508f
C5034 X2.X2.X1.X1.X2.X2.X3.vin2 d4 0.0265f
C5035 X2.X1.X3.vin1 X2.X1.X2.X1.X3.vin1 0.00304f
C5036 a_2582_23258# d1 0.00148f
C5037 a_8186_18358# a_8872_16452# 3.08e-19
C5038 X2.X2.X2.X2.X2.X1.X1.vin1 d3 6.34e-20
C5039 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X1.vin2 3.94e-19
C5040 X2.X1.X1.X1.X2.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin1 0.267f
C5041 a_2582_8010# a_4696_7064# 2.95e-20
C5042 a_2582_6104# d1 3.41e-19
C5043 a_52492_25982# a_54606_25076# 4.72e-20
C5044 a_25326_25076# a_25712_25076# 0.419f
C5045 d0 X2.X1.X2.X1.X1.X1.X1.vin1 0.269f
C5046 a_25326_6016# X1.X2.X2.X1.X1.X1.X2.vin1 0.402f
C5047 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X3.vin1 0.00118f
C5048 d3 a_48702_31882# 3.23e-19
C5049 X1.X2.X1.X1.X2.X2.X1.vin2 a_16836_19446# 1.78e-19
C5050 X2.X1.X2.X2.X1.X2.vout d1 0.033f
C5051 d2 X2.X1.X2.X1.X2.X2.X1.vin1 0.0106f
C5052 a_17222_25164# X1.X2.X1.X1.X2.X1.X1.vin1 0.417f
C5053 X1.X1.X2.X1.X2.X2.X1.vin1 X1.X2.X1.X2.X1.X2.vrefh 0.00437f
C5054 a_16836_25164# X1.X2.X1.X1.X2.X1.X3.vin1 0.354f
C5055 d3 a_17222_9916# 0.00112f
C5056 a_10686_17452# X1.X1.X2.X1.X2.X2.X3.vin2 0.567f
C5057 d4 a_34362_18540# 0.257f
C5058 X1.X1.X2.X1.X1.X2.vout d1 0.033f
C5059 X2.X1.X1.X1.X2.X2.X3.vin2 d4 0.0265f
C5060 X1.X1.X2.X3.vin2 X1.X1.X2.X3.vin1 0.559f
C5061 a_52406_12640# vdd 0.561f
C5062 X2.X2.X1.X1.X1.X2.X3.vin2 a_46502_27070# 0.567f
C5063 X2.X1.X1.X1.X1.X1.X3.vin1 a_34062_31882# 0.428f
C5064 a_8486_31700# a_8872_31700# 0.419f
C5065 a_22826_29834# vdd 0.477f
C5066 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.X1.X3.vin2 2.23e-19
C5067 a_54992_26982# X2.X2.X2.X2.X2.X1.X2.vin1 1.78e-19
C5068 a_33976_22312# a_34062_20446# 3.38e-19
C5069 a_34362_22312# a_33676_20446# 3.31e-19
C5070 X1.X2.X1.X2.X1.X2.vrefh a_17222_13728# 8.22e-20
C5071 d3 d1 0.373f
C5072 d0 a_31476_11822# 0.515f
C5073 d3 X2.X1.X2.X2.X2.X2.vout 0.222f
C5074 d2 a_8486_8828# 0.00138f
C5075 a_4782_28070# X1.X1.X1.X1.X1.X2.X3.vin2 0.277f
C5076 X2.X1.X2.X2.X1.X2.vrefh vdd 0.414f
C5077 a_8186_10734# a_8486_8828# 4.41e-20
C5078 a_16836_32788# d1 2.25e-20
C5079 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin2 7.84e-19
C5080 X1.X2.X2.X1.X1.X1.vout vdd 0.78f
C5081 d2 a_31862_8010# 0.00665f
C5082 X1.X2.X2.X2.X1.X2.X1.vin1 d2 0.0114f
C5083 a_39966_32700# d4 8.99e-20
C5084 X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.vout 3.38e-19
C5085 a_25712_32700# d2 3.9e-19
C5086 X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X1.X1.vin1 0.267f
C5087 a_5082_29936# X1.X1.X1.X1.X3.vin1 0.434f
C5088 d3 X2.X2.X1.X1.X1.X1.X3.vin1 0.0103f
C5089 X2.X2.X2.X2.X2.X2.vout d1 0.033f
C5090 X1.X2.X1.X1.X2.X2.X3.vin2 d4 0.0265f
C5091 X1.X2.X2.vrefh X1.X3.vin2 4.75e-20
C5092 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X2.X1.X1.X2.X2.vrefh 0.00437f
C5093 X1.X1.X3.vin2 a_5082_14688# 2.04e-19
C5094 X2.X2.X1.X2.X1.X2.X1.vin1 d1 0.0118f
C5095 d0 a_11072_4110# 0.518f
C5096 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X1.X3.vin1 0.0425f
C5097 a_40352_6016# a_40352_4110# 0.00396f
C5098 d0 a_31862_15634# 0.0489f
C5099 X2.X2.X2.X2.X2.X1.X3.vin2 d1 0.15f
C5100 X2.X1.X1.X1.X2.X2.vrefh d0 0.848f
C5101 d2 a_52406_31700# 0.00157f
C5102 a_52406_31700# a_54606_32700# 4.77e-21
C5103 a_19336_18540# vdd 1.05f
C5104 d1 a_14082_892# 2.34e-19
C5105 X2.X1.X1.X1.X1.X1.X3.vin2 a_31476_30882# 0.354f
C5106 X2.X1.X2.X3.vin2 d1 0.0129f
C5107 a_2582_25164# d2 0.00328f
C5108 d0 X1.X1.X1.X2.X2.X2.vrefh 0.844f
C5109 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 0.049f
C5110 a_23126_16452# a_22826_14586# 5.55e-20
C5111 a_5082_26164# X1.X1.X1.X1.X2.X1.X3.vin1 0.00837f
C5112 X2.X1.X2.X2.X2.X1.X3.vin2 X2.X1.X2.X2.X2.X2.X3.vin1 1.22e-19
C5113 X1.X1.X2.X1.X3.vin2 a_8486_12640# 0.00101f
C5114 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X1.X2.X1.vin2 0.076f
C5115 d2 X2.X1.X2.X2.X2.X2.X1.vin1 9.24e-20
C5116 a_38152_27888# X2.X1.X2.X2.X2.X1.X3.vin2 0.1f
C5117 a_8872_8828# a_8572_6962# 6.71e-19
C5118 a_54992_6016# vdd 1.05f
C5119 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X1.vin2 0.668f
C5120 X1.X1.X3.vin2 a_5646_892# 0.0927f
C5121 X1.X2.X3.vin1 X1.X2.X3.vin2 3.25f
C5122 X2.X2.X1.X1.X2.X1.X1.vin2 vdd 0.36f
C5123 X1.X2.X1.X3.vin2 X1.X2.X2.X3.vin1 1.22e-19
C5124 d0 X1.X1.X2.X1.X2.X1.X1.vin2 0.276f
C5125 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X3.vin1 0.00117f
C5126 a_17222_23258# d0 0.0489f
C5127 X2.X2.X2.X2.X1.X2.X3.vin2 a_52406_24076# 0.277f
C5128 d1 X1.X1.X2.vrefh 0.257f
C5129 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X1.X2.vout 0.075f
C5130 a_34062_28070# a_31862_28976# 4.2e-20
C5131 X2.X1.X1.X1.X1.X2.X2.vin1 X2.X1.X1.X1.X1.X2.X3.vin1 0.00117f
C5132 a_17222_17540# a_19422_16634# 4.2e-20
C5133 X2.X1.X2.X1.X1.X1.X3.vin2 vdd 0.937f
C5134 X1.X1.X1.X1.X1.X1.X1.vin2 a_2582_30882# 8.88e-20
C5135 d3 X2.X2.X3.vin2 0.77f
C5136 d3 X1.X1.X2.X2.X2.X1.vout 0.0421f
C5137 X2.X1.X1.X1.X2.X1.X3.vin1 vdd 0.997f
C5138 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X1.vin2 0.076f
C5139 d2 a_19422_9010# 7.51e-19
C5140 X2.X2.X2.X1.X1.X2.X1.vin1 a_54992_6016# 1.64e-19
C5141 d2 X2.X2.X2.X1.X2.X2.X3.vin2 0.113f
C5142 a_34362_22312# X2.X1.X1.X1.X2.X2.X3.vin1 0.00874f
C5143 d3 a_23126_24076# 0.00122f
C5144 X1.X1.X2.X2.X2.X2.X3.vin2 d0 4.34e-19
C5145 a_49002_29936# X2.X2.X1.X1.X1.X2.X3.vin1 0.00874f
C5146 d2 X2.X2.X2.X1.X2.X1.vout 0.00174f
C5147 X2.X1.X2.X1.X1.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin2 0.0128f
C5148 X2.X2.X2.X2.X1.X1.X3.vin2 X2.X2.X2.X2.X1.X1.X3.vin1 0.581f
C5149 a_8186_25982# X1.X1.X2.X3.vin2 0.452f
C5150 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X1.X2.X2.X1.X2.vrefh 0.1f
C5151 a_19422_28070# d1 0.0749f
C5152 X1.X2.X2.X2.X1.X1.vout d1 0.0238f
C5153 d0 a_42976_892# 2.73e-19
C5154 X2.X2.X2.X2.X1.X1.X1.vin1 a_54992_17452# 1.64e-19
C5155 a_16836_27070# d2 0.00533f
C5156 a_8186_29834# a_8872_27888# 2.86e-19
C5157 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X2.X1.X2.X2.vrefh 0.0128f
C5158 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.X3.vin2 1.22e-19
C5159 d0 a_39966_13640# 0.0489f
C5160 X1.X2.X1.X2.X2.X1.X1.vin2 vdd 0.36f
C5161 d2 X2.X2.vrefh 0.0108f
C5162 a_16836_6104# X1.X2.X1.X2.X2.X2.X1.vin2 0.12f
C5163 X1.X2.X1.X2.X2.X2.X1.vin2 X1.X2.X1.X2.X2.X2.X2.vin1 0.242f
C5164 a_33676_16634# X2.X1.X1.X2.X1.X1.X3.vin2 0.1f
C5165 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X3.vin1 0.00789f
C5166 d3 X2.X2.X2.X1.X1.X2.vout 6.06e-19
C5167 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 0.0903f
C5168 a_31862_30882# d0 0.0489f
C5169 a_31862_32788# X2.X1.X1.X1.X1.X1.X1.vin1 0.42f
C5170 a_31476_32788# X2.X1.X1.X1.X1.X1.X3.vin1 0.354f
C5171 X1.X1.X1.X2.X2.X1.X3.vin1 vdd 0.997f
C5172 d2 a_19422_31882# 9.83e-19
C5173 a_10686_25076# X1.X1.X2.X2.X1.X2.X1.vin2 8.88e-20
C5174 a_46502_28976# d0 0.0675f
C5175 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X3.vin2 0.552f
C5176 X1.X2.X1.X1.X3.vin1 d1 0.00179f
C5177 d3 a_5082_18540# 0.0469f
C5178 a_11072_26982# a_11072_28888# 0.00396f
C5179 a_25712_21264# vdd 1.05f
C5180 d2 a_49002_7064# 0.254f
C5181 X2.X2.X1.X3.vin2 a_49002_10916# 0.452f
C5182 X1.X1.X1.X2.X3.vin1 a_5082_10916# 0.372f
C5183 a_25326_32700# X2.vrefh 0.3f
C5184 X1.X2.X2.X2.X2.X2.X2.vin1 a_25712_32700# 0.197f
C5185 X1.X1.X2.X2.X2.X2.X1.vin1 X1.X2.X1.X1.X1.X2.vrefh 0.00437f
C5186 a_19722_22312# X1.X2.X1.X1.X2.X2.vout 0.263f
C5187 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X2.vin1 0.564f
C5188 X2.X1.X2.X1.X2.X1.X3.vin1 d1 0.151f
C5189 a_46116_4198# vdd 1.05f
C5190 X1.X1.X2.X2.X1.X1.X3.vin2 vdd 0.905f
C5191 X2.X2.X1.X1.X2.X2.vout X2.X2.X1.X1.X2.X2.X3.vin2 0.08f
C5192 a_39966_19358# X2.X1.X2.X1.X2.X2.X3.vin2 8.07e-19
C5193 a_5646_892# a_6032_892# 0.419f
C5194 a_8572_25982# vdd 1.05f
C5195 d3 a_8486_12640# 0.00195f
C5196 X2.X2.X2.vrefh vdd 0.702f
C5197 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.X1.vin2 0.216f
C5198 X1.X2.X2.X1.X2.X2.X3.vin1 a_25326_15546# 0.52f
C5199 X2.X2.X2.X2.X2.X2.X2.vin1 vdd 0.578f
C5200 a_17222_32788# X1.X2.X1.X1.X1.X1.X3.vin1 0.52f
C5201 a_23512_24076# d2 6.04e-19
C5202 d0 X2.X1.X1.X2.X1.X1.X1.vin1 0.267f
C5203 X1.X1.X2.X1.X3.vin1 vdd 0.805f
C5204 a_52106_22210# vdd 0.477f
C5205 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X3.vin2 0.161f
C5206 X1.X2.X1.X2.X1.X1.X2.vin1 a_16836_15634# 0.197f
C5207 d2 X2.X1.X1.X2.X1.X2.X3.vin2 0.121f
C5208 X1.X2.X2.X1.X2.X2.vout a_23512_16452# 0.36f
C5209 a_39966_11734# X2.X1.X2.X1.X2.vrefh 8.22e-20
C5210 d4 X2.X2.X2.X3.vin1 0.0865f
C5211 a_46116_17540# X2.X2.X1.X2.X1.X1.X2.vin1 1.78e-19
C5212 d2 a_54992_7922# 0.00351f
C5213 d3 X1.X1.X2.X2.X1.X2.X3.vin2 0.0247f
C5214 d3 X1.X1.X1.X1.X2.vrefh 6.65e-20
C5215 X2.X1.X1.X2.X2.X1.X1.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 2.23e-19
C5216 X2.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.vout 0.399f
C5217 a_48616_29936# vdd 1.05f
C5218 X2.X2.X1.X1.X1.X2.X3.vin2 d3 0.103f
C5219 X1.X2.X2.X2.X1.X2.X3.vin1 a_22826_22210# 0.00874f
C5220 X2.X2.X1.X1.X2.X2.X2.vin1 X2.X2.X1.X2.vrefh 0.564f
C5221 a_52492_6962# a_52792_5016# 6.1e-19
C5222 d0 X2.X1.X1.X2.X2.X2.X3.vin2 4.34e-19
C5223 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X2.vrefh 0.00118f
C5224 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X2.vin1 0.242f
C5225 d3 a_52492_10734# 0.621f
C5226 X2.X2.X2.X2.X2.X1.X1.vin2 a_54992_28888# 1.78e-19
C5227 d0 a_54992_15546# 0.518f
C5228 a_2196_17540# a_2582_17540# 0.419f
C5229 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X2.vin1 0.564f
C5230 a_19336_18540# X1.X2.X1.X2.X1.X1.X3.vin1 0.00232f
C5231 X1.X2.X1.X2.X2.X2.vrefh a_17222_8010# 0.3f
C5232 a_23512_8828# a_25326_7922# 1.06e-19
C5233 X2.X2.X2.X2.X1.X1.X3.vin2 a_54992_21264# 0.354f
C5234 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X1.vout 0.033f
C5235 a_16836_4198# vdd 1.05f
C5236 a_19336_7064# X1.X2.X1.X2.X2.X2.vout 0.0929f
C5237 d4 a_37766_16452# 8.66e-19
C5238 a_52492_18358# a_52406_16452# 3.3e-19
C5239 X1.X2.X2.X2.X1.X2.vout a_23512_24076# 0.36f
C5240 X1.X2.X2.vrefh vdd 0.707f
C5241 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X3.vin1 0.206f
C5242 X1.X2.X2.vrefh a_28096_892# 4.63e-19
C5243 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.vout 0.075f
C5244 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.X2.vin1 0.00117f
C5245 X1.X1.X1.X1.X1.X1.X1.vin1 d1 1.51e-19
C5246 a_37466_18358# vdd 0.476f
C5247 X2.X2.X1.X2.X1.X1.X3.vin2 vdd 0.905f
C5248 a_25712_11734# X1.X2.X2.X1.X2.vrefh 1.64e-19
C5249 X2.X1.X2.X2.X1.X2.X1.vin1 d0 0.267f
C5250 X1.X1.X1.X1.X2.X1.vout X1.X1.X1.X1.X2.X2.vout 0.514f
C5251 d2 a_34062_9010# 7.51e-19
C5252 d3 a_4696_26164# 0.621f
C5253 a_23212_10734# a_25326_9828# 4.72e-20
C5254 a_31476_13728# d1 2.25e-20
C5255 X1.X1.X1.X1.X2.X2.vrefh vdd 0.415f
C5256 a_2196_15634# a_2196_13728# 0.00396f
C5257 a_34362_18540# X2.X1.X1.X3.vin2 0.233f
C5258 a_16836_27070# a_16836_25164# 0.00396f
C5259 X2.X2.X2.X1.X1.X1.vout vdd 0.78f
C5260 a_49002_10916# X2.X2.X1.X2.X3.vin2 0.263f
C5261 d2 a_40352_13640# 0.00464f
C5262 X1.X2.X1.X1.X2.vrefh a_17222_25164# 8.22e-20
C5263 a_23512_12640# vdd 1.05f
C5264 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X2.vrefh 0.00118f
C5265 a_39966_28888# d1 0.00148f
C5266 X1.X2.X2.X1.X2.X1.X1.vin2 X1.X2.X2.X1.X2.X1.X1.vin1 0.668f
C5267 X2.X1.X1.X1.X2.X1.X3.vin2 vdd 0.903f
C5268 X2.X1.X2.X1.X1.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X3.vin1 0.581f
C5269 a_40352_26982# d2 0.00272f
C5270 d2 X2.X2.X1.X1.X1.X2.X1.vin2 0.226f
C5271 X2.X1.X2.X1.X2.X2.X1.vin2 a_39966_15546# 0.273f
C5272 d2 X1.X2.X2.X1.X2.X1.X3.vin2 0.171f
C5273 X1.X2.X1.X2.X1.X1.vout X1.X2.X1.X2.X3.vin1 0.131f
C5274 X2.X2.X1.X2.X1.X2.X3.vin2 a_46502_9916# 8.07e-19
C5275 a_2582_6104# X1.X1.X1.X2.X2.X2.X1.vin2 0.273f
C5276 X1.X1.X1.X2.X2.X1.X3.vin2 vdd 0.903f
C5277 X2.X2.X2.X1.X3.vin2 d1 0.00807f
C5278 a_33676_31882# X2.X1.X1.X1.X1.X1.X3.vin2 0.1f
C5279 X2.X1.X2.X2.X2.X2.X1.vin1 X2.X1.X2.X2.X2.X2.X3.vin2 2.23e-19
C5280 a_52106_25982# d4 7.15e-19
C5281 X2.X2.X1.X2.X2.X1.X3.vin2 a_46502_8010# 0.567f
C5282 a_34062_28070# X2.X1.X1.X1.X1.X2.X3.vin2 0.277f
C5283 X1.X2.X2.X2.X2.X2.X3.vin2 vdd 0.738f
C5284 a_54992_30794# d0 0.518f
C5285 d2 X2.X1.X1.X1.X1.X2.X3.vin1 0.158f
C5286 X1.X1.X2.X2.X3.vin1 d1 0.00179f
C5287 a_4696_22312# a_4396_20446# 6.71e-19
C5288 d2 a_34362_10916# 7.13e-19
C5289 X1.X2.X2.X2.X2.X1.X3.vin2 a_25326_30794# 8.07e-19
C5290 X1.X2.X2.X1.X2.X2.X2.vin1 d1 1.03e-19
C5291 d2 a_8872_5016# 0.00251f
C5292 a_25326_6016# vdd 0.541f
C5293 X1.X2.X1.X1.X2.X2.X3.vin1 d4 2.08e-19
C5294 a_46502_8010# a_46502_6104# 0.00198f
C5295 a_54606_21264# a_52792_20264# 1.15e-20
C5296 a_17222_25164# vdd 0.553f
C5297 a_46116_8010# X2.X2.X1.X2.X2.X2.X1.vin1 1.64e-19
C5298 X1.X1.X3.vin1 X1.X1.X2.X3.vin1 3.45e-19
C5299 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X1.X2.X2.X2.X2.vrefh 0.00437f
C5300 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X1.vin2 8.93e-19
C5301 X2.X1.X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X1.vin2 8.93e-19
C5302 X1.X1.X1.X1.X2.X2.X2.vin1 d0 0.262f
C5303 X2.X1.X2.X2.X1.X2.X2.vin1 a_39966_23170# 8.88e-20
C5304 d2 a_39966_17452# 0.00583f
C5305 X2.X1.X2.X1.X2.X1.X2.vin1 a_39966_11734# 8.88e-20
C5306 d3 X1.X2.X2.X3.vin1 0.676f
C5307 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.vout 0.08f
C5308 X2.X2.X1.X1.X1.X1.X3.vin2 vdd 0.939f
C5309 a_37466_14586# a_37852_14586# 0.419f
C5310 a_4782_28070# vdd 0.47f
C5311 a_46502_21352# X2.X2.X1.X1.X2.X2.X2.vin1 8.88e-20
C5312 a_2582_28976# X1.X1.X1.X1.X1.X2.X1.vin2 0.273f
C5313 X1.X2.X2.X2.X2.X2.X3.vin1 a_25326_30794# 0.52f
C5314 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X1.X3.vin2 0.0523f
C5315 a_46502_19446# a_46502_17540# 0.00198f
C5316 a_23126_27888# a_25326_26982# 4.2e-20
C5317 a_5082_14688# d1 0.0422f
C5318 a_46116_19446# X2.X2.X1.X2.X1.X1.X1.vin1 1.64e-19
C5319 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X1.X1.vin2 0.216f
C5320 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X2.X1.X3.vin1 0.0131f
C5321 X1.X1.X2.X1.X2.X1.X1.vin1 a_11072_11734# 0.195f
C5322 X2.X1.X2.X2.X2.X2.X3.vin2 X2.X2.vrefh 0.183f
C5323 X1.X2.X2.X2.X2.X2.vout a_23512_31700# 0.36f
C5324 X1.X2.X1.X1.X1.X1.X2.vin1 a_16836_30882# 0.197f
C5325 X1.X2.X2.X2.X1.X2.X1.vin2 a_25326_23170# 0.273f
C5326 a_52492_18358# X2.X2.X2.X1.X2.X2.X3.vin2 0.00517f
C5327 X2.X2.X1.X1.X3.vin1 X2.X2.X2.X2.X3.vin2 0.0604f
C5328 a_39966_15546# X2.X1.X2.X1.X2.X1.X3.vin2 8.07e-19
C5329 a_46502_9916# X2.X2.X1.X2.X2.X1.X2.vin1 8.88e-20
C5330 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X3.vin2 0.161f
C5331 a_25712_28888# d0 0.515f
C5332 d0 X1.X1.X1.X2.X1.X2.X1.vin1 0.267f
C5333 X2.X2.X3.vin2 X2.X2.X2.X1.X3.vin2 0.039f
C5334 a_39966_21264# X2.X1.X2.X2.X1.X1.X3.vin1 0.00207f
C5335 a_4396_12822# a_2582_11822# 1.15e-20
C5336 d2 a_8572_29834# 0.627f
C5337 X1.X2.X2.X1.X2.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin1 0.00437f
C5338 X1.X1.X2.X2.X2.X1.X3.vin2 d0 4.34e-19
C5339 a_48316_12822# a_46502_11822# 1.15e-20
C5340 d2 X2.X1.X2.X1.X2.X2.vrefh 0.168f
C5341 X1.X2.X1.X1.X2.X1.X1.vin2 a_16836_23258# 1.78e-19
C5342 X2.X1.X3.vin1 d1 0.0876f
C5343 X2.X1.X1.X1.X3.vin2 a_34062_20446# 9.7e-20
C5344 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.X3.vin1 1.22e-19
C5345 X2.X2.X2.X2.X1.X2.vout a_52106_22210# 0.254f
C5346 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X1.vout 0.13f
C5347 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.vrefh 0.161f
C5348 d1 a_2196_4198# 2.92e-22
C5349 X1.X1.X2.X2.X1.X1.X3.vin1 a_10686_19358# 0.52f
C5350 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X2.vin1 0.564f
C5351 X1.X2.X2.X1.X1.X2.X1.vin1 X2.X1.X1.X2.X2.X2.vrefh 0.00437f
C5352 X2.X1.X2.X1.X1.X2.X2.vin1 a_40352_9828# 0.197f
C5353 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X1.X3.vin2 0.0943f
C5354 a_23212_14586# vdd 1.05f
C5355 X1.X1.X2.X1.X1.X1.X3.vin2 a_8872_5016# 0.1f
C5356 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X2.vrefh 0.076f
C5357 X1.X2.X1.X2.X1.X2.X1.vin1 X1.X2.X1.X2.X1.X2.X2.vin1 0.0689f
C5358 a_17222_13728# a_19036_12822# 1.06e-19
C5359 X2.X1.X2.X2.X2.X2.X2.vin1 d1 7.58e-19
C5360 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin1 0.52f
C5361 a_34362_26164# a_34062_24258# 5.25e-20
C5362 a_19722_22312# vdd 0.567f
C5363 a_33976_26164# X2.X1.X1.X1.X2.X1.vout 1.64e-19
C5364 X1.X1.X2.X2.X2.X1.X1.vin1 d0 0.267f
C5365 a_33976_14688# a_33676_12822# 6.71e-19
C5366 a_33976_7064# a_34062_5198# 3.38e-19
C5367 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.X2.vin1 0.00117f
C5368 a_34362_7064# a_33676_5198# 3.31e-19
C5369 a_2582_6104# a_4782_5198# 4.2e-20
C5370 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X1.X2.X1.vin2 0.216f
C5371 a_46502_19446# a_48616_18540# 4.72e-20
C5372 X2.X2.X1.X2.vrefh d0 0.848f
C5373 a_25712_9828# a_25712_7922# 0.00396f
C5374 a_52792_20264# a_52106_18358# 2.97e-19
C5375 a_39966_17452# a_38152_16452# 1.15e-20
C5376 X2.X2.X2.X1.X1.X1.X3.vin2 X2.X2.X2.X1.X1.X1.X1.vin1 2.23e-19
C5377 X2.X2.X2.X1.X1.X1.X2.vin1 a_54992_4110# 1.78e-19
C5378 a_25326_19358# a_25326_17452# 0.00198f
C5379 X1.X1.X2.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X3.vin1 0.581f
C5380 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X2.vrefh 0.00118f
C5381 a_8186_29834# X1.X1.X2.X2.X2.X2.vout 0.263f
C5382 a_2196_17540# vdd 1.05f
C5383 a_52792_27888# a_52492_25982# 6.2e-19
C5384 a_46502_27070# a_48616_26164# 4.72e-20
C5385 X2.X2.X1.X2.X2.X1.X3.vin1 d1 0.151f
C5386 X2.X2.X2.X1.X2.X2.X3.vin1 a_54992_15546# 0.354f
C5387 a_46116_27070# a_46116_28976# 0.00396f
C5388 d3 a_22826_25982# 0.29f
C5389 X2.X1.X1.X2.X1.X2.X3.vin2 a_31862_11822# 0.567f
C5390 X2.X1.X1.X2.X1.X1.vout a_34362_14688# 0.387f
C5391 a_34062_16634# X2.X1.X1.X2.X3.vin1 1.52e-19
C5392 d3 a_22826_10734# 0.284f
C5393 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin2 0.12f
C5394 a_54992_30794# a_54992_32700# 0.00396f
C5395 a_52406_27888# a_54606_28888# 4.77e-21
C5396 X2.X1.X2.X2.X2.X2.X1.vin2 a_39966_30794# 0.273f
C5397 a_48316_16634# a_46502_15634# 1.15e-20
C5398 d5 a_49566_892# 0.505f
C5399 a_48702_24258# X2.X2.X1.X1.X2.X1.X3.vin2 0.267f
C5400 a_10686_21264# a_8486_20264# 4.77e-21
C5401 a_39966_21264# X2.X1.X2.X2.X1.X1.X3.vin2 0.567f
C5402 X2.X2.X2.X2.X1.X1.X3.vin2 d1 0.15f
C5403 d2 X2.X1.X2.X2.X2.X2.vrefh 0.168f
C5404 d3 X2.X2.X2.X2.X2.X1.vout 0.0015f
C5405 d2 a_2196_27070# 0.00533f
C5406 X2.X1.X2.X1.X2.X2.X1.vin2 vdd 0.36f
C5407 X1.X2.X2.X2.X2.X1.X3.vin1 d3 0.0195f
C5408 d1 a_23512_8828# 0.521f
C5409 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 0.581f
C5410 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X2.X3.vin2 0.0565f
C5411 X1.X3.vin1 d6 0.0237f
C5412 d3 a_19336_14688# 7.7e-20
C5413 X1.X1.X1.X3.vin2 vdd 0.716f
C5414 a_34362_26164# d1 0.0318f
C5415 a_39966_6016# a_38152_5016# 1.15e-20
C5416 a_31476_28976# X2.X1.X1.X1.X1.X2.vrefh 1.64e-19
C5417 X2.X2.X2.X1.X3.vin2 a_52492_10734# 0.0927f
C5418 X2.X2.X2.X2.X2.X1.vout X2.X2.X2.X2.X2.X2.vout 0.514f
C5419 X1.X1.X2.X2.X1.X1.vout a_8872_20264# 0.359f
C5420 a_31476_32788# d0 0.511f
C5421 X2.X1.X1.X2.X1.X2.vout X2.X1.X1.X2.X1.X2.X3.vin1 0.326f
C5422 X1.X1.X2.X1.X2.X1.X1.vin1 vdd 0.592f
C5423 a_54606_17452# X2.X2.X2.X1.X2.X2.X2.vin1 0.402f
C5424 X1.X2.X2.X2.X1.X2.X1.vin2 vdd 0.361f
C5425 a_31862_6104# X2.X1.X1.X2.X2.X2.X2.vin1 8.88e-20
C5426 a_37852_22210# X2.X1.X2.X2.X1.X1.X3.vin2 0.00546f
C5427 X2.X1.X2.X2.X2.X2.X1.vin2 a_40352_32700# 1.78e-19
C5428 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X1.vin1 0.206f
C5429 a_19722_18540# X1.X2.X3.vin1 0.47f
C5430 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X1.vin1 0.0689f
C5431 X2.X2.X2.X2.X1.X1.X3.vin2 a_54606_19358# 7.84e-19
C5432 d2 a_10686_13640# 0.00665f
C5433 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X1.vin2 0.1f
C5434 X2.X2.X2.X2.X2.vrefh d0 0.844f
C5435 X2.X2.X2.X1.X2.X2.vrefh a_54992_13640# 0.118f
C5436 X2.X2.X2.X2.X2.X1.vout X2.X2.X2.X2.X2.X1.X3.vin2 0.326f
C5437 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X2.X1.X3.vin2 8.93e-19
C5438 a_48616_26164# X2.X2.X1.X1.X1.X2.vout 7.93e-20
C5439 X1.X1.X1.X1.X1.X2.X1.vin1 d1 0.0118f
C5440 a_25326_26982# X1.X2.X2.X2.X2.X1.X2.vin1 8.88e-20
C5441 X2.X1.X1.X1.X2.X1.X2.vin1 a_31862_23258# 0.402f
C5442 d3 a_49002_18540# 0.0469f
C5443 d0 X2.X1.X2.X1.X1.X2.X2.vin1 0.262f
C5444 d3 X2.X2.X1.X1.X2.X1.X3.vin2 2.81e-19
C5445 X1.X1.X2.X1.X2.X2.X2.vin1 a_10686_15546# 8.88e-20
C5446 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.X1.vin2 8.93e-19
C5447 d2 a_17222_28976# 0.00479f
C5448 X1.X2.X2.X1.X2.X1.vout d1 0.0238f
C5449 a_46502_11822# d1 0.00151f
C5450 a_54992_13640# vdd 1.05f
C5451 a_48316_9010# X2.X2.X1.X2.X2.X1.X3.vin2 0.1f
C5452 X1.X2.X1.X2.X1.X1.X2.vin1 vdd 0.576f
C5453 a_2582_32788# a_4782_31882# 4.2e-20
C5454 X2.X3.vin2 vdd 0.665f
C5455 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.vout 0.335f
C5456 X1.X2.X1.X1.X3.vin2 d4 0.00419f
C5457 X1.X2.X2.X2.X3.vin1 a_22826_22210# 0.436f
C5458 a_4696_10916# X1.X1.X1.X2.X3.vin2 0.0927f
C5459 X2.X2.X1.X2.X1.X2.vrefh a_46502_13728# 8.22e-20
C5460 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 0.0565f
C5461 a_52492_25982# vdd 1.05f
C5462 X2.X1.X2.X1.X2.X1.X3.vin2 vdd 0.903f
C5463 X2.X1.X2.X2.X1.X1.vout d2 0.00169f
C5464 a_4782_16634# a_4696_14688# 3.14e-19
C5465 a_4396_16634# a_5082_14688# 2.86e-19
C5466 a_46502_21352# d0 0.0675f
C5467 d4 a_46116_32788# 1.8e-19
C5468 a_54606_25076# X2.X2.X2.X2.X1.X2.X2.vin1 0.402f
C5469 X2.X1.X2.X2.X2.X2.X1.vin2 vdd 0.387f
C5470 a_54606_9828# a_52406_8828# 4.77e-21
C5471 X1.X2.X2.X1.X1.X2.vout a_23212_6962# 0.0929f
C5472 X2.X2.X1.X1.X1.X2.X3.vin1 vdd 0.96f
C5473 a_46116_15634# d1 2.92e-22
C5474 a_22826_14586# X1.X2.X2.X1.X3.vin2 0.423f
C5475 a_49002_26164# a_48316_24258# 2.97e-19
C5476 a_48616_26164# a_48702_24258# 3.21e-19
C5477 a_48616_14688# a_48702_12822# 3.38e-19
C5478 a_49002_14688# a_48316_12822# 3.31e-19
C5479 X2.X1.X2.X1.X1.X2.X3.vin1 a_39966_7922# 0.52f
C5480 a_46502_19446# d4 1.89e-19
C5481 d1 a_19336_7064# 0.00613f
C5482 d3 a_2582_11822# 1.89e-19
C5483 X1.X2.X1.X2.X2.X1.X2.vin1 vdd 0.576f
C5484 a_54606_17452# vdd 0.541f
C5485 a_48316_20446# d2 6.04e-19
C5486 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin2 0.12f
C5487 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.vout 0.118f
C5488 X1.X1.X2.X1.X1.X1.X3.vin1 vdd 1.03f
C5489 X2.X1.X2.X1.X1.X2.vout a_38152_8828# 0.36f
C5490 X2.X1.X1.X2.X2.X1.X2.vin1 a_31476_8010# 0.197f
C5491 d4 a_10686_17452# 1.89e-19
C5492 a_22826_29834# a_23512_31700# 3.31e-19
C5493 X1.X2.X2.X1.X2.X1.X1.vin2 d1 4.01e-19
C5494 a_52406_12640# a_52792_12640# 0.419f
C5495 a_19336_26164# a_19036_24258# 6.2e-19
C5496 X1.X2.X1.X1.X2.X1.vout d2 0.00174f
C5497 X2.X2.X2.X1.X2.vrefh vdd 0.426f
C5498 d3 a_10686_32700# 1.28e-19
C5499 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X3.vin1 0.00118f
C5500 a_48702_16634# a_49002_14688# 4.19e-20
C5501 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X3.vin2 0.418f
C5502 X2.X2.X1.X2.X1.X1.vout a_48616_14688# 0.169f
C5503 X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.vout 3.2e-19
C5504 X2.X2.X2.X2.X2.X2.X3.vin1 a_54992_30794# 0.354f
C5505 X1.X1.X2.vrefh a_10686_4110# 4.89e-19
C5506 a_23212_18358# d2 0.0113f
C5507 a_33676_20446# d2 6.04e-19
C5508 X2.X1.X2.X1.X2.X2.X3.vin1 d1 0.146f
C5509 X1.X2.X1.X3.vin1 a_19336_18540# 0.17f
C5510 a_54606_23170# a_54992_23170# 0.419f
C5511 a_48316_31882# a_46502_30882# 1.15e-20
C5512 X1.X2.X1.X1.X1.X1.X2.vin1 vdd 0.578f
C5513 X2.X1.X1.X1.X1.X2.vout vdd 0.696f
C5514 d3 a_48616_26164# 0.621f
C5515 a_8186_25982# a_8872_24076# 3.08e-19
C5516 a_22826_18358# X1.X2.X2.X1.X2.X2.X3.vin2 0.00846f
C5517 a_25712_15546# d1 2.25e-20
C5518 a_37852_6962# vdd 1.05f
C5519 a_25326_9828# X1.X2.X2.X1.X1.X2.X2.vin1 0.402f
C5520 a_54992_6016# X2.X2.X2.X1.X1.X1.X1.vin2 1.78e-19
C5521 d3 X1.X2.X2.X1.X1.X2.X3.vin1 2.1e-19
C5522 X1.X1.X2.X2.X3.vin2 a_8572_29834# 0.363f
C5523 X2.X1.X2.X2.X1.X2.vrefh d0 0.848f
C5524 X2.X1.X2.X1.X2.X1.X2.vin1 a_40352_13640# 0.197f
C5525 d2 X2.X1.X1.X2.X1.X1.X3.vin2 0.169f
C5526 a_10686_13640# a_8872_12640# 1.15e-20
C5527 d3 X1.X2.X2.X2.X2.X1.X3.vin2 7.71e-19
C5528 a_46116_30882# d1 2.92e-22
C5529 X2.X2.X2.X2.X1.X2.X3.vin2 a_52106_22210# 3.85e-19
C5530 a_19036_20446# d2 6.04e-19
C5531 a_31862_13728# X2.X1.X1.X2.X1.X2.X3.vin1 0.52f
C5532 a_4696_10916# a_4782_9010# 3.21e-19
C5533 a_22826_14586# a_23126_12640# 4.19e-20
C5534 X2.X1.X3.vin1 a_37466_6962# 6.45e-19
C5535 a_2582_13728# X1.X1.X1.X2.X1.X2.X2.vin1 8.88e-20
C5536 a_5082_10916# a_4396_9010# 2.97e-19
C5537 a_31862_9916# d1 3.95e-19
C5538 a_33676_12822# vdd 1.05f
C5539 a_4782_16634# a_2582_15634# 4.77e-21
C5540 a_54606_7922# vdd 0.553f
C5541 d3 a_37466_14586# 9.23e-19
C5542 d2 a_46116_9916# 0.00272f
C5543 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X2.X2.vrefh 0.076f
C5544 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X2.X1.vin2 0.668f
C5545 X2.X1.X1.X2.X1.X2.X2.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 0.234f
C5546 d3 X2.X2.X2.X1.X2.X1.X1.vin1 6.34e-20
C5547 X2.X2.X2.X2.X3.vin1 d1 0.00179f
C5548 a_17222_32788# d4 8.99e-20
C5549 a_33676_12822# a_34062_12822# 0.419f
C5550 X1.X1.X1.X1.X3.vin2 a_4782_20446# 9.7e-20
C5551 X1.X2.X2.X2.X1.X1.X2.vin1 X2.X1.X1.X1.X2.X2.X1.vin2 0.00232f
C5552 a_31476_21352# a_31862_21352# 0.419f
C5553 X1.X1.X2.X2.X2.X1.X3.vin2 a_8486_27888# 0.267f
C5554 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X1.X2.X2.X2.X1.X3.vin1 0.00117f
C5555 X2.X2.X2.X1.X1.X2.X1.vin2 a_54992_7922# 0.12f
C5556 a_54606_7922# X2.X2.X2.X1.X1.X2.X1.vin1 0.417f
C5557 a_39966_21264# d1 0.00148f
C5558 X2.X2.X1.X1.X2.X2.X1.vin2 d2 0.231f
C5559 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.X2.vin1 0.00117f
C5560 X2.X1.X2.X2.X2.X2.X3.vin1 d1 0.147f
C5561 a_25326_28888# X1.X2.X2.X2.X2.X2.vrefh 0.3f
C5562 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.vout 0.335f
C5563 d0 a_54992_6016# 0.515f
C5564 X2.X2.X2.X2.X3.vin2 a_52406_31700# 9.7e-20
C5565 X2.X2.X1.X1.X2.X1.X1.vin2 d0 0.276f
C5566 a_38152_27888# d1 0.521f
C5567 a_8572_22210# a_8486_20264# 3.14e-19
C5568 X1.X1.X1.X2.X2.X2.X1.vin2 a_2196_4198# 1.78e-19
C5569 X1.X1.X1.X2.X1.X2.vout a_4396_12822# 0.36f
C5570 X2.X1.X1.X1.X2.X2.X3.vin1 d2 0.153f
C5571 a_25712_30794# d1 2.25e-20
C5572 d0 X2.X1.X2.X1.X1.X1.X3.vin2 4.34e-19
C5573 X2.X1.X1.X1.X2.X2.vrefh X1.X2.X2.X2.X1.X2.vrefh 0.117f
C5574 X2.X1.X1.X1.X2.X1.X3.vin1 d0 4.36e-19
C5575 a_49002_14688# d1 0.0422f
C5576 a_4782_24258# a_2582_23258# 4.77e-21
C5577 a_39966_11734# X2.X1.X2.X1.X1.X2.X3.vin2 8.07e-19
C5578 a_10686_26982# X1.X1.X2.X2.X2.X1.X3.vin1 0.52f
C5579 a_19336_26164# a_19722_26164# 0.414f
C5580 a_4696_10916# d1 0.0126f
C5581 d2 X2.X1.X1.X1.X1.X1.X3.vin2 0.0661f
C5582 a_37766_27888# d2 0.00123f
C5583 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X3.vin1 0.00117f
C5584 X2.X2.X2.vrefh X2.X2.X2.X1.X1.X1.X1.vin2 0.096f
C5585 X1.X1.X2.X2.X2.X2.X3.vin2 a_8486_31700# 0.277f
C5586 a_11072_32700# vdd 1.05f
C5587 a_8486_5016# a_8872_5016# 0.419f
C5588 a_37852_22210# d1 0.00613f
C5589 X1.X1.X2.X1.X2.X2.vout a_8572_14586# 0.0929f
C5590 X2.X1.X1.X2.X2.X1.X2.vin1 vdd 0.576f
C5591 a_4782_20446# vdd 0.471f
C5592 d0 X1.X2.X1.X2.X2.X1.X1.vin2 0.276f
C5593 a_17222_25164# a_19422_24258# 4.2e-20
C5594 d2 a_52492_29834# 0.627f
C5595 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X2.vin1 0.00117f
C5596 a_37766_27888# a_37852_29834# 3.14e-19
C5597 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X2.vin1 0.564f
C5598 X2.X2.X2.X3.vin2 X2.X2.X2.X3.vin1 0.559f
C5599 a_33976_26164# X2.X1.X1.X1.X3.vin1 0.169f
C5600 a_52492_25982# X2.X2.X2.X2.X1.X2.vout 7.93e-20
C5601 d0 X1.X1.X1.X2.X2.X1.X3.vin1 4.36e-19
C5602 a_25326_13640# vdd 0.541f
C5603 a_39966_26982# vdd 0.553f
C5604 a_54606_23170# d1 3.41e-19
C5605 a_39966_21264# X2.X1.X2.X2.X1.X1.X1.vin2 8.88e-20
C5606 d3 a_4782_24258# 0.00195f
C5607 a_23212_29834# a_25326_28888# 2.95e-20
C5608 a_25712_21264# d0 0.515f
C5609 a_11072_6016# X1.X1.X2.X1.X1.X2.vrefh 0.118f
C5610 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.X1.X1.X3.vin1 1.22e-19
C5611 X1.X1.X1.X1.X2.X2.vout d2 0.00117f
C5612 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X2.vrefh 2.33e-19
C5613 X1.X2.X2.X3.vin2 vdd 0.716f
C5614 a_49002_29936# X2.X2.X1.X1.X3.vin1 0.434f
C5615 a_31862_28976# vdd 0.553f
C5616 d0 a_46116_4198# 0.515f
C5617 X1.X1.X2.X2.X1.X1.X3.vin2 d0 4.34e-19
C5618 X1.X2.X1.X1.X2.X1.X3.vin2 d1 0.15f
C5619 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin2 0.1f
C5620 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin2 0.1f
C5621 a_23212_10734# vdd 1.05f
C5622 d0 X2.X2.X2.vrefh 4.73f
C5623 d3 X2.X2.X2.X1.X1.X2.X2.vin1 8.68e-20
C5624 d0 X2.X2.X2.X2.X2.X2.X2.vin1 0.199f
C5625 X2.X2.X3.vin2 a_49002_14688# 2.04e-19
C5626 a_39966_9828# X2.X1.X2.X1.X1.X2.X1.vin2 8.88e-20
C5627 d3 X2.X1.X2.X1.X1.X2.X3.vin1 2.1e-19
C5628 X2.X2.X1.X2.X1.X1.X2.vin1 d1 1.03e-19
C5629 X1.X1.X2.X1.X1.X1.vout X1.X1.X2.X1.X1.X1.X3.vin1 0.118f
C5630 a_33676_12822# a_33976_10916# 6.48e-19
C5631 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X3.vin1 0.546f
C5632 a_8186_14586# X1.X1.X2.X1.X2.X1.vout 0.383f
C5633 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X1.X2.vout 0.075f
C5634 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X2.X1.X1.vin1 0.668f
C5635 X2.X2.X1.X1.X2.X1.vout X2.X2.X1.X1.X2.X2.vout 0.514f
C5636 X1.X1.X2.X2.X1.X2.vout d1 0.033f
C5637 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X1.vin1 5.19e-19
C5638 a_11072_32700# X1.X2.vrefh 0.118f
C5639 X1.X2.X1.X2.X1.X1.X1.vin1 vdd 0.592f
C5640 X2.X1.X2.X1.X2.X1.vout a_37766_12640# 0.422f
C5641 X1.X2.X2.X2.vrefh a_25326_17452# 0.3f
C5642 d1 X2.X2.X2.X1.X1.X2.X3.vin1 0.146f
C5643 a_19422_12822# d1 0.0749f
C5644 d2 a_16836_11822# 0.00533f
C5645 X2.X1.X1.X1.X2.X1.X2.vin1 d1 1.03e-19
C5646 a_4396_5198# a_2582_4198# 1.15e-20
C5647 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.X1.vin2 0.23f
C5648 a_4782_20446# X1.X1.X1.X1.X2.X2.X3.vin2 0.277f
C5649 d1 a_40352_7922# 2.25e-20
C5650 X2.X2.X2.X2.X2.X1.X3.vin2 a_54606_30794# 8.07e-19
C5651 a_37766_5016# vdd 0.562f
C5652 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X1.vin2 0.242f
C5653 a_4782_31882# a_2582_30882# 4.77e-21
C5654 a_10686_13640# a_10686_11734# 0.00198f
C5655 a_19422_24258# a_19722_22312# 4.19e-20
C5656 X1.X2.X1.X1.X2.X1.vout a_19336_22312# 0.169f
C5657 X1.X1.X1.X2.X2.X1.X2.vin1 d1 1.03e-19
C5658 d2 X2.X2.X1.X2.X2.X1.X3.vin2 0.175f
C5659 a_40352_25076# d1 2.92e-22
C5660 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.vout 0.038f
C5661 X1.X2.X2.X1.X1.X1.vout a_23212_6962# 0.169f
C5662 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X1.X2.X2.X2.X2.vrefh 0.00437f
C5663 d0 a_16836_4198# 0.515f
C5664 X1.X1.X1.X2.X1.X2.X3.vin2 d1 0.171f
C5665 d1 X2.X1.X1.X2.X2.X2.X1.vin1 0.0118f
C5666 X1.X2.X2.vrefh X1.X2.X2.X1.X1.X1.X1.vin2 0.096f
C5667 a_46116_6104# a_46116_4198# 0.00396f
C5668 X1.X2.X1.X2.X1.X1.X3.vin2 a_17222_13728# 8.07e-19
C5669 X1.X1.X1.X1.X1.X2.vout X1.X1.X1.X1.X1.X1.vout 0.507f
C5670 X1.X2.X2.X2.X1.X2.X3.vin2 d1 0.171f
C5671 d0 X1.X2.X2.vrefh 4.78f
C5672 a_52106_25982# X2.X2.X2.X3.vin2 0.452f
C5673 X2.X2.X2.X2.X2.X1.X1.vin2 d1 4.01e-19
C5674 d2 X1.X2.X2.X1.X2.X2.X1.vin2 0.231f
C5675 X2.X2.X1.X3.vin2 vdd 0.716f
C5676 d2 a_46502_6104# 6.36e-19
C5677 X1.X1.X1.X1.X3.vin1 vdd 0.805f
C5678 a_8186_6962# vdd 0.477f
C5679 d0 X2.X2.X1.X2.X1.X1.X3.vin2 4.34e-19
C5680 X2.X1.X2.X2.X1.X2.X2.vin1 d2 0.0329f
C5681 d1 a_49566_892# 4.67e-19
C5682 X2.X1.X2.X2.X2.X1.X1.vin2 a_40352_26982# 0.12f
C5683 a_19336_26164# X1.X2.X1.X1.X2.X1.X3.vin1 0.00251f
C5684 a_39966_26982# X2.X1.X2.X2.X2.X1.X1.vin1 0.417f
C5685 X2.X2.X1.X1.X1.X1.X2.vin1 d1 0.0144f
C5686 a_25326_13640# X1.X2.X2.X1.X2.X1.X2.vin1 0.402f
C5687 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X2.vrefh 0.076f
C5688 X1.X2.X2.X2.X2.X2.X3.vin2 a_23512_31700# 0.101f
C5689 X2.X2.X1.X2.X2.X1.vout a_49002_7064# 0.383f
C5690 X1.X1.X1.X1.X2.X2.vrefh d0 0.844f
C5691 a_11072_9828# d1 2.92e-22
C5692 X1.X2.X1.X2.X2.X1.X3.vin2 X1.X2.X1.X2.X2.X2.vrefh 0.161f
C5693 a_10686_6016# a_8572_6962# 2.95e-20
C5694 a_19336_22312# a_19036_20446# 6.71e-19
C5695 a_23512_16452# a_23212_14586# 6.71e-19
C5696 X1.X2.X2.X1.X2.X2.X3.vin2 a_23126_16452# 0.277f
C5697 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X3.vin1 0.00117f
C5698 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X3.vin1 0.00836f
C5699 X2.X1.X2.X2.X1.X2.X3.vin1 X2.X1.X2.X2.X1.X2.vrefh 2.33e-19
C5700 a_19722_10916# X1.X2.X1.X2.X2.X1.X3.vin1 0.00837f
C5701 d4 X1.X2.X1.X2.X1.X1.X3.vin2 4.77e-19
C5702 a_39966_28888# a_40352_28888# 0.419f
C5703 X1.X2.X3.vin1 X1.X3.vin2 0.12f
C5704 X2.X2.X1.X1.X1.X1.X2.vin1 X2.X2.X1.X1.X1.X1.X3.vin1 0.00117f
C5705 a_22826_10734# a_23512_8828# 3.08e-19
C5706 X2.X1.X1.X1.X2.X1.X3.vin2 d0 4.34e-19
C5707 X1.X1.X1.X1.X1.X1.X3.vin1 d4 0.00851f
C5708 a_48702_31882# a_46502_32788# 4.2e-20
C5709 X1.X1.X2.X2.X2.X1.X1.vin2 d3 3.99e-21
C5710 d3 X2.X2.X1.X2.X1.X2.X3.vin2 0.0247f
C5711 d2 X1.X1.X2.X1.X1.X2.X2.vin1 0.0329f
C5712 d3 X1.X1.X1.X2.X1.X2.vout 0.0232f
C5713 X2.X2.X1.X1.X2.X1.X1.vin2 a_46116_23258# 1.78e-19
C5714 a_31862_28976# X2.X1.X1.X1.X1.X2.X1.vin1 0.417f
C5715 a_31476_28976# X2.X1.X1.X1.X1.X2.X3.vin1 0.354f
C5716 a_2196_28976# X1.X1.X1.X1.X1.X2.X2.vin1 1.78e-19
C5717 X2.X1.X1.X1.X1.X1.X1.vin1 vdd 0.596f
C5718 d0 X1.X1.X1.X2.X2.X1.X3.vin2 4.34e-19
C5719 X1.X1.X1.X1.X2.X2.X1.vin1 d1 0.0118f
C5720 X1.X2.X2.X2.X2.X2.X3.vin2 d0 4.34e-19
C5721 X2.X2.X2.X1.X1.X2.vrefh X2.X2.X2.X1.X1.X1.X3.vin2 0.165f
C5722 X1.X2.X2.X2.X2.X1.X1.vin1 d1 0.0118f
C5723 d4 X1.X1.X2.X1.X2.X2.vout 6.95e-19
C5724 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X3.vin2 2.23e-19
C5725 X2.X2.X1.X2.X1.X2.X3.vin1 a_48702_12822# 0.42f
C5726 X2.X2.X1.X1.X2.X1.X3.vin1 a_48702_24258# 0.428f
C5727 a_25326_6016# X1.X2.X2.X1.X1.X1.X1.vin2 8.88e-20
C5728 a_17222_21352# d2 0.00393f
C5729 a_46502_32788# d1 2.7e-19
C5730 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X2.vout 0.326f
C5731 d0 a_25326_6016# 0.0489f
C5732 a_54606_32700# vrefl 0.3f
C5733 X2.X2.X2.X2.X2.X2.X2.vin1 a_54992_32700# 0.197f
C5734 a_17222_25164# d0 0.0675f
C5735 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X3.vin1 0.00117f
C5736 X2.X2.X3.vin2 a_49566_892# 0.0912f
C5737 a_23126_20264# a_22826_18358# 5.25e-20
C5738 a_54992_9828# a_54992_7922# 0.00396f
C5739 X1.X2.X2.X2.X1.X2.X3.vin2 a_23126_24076# 0.277f
C5740 d2 X1.X2.X2.X2.X2.X2.X1.vin2 7.2e-20
C5741 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X3.vin2 0.161f
C5742 X2.X2.X1.X2.X2.X2.X2.vin1 a_46116_4198# 0.197f
C5743 X2.X2.X1.X1.X1.X1.X3.vin2 d0 4.34e-19
C5744 a_46502_32788# X2.X2.X1.X1.X1.X1.X3.vin1 0.52f
C5745 d2 a_48316_5198# 0.00393f
C5746 X1.X1.X2.X1.X1.X2.vrefh vdd 0.43f
C5747 X2.X2.X1.X3.vin1 a_48702_20446# 5.31e-19
C5748 X2.X2.X1.X2.X2.X2.X2.vin1 X2.X2.X2.vrefh 0.564f
C5749 a_8186_22210# d1 0.0422f
C5750 X1.X2.X2.X1.X2.X2.X3.vin2 a_25712_17452# 0.354f
C5751 X1.X2.X1.X3.vin1 a_19722_22312# 7.98e-19
C5752 X2.X2.X1.X2.X3.vin2 a_48616_7064# 0.363f
C5753 X2.X2.X1.X1.X2.X2.X3.vin1 vdd 0.962f
C5754 d4 X1.X2.X2.X1.X2.X2.X3.vin2 0.0264f
C5755 d6 a_42976_892# 0.506f
C5756 X1.X1.X2.X1.X2.X2.X2.vin1 d1 1.03e-19
C5757 X2.X2.X2.X1.X2.X1.vout X2.X2.X2.X1.X2.X1.X3.vin1 0.118f
C5758 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X3.vin1 0.206f
C5759 X3.vin1 d7 0.0163f
C5760 a_19336_18540# X1.X2.X1.X2.X1.X1.vout 1.64e-19
C5761 a_19722_18540# a_19422_16634# 5.25e-20
C5762 X1.X1.X3.vin1 a_4782_12822# 2.12e-19
C5763 a_39966_7922# a_39966_6016# 0.00198f
C5764 X2.X2.X1.X2.X3.vin2 vdd 1.29f
C5765 d3 X2.X2.X1.X1.X2.X1.X3.vin1 0.0195f
C5766 d2 X1.X2.X2.X2.X3.vin2 0.0685f
C5767 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.vout 0.075f
C5768 a_31862_19446# d1 0.00148f
C5769 a_16836_15634# a_17222_15634# 0.419f
C5770 X2.X1.X1.X1.X1.X2.X3.vin2 vdd 0.787f
C5771 a_46502_17540# a_46502_15634# 0.00198f
C5772 d2 a_40352_11734# 0.00272f
C5773 a_46502_23258# d2 0.00665f
C5774 d2 a_33976_7064# 0.608f
C5775 d1 a_23126_5016# 0.0752f
C5776 a_11072_28888# vdd 1.05f
C5777 a_31862_6104# X2.X1.X1.X2.X2.X2.X1.vin2 0.273f
C5778 X1.X1.X2.X2.X1.X2.X1.vin2 d1 0.00406f
C5779 X2.X1.X2.X1.X3.vin2 vdd 1.32f
C5780 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin2 0.1f
C5781 d4 X1.X1.X2.X2.X2.X2.vout 1.45e-19
C5782 X2.X1.X1.X2.X2.X2.X2.vin1 a_31476_4198# 0.197f
C5783 X1.X2.X2.X2.X1.X2.X3.vin2 a_25712_25076# 0.354f
C5784 a_52492_25982# X2.X2.X2.X2.X1.X2.X3.vin2 0.00535f
C5785 d3 X2.X1.X1.X2.X2.X1.X1.vin2 3.99e-21
C5786 X1.X1.X1.X2.X2.X2.X3.vin1 d1 0.149f
C5787 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X3.vin2 0.234f
C5788 d2 a_19422_5198# 0.00202f
C5789 X2.X1.X1.X2.X2.X2.X2.vin1 X2.X1.X2.vrefh 0.564f
C5790 X1.X2.X2.X1.X2.X2.vrefh d1 0.0124f
C5791 a_37766_5016# X2.X1.X2.X1.X1.X1.X3.vin1 0.428f
C5792 X1.X2.X1.X2.X2.X2.X1.vin1 d2 9.24e-20
C5793 X2.X1.X1.X1.X1.X1.X1.vin2 a_31862_30882# 8.88e-20
C5794 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X3.vin1 0.206f
C5795 a_17222_19446# d1 0.00148f
C5796 d3 X1.X2.X1.X2.X2.X1.X3.vin1 0.0195f
C5797 X2.X1.X3.vin1 a_37466_14586# 2.24e-19
C5798 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.vout 0.197f
C5799 X2.X1.X1.X1.X2.X2.X3.vin2 a_31862_17540# 8.07e-19
C5800 a_25712_23170# a_25712_21264# 0.00396f
C5801 X2.X1.X1.X1.X2.X2.vout a_33976_18540# 7.93e-20
C5802 X2.X1.X1.X1.X2.X2.vout a_34062_20446# 0.418f
C5803 a_34362_22312# X2.X1.X1.X1.X2.X2.X3.vin2 3.85e-19
C5804 X1.X1.X1.X2.X2.X2.vrefh a_2196_8010# 0.118f
C5805 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X1.X3.vin2 0.0533f
C5806 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X3.vin1 2.33e-19
C5807 X1.X2.X2.X2.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin1 0.00437f
C5808 d3 X2.X1.X1.X1.X3.vin2 0.387f
C5809 X1.X1.X2.X2.X1.X2.vrefh d1 0.0071f
C5810 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X2.X2.vrefh 0.076f
C5811 a_2196_17540# d0 0.518f
C5812 X1.X2.X1.X1.X1.X1.X1.vin1 d1 1.51e-19
C5813 X1.X1.X2.X1.X2.X2.X1.vin2 X1.X1.X2.X1.X2.X2.X1.vin1 0.668f
C5814 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.X3.vin1 0.0174f
C5815 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 0.581f
C5816 a_2582_19446# d1 0.00148f
C5817 d2 X2.X1.X2.X1.X1.X2.X1.vin2 0.226f
C5818 X2.X1.X1.X2.X2.vrefh X1.X2.X2.X1.X2.vrefh 0.117f
C5819 X2.X2.X2.X1.X2.X1.X3.vin2 a_52106_10734# 3.49e-19
C5820 X2.X2.X3.vin1 X2.X2.X2.X3.vin1 3.45e-19
C5821 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 0.242f
C5822 a_25326_32700# a_25326_30794# 0.00198f
C5823 X1.X1.X2.X2.X1.X2.X3.vin1 a_8572_22210# 0.00329f
C5824 a_19036_24258# vdd 1.05f
C5825 X1.X2.X1.X2.X2.X2.X2.vin1 a_17222_4198# 0.402f
C5826 a_8186_6962# X1.X1.X2.X1.X1.X1.vout 0.386f
C5827 X1.X1.X2.X1.X2.X2.X1.vin1 a_11072_13640# 1.64e-19
C5828 a_10686_25076# d1 0.00151f
C5829 X1.X2.X2.X2.X2.X1.X1.vin1 a_25712_25076# 1.64e-19
C5830 X1.X2.X2.X2.X1.X1.vout a_23512_20264# 0.359f
C5831 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X3.vin1 0.00118f
C5832 d2 X1.X1.X1.X2.X1.X2.X2.vin1 0.0329f
C5833 d0 X2.X1.X2.X1.X2.X2.X1.vin2 0.276f
C5834 X1.X2.X1.X1.X2.X1.X1.vin2 d2 0.231f
C5835 a_46116_27070# d2 0.00533f
C5836 X1.X2.X2.X1.X1.X2.X3.vin1 a_23512_8828# 0.199f
C5837 a_48316_28070# d1 0.521f
C5838 X2.X1.X2.X2.X1.X1.X3.vin1 a_37852_18358# 0.00255f
C5839 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.X2.vin1 0.00117f
C5840 a_52406_31700# X2.X2.X2.X2.X2.X2.X3.vin2 0.277f
C5841 X1.X2.X3.vin1 vdd 0.858f
C5842 X2.X1.X1.X1.X3.vin2 X2.X1.X2.X3.vin2 7.46e-20
C5843 a_8572_25982# a_8486_27888# 3.21e-19
C5844 a_37466_25982# X2.X1.X2.X2.X3.vin1 0.372f
C5845 a_31862_27070# X2.X1.X1.X1.X1.X2.X1.vin2 8.88e-20
C5846 d2 X1.X1.X2.X2.X2.X1.X3.vin1 0.104f
C5847 X1.X1.X1.X1.X2.X1.X3.vin1 d2 0.104f
C5848 X1.X2.X2.X2.X2.X2.vrefh d1 0.0124f
C5849 a_8872_20264# d4 0.00161f
C5850 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X2.X1.X2.X2.X2.vrefh 0.0128f
C5851 X1.X1.X1.X1.X2.X1.X3.vin2 vdd 0.903f
C5852 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X1.X2.X2.X1.X2.X1.vin1 0.668f
C5853 X1.X2.X3.vin2 a_23212_18358# 0.355f
C5854 X2.X2.X2.X2.X2.X2.vrefh a_54992_28888# 0.118f
C5855 d0 X1.X1.X2.X1.X2.X1.X1.vin1 0.267f
C5856 X2.X2.X2.X2.X1.X2.X2.vin1 vdd 0.576f
C5857 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X1.X2.X1.vin1 2.23e-19
C5858 a_10686_19358# a_10686_17452# 0.00198f
C5859 a_34062_28070# X2.X1.X1.X1.X1.X2.X3.vin1 0.42f
C5860 X1.X2.X2.X2.X1.X2.X1.vin2 d0 0.276f
C5861 X1.X2.X2.X2.X2.vrefh d2 0.158f
C5862 X1.X1.X2.X2.X1.X2.X3.vin2 a_8186_22210# 3.85e-19
C5863 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X3.vin1 0.00789f
C5864 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X1.X2.X2.vin1 0.242f
C5865 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X2.vin1 0.242f
C5866 X1.X1.X2.X1.X1.X2.X1.vin2 X1.X1.X2.X1.X1.X2.X1.vin1 0.668f
C5867 a_33976_18540# a_34062_16634# 3.21e-19
C5868 a_34362_18540# a_33676_16634# 2.97e-19
C5869 a_23212_6962# a_25326_6016# 2.95e-20
C5870 X2.X1.X1.X3.vin1 d4 1f
C5871 a_2582_21352# X1.X1.X1.X1.X2.X2.X1.vin2 0.273f
C5872 d0 a_54992_13640# 0.515f
C5873 d0 X1.X2.X1.X2.X1.X1.X2.vin1 0.262f
C5874 d2 a_19336_10916# 0.0057f
C5875 d0 X2.X3.vin2 0.00479f
C5876 a_23512_27888# a_23212_25982# 6.2e-19
C5877 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X2.vrefh 0.267f
C5878 X1.X1.X2.X1.X3.vin1 a_8572_10734# 0.169f
C5879 X1.X2.X2.X2.X1.X1.vout X1.X2.X2.X2.X1.X1.X3.vin2 0.342f
C5880 X2.X1.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X1.X3.vin2 0.0533f
C5881 a_52492_22210# d2 0.526f
C5882 a_16836_30882# a_17222_30882# 0.419f
C5883 d0 X2.X1.X2.X1.X2.X1.X3.vin2 4.34e-19
C5884 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X2.X1.X2.X2.vrefh 0.00437f
C5885 X2.X1.X1.X2.X2.vrefh a_31476_9916# 1.64e-19
C5886 X1.X2.X2.X1.X1.X2.X2.vin1 vdd 0.576f
C5887 X2.X1.X1.X2.X1.X1.vout X2.X1.X1.X2.X1.X1.X3.vin2 0.342f
C5888 a_19336_22312# a_17222_21352# 2.68e-20
C5889 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X1.vin2 0.668f
C5890 d4 X1.X1.X1.X1.X1.X2.X3.vin1 0.00851f
C5891 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X3.vin1 0.206f
C5892 X2.X1.X2.X2.X2.X2.X1.vin2 d0 0.253f
C5893 a_23212_29834# d1 0.00613f
C5894 X2.X2.X1.X1.X1.X2.X3.vin1 d0 4.36e-19
C5895 X1.X1.X2.X2.X1.X2.X2.vin1 a_10686_23170# 8.88e-20
C5896 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X1.vin2 8.93e-19
C5897 d3 X1.X2.X2.X1.X2.X1.X3.vin1 0.0195f
C5898 a_4696_14688# a_2582_13728# 2.68e-20
C5899 a_33976_14688# a_34362_14688# 0.419f
C5900 a_31862_21352# vdd 0.553f
C5901 X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin1 0.00304f
C5902 X1.X2.X2.X2.X2.X2.X3.vin2 X2.vrefh 0.183f
C5903 d0 X1.X2.X1.X2.X2.X1.X2.vin1 0.262f
C5904 d0 a_54606_17452# 0.0489f
C5905 X1.X1.X1.X1.X3.vin2 a_4696_22312# 0.363f
C5906 X1.X3.vin1 a_14082_892# 0.413f
C5907 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X1.vin2 0.076f
C5908 a_37766_12640# a_37852_10734# 3.21e-19
C5909 a_19722_26164# vdd 0.489f
C5910 d0 X1.X1.X2.X1.X1.X1.X3.vin1 4.36e-19
C5911 a_52406_20264# d4 0.00154f
C5912 X1.X2.X2.X1.X2.X2.X3.vin1 a_25712_15546# 0.354f
C5913 d3 a_31862_25164# 0.00112f
C5914 X1.X1.X2.vrefh X1.X3.vin1 0.0451f
C5915 d0 X2.X2.X2.X1.X2.vrefh 0.844f
C5916 X1.X1.X2.X2.X2.X2.X1.vin2 X1.X1.X2.X2.X2.X2.X1.vin1 0.668f
C5917 a_46502_17540# a_48316_16634# 1.06e-19
C5918 a_19036_16634# a_17222_15634# 1.15e-20
C5919 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X2.vin1 0.0689f
C5920 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 0.049f
C5921 a_40352_11734# X2.X1.X2.X1.X2.vrefh 1.64e-19
C5922 X2.X1.X3.vin2 d2 0.1f
C5923 a_48316_24258# d2 3.82e-19
C5924 a_37466_25982# a_37766_24076# 4.41e-20
C5925 X1.X1.X3.vin2 d5 0.0378f
C5926 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X1.X2.X1.X1.X2.X3.vin2 3.94e-19
C5927 X1.X1.X2.X1.X2.X1.X1.vin1 a_10686_9828# 8.22e-20
C5928 a_5082_14688# X1.X1.X1.X2.X1.X2.vout 0.254f
C5929 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin2 0.12f
C5930 X2.X2.X1.X1.X3.vin1 vdd 0.805f
C5931 a_2196_23258# d2 0.00464f
C5932 X1.X2.X1.X1.X1.X1.X2.vin1 d0 0.262f
C5933 a_10686_17452# a_11072_17452# 0.419f
C5934 a_37766_20264# d4 0.0013f
C5935 X1.X1.X2.X1.X2.X1.vout vdd 0.805f
C5936 a_10686_25076# X1.X1.X2.X2.X1.X2.X3.vin2 0.567f
C5937 X2.X1.X1.X1.X1.X1.X1.vin2 a_34062_31882# 0.00743f
C5938 d3 a_2582_9916# 0.00112f
C5939 X2.X1.X2.X1.X2.X1.X1.vin2 a_39966_11734# 0.273f
C5940 a_4696_22312# vdd 1.05f
C5941 d3 X1.X1.X1.X2.X1.X1.vout 0.00883f
C5942 a_2196_17540# X1.X1.X1.X2.X1.X1.X3.vin1 0.354f
C5943 a_2582_17540# X1.X1.X1.X2.X1.X1.X1.vin1 0.417f
C5944 a_17222_23258# X1.X2.X1.X1.X2.X2.X1.vin1 8.22e-20
C5945 a_2582_25164# X1.X1.X1.X1.X1.X2.X3.vin2 8.07e-19
C5946 X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.vout 3.08e-19
C5947 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X3.vin1 0.449f
C5948 X2.X1.X2.X1.X2.X2.X3.vin1 a_37466_14586# 0.00874f
C5949 a_37466_10734# a_37766_8828# 4.41e-20
C5950 a_48316_28070# X2.X2.X1.X1.X1.X2.X3.vin2 0.101f
C5951 d3 X2.X2.X1.X2.X1.X2.vout 0.0232f
C5952 a_22826_25982# X1.X2.X2.X2.X1.X2.X3.vin2 0.00846f
C5953 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X3.vin1 1.42e-20
C5954 a_2582_11822# a_4696_10916# 4.72e-20
C5955 X1.X1.X1.X1.X2.X2.X1.vin2 a_2196_19446# 1.78e-19
C5956 a_23126_20264# d4 0.00154f
C5957 d3 X2.X2.X1.X1.X1.X1.X1.vin2 1.14e-19
C5958 d0 a_54606_7922# 0.0675f
C5959 d3 X1.X1.X1.X3.vin1 0.675f
C5960 a_19336_14688# a_19422_12822# 3.38e-19
C5961 a_19722_14688# a_19036_12822# 3.31e-19
C5962 a_23212_22210# a_23126_20264# 3.14e-19
C5963 X1.X2.X1.X2.X2.X1.X1.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 2.23e-19
C5964 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X1.vin2 0.076f
C5965 a_48616_18540# a_48316_16634# 6.2e-19
C5966 a_23212_10734# X1.X2.X2.X1.X1.X2.X3.vin2 0.00535f
C5967 X2.X1.X1.X2.X1.X2.X1.vin1 d1 0.0118f
C5968 a_2582_15634# a_2582_13728# 0.00198f
C5969 a_54992_28888# d1 2.92e-22
C5970 a_17222_27070# a_17222_25164# 0.00198f
C5971 a_16836_27070# X1.X2.X1.X1.X2.X1.X1.vin1 1.64e-19
C5972 a_2196_15634# X1.X1.X1.X2.X1.X2.X1.vin1 1.64e-19
C5973 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X1.X3.vin1 0.0425f
C5974 d2 a_46502_13728# 0.00479f
C5975 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 1.22e-19
C5976 a_31862_27070# a_33976_26164# 4.72e-20
C5977 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X3.vin1 2.33e-19
C5978 X2.X1.X1.X2.X1.X2.vrefh vdd 0.414f
C5979 d5 a_6032_892# 0.04f
C5980 X2.X2.X3.vin1 a_52406_8828# 8.66e-20
C5981 a_37852_14586# a_39966_13640# 2.95e-20
C5982 X2.X1.X2.X2.X2.X1.X3.vin2 d1 0.15f
C5983 a_25326_11734# a_25712_11734# 0.419f
C5984 a_37852_18358# X2.X1.X2.X1.X2.X2.vout 7.93e-20
C5985 X2.X1.X2.X1.X2.X2.X1.vin2 a_40352_15546# 0.12f
C5986 a_39966_15546# X2.X1.X2.X1.X2.X2.X1.vin1 0.417f
C5987 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X3.vin1 1.22e-19
C5988 d2 X2.X2.X2.X2.X2.X1.X2.vin1 0.0318f
C5989 d2 X1.X1.X2.X1.X2.X2.X3.vin1 0.153f
C5990 a_38152_8828# a_37852_6962# 6.71e-19
C5991 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.X1.vin2 0.22f
C5992 X2.X1.X1.X1.X1.X2.X2.vin1 X2.X1.X1.X1.X1.X2.X1.vin2 0.242f
C5993 X2.X1.X1.X1.X1.X1.vout X2.X1.X1.X1.X1.X1.X3.vin2 0.342f
C5994 X1.X2.X1.X3.vin1 X1.X2.X2.X3.vin2 1.22e-19
C5995 a_46116_17540# d1 2.25e-20
C5996 a_5082_22312# a_4782_20446# 5.55e-20
C5997 a_17222_15634# vdd 0.541f
C5998 a_40352_6016# vdd 1.05f
C5999 X1.X1.X1.X1.X2.X2.vout a_4396_20446# 0.36f
C6000 X1.X1.X1.X2.X2.vrefh vdd 0.426f
C6001 X2.X2.X2.X1.X1.X1.vout a_52492_6962# 0.169f
C6002 d2 a_54992_17452# 0.00441f
C6003 X2.X1.X1.X1.X2.X1.X1.vin2 vdd 0.36f
C6004 a_4396_9010# a_4696_7064# 6.1e-19
C6005 X1.X2.X1.X2.X3.vin2 X1.X2.X2.X1.X3.vin1 0.0604f
C6006 d1 X1.X1.X1.X2.X2.X2.X2.vin1 0.0144f
C6007 a_11072_32700# d0 0.515f
C6008 X1.X1.X2.X3.vin1 a_8572_18358# 0.17f
C6009 X1.X2.X2.X1.X1.X1.X3.vin2 vdd 0.937f
C6010 X2.X2.X2.X2.X1.X1.X3.vin2 a_52792_20264# 0.1f
C6011 d0 X2.X1.X1.X2.X2.X1.X2.vin1 0.262f
C6012 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X2.vin1 0.564f
C6013 X1.X2.X1.X1.X2.X1.X3.vin1 vdd 0.997f
C6014 d2 X2.X1.X2.X1.X2.X2.X3.vin2 0.113f
C6015 X2.X1.X2.X1.X2.X1.X2.vin1 a_40352_11734# 1.78e-19
C6016 X2.X1.X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X1.vin1 2.23e-19
C6017 X2.X1.X2.X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X2.X1.vin1 2.23e-19
C6018 X2.X1.X2.X2.X1.X2.X2.vin1 a_40352_23170# 1.78e-19
C6019 d1 a_31862_4198# 0.0015f
C6020 X1.X1.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X1.X3.vin1 0.0321f
C6021 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X1.X2.X2.X2.vin1 0.00117f
C6022 a_46502_21352# a_48702_20446# 4.2e-20
C6023 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X2.X1.vin2 0.216f
C6024 X1.X2.X2.X2.X2.X2.X3.vin1 a_25712_30794# 0.354f
C6025 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X1.X1.vin1 0.206f
C6026 a_39966_26982# d0 0.0675f
C6027 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin2 0.12f
C6028 X1.X2.X1.X2.X3.vin1 a_19722_10916# 0.372f
C6029 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X2.X1.X2.X1.X2.X2.vin1 0.00232f
C6030 d0 a_25326_13640# 0.0489f
C6031 X1.X1.X1.X2.X2.X1.X1.vin2 vdd 0.36f
C6032 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 2.23e-19
C6033 a_19036_28070# d2 0.00393f
C6034 a_22826_22210# d2 0.0191f
C6035 X2.X2.X2.X2.X3.vin2 a_52492_29834# 0.363f
C6036 X1.X2.X2.X2.X1.X2.X1.vin2 a_25712_23170# 0.12f
C6037 a_25326_23170# X1.X2.X2.X2.X1.X2.X1.vin1 0.417f
C6038 a_19036_31882# a_17222_30882# 1.15e-20
C6039 X2.X1.X2.X2.X3.vin1 vdd 0.804f
C6040 X1.X1.X2.X2.X1.X1.X3.vin1 a_8572_18358# 0.00255f
C6041 a_31476_8010# a_31862_8010# 0.419f
C6042 X2.X1.X1.X1.X1.X2.vrefh vdd 0.43f
C6043 a_46502_9916# a_48702_9010# 4.2e-20
C6044 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.X2.vin1 0.00117f
C6045 d5 X3.vin2 0.00102f
C6046 a_31862_28976# d0 0.0675f
C6047 d5 a_20672_892# 0.033f
C6048 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X2.vrefh 0.00118f
C6049 X2.X1.X2.X2.X1.X1.X3.vin2 X2.X1.X2.X2.X1.X1.X3.vin1 0.581f
C6050 a_38152_12640# d1 0.521f
C6051 a_37852_18358# d1 0.00638f
C6052 a_11072_21264# vdd 1.05f
C6053 d3 a_25326_32700# 1.28e-19
C6054 d2 a_19722_29936# 0.254f
C6055 d2 X1.X1.X2.X2.X2.X2.X3.vin1 0.0571f
C6056 X1.X1.X1.X2.X1.X2.X3.vin2 a_2582_11822# 0.567f
C6057 a_54606_17452# X2.X2.X2.X1.X2.X2.X3.vin1 0.00207f
C6058 X2.X1.X1.X3.vin1 X2.X1.X1.X3.vin2 0.552f
C6059 X1.X2.X1.X2.X1.X2.X1.vin2 a_16836_11822# 1.78e-19
C6060 X2.X2.X1.X2.X1.X2.X3.vin2 a_46502_11822# 0.567f
C6061 a_17222_32788# X1.X2.X1.X1.X1.X1.X1.vin2 0.273f
C6062 a_17222_30882# vdd 0.541f
C6063 X1.X1.X2.X2.X1.X1.X3.vin1 a_11072_19358# 0.354f
C6064 a_52406_16452# a_52106_14586# 5.55e-20
C6065 X1.X2.X2.X2.X1.X2.vrefh a_25712_21264# 0.118f
C6066 d3 X2.X2.X2.X1.X2.X1.X3.vin2 2.81e-19
C6067 d0 X1.X2.X1.X2.X1.X1.X1.vin1 0.267f
C6068 X1.X1.X3.vin2 a_6032_892# 0.268f
C6069 a_34362_14688# vdd 0.477f
C6070 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin2 7.84e-19
C6071 X1.X2.X1.X2.X1.X2.X3.vin1 a_19036_12822# 0.199f
C6072 a_52406_27888# d3 0.00148f
C6073 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X2.X1.vout 0.038f
C6074 d3 X1.X1.X1.X1.X1.X2.X2.vin1 8.68e-20
C6075 a_34362_14688# a_34062_12822# 5.55e-20
C6076 X1.X2.X2.X2.X1.X2.vout a_22826_22210# 0.254f
C6077 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 2.23e-19
C6078 X1.X1.X2.X2.X1.X1.X3.vin2 a_8186_18358# 3.49e-19
C6079 a_19036_16634# a_19422_16634# 0.419f
C6080 X2.X1.X1.X2.X2.X2.vout a_34062_5198# 0.418f
C6081 X1.X1.X1.X2.X2.X2.X3.vin1 a_4782_5198# 0.42f
C6082 a_34362_7064# X2.X1.X1.X2.X2.X2.X3.vin2 3.85e-19
C6083 d4 a_48316_16634# 0.00176f
C6084 a_39966_26982# a_39966_25076# 0.00198f
C6085 X1.X2.X2.X1.X1.X2.X1.vin2 X1.X2.X2.X1.X1.X2.X1.vin1 0.668f
C6086 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X2.vrefh 0.076f
C6087 X2.X1.X2.X1.X2.X2.X3.vin2 a_38152_16452# 0.101f
C6088 X1.X1.X2.X3.vin1 d2 6.42e-19
C6089 a_31862_32788# X2.X1.X1.X1.X1.X1.X3.vin2 7.84e-19
C6090 X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin2 0.00254f
C6091 X1.X1.X2.X3.vin1 a_8186_10734# 0.509f
C6092 X2.X2.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 0.0565f
C6093 a_25326_19358# X1.X2.X2.X1.X2.X2.X3.vin2 8.07e-19
C6094 a_39966_11734# vdd 0.553f
C6095 a_2196_25164# a_2582_25164# 0.419f
C6096 X1.X1.X1.X2.X1.X1.X1.vin1 vdd 0.592f
C6097 a_46502_27070# a_46502_28976# 0.00198f
C6098 a_48616_10916# a_46502_9916# 5.36e-21
C6099 a_52406_27888# X2.X2.X2.X2.X2.X1.X3.vin2 0.267f
C6100 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X3.vin1 0.00118f
C6101 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X1.vin2 0.668f
C6102 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X2.X1.X2.vin1 0.00117f
C6103 a_4696_29936# X1.X1.X1.X1.X1.X2.vout 0.0929f
C6104 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X2.vin1 0.242f
C6105 X2.X1.X2.X2.X2.X2.X1.vin2 a_40352_30794# 0.12f
C6106 a_39966_30794# X2.X1.X2.X2.X2.X2.X1.vin1 0.417f
C6107 a_52406_16452# vdd 0.471f
C6108 X1.X2.X1.X2.X2.X2.X2.vin1 vdd 0.578f
C6109 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X1.X2.X2.X1.X1.X3.vin1 0.00117f
C6110 X1.X1.X2.X2.X1.X1.X3.vin2 a_8486_20264# 0.267f
C6111 a_19036_24258# a_19422_24258# 0.419f
C6112 a_16836_6104# vdd 1.05f
C6113 X1.X2.X1.X2.X1.X1.X3.vin1 a_17222_15634# 0.00207f
C6114 a_10686_15546# d1 3.41e-19
C6115 X1.X1.X3.vin1 X1.X1.X1.X2.X3.vin1 7.18e-19
C6116 X2.X1.X2.X1.X2.X2.X1.vin1 vdd 0.592f
C6117 X1.X1.X2.X2.X1.X1.X3.vin1 d2 0.104f
C6118 X1.X1.X2.X2.vrefh a_10686_17452# 0.3f
C6119 X2.X1.X1.X2.X2.X2.X1.vin2 a_31476_4198# 1.78e-19
C6120 a_5646_892# X1.X3.vin1 0.354f
C6121 d3 X1.X2.X1.X2.X3.vin1 0.375f
C6122 a_11072_9828# a_11072_7922# 0.00396f
C6123 X1.X1.X1.X2.X2.X2.X3.vin1 a_5082_7064# 0.00874f
C6124 d3 a_8572_22210# 7.7e-20
C6125 a_16836_13728# d1 2.25e-20
C6126 X2.X1.X2.X1.X1.X1.X3.vin2 a_38152_5016# 0.1f
C6127 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X2.vrefh 0.076f
C6128 a_34362_26164# X2.X1.X1.X1.X3.vin2 0.241f
C6129 a_37766_24076# vdd 0.47f
C6130 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X2.vrefh 0.267f
C6131 X2.X1.X2.X1.X3.vin1 d1 0.00179f
C6132 d1 d5 9.06f
C6133 d2 a_25712_13640# 0.00464f
C6134 X2.X1.X1.X1.X1.X1.X1.vin1 d0 0.0488f
C6135 a_19036_9010# a_19422_9010# 0.419f
C6136 a_8486_8828# vdd 0.47f
C6137 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X1.X2.X2.X2.X2.vin1 0.00117f
C6138 a_31862_6104# a_34062_5198# 4.2e-20
C6139 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 0.234f
C6140 X1.X2.X2.X2.X1.X2.X1.vin1 vdd 0.592f
C6141 a_23512_24076# a_25326_23170# 1.06e-19
C6142 a_10686_7922# d1 3.41e-19
C6143 X1.X2.X1.X1.X2.X2.vrefh a_17222_23258# 0.3f
C6144 a_31862_8010# vdd 0.541f
C6145 a_25326_28888# d1 0.00148f
C6146 d2 X1.X1.X2.X1.X2.X1.X3.vin2 0.171f
C6147 X2.X2.X2.X1.X2.X2.X3.vin2 a_52106_14586# 3.85e-19
C6148 a_25712_32700# vdd 1.05f
C6149 X1.X1.X2.X1.X2.X1.X3.vin2 a_8186_10734# 3.49e-19
C6150 d2 X2.X1.X1.X1.X1.X2.X1.vin2 0.226f
C6151 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X3.vin1 0.546f
C6152 a_34062_24258# a_31862_23258# 4.77e-21
C6153 a_2582_6104# X1.X1.X1.X2.X2.X2.vrefh 8.22e-20
C6154 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.X1.X3.vin2 2.23e-19
C6155 a_52106_14586# X2.X2.X2.X1.X2.X1.vout 0.383f
C6156 a_25712_26982# X1.X2.X2.X2.X2.X1.X2.vin1 1.78e-19
C6157 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X2.vrefh 0.00118f
C6158 X1.X1.X1.X1.X2.X2.X3.vin2 X1.X1.X1.X2.X1.X1.X1.vin1 5.19e-19
C6159 X1.X1.X2.X1.X2.X2.X3.vin2 X1.X1.X2.X1.X2.X2.X1.vin1 2.23e-19
C6160 a_54992_23170# a_54992_21264# 0.00396f
C6161 X1.X1.X2.X1.X2.X2.X2.vin1 a_11072_15546# 1.78e-19
C6162 d2 X1.X2.X1.X1.X1.X2.X3.vin1 0.158f
C6163 X2.X2.X2.X1.X2.X1.X1.vin2 d1 4.01e-19
C6164 X2.X2.X1.X2.X2.X1.vout X2.X2.X1.X2.X2.X1.X3.vin2 0.326f
C6165 X1.X1.X1.X1.X1.X1.X3.vin1 a_4782_31882# 0.428f
C6166 a_40352_25076# X2.X1.X2.X2.X1.X2.X1.vin2 1.78e-19
C6167 a_40352_13640# X2.X1.X2.X1.X2.X1.X1.vin2 1.78e-19
C6168 a_19422_16634# vdd 0.561f
C6169 a_8186_25982# d2 7.13e-19
C6170 a_19036_20446# a_19722_18540# 3.08e-19
C6171 a_19422_20446# a_19336_18540# 3.3e-19
C6172 a_52406_31700# vdd 0.471f
C6173 X1.X1.X1.X1.X2.X2.X3.vin1 d4 2.08e-19
C6174 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X3.vin1 2.33e-19
C6175 d0 X1.X1.X2.X1.X1.X2.vrefh 0.848f
C6176 a_4782_16634# X1.X1.X1.X2.X3.vin1 1.52e-19
C6177 d2 a_25326_17452# 0.00583f
C6178 X1.X1.X1.X2.X1.X1.vout a_5082_14688# 0.387f
C6179 a_2582_25164# vdd 0.553f
C6180 X2.X2.X1.X1.X2.X2.X3.vin1 d0 4.36e-19
C6181 d4 X2.X2.X1.X1.X1.X1.X1.vin1 0.00332f
C6182 a_48616_22312# X2.X2.X1.X1.X2.X2.vout 0.0929f
C6183 a_10686_30794# d1 3.41e-19
C6184 X2.X2.X2.X2.X1.X2.X2.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 0.234f
C6185 X2.X1.X2.X2.X2.X2.X1.vin1 vdd 0.592f
C6186 X2.X2.X2.X1.X1.X2.X2.vin1 X2.X2.X2.X1.X1.X2.X3.vin1 0.00117f
C6187 X1.X2.X1.X1.X2.vrefh a_16836_27070# 0.118f
C6188 X2.X2.X2.X1.X1.X2.X3.vin2 a_52406_8828# 0.277f
C6189 a_40352_32700# X2.X2.vrefh 0.118f
C6190 X2.X2.X2.X2.X1.X1.X3.vin1 d1 0.146f
C6191 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.vrefh 2.33e-19
C6192 d2 X2.X1.X2.X2.X2.X1.vout 0.115f
C6193 X2.X2.X2.X2.X1.X1.X1.vin2 d4 3.99e-21
C6194 X2.X2.X1.X3.vin1 a_48702_24258# 5.28e-19
C6195 X2.X2.X1.X2.X3.vin1 a_48702_12822# 9.54e-19
C6196 a_49002_14688# X2.X2.X1.X2.X1.X2.X3.vin2 3.85e-19
C6197 X2.X2.X2.X2.X2.vrefh a_54992_25076# 0.118f
C6198 a_19422_9010# vdd 0.561f
C6199 d2 a_4696_14688# 0.526f
C6200 X2.X1.X2.X1.X1.X2.X3.vin1 a_40352_7922# 0.354f
C6201 d3 X1.X1.X2.X1.X2.X1.X1.vin2 3.99e-21
C6202 d1 X1.X2.X1.X2.X2.X2.vout 0.0331f
C6203 a_39966_21264# a_38152_20264# 1.15e-20
C6204 X2.X1.X1.X1.X1.X2.X3.vin2 d0 4.34e-19
C6205 X1.X1.X2.X2.X1.X1.vout d4 0.00132f
C6206 X1.X1.X1.X2.X1.X2.vout a_4696_10916# 7.93e-20
C6207 X2.X2.X2.X1.X2.X2.X3.vin2 vdd 0.761f
C6208 X2.X2.X1.X1.X2.X2.X3.vin2 d2 0.113f
C6209 a_19036_31882# a_19422_31882# 0.419f
C6210 X2.X2.X2.X1.X2.X1.vout vdd 0.805f
C6211 d4 X1.X1.X2.X1.X2.X2.X3.vin2 0.0264f
C6212 a_33676_9010# a_31862_8010# 1.15e-20
C6213 a_11072_28888# d0 0.515f
C6214 X2.X1.X2.X2.X2.X1.vout a_37852_29834# 0.169f
C6215 X2.X1.X2.X2.X1.X1.X3.vin1 d1 0.146f
C6216 a_31862_21352# X2.X1.X1.X1.X2.X2.X2.vin1 8.88e-20
C6217 a_19722_26164# a_19422_24258# 5.25e-20
C6218 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.X1.vin2 3.94e-19
C6219 X1.X2.X2.X1.X2.X1.X1.vin1 d1 0.0118f
C6220 a_19336_26164# X1.X2.X1.X1.X2.X1.vout 1.64e-19
C6221 X1.X1.X1.X2.vrefh a_2582_19446# 0.3f
C6222 a_8872_20264# a_10686_19358# 1.06e-19
C6223 a_31862_23258# d1 0.00148f
C6224 d3 X1.X1.X2.X2.X2.X2.X3.vin2 0.109f
C6225 X2.X2.X2.X2.X1.X2.X3.vin1 a_52492_22210# 0.00329f
C6226 a_16836_27070# vdd 1.05f
C6227 X2.X2.X2.X2.X1.X1.X3.vin1 a_54606_19358# 0.52f
C6228 X1.X1.X2.vrefh a_11072_4110# 9.79e-19
C6229 d4 a_8186_29834# 5.68e-19
C6230 X2.X2.vrefh vdd 0.419f
C6231 X2.X2.X1.X2.X1.X1.vout X2.X2.X1.X2.X3.vin1 0.131f
C6232 X1.X1.X3.vin2 d1 0.0461f
C6233 a_49002_10916# X2.X2.X1.X2.X2.X1.X3.vin2 3.49e-19
C6234 a_34362_18540# d2 0.00132f
C6235 a_39966_17452# a_39966_15546# 0.00198f
C6236 X1.X2.X1.X3.vin1 X1.X2.X3.vin1 0.188f
C6237 X2.X1.X1.X1.X2.X2.X3.vin2 d2 0.113f
C6238 a_48616_7064# a_49002_7064# 0.419f
C6239 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 0.242f
C6240 a_19422_31882# vdd 0.565f
C6241 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X2.vrefh 0.00118f
C6242 X2.X2.X2.X2.X1.X2.X1.vin2 X2.X2.X2.X2.X1.X2.vrefh 0.1f
C6243 a_37852_22210# a_38152_20264# 6.1e-19
C6244 a_31862_9916# X2.X1.X1.X2.X2.X1.X1.vin2 0.273f
C6245 X1.X1.X1.X1.X2.X1.X2.vin1 d1 1.03e-19
C6246 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.X2.vin1 0.242f
C6247 X1.X2.X2.X2.X1.X1.X3.vin1 d1 0.146f
C6248 d3 X2.X2.X1.X3.vin1 0.702f
C6249 a_25326_21264# X1.X2.X2.X2.X1.X1.X3.vin1 0.00207f
C6250 X1.X1.X1.X1.X1.X2.X3.vin2 a_2196_27070# 0.354f
C6251 a_49002_7064# vdd 0.477f
C6252 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 0.234f
C6253 a_39966_32700# d2 1.95e-19
C6254 X1.X1.X2.X1.X2.X1.X3.vin2 a_8872_12640# 0.1f
C6255 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X2.X1.X1.X1.X1.X1.vin2 0.00232f
C6256 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X2.vrefh 0.076f
C6257 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X1.vin2 0.076f
C6258 X2.X2.X1.X2.X2.X1.X1.vin2 d1 4.01e-19
C6259 d4 a_4696_18540# 0.63f
C6260 a_28096_892# a_28482_892# 0.419f
C6261 a_23512_24076# vdd 1.05f
C6262 X1.X2.X1.X1.X2.X2.X3.vin2 d2 0.113f
C6263 a_28482_892# vdd 0.473f
C6264 a_2582_13728# a_4782_12822# 4.2e-20
C6265 X1.X2.X2.X1.X2.X1.vout X1.X2.X2.X1.X2.X1.X3.vin1 0.118f
C6266 X1.X1.X1.X2.X3.vin2 a_4782_9010# 0.00101f
C6267 X1.X1.X1.X2.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X2.vin1 0.00117f
C6268 X2.X1.X1.X2.X2.X1.X3.vin1 d1 0.151f
C6269 a_48316_28070# a_48616_26164# 6.48e-19
C6270 X2.X1.X1.X2.X1.X2.X3.vin2 vdd 0.787f
C6271 d1 a_25326_7922# 3.41e-19
C6272 d2 X1.X2.X1.X2.X1.X2.vrefh 0.177f
C6273 X2.X2.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X3.vin2 0.0533f
C6274 a_37766_20264# a_39966_19358# 4.2e-20
C6275 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X2.X1.X1.X1.vin2 0.216f
C6276 X1.X1.X1.X1.X2.X1.X3.vin2 a_5082_22312# 0.00815f
C6277 d2 X2.X2.X1.X2.X2.X1.X1.vin1 0.0105f
C6278 a_54992_21264# d1 2.92e-22
C6279 a_39966_21264# a_40352_21264# 0.419f
C6280 a_54992_7922# vdd 1.05f
C6281 X2.X2.X1.X1.X1.X2.X2.vin1 a_46116_28976# 1.78e-19
C6282 a_39966_15546# X2.X1.X2.X1.X2.X2.vrefh 8.22e-20
C6283 a_34062_12822# X2.X1.X1.X2.X1.X2.X3.vin2 0.277f
C6284 X1.X2.X3.vin1 d0 0.04f
C6285 a_23512_27888# d3 0.00178f
C6286 a_48316_16634# X2.X2.X1.X2.X1.X1.vout 0.359f
C6287 d3 X2.X1.X1.X1.X2.X2.vout 8.47e-19
C6288 X2.X1.X2.X2.X1.X1.X3.vin2 d1 0.15f
C6289 a_31476_21352# X2.X1.X1.X1.X2.X2.X3.vin1 0.354f
C6290 a_2196_21352# X1.X1.X1.X1.X2.X2.X2.vin1 1.78e-19
C6291 a_31862_21352# X2.X1.X1.X1.X2.X2.X1.vin1 0.417f
C6292 X1.X2.X1.X1.X1.X1.X1.vin2 X1.X2.X1.X1.X1.X1.X3.vin2 8.93e-19
C6293 X1.X1.X1.X1.X2.X1.X3.vin2 d0 4.34e-19
C6294 X1.X2.X1.X1.X2.X2.X3.vin2 a_17222_17540# 8.07e-19
C6295 X2.X2.X2.X1.X1.X2.X1.vin1 a_54992_7922# 0.195f
C6296 d2 a_2582_15634# 0.0059f
C6297 X2.X2.X2.X2.X1.X1.X2.vin1 d2 0.031f
C6298 X1.X2.X2.X2.X2.X1.X3.vin2 X1.X2.X2.X2.X2.X2.vrefh 0.161f
C6299 X1.X2.X1.X2.X1.X1.X3.vin1 a_19422_16634# 0.428f
C6300 X1.X2.X1.X2.X1.X1.X3.vin2 a_19722_14688# 0.00815f
C6301 X2.X2.X2.X2.X1.X2.X2.vin1 d0 0.262f
C6302 a_52492_6962# a_54606_7922# 2.68e-20
C6303 X1.X1.X1.X2.X1.X2.vout X1.X1.X1.X2.X1.X2.X3.vin2 0.075f
C6304 X1.X1.X2.X1.X1.X2.X3.vin1 a_8186_6962# 0.00874f
C6305 a_33976_26164# d2 0.0057f
C6306 a_11072_26982# X1.X1.X2.X2.X2.X1.X3.vin1 0.354f
C6307 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X2.X1.X1.vin2 0.216f
C6308 a_23126_12640# a_25326_11734# 4.2e-20
C6309 X2.X2.X2.X2.X2.X2.vrefh d1 0.0124f
C6310 a_46116_17540# X2.X2.X1.X2.X1.X1.X1.vin1 0.195f
C6311 X1.X1.X1.X2.X3.vin2 d1 0.00807f
C6312 X2.X2.X2.vrefh X2.X2.X2.X1.X1.X1.X1.vin1 0.142f
C6313 a_19722_26164# X1.X2.X1.X3.vin1 0.509f
C6314 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.vrefh 2.33e-19
C6315 a_49002_22312# d1 0.0422f
C6316 X2.X1.X2.X2.X3.vin1 a_37466_22210# 0.436f
C6317 X1.X2.X2.X2.X2.X1.X1.vin2 a_25712_28888# 1.78e-19
C6318 d3 a_52406_24076# 0.00122f
C6319 a_34062_9010# vdd 0.561f
C6320 a_11072_17452# X1.X1.X2.X1.X2.X2.X1.vin2 1.78e-19
C6321 a_5082_18540# X1.X1.X3.vin2 6.58e-20
C6322 d2 a_2582_8010# 0.00665f
C6323 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X2.X1.X1.X1.vin2 0.216f
C6324 a_23126_20264# a_25326_19358# 4.2e-20
C6325 X1.X2.X2.X2.X1.X2.X1.vin2 X1.X2.X2.X2.X1.X2.vrefh 0.1f
C6326 X2.X2.X2.X3.vin2 a_52406_20264# 5.21e-19
C6327 d0 X1.X2.X2.X1.X1.X2.X2.vin1 0.262f
C6328 X2.X1.X2.X2.X3.vin2 X2.X1.X2.X2.X2.X2.vout 0.0866f
C6329 X2.X2.X2.X1.X1.X2.X3.vin1 X2.X2.X2.X1.X1.X1.X3.vin2 1.22e-19
C6330 X1.X2.X1.X1.X2.X1.X3.vin1 a_19422_24258# 0.428f
C6331 a_52406_12640# a_52106_10734# 5.25e-20
C6332 d2 X1.X2.X1.X1.X1.X2.vrefh 6.65e-20
C6333 a_46502_23258# X2.X2.X1.X1.X2.X2.X1.vin1 8.22e-20
C6334 a_33676_24258# X2.X1.X1.X1.X2.X1.vout 0.359f
C6335 d2 a_2582_28976# 0.00479f
C6336 X2.X1.X2.X2.X3.vin2 d1 0.00807f
C6337 a_40352_13640# vdd 1.05f
C6338 X2.X1.X1.X3.vin1 X2.X1.X1.X1.X3.vin1 0.199f
C6339 a_31476_13728# a_31476_11822# 0.00396f
C6340 a_31476_25164# a_31476_23258# 0.00396f
C6341 d2 a_46116_11822# 0.00533f
C6342 d2 a_22826_14586# 0.0191f
C6343 a_48316_12822# d1 0.521f
C6344 a_2582_27070# d1 0.00151f
C6345 X1.X2.X2.X1.X2.X1.X3.vin2 vdd 0.903f
C6346 a_40352_26982# vdd 1.05f
C6347 X2.X1.X2.X2.X1.X1.X3.vin2 X2.X1.X2.X2.X1.X1.X1.vin2 8.93e-19
C6348 a_39966_13640# X2.X1.X2.X1.X2.X1.X3.vin1 0.00207f
C6349 X1.X1.X3.vin2 a_8486_12640# 2.33e-19
C6350 a_54992_23170# d1 2.25e-20
C6351 X2.X1.X2.X2.X1.X1.X2.vin1 a_39966_19358# 8.88e-20
C6352 a_22826_18358# a_23126_16452# 4.41e-20
C6353 a_23212_29834# X1.X2.X2.X2.X2.X1.X3.vin2 0.00546f
C6354 X2.X1.X2.X1.X3.vin1 a_37466_6962# 0.436f
C6355 X2.X2.X1.X1.X1.X2.X1.vin2 vdd 0.361f
C6356 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X1.vout 0.0524f
C6357 a_4396_9010# X1.X1.X1.X2.X2.X1.vout 0.359f
C6358 X1.X1.X2.X2.X3.vin1 a_8572_22210# 0.363f
C6359 a_31862_21352# d0 0.0675f
C6360 X2.vrefh X2.X1.X1.X1.X1.X1.X1.vin1 0.108f
C6361 a_46116_25164# X2.X2.X1.X1.X2.X1.X1.vin1 0.195f
C6362 d3 a_34062_16634# 4.67e-19
C6363 d2 a_2582_30882# 4.64e-19
C6364 d1 X3.vin2 3.83e-19
C6365 X2.X1.X1.X1.X1.X2.X3.vin1 vdd 0.96f
C6366 d1 a_20672_892# 5.18e-19
C6367 a_34362_10916# vdd 0.487f
C6368 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.X1.vin2 8.93e-19
C6369 X2.X1.X2.X1.X1.X2.X2.vin1 a_39966_7922# 8.88e-20
C6370 X2.X1.X2.vrefh a_39966_4110# 4.89e-19
C6371 a_8872_5016# vdd 1.05f
C6372 a_8186_25982# X1.X1.X2.X2.X3.vin2 0.263f
C6373 d2 X1.X2.X2.X1.X2.vrefh 0.158f
C6374 a_48702_16634# d1 0.0749f
C6375 a_23212_29834# X1.X2.X2.X2.X2.X2.X3.vin1 0.00329f
C6376 X2.X1.X1.X2.X1.X2.X3.vin2 a_33976_10916# 0.00535f
C6377 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.X1.vin1 5.19e-19
C6378 X2.X2.X2.X3.vin1 d2 6.42e-19
C6379 a_48616_18540# a_46502_17540# 5.36e-21
C6380 a_39966_17452# vdd 0.541f
C6381 a_52792_24076# d2 6.04e-19
C6382 a_34062_12822# a_34362_10916# 4.41e-20
C6383 d3 X1.X2.X2.X1.X2.X2.vout 8.47e-19
C6384 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.vrefh 2.33e-19
C6385 d2 a_8572_6962# 0.625f
C6386 X2.X2.X1.X2.vrefh a_46116_19446# 0.118f
C6387 a_54606_26982# a_54992_26982# 0.419f
C6388 a_4696_7064# a_4396_5198# 6.71e-19
C6389 a_4696_22312# a_5082_22312# 0.419f
C6390 a_33676_9010# a_34062_9010# 0.419f
C6391 X1.X2.X2.X2.vrefh X1.X2.X2.X1.X2.X2.X3.vin2 0.161f
C6392 X2.X2.X1.X2.X2.X2.vout d1 0.0331f
C6393 X2.X1.X2.X1.X2.X2.vout d1 0.033f
C6394 X1.X2.X2.X2.X2.X1.vout X1.X2.X2.X2.X3.vin2 0.399f
C6395 X1.X1.X1.X2.X2.X2.X3.vin2 a_2582_4198# 0.567f
C6396 X1.X1.X2.X2.X1.X2.X3.vin1 X1.X1.X2.X2.X1.X1.X3.vin2 1.22e-19
C6397 a_34062_24258# d1 0.0749f
C6398 a_39966_32700# a_38152_31700# 1.15e-20
C6399 X1.X2.X1.X1.X2.X1.vout X1.X2.X1.X1.X2.X2.vout 0.514f
C6400 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X1.vin1 0.0689f
C6401 X1.X1.X2.X1.X2.X1.X3.vin2 a_10686_11734# 7.84e-19
C6402 d4 a_22826_18358# 0.281f
C6403 a_4782_9010# d1 0.0749f
C6404 a_2196_25164# a_2196_27070# 0.00396f
C6405 d1 a_54606_6016# 0.00148f
C6406 a_46502_25164# d1 3.95e-19
C6407 a_39966_30794# X2.X1.X2.X2.X2.X2.vrefh 8.22e-20
C6408 X1.X2.X1.X2.X2.X1.X1.vin2 a_16836_8010# 1.78e-19
C6409 d3 X1.X2.X2.X1.X1.X2.vout 6.06e-19
C6410 X1.X1.X3.vin1 a_5082_10916# 6.09e-19
C6411 a_48316_31882# X2.X2.X1.X1.X1.X1.vout 0.359f
C6412 a_46502_6104# a_46502_4198# 0.00198f
C6413 a_8572_29834# vdd 1.05f
C6414 X1.X2.X2.vrefh X1.X2.X2.X1.X1.X1.X1.vin1 0.142f
C6415 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X3.vin1 1.22e-19
C6416 X1.X1.X1.X2.X2.X1.X3.vin2 a_2196_8010# 0.354f
C6417 a_37766_24076# a_37466_22210# 5.55e-20
C6418 a_16836_9916# X1.X2.X1.X2.X2.X1.X1.vin1 0.195f
C6419 X2.X1.X2.X1.X2.X2.vrefh vdd 0.415f
C6420 a_54606_6016# X2.X2.X2.X1.X1.X1.X3.vin1 0.00207f
C6421 X2.X1.X1.X2.X1.X1.X3.vin2 a_33976_14688# 0.00546f
C6422 d2 X1.X2.X2.X1.X2.X2.X1.vin1 0.0106f
C6423 d2 X2.X2.X1.X2.X2.X2.X3.vin1 0.0577f
C6424 X2.X2.X2.X2.X2.X1.X1.vin1 d1 0.0118f
C6425 a_31862_13728# X2.X1.X1.X2.X1.X2.X1.vin2 0.273f
C6426 a_39966_32700# X2.X1.X2.X2.X2.X2.X3.vin2 0.567f
C6427 a_33976_10916# a_34062_9010# 3.21e-19
C6428 d2 X2.X1.X1.X2.X2.X2.vrefh 0.168f
C6429 a_34362_10916# a_33676_9010# 2.97e-19
C6430 d3 X1.X1.X2.X2.X2.X1.X3.vin2 0.0952f
C6431 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X3.vin1 0.0131f
C6432 X2.X1.X2.X2.X2.X1.X1.vin1 a_40352_26982# 0.195f
C6433 X1.X2.X2.X1.X2.X1.X2.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 0.234f
C6434 a_46116_30882# X2.X2.X1.X1.X1.X1.X1.vin2 1.78e-19
C6435 a_48702_31882# d1 0.0394f
C6436 a_17222_9916# d1 3.95e-19
C6437 X1.X1.X2.X1.X1.X1.X3.vin2 a_8572_6962# 0.00546f
C6438 X1.X2.X1.X1.X2.X2.vout a_19036_20446# 0.36f
C6439 d3 X1.X2.X2.X2.X2.X2.vout 1.05e-19
C6440 a_19722_22312# a_19422_20446# 5.55e-20
C6441 d2 a_31476_9916# 0.00272f
C6442 d0 X2.X1.X1.X2.X1.X2.vrefh 0.848f
C6443 X2.X1.X2.X2.X2.X1.X3.vin2 a_40352_28888# 0.354f
C6444 d2 a_17222_8010# 0.00665f
C6445 X2.X2.X3.vin2 X2.X2.X1.X2.X2.X2.vout 1.5e-19
C6446 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X2.vin1 0.564f
C6447 a_48702_31882# X2.X2.X1.X1.X1.X1.X3.vin1 0.428f
C6448 X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin1 0.00437f
C6449 X1.X1.X2.X2.X2.X1.X1.vin1 d3 6.34e-20
C6450 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X2.vin1 0.242f
C6451 a_52106_29834# a_52792_31700# 3.31e-19
C6452 a_37766_27888# a_37466_25982# 5.25e-20
C6453 a_52106_25982# d2 7.13e-19
C6454 X2.X1.X2.X2.X2.X2.vout d1 0.033f
C6455 a_25326_21264# d1 0.00148f
C6456 a_54606_13640# X2.X2.X2.X1.X2.X1.X1.vin2 8.88e-20
C6457 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 0.0565f
C6458 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X2.vin1 0.0689f
C6459 a_2582_28976# a_4396_28070# 1.06e-19
C6460 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X2.X3.vin1 0.206f
C6461 d2 X2.X2.X2.X1.X3.vin1 0.0619f
C6462 X2.X1.X1.X1.X2.X2.X1.vin2 d2 0.231f
C6463 a_33976_10916# a_34362_10916# 0.414f
C6464 d0 a_17222_15634# 0.0489f
C6465 d0 a_40352_6016# 0.515f
C6466 a_19336_18540# X1.X2.X1.X3.vin2 0.0927f
C6467 d0 X1.X1.X1.X2.X2.vrefh 0.844f
C6468 a_4696_10916# a_2582_9916# 5.36e-21
C6469 X2.X1.X1.X1.X2.X1.X1.vin2 d0 0.276f
C6470 X1.X2.X1.X1.X2.X2.X3.vin1 d2 0.153f
C6471 X2.X2.X1.X1.X1.X1.X3.vin1 d1 0.0296f
C6472 d2 a_37766_31700# 0.00166f
C6473 a_2582_27070# X1.X1.X1.X1.X2.vrefh 0.3f
C6474 a_10686_26982# a_8872_27888# 1.06e-19
C6475 X1.X2.X2.X1.X1.X1.X2.vin1 a_25326_4110# 8.88e-20
C6476 d1 X2.X2.X2.X1.X1.X1.X3.vin1 0.16f
C6477 X1.X2.X2.X1.X1.X1.X3.vin2 X1.X2.X2.X1.X1.X1.X1.vin2 8.93e-19
C6478 d0 X1.X2.X2.X1.X1.X1.X3.vin2 4.34e-19
C6479 X2.X2.X2.X2.X2.X2.X3.vin2 vrefl 0.183f
C6480 X1.X2.X1.X1.X2.X1.X3.vin1 d0 4.36e-19
C6481 X2.X1.X2.X2.X2.X2.vrefh vdd 0.415f
C6482 d2 X1.X2.X2.X2.X2.X2.X1.vin1 9.24e-20
C6483 a_49002_14688# X2.X2.X1.X2.X1.X2.vout 0.254f
C6484 a_37766_16452# a_38152_16452# 0.419f
C6485 a_48316_5198# a_46502_4198# 1.15e-20
C6486 d2 a_48616_14688# 0.526f
C6487 a_2196_27070# vdd 1.05f
C6488 a_54606_19358# d1 3.95e-19
C6489 a_16836_27070# a_16836_28976# 0.00396f
C6490 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X2.X3.vin2 0.0523f
C6491 d2 X2.X2.X1.X2.X2.X2.X3.vin2 8.42e-19
C6492 a_37852_29834# a_37766_31700# 3.38e-19
C6493 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X2.vin1 0.242f
C6494 d4 a_46502_17540# 0.00112f
C6495 a_2196_17540# a_2196_15634# 0.00396f
C6496 X1.X2.X2.X2.X2.X1.X3.vin1 a_25326_28888# 0.00207f
C6497 X1.X1.X1.X1.X1.X2.vout a_4782_28070# 0.418f
C6498 d0 X1.X1.X1.X2.X2.X1.X1.vin2 0.276f
C6499 d6 X2.X3.vin2 0.00878f
C6500 d3 a_48702_9010# 0.00148f
C6501 X2.X1.X1.X1.X1.X2.vrefh d0 0.848f
C6502 X1.X2.X3.vin1 X1.X2.X1.X2.X1.X1.vout 2.91e-19
C6503 d4 a_52106_29834# 0.00116f
C6504 a_23126_27888# d4 2.4e-19
C6505 a_39966_7922# X2.X1.X2.X1.X1.X1.X3.vin2 8.07e-19
C6506 X2.X2.X3.vin2 d1 0.0892f
C6507 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.X1.X1.X1.vin2 3.94e-19
C6508 X1.X1.X2.X2.X2.X1.vout d1 0.0238f
C6509 d3 a_31476_32788# 2.56e-19
C6510 a_31862_25164# X2.X1.X1.X1.X2.X1.X2.vin1 8.88e-20
C6511 X2.X1.X2.X2.X1.X1.X1.vin2 d1 1.49e-19
C6512 a_10686_13640# vdd 0.541f
C6513 a_11072_21264# d0 0.515f
C6514 X2.X2.X1.X2.X1.X1.X3.vin1 a_46502_15634# 0.00207f
C6515 X2.X2.X2.X2.X1.X2.X1.vin2 d2 0.226f
C6516 X2.X2.X2.X2.X1.X1.X1.vin2 X2.X2.X2.X2.X1.X1.X1.vin1 0.668f
C6517 a_2582_27070# a_4696_26164# 4.72e-20
C6518 a_23126_24076# d1 0.0749f
C6519 d2 X2.X1.X1.X2.X2.X2.vout 0.11f
C6520 X1.X2.X2.X1.X1.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin1 0.00437f
C6521 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 2.23e-19
C6522 a_17222_28976# vdd 0.553f
C6523 X2.X1.X1.X2.X2.X2.X3.vin1 X2.X1.X1.X2.X2.X2.X1.vin2 0.22f
C6524 X2.X2.X2.X2.X2.vrefh d3 6.65e-20
C6525 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X1.vin2 0.076f
C6526 d3 X2.X1.X2.X1.X1.X2.vout 6.06e-19
C6527 a_17222_30882# d0 0.0489f
C6528 X1.X1.X2.X2.X1.X2.X1.vin1 d1 0.0118f
C6529 X1.X1.X2.X1.X1.X1.vout a_8872_5016# 0.359f
C6530 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X1.X3.vin1 0.00836f
C6531 d3 X2.X1.X2.X1.X1.X2.X2.vin1 8.68e-20
C6532 a_33676_5198# a_31862_4198# 1.15e-20
C6533 a_52106_6962# X2.X2.X2.X1.X3.vin1 0.436f
C6534 a_37852_25982# a_38152_24076# 6.48e-19
C6535 X2.X1.X2.X2.X1.X1.vout vdd 0.78f
C6536 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X1.vout 0.0215f
C6537 X1.X2.X2.X2.X1.X1.X1.vin2 d1 1.49e-19
C6538 X2.X2.X1.X1.X1.X2.X3.vin2 a_46502_25164# 8.07e-19
C6539 a_25326_21264# X1.X2.X2.X2.X1.X1.X1.vin2 8.88e-20
C6540 a_37466_14586# a_38152_12640# 2.86e-19
C6541 d4 a_52792_16452# 0.00119f
C6542 a_37852_6962# a_38152_5016# 6.1e-19
C6543 d1 X2.X2.X2.X1.X1.X2.vout 0.033f
C6544 d4 a_48616_18540# 0.63f
C6545 a_34362_18540# X2.X1.X1.X2.X1.X1.X3.vin1 0.00837f
C6546 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.X1.X1.X3.vin1 1.22e-19
C6547 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X1.vin2 0.076f
C6548 a_5082_18540# d1 0.0424f
C6549 a_2582_9916# X1.X1.X1.X2.X2.X1.X2.vin1 8.88e-20
C6550 d2 a_52406_8828# 0.00138f
C6551 X2.X3.vin1 a_43362_892# 0.413f
C6552 X1.X1.X1.X2.X1.X2.X3.vin2 a_2582_9916# 8.07e-19
C6553 X1.X2.X2.X2.X3.vin1 a_23126_20264# 1.52e-19
C6554 d0 a_39966_11734# 0.0675f
C6555 a_10686_15546# a_11072_15546# 0.419f
C6556 d3 a_48616_10916# 0.621f
C6557 X1.X1.X1.X2.X1.X1.X1.vin1 d0 0.267f
C6558 d2 a_19036_12822# 6.04e-19
C6559 a_48316_20446# vdd 1.05f
C6560 X2.X2.X2.X3.vin1 a_52492_18358# 0.17f
C6561 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X2.vrefh 2.33e-19
C6562 X1.X1.X2.X2.X1.X1.X1.vin2 d1 1.49e-19
C6563 a_8486_12640# d1 0.0749f
C6564 d2 X2.X1.X2.X1.X1.X2.X1.vin1 0.0114f
C6565 X2.X2.X1.X2.X1.X2.vrefh a_46502_15634# 0.3f
C6566 X2.X2.X2.X2.X2.X1.X3.vin1 a_52106_25982# 0.00837f
C6567 a_25712_25076# d1 2.92e-22
C6568 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 0.049f
C6569 a_33676_28070# d3 0.00108f
C6570 X1.X2.X2.X2.X2.X2.X3.vin2 a_25326_30794# 7.84e-19
C6571 X1.X2.X2.X2.X2.X2.X2.vin1 X1.X2.X2.X2.X2.X2.X1.vin1 0.0689f
C6572 X1.X2.X1.X1.X2.X1.vout vdd 0.805f
C6573 a_19422_5198# a_17222_4198# 4.77e-21
C6574 X1.X2.X1.X2.X2.X2.X3.vin2 a_16836_4198# 0.354f
C6575 X1.X1.X2.X2.X1.X2.X3.vin2 d1 0.171f
C6576 X1.X1.X1.X1.X2.vrefh d1 0.00745f
C6577 d0 X1.X2.X1.X2.X2.X2.X2.vin1 0.262f
C6578 a_25326_15546# a_23212_14586# 2.68e-20
C6579 X1.X2.X1.X2.X2.X2.X3.vin2 X1.X2.X2.vrefh 0.172f
C6580 a_16836_6104# d0 0.518f
C6581 d2 a_31862_6104# 6.36e-19
C6582 X1.X2.X2.X2.X1.X2.X2.vin1 d2 0.0329f
C6583 a_23212_18358# vdd 1.05f
C6584 a_8572_18358# a_10686_17452# 4.72e-20
C6585 d0 X2.X1.X2.X1.X2.X2.X1.vin1 0.267f
C6586 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X2.vrefh 0.00118f
C6587 a_33676_20446# vdd 1.05f
C6588 X2.X2.X1.X1.X1.X2.X3.vin2 d1 0.171f
C6589 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X2.vout 0.0898f
C6590 X1.X1.X2.X1.X1.X2.X1.vin1 X1.X2.X1.X2.X2.X2.vrefh 0.00437f
C6591 a_16836_13728# X1.X2.X1.X2.X1.X2.X1.vin1 0.195f
C6592 d4 a_23126_16452# 8.66e-19
C6593 a_52492_10734# d1 0.0126f
C6594 a_10686_23170# a_11072_23170# 0.419f
C6595 X2.X2.X1.X1.X1.X1.X2.vin1 X2.X2.X1.X1.X1.X1.X1.vin2 0.242f
C6596 a_4396_16634# d1 0.521f
C6597 d3 a_52406_12640# 0.00195f
C6598 a_52792_27888# a_52492_29834# 6.1e-19
C6599 X2.X1.X1.X2.X1.X1.X3.vin2 vdd 0.905f
C6600 a_37766_31700# a_38152_31700# 0.419f
C6601 X1.X1.X3.vin2 a_5082_7064# 5.84e-19
C6602 a_10686_19358# X1.X1.X2.X1.X2.X2.X3.vin2 8.07e-19
C6603 X1.X2.X2.X2.X1.X2.X1.vin1 d0 0.267f
C6604 a_31476_28976# X2.X1.X1.X1.X1.X2.X1.vin2 0.12f
C6605 d0 a_31862_8010# 0.0489f
C6606 d3 a_22826_29834# 2.73e-19
C6607 a_25712_32700# d0 0.515f
C6608 a_19036_20446# vdd 1.05f
C6609 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X1.vin2 0.242f
C6610 a_10686_32700# a_10686_30794# 0.00198f
C6611 X2.X2.X2.X1.X1.X2.vrefh a_54992_6016# 0.118f
C6612 a_25326_28888# X1.X2.X2.X2.X2.X1.X3.vin2 0.567f
C6613 X2.X1.X3.vin1 a_34062_16634# 2.92e-19
C6614 a_10686_7922# a_11072_7922# 0.419f
C6615 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X3.vin1 0.00118f
C6616 a_23212_6962# X1.X2.X2.X1.X1.X1.X3.vin2 0.00546f
C6617 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.vrefh 0.161f
C6618 a_52106_6962# a_52406_8828# 5.55e-20
C6619 a_4696_26164# d1 0.0126f
C6620 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X1.X2.X2.X1.vin2 0.216f
C6621 X1.X2.X1.X1.X3.vin2 d2 0.00194f
C6622 a_46116_9916# vdd 1.05f
C6623 d2 X1.X2.X1.X2.X3.vin2 0.0501f
C6624 a_37766_31700# X2.X1.X2.X2.X2.X2.X3.vin2 0.277f
C6625 X2.X1.X1.X3.vin1 a_34362_22312# 7.98e-19
C6626 a_2582_21352# d2 0.00393f
C6627 X2.X2.X2.X2.vrefh a_54992_17452# 0.118f
C6628 a_25326_26982# d2 0.00328f
C6629 X2.X1.X1.X2.X2.vrefh X2.X1.X1.X2.X2.X1.X1.vin1 0.267f
C6630 X1.X1.X1.X2.X3.vin2 a_4782_5198# 9.7e-20
C6631 a_4696_18540# X1.X1.X3.vin1 0.354f
C6632 a_46502_32788# X2.X2.X1.X1.X1.X1.X1.vin2 0.273f
C6633 X2.X2.X2.X2.X1.X1.vout a_52492_22210# 0.169f
C6634 d2 a_46116_32788# 3.9e-19
C6635 X2.X2.X1.X2.X2.X2.vrefh a_46502_6104# 8.22e-20
C6636 a_2582_25164# d0 0.0675f
C6637 a_34926_892# vdd 1.05f
C6638 a_19336_22312# X1.X2.X1.X1.X2.X2.X3.vin1 0.00329f
C6639 X2.X1.X2.X2.X2.X2.X1.vin1 d0 0.267f
C6640 X2.X2.X1.X1.X2.X2.X1.vin2 vdd 0.36f
C6641 a_34362_29936# d1 0.0422f
C6642 d3 a_19336_18540# 7.7e-20
C6643 a_39966_25076# a_37766_24076# 4.77e-21
C6644 X1.X1.X2.X2.X1.X2.X2.vin1 a_11072_23170# 1.78e-19
C6645 a_34362_14688# X2.X1.X1.X2.X3.vin1 0.436f
C6646 a_4696_14688# X1.X1.X1.X2.X1.X2.X3.vin1 0.00329f
C6647 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X1.vin1 2.23e-19
C6648 X2.X2.X2.X1.X2.X1.vout a_52792_12640# 0.359f
C6649 a_46502_19446# d2 0.00583f
C6650 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X1.vin2 0.668f
C6651 X2.X1.X1.X1.X2.X2.X3.vin1 vdd 0.962f
C6652 d1 a_37466_6962# 0.0422f
C6653 X2.X2.X2.X1.X2.X1.X1.vin2 X2.X2.X2.X1.X2.X1.X1.vin1 0.668f
C6654 d4 a_23126_31700# 2.4e-19
C6655 X1.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X3.vin1 0.546f
C6656 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X3.vin1 0.0131f
C6657 X1.X1.X2.X1.X2.X1.vout a_8572_10734# 1.64e-19
C6658 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X2.vout 0.0866f
C6659 d3 X2.X2.X1.X1.X2.X1.X1.vin2 3.99e-21
C6660 d0 X2.X2.X2.X1.X2.X2.X3.vin2 4.34e-19
C6661 a_4396_31882# d1 0.511f
C6662 a_48616_29936# X2.X2.X1.X1.X1.X2.vout 0.0929f
C6663 X2.X1.X1.X1.X1.X1.X3.vin2 vdd 0.939f
C6664 a_54606_4110# vdd 0.553f
C6665 a_37766_27888# vdd 0.561f
C6666 a_10686_17452# d2 0.00583f
C6667 a_52792_16452# a_52492_14586# 6.71e-19
C6668 d3 X2.X1.X1.X1.X2.X1.X3.vin1 0.0195f
C6669 X2.X2.X3.vin1 X2.X2.X1.X2.X3.vin1 7.18e-19
C6670 a_16836_27070# d0 0.515f
C6671 a_8572_6962# a_8486_5016# 3.14e-19
C6672 d4 X1.X2.X1.X1.X1.X2.vout 1.45e-19
C6673 X1.X2.X2.X3.vin1 d1 0.00955f
C6674 X1.X1.X1.X2.X2.X2.X1.vin2 d1 0.0985f
C6675 a_52492_10734# X2.X2.X2.X1.X1.X2.vout 7.93e-20
C6676 a_31476_19446# d2 0.00441f
C6677 X2.X2.X1.X2.X1.X1.X3.vin1 a_48316_16634# 0.199f
C6678 X2.X2.X1.X1.X2.X1.vout d2 0.00174f
C6679 d0 X2.X2.vrefh 0.0263f
C6680 a_10686_30794# a_11072_30794# 0.419f
C6681 X1.X1.X1.X2.X3.vin2 a_5082_7064# 0.422f
C6682 X2.X2.X1.X1.X2.X2.vout a_48616_18540# 7.93e-20
C6683 a_37766_5016# a_38152_5016# 0.419f
C6684 a_52492_29834# vdd 1.05f
C6685 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X3.vin1 0.0174f
C6686 X1.X2.X2.X1.X1.X1.X2.vin1 a_25712_6016# 0.197f
C6687 X2.X2.X1.X1.X1.X2.vrefh a_46502_30882# 0.3f
C6688 X1.X1.X2.X1.X2.X1.X1.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 5.19e-19
C6689 a_10686_9828# a_8486_8828# 4.77e-21
C6690 X2.X2.X1.X1.X2.X1.X3.vin2 a_49002_22312# 0.00815f
C6691 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X1.vin2 0.668f
C6692 d3 X1.X2.X1.X2.X2.X1.X1.vin2 3.99e-21
C6693 X1.X1.X2.X1.X2.X2.X3.vin2 a_11072_17452# 0.354f
C6694 a_4696_18540# a_4782_16634# 3.21e-19
C6695 a_5082_18540# a_4396_16634# 2.97e-19
C6696 X1.X1.X1.X1.X2.X2.vrefh a_2196_21352# 1.64e-19
C6697 X1.X1.X1.X2.X2.X2.X1.vin1 d2 9.24e-20
C6698 d3 X1.X1.X1.X2.X2.X1.X3.vin1 0.0195f
C6699 X1.X1.X1.X1.X2.X2.vout vdd 0.865f
C6700 a_39966_11734# X2.X1.X2.X1.X2.X1.X1.vin1 0.417f
C6701 X2.X1.X2.X1.X2.X1.X1.vin2 a_40352_11734# 0.12f
C6702 a_16836_19446# d2 0.00441f
C6703 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X3.vin1 0.206f
C6704 X1.X2.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin2 0.1f
C6705 a_31862_23258# a_33976_22312# 2.95e-20
C6706 X1.X2.X3.vin2 a_22826_14586# 3.67e-19
C6707 X2.X1.X1.X2.X1.X1.X1.vin2 X2.X1.X1.X2.X1.X1.X3.vin2 8.93e-19
C6708 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 1.22e-19
C6709 a_25326_4110# vdd 0.553f
C6710 X1.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.vout 0.398f
C6711 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.X3.vin1 0.0174f
C6712 d0 a_28482_892# 1.37e-19
C6713 X1.X1.X2.X2.X1.X2.vrefh a_10686_21264# 0.3f
C6714 a_8872_16452# a_10686_15546# 1.06e-19
C6715 X1.X1.X1.X2.X1.X2.vrefh a_2582_15634# 0.3f
C6716 X2.X2.X2.X2.X1.X2.X3.vin1 a_52792_24076# 0.199f
C6717 X1.X1.X2.X2.X1.X2.vout a_8572_22210# 0.0929f
C6718 X1.X2.X2.X1.X1.X2.X3.vin1 a_25326_7922# 0.52f
C6719 d3 a_8572_25982# 0.621f
C6720 d0 X2.X1.X1.X2.X1.X2.X3.vin2 4.34e-19
C6721 a_54606_13640# d1 0.00148f
C6722 X1.X2.X1.X2.X3.vin1 a_19422_12822# 9.54e-19
C6723 a_19722_14688# X1.X2.X1.X2.X1.X2.X3.vin2 3.85e-19
C6724 d3 X1.X1.X2.X1.X3.vin1 0.0869f
C6725 d3 a_52106_22210# 0.0474f
C6726 d0 a_54992_7922# 0.518f
C6727 a_17222_32788# d2 1.95e-19
C6728 a_2196_19446# d2 0.00441f
C6729 X1.X2.X2.X1.X1.X1.X3.vin1 a_23512_5016# 0.199f
C6730 a_52406_16452# X2.X2.X2.X1.X2.X2.X3.vin1 0.42f
C6731 X1.X2.X2.X1.X1.X2.vout a_23512_8828# 0.36f
C6732 X2.X1.X2.X3.vin1 X2.X1.X3.vin2 1.16f
C6733 a_48616_18540# X2.X2.X1.X2.X1.X1.vout 1.64e-19
C6734 X1.X2.X1.X2.X2.X1.X2.vin1 a_16836_8010# 0.197f
C6735 a_49002_18540# a_48702_16634# 5.25e-20
C6736 a_38152_20264# a_37852_18358# 6.2e-19
C6737 X2.X2.X1.X2.X2.X1.X3.vin2 a_48616_7064# 0.00546f
C6738 a_16836_11822# vdd 1.05f
C6739 a_54606_11734# a_54606_9828# 0.00198f
C6740 d2 X2.X2.X1.X2.X1.X2.X3.vin1 0.155f
C6741 a_17222_6104# X1.X2.X1.X2.X2.X2.X2.vin1 8.88e-20
C6742 d2 a_8872_27888# 0.00251f
C6743 X1.X1.X1.X1.X2.X1.X1.vin2 d2 0.231f
C6744 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.vrefh 0.161f
C6745 X2.X1.X2.X2.X2.X1.X3.vin1 a_39966_26982# 0.52f
C6746 a_37852_14586# X2.X1.X2.X1.X2.X1.X3.vin2 0.00546f
C6747 a_16836_6104# a_17222_6104# 0.419f
C6748 X1.X2.X2.X1.X2.X2.vout X1.X2.X2.X1.X2.X1.vout 0.514f
C6749 a_8486_24076# vdd 0.47f
C6750 X2.X2.X1.X2.X2.X1.X3.vin2 vdd 0.903f
C6751 X2.X1.X2.X1.X2.X2.X1.vin1 a_40352_15546# 0.195f
C6752 a_48616_7064# a_46502_6104# 2.68e-20
C6753 X2.X2.X1.X1.X1.X2.X2.vin1 d2 0.0329f
C6754 X1.X2.X2.X3.vin2 a_23212_25982# 0.355f
C6755 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 5.19e-19
C6756 a_8872_24076# a_10686_23170# 1.06e-19
C6757 X1.X1.X1.X1.X2.X2.vrefh a_2582_23258# 0.3f
C6758 a_22826_25982# d1 0.0316f
C6759 X2.X2.X1.X2.X1.X1.X1.vin1 d1 0.011f
C6760 a_22826_10734# d1 0.0318f
C6761 X1.X2.X2.X1.X2.X2.X1.vin2 vdd 0.36f
C6762 a_46502_6104# vdd 0.553f
C6763 X1.X1.X1.X1.X2.X2.vout X1.X1.X1.X1.X2.X2.X3.vin2 0.08f
C6764 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin2 7.84e-19
C6765 X1.X1.X1.X2.X2.X1.vout a_4696_7064# 0.169f
C6766 X1.X2.X1.X1.X2.X1.X3.vin2 a_17222_23258# 0.567f
C6767 a_4782_9010# a_5082_7064# 4.19e-20
C6768 X2.X1.X2.X2.X1.X2.X2.vin1 vdd 0.576f
C6769 d1 a_4782_5198# 0.0751f
C6770 a_52406_8828# a_52792_8828# 0.419f
C6771 X1.X1.X2.X2.X2.X1.X2.vin1 X1.X2.X1.X1.X1.X2.X1.vin2 0.00232f
C6772 a_16836_28976# a_17222_28976# 0.419f
C6773 a_37766_24076# X2.X1.X2.X2.X1.X2.X3.vin1 0.42f
C6774 d3 a_37466_18358# 0.0469f
C6775 X2.X2.X2.X2.X2.X1.vout d1 0.0238f
C6776 a_2582_6104# X1.X1.X1.X2.X2.X1.X3.vin2 8.07e-19
C6777 X2.X1.X1.X1.X2.X1.X2.vin1 X2.X1.X1.X1.X2.X2.vrefh 0.564f
C6778 X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.vout 1.71e-19
C6779 X1.X2.X2.X2.X2.X1.X3.vin1 d1 0.151f
C6780 d1 X2.X1.X2.X1.X1.X1.X1.vin2 0.0985f
C6781 X1.X1.X2.X1.X2.X2.X3.vin1 a_8186_14586# 0.00874f
C6782 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X2.X1.X2.X2.X2.vrefh 0.0128f
C6783 d0 a_40352_13640# 0.515f
C6784 X2.X2.X3.vin1 a_49952_892# 0.386f
C6785 X2.X2.X1.X1.X2.X2.X3.vin1 a_48702_20446# 0.42f
C6786 X2.X2.X1.X1.X2.X2.X1.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 2.23e-19
C6787 d2 X2.X1.X1.X2.X1.X2.vout 0.00124f
C6788 X2.X2.X1.X2.X2.X1.X1.vin2 a_46116_8010# 1.78e-19
C6789 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X2.vin1 0.564f
C6790 a_19336_14688# d1 0.00613f
C6791 X2.X1.X2.X2.vrefh d1 0.00964f
C6792 X1.X1.X2.X3.vin2 d4 0.535f
C6793 X2.X2.X1.X2.X1.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X1.vin1 5.19e-19
C6794 X1.X2.X1.X1.X3.vin2 a_19336_22312# 0.363f
C6795 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X1.vin2 0.696f
C6796 a_40352_26982# d0 0.518f
C6797 a_8486_8828# X1.X1.X2.X1.X1.X2.X3.vin1 0.42f
C6798 X1.X1.X1.X2.X2.X1.X2.vin1 X1.X1.X1.X2.X2.X2.vrefh 0.564f
C6799 X2.X2.X1.X1.X2.X2.vout d4 6.02e-19
C6800 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.vrefh 0.161f
C6801 X1.X1.X2.X1.X1.X2.X2.vin1 vdd 0.576f
C6802 d0 X1.X2.X2.X1.X2.X1.X3.vin2 4.34e-19
C6803 a_19036_28070# a_19336_26164# 6.48e-19
C6804 X1.X2.X1.X1.X1.X2.X3.vin2 d2 0.122f
C6805 d3 a_23512_12640# 0.00178f
C6806 a_11072_25076# X1.X1.X2.X2.X1.X2.X1.vin2 1.78e-19
C6807 X2.X2.X1.X1.X1.X2.X1.vin2 d0 0.276f
C6808 X2.X2.X2.X2.X3.vin1 a_52406_24076# 9.54e-19
C6809 a_37466_22210# X2.X1.X2.X2.X1.X1.vout 0.387f
C6810 d3 X2.X1.X1.X1.X2.X1.X3.vin2 2.81e-19
C6811 X2.X2.X2.X1.X3.vin2 a_52406_12640# 0.00101f
C6812 X1.X2.X2.X2.X1.X2.X1.vin1 a_25712_23170# 0.195f
C6813 X1.X2.X2.vrefh a_14082_892# 2.22e-19
C6814 X2.X2.X1.X2.X2.X1.X3.vin1 a_48702_9010# 0.428f
C6815 X2.X1.X1.X1.X1.X2.X3.vin1 d0 4.36e-19
C6816 a_10686_28888# a_10686_30794# 0.00198f
C6817 d3 X1.X1.X1.X2.X2.X1.X3.vin2 7.71e-19
C6818 a_25712_32700# X2.vrefh 0.118f
C6819 a_17222_21352# vdd 0.553f
C6820 X2.X1.X2.X3.vin2 a_37466_18358# 0.263f
C6821 a_49002_18540# d1 0.0424f
C6822 d3 X1.X2.X2.X2.X2.X2.X3.vin2 0.0028f
C6823 d1 a_5082_7064# 0.0422f
C6824 X2.X1.X2.X2.X1.X2.X1.vin1 a_39966_21264# 8.22e-20
C6825 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X1.X2.X2.X1.X1.X3.vin2 3.94e-19
C6826 X2.X2.X1.X1.X2.X1.X3.vin2 d1 0.15f
C6827 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.X1.vin2 0.23f
C6828 a_40352_19358# a_40352_17452# 0.00396f
C6829 a_2582_28976# X1.X1.X1.X1.X1.X2.vrefh 8.22e-20
C6830 a_22826_25982# a_23126_24076# 4.41e-20
C6831 a_25326_25076# X1.X2.X2.X2.X1.X2.X1.vin2 8.88e-20
C6832 vrefl vdd 0.418f
C6833 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X3.vin1 0.587f
C6834 a_48616_7064# a_48316_5198# 6.71e-19
C6835 X1.X1.X2.vrefh X1.X2.X2.vrefh 0.0959f
C6836 d0 a_39966_17452# 0.0489f
C6837 X1.X2.X2.X2.X2.X2.X1.vin2 vdd 0.387f
C6838 a_8186_22210# a_8572_22210# 0.419f
C6839 a_8572_18358# X1.X1.X2.X1.X2.X2.vout 7.93e-20
C6840 d1 a_10686_4110# 0.00107f
C6841 X2.X2.X3.vin1 a_52406_5016# 8.66e-20
C6842 a_48316_5198# vdd 1.05f
C6843 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 0.139f
C6844 d3 a_17222_25164# 0.00112f
C6845 a_33976_29936# X2.X1.X1.X1.X3.vin1 0.363f
C6846 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 0.587f
C6847 d3 X2.X2.X1.X1.X1.X1.X3.vin2 0.0678f
C6848 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 0.0565f
C6849 a_10686_15546# X1.X1.X2.X1.X2.X2.vrefh 8.22e-20
C6850 a_8872_31700# a_10686_30794# 1.06e-19
C6851 X2.X2.X2.X2.X1.X1.X3.vin1 a_52792_20264# 0.199f
C6852 X1.X1.X1.X1.X1.X2.vrefh a_2582_30882# 0.3f
C6853 d3 a_4782_28070# 7.51e-19
C6854 a_25326_15546# a_25326_13640# 0.00198f
C6855 d2 X2.X1.X2.X1.X1.X2.vrefh 6.65e-20
C6856 a_19422_16634# X1.X2.X1.X2.X1.X1.vout 0.422f
C6857 d4 X2.X2.X1.X2.X1.X1.vout 0.00145f
C6858 a_48616_26164# a_46502_25164# 5.36e-21
C6859 d4 X2.X1.X1.X3.vin2 0.134f
C6860 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X1.X2.X2.vrefh 0.1f
C6861 a_39966_26982# X2.X1.X2.X2.X1.X2.X3.vin2 8.07e-19
C6862 a_25326_7922# a_25712_7922# 0.419f
C6863 a_10686_25076# a_11072_25076# 0.419f
C6864 X2.X1.X1.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 0.581f
C6865 a_52406_31700# X2.X2.X2.X2.X2.X2.X3.vin1 0.42f
C6866 a_2196_17540# X1.X1.X1.X2.X1.X1.X1.vin2 0.12f
C6867 a_2582_11822# d1 0.00151f
C6868 X1.X2.X2.X2.X3.vin2 vdd 1.29f
C6869 a_40352_11734# vdd 1.05f
C6870 a_2196_25164# X1.X1.X1.X1.X2.X1.X3.vin1 0.354f
C6871 X2.X1.X2.X1.X2.X2.vout a_37466_14586# 0.263f
C6872 a_2582_25164# X1.X1.X1.X1.X2.X1.X1.vin1 0.417f
C6873 a_46502_23258# vdd 0.541f
C6874 a_46502_27070# X2.X2.X1.X1.X1.X2.X3.vin1 0.00207f
C6875 a_33976_7064# vdd 1.05f
C6876 a_52406_24076# a_54606_23170# 4.2e-20
C6877 a_48616_10916# X2.X2.X1.X2.X2.X1.X3.vin1 0.00251f
C6878 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X1.vin2 0.216f
C6879 d0 X2.X1.X2.X1.X2.X2.vrefh 0.848f
C6880 a_8572_10734# a_8486_8828# 3.3e-19
C6881 X1.X1.X1.X2.vrefh d1 0.00964f
C6882 X2.X1.X1.X1.X2.X1.vout d4 3.29e-19
C6883 a_49002_18540# X2.X2.X3.vin2 6.58e-20
C6884 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.vout 0.398f
C6885 X1.X2.X2.X1.X2.X2.X3.vin1 d1 0.146f
C6886 a_33676_24258# a_34362_22312# 2.86e-19
C6887 a_10686_32700# d1 0.00148f
C6888 X2.X1.X2.X2.X2.X2.X1.vin1 a_40352_30794# 0.195f
C6889 a_34062_24258# a_33976_22312# 3.14e-19
C6890 X2.X2.X2.X2.X2.X2.vrefh a_54606_30794# 8.22e-20
C6891 X1.X1.X1.X3.vin2 X1.X1.X2.X1.X3.vin2 7.46e-20
C6892 a_19422_5198# vdd 0.47f
C6893 X1.X1.X2.X3.vin1 a_8186_14586# 7.98e-19
C6894 a_19422_24258# X1.X2.X1.X1.X2.X1.vout 0.422f
C6895 a_11072_15546# d1 2.25e-20
C6896 X1.X2.X1.X2.X2.X2.X1.vin1 vdd 0.592f
C6897 X2.X1.X2.X3.vin1 a_37766_12640# 5.28e-19
C6898 X1.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X2.X3.vin2 0.161f
C6899 d2 X1.X2.X1.X2.X1.X1.X3.vin2 0.169f
C6900 X1.X1.X1.X1.X1.X1.X3.vin1 d2 1.69e-19
C6901 a_48616_26164# d1 0.0126f
C6902 X2.X1.X2.X2.X1.X1.X3.vin1 a_38152_20264# 0.199f
C6903 d3 a_19722_22312# 9.23e-19
C6904 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin2 0.1f
C6905 a_39966_7922# a_37852_6962# 2.68e-20
C6906 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X1.X3.vin1 0.0321f
C6907 a_23126_16452# X1.X2.X2.X1.X3.vin2 9.7e-20
C6908 X1.X2.X1.X2.X1.X2.X1.vin1 d1 0.0118f
C6909 X1.X2.X2.X1.X1.X2.X3.vin1 d1 0.146f
C6910 a_40352_28888# d1 2.92e-22
C6911 d2 a_31862_13728# 0.00479f
C6912 d4 X2.X2.X1.X1.X1.X1.vout 4.78e-20
C6913 a_37466_10734# a_37852_10734# 0.414f
C6914 a_19422_9010# X1.X2.X1.X2.X2.X1.vout 0.422f
C6915 X2.X2.X1.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X1.vin2 3.94e-19
C6916 X2.X1.X1.X2.X2.X2.X3.vin1 a_34062_5198# 0.42f
C6917 d2 X1.X1.X2.X1.X2.X2.vout 0.00117f
C6918 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X3.vin2 2.23e-19
C6919 a_34062_28070# a_33976_26164# 3.3e-19
C6920 X1.X2.X2.X2.X2.X1.X3.vin2 d1 0.15f
C6921 X2.X1.X2.X1.X1.X2.X1.vin2 vdd 0.361f
C6922 a_33676_28070# a_34362_26164# 3.08e-19
C6923 a_11072_7922# d1 2.25e-20
C6924 a_52106_25982# X2.X2.X2.X2.X3.vin2 0.263f
C6925 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin2 7.84e-19
C6926 d2 X1.X2.X1.X2.X2.X1.X3.vin2 0.175f
C6927 d2 X2.X1.X2.X2.X2.X1.X2.vin1 0.0318f
C6928 a_19336_10916# a_19036_9010# 6.2e-19
C6929 a_25712_28888# a_25712_30794# 0.00396f
C6930 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X2.vrefh 2.33e-19
C6931 a_33676_9010# a_33976_7064# 6.1e-19
C6932 X2.X1.X2.X2.X2.X2.vrefh d0 0.848f
C6933 X2.X2.X1.X1.X1.X2.vout X2.X2.X1.X1.X1.X2.X3.vin1 0.326f
C6934 a_31476_17540# d1 2.25e-20
C6935 a_37466_14586# d1 0.0422f
C6936 a_25712_6016# vdd 1.05f
C6937 X1.X1.X1.X2.X1.X2.X2.vin1 vdd 0.576f
C6938 X2.X1.X1.X2.X3.vin1 a_34362_10916# 0.372f
C6939 X2.X2.X2.X1.X2.X1.X1.vin1 d1 0.0118f
C6940 X1.X2.X1.X1.X2.X1.X1.vin2 vdd 0.36f
C6941 a_2196_27070# d0 0.515f
C6942 d2 a_40352_17452# 0.00441f
C6943 X1.X1.X2.X2.X3.vin1 a_8572_25982# 0.17f
C6944 a_46502_11822# a_48616_10916# 4.72e-20
C6945 a_46116_27070# vdd 1.05f
C6946 X1.X2.X2.X2.X2.X2.X3.vin1 d1 0.147f
C6947 a_33976_22312# d1 0.00613f
C6948 a_19422_20446# X1.X2.X3.vin1 1.64e-19
C6949 X1.X2.X1.X1.X2.X2.X3.vin2 a_19722_18540# 0.00846f
C6950 X2.X2.X1.X1.X2.X2.X1.vin2 X2.X2.X1.X1.X2.X2.X2.vin1 0.242f
C6951 X1.X1.X2.X2.X2.X1.X3.vin1 vdd 0.997f
C6952 a_16836_27070# a_17222_27070# 0.419f
C6953 d2 X1.X2.X2.X1.X2.X2.X3.vin2 0.113f
C6954 a_8186_14586# X1.X1.X2.X1.X2.X1.X3.vin2 0.00815f
C6955 X1.X1.X1.X1.X2.X1.X3.vin1 vdd 0.997f
C6956 a_23212_18358# a_23512_16452# 6.48e-19
C6957 a_11072_30794# d1 2.25e-20
C6958 d2 X1.X2.X1.X1.X1.X1.X3.vin2 0.0661f
C6959 X1.X2.X2.X2.X1.X1.X3.vin1 a_23512_20264# 0.199f
C6960 X2.X2.X1.X1.X2.X2.vrefh a_46116_21352# 1.64e-19
C6961 X1.X1.X2.X1.X1.X2.X3.vin2 a_8186_6962# 3.85e-19
C6962 d1 a_33676_5198# 0.522f
C6963 d3 X1.X1.X1.X3.vin2 0.482f
C6964 a_8872_20264# a_8572_18358# 6.2e-19
C6965 a_40352_15546# a_40352_13640# 0.00396f
C6966 a_54606_15546# d1 3.41e-19
C6967 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X2.vin1 0.242f
C6968 X2.X2.X2.X2.X1.X1.X1.vin1 d4 6.34e-20
C6969 d0 a_10686_13640# 0.0489f
C6970 X1.X2.X2.X2.X2.vrefh vdd 0.426f
C6971 a_13696_892# X1.X3.vin2 0.0927f
C6972 d3 X1.X1.X2.X1.X2.X1.X1.vin1 6.34e-20
C6973 a_2196_25164# a_2196_23258# 0.00396f
C6974 d2 X1.X1.X1.X2.X3.vin1 0.0014f
C6975 a_10686_30794# X1.X1.X2.X2.X2.X2.vrefh 8.22e-20
C6976 X2.X1.X2.X2.X1.X1.X3.vin2 a_38152_20264# 0.1f
C6977 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X2.vrefh 0.076f
C6978 a_19422_31882# X1.X2.X1.X1.X1.X1.vout 0.422f
C6979 d2 X1.X1.X2.X2.X2.X2.vout 0.102f
C6980 a_17222_28976# d0 0.0675f
C6981 a_19336_29936# a_17222_30882# 2.95e-20
C6982 a_31862_21352# a_34062_20446# 4.2e-20
C6983 d5 X1.X3.vin1 0.0932f
C6984 X2.X1.X1.X1.X2.X2.X3.vin1 X2.X1.X1.X1.X2.X2.X2.vin1 0.00117f
C6985 a_19336_10916# vdd 1.05f
C6986 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.vout 0.038f
C6987 a_52492_22210# vdd 1.05f
C6988 d1 a_46116_8010# 2.92e-22
C6989 X2.X1.X2.X2.X1.X2.X1.vin2 d1 0.00406f
C6990 X2.X2.X2.X2.X1.X1.X3.vin1 a_54992_19358# 0.354f
C6991 a_31862_19446# X2.X1.X1.X2.X1.X1.X1.vin1 8.22e-20
C6992 a_39966_19358# d4 0.00112f
C6993 X1.X2.X2.X3.vin1 a_22826_10734# 0.509f
C6994 a_48316_12822# X2.X2.X1.X2.X1.X2.X3.vin2 0.101f
C6995 X1.X2.X3.vin2 X1.X2.X1.X2.X3.vin2 0.00254f
C6996 d3 X2.X1.X2.X1.X2.X1.X3.vin2 2.81e-19
C6997 X2.X1.X2.X1.X2.X2.X3.vin2 a_39966_15546# 7.84e-19
C6998 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X1.vin1 0.0689f
C6999 X1.X2.X2.X2.X1.X2.X3.vin1 a_23212_22210# 0.00329f
C7000 d3 a_52492_25982# 0.621f
C7001 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X1.vin2 0.216f
C7002 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X2.vrefh 0.267f
C7003 a_4782_24258# d1 0.0749f
C7004 a_2196_11822# a_2196_9916# 0.00396f
C7005 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X1.X3.vin1 0.0131f
C7006 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X2.vrefh 0.00118f
C7007 X1.X2.X2.X2.X1.X1.X3.vin2 X1.X2.X2.X2.X1.X1.X3.vin1 0.581f
C7008 X2.X1.X1.X2.X1.X1.X2.vin1 d1 1.03e-19
C7009 d3 X2.X2.X1.X1.X1.X2.X3.vin1 0.0105f
C7010 a_25326_19358# d4 0.00112f
C7011 X2.X2.X2.X1.X1.X2.X2.vin1 d1 1.03e-19
C7012 a_34362_26164# X2.X1.X1.X1.X2.X1.X3.vin1 0.00837f
C7013 a_54606_30794# d1 3.41e-19
C7014 d1 X2.X1.X2.X1.X1.X2.X3.vin1 0.146f
C7015 d4 X1.X1.X3.vin1 0.287f
C7016 X1.X1.X1.X2.X1.X2.X1.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 2.23e-19
C7017 X1.X1.X1.X2.X1.X2.X3.vin1 a_4782_12822# 0.42f
C7018 a_28482_892# vout 0.399f
C7019 X1.X2.X1.X2.X2.X1.X3.vin2 X1.X2.X1.X2.X2.X2.X1.vin2 3.94e-19
C7020 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X1.X2.X1.vin2 0.076f
C7021 a_48702_28070# a_49002_26164# 4.41e-20
C7022 X2.X1.X3.vin2 vdd 0.834f
C7023 d1 a_25712_7922# 2.25e-20
C7024 X2.X2.X1.X1.X1.X2.X3.vin2 a_48616_26164# 0.00535f
C7025 a_48316_24258# vdd 1.05f
C7026 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X2.X1.X1.X1.vin1 0.206f
C7027 X2.X1.X2.X2.X1.X1.X3.vin2 a_40352_21264# 0.354f
C7028 X2.X2.X1.X1.X1.X2.X2.vin1 X2.X2.X1.X1.X1.X2.X1.vin1 0.0689f
C7029 a_48316_28070# a_46502_28976# 1.06e-19
C7030 a_40352_15546# X2.X1.X2.X1.X2.X2.vrefh 1.64e-19
C7031 X1.X2.X1.X2.X1.X1.X1.vin2 a_17222_15634# 8.88e-20
C7032 d3 X2.X2.X2.X1.X2.vrefh 6.65e-20
C7033 d2 X2.X1.X1.X2.X2.X1.X3.vin2 0.175f
C7034 a_10686_19358# d4 0.00112f
C7035 a_8872_20264# d2 3.82e-19
C7036 a_2196_23258# vdd 1.05f
C7037 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X3.vin1 0.206f
C7038 a_2196_6104# vdd 1.05f
C7039 X1.X1.X1.X1.X2.X2.X1.vin1 X1.X1.X1.X1.X2.X2.X2.vin1 0.0689f
C7040 X2.X1.X3.vin1 a_37466_18358# 5.87e-20
C7041 a_2582_21352# a_4396_20446# 1.06e-19
C7042 a_54606_7922# X2.X2.X2.X1.X1.X2.vrefh 8.22e-20
C7043 a_8872_16452# d1 0.521f
C7044 a_31476_27070# d1 2.92e-22
C7045 d2 X1.X1.X2.X1.X2.X2.X1.vin2 0.231f
C7046 a_16836_32788# X1.X2.X1.X1.X1.X1.X2.vin1 1.78e-19
C7047 d3 X2.X1.X1.X1.X1.X2.vout 6.83e-19
C7048 d0 X2.X1.X1.X2.X1.X1.X3.vin2 4.34e-19
C7049 a_52106_22210# X2.X2.X2.X2.X1.X1.X3.vin2 0.00815f
C7050 a_10686_6016# X1.X1.X2.X1.X1.X1.X1.vin2 8.88e-20
C7051 a_54606_25076# a_52792_24076# 1.15e-20
C7052 X2.X2.X2.X1.X2.X2.X2.vin1 a_54992_17452# 0.197f
C7053 X2.X1.X1.X2.X2.X2.X1.vin2 X2.X1.X1.X2.X2.X2.X2.vin1 0.242f
C7054 a_2196_13728# d1 2.25e-20
C7055 X1.X1.X3.vin2 X1.X3.vin1 0.238f
C7056 X2.X2.X2.X3.vin2 d4 1.03f
C7057 X2.X1.X1.X1.X1.X1.X2.vin1 d1 0.0144f
C7058 a_54992_21264# a_54992_19358# 0.00396f
C7059 X1.X2.X2.X1.X2.X1.X3.vin1 X1.X2.X2.X1.X2.X1.X1.vin1 0.206f
C7060 X2.X2.X2.X1.X1.X1.X1.vin2 a_54606_4110# 0.273f
C7061 d2 a_11072_13640# 0.00464f
C7062 X2.X1.X1.X3.vin1 d2 6.42e-19
C7063 a_46502_17540# X2.X2.X1.X2.X1.X1.X3.vin1 0.52f
C7064 X2.X2.X1.X2.X3.vin2 a_48702_5198# 9.7e-20
C7065 d2 a_37466_10734# 7.13e-19
C7066 a_10686_28888# d1 0.00148f
C7067 d0 a_46116_9916# 0.518f
C7068 d4 a_4782_16634# 0.00142f
C7069 d2 X1.X2.X1.X1.X1.X2.X1.vin2 0.226f
C7070 d2 X1.X1.X2.X1.X1.X2.X1.vin2 0.226f
C7071 X1.X2.X1.X1.X1.X2.X1.vin1 a_17222_30882# 8.22e-20
C7072 X1.X1.X1.X1.X1.X1.X1.vin2 a_4782_31882# 0.00743f
C7073 d3 a_33676_12822# 0.00108f
C7074 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X2.vrefh 0.267f
C7075 X1.X2.X2.X2.X1.X1.X3.vin1 X1.X2.X2.X2.X1.X1.X1.vin1 0.206f
C7076 X2.X1.X2.X1.X3.vin2 a_37852_14586# 0.363f
C7077 X2.X2.X1.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin2 0.1f
C7078 a_8572_29834# a_8486_27888# 3.14e-19
C7079 a_4396_5198# X1.X1.X1.X2.X2.X2.X3.vin2 0.101f
C7080 a_46502_13728# vdd 0.553f
C7081 X1.X2.X2.X1.X2.vrefh a_25326_9828# 0.3f
C7082 d2 X1.X1.X1.X1.X1.X2.X3.vin1 0.158f
C7083 d0 a_34926_892# 2.73e-19
C7084 X1.X2.X2.X2.X2.X1.X3.vin1 a_22826_25982# 0.00837f
C7085 a_31862_13728# a_31862_11822# 0.00198f
C7086 a_31862_25164# a_31862_23258# 0.00198f
C7087 X2.X2.X1.X1.X2.X2.X1.vin2 d0 0.276f
C7088 X1.X1.X2.X2.X2.X1.X1.vin2 d1 4.01e-19
C7089 X2.X1.X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X3.vin1 0.581f
C7090 X1.X2.X1.X2.X1.X2.vout a_19336_10916# 7.93e-20
C7091 X2.X2.X1.X2.X1.X2.X3.vin2 d1 0.171f
C7092 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X2.vrefh 0.00118f
C7093 X2.X2.X2.X2.X1.X2.X2.vin1 a_54992_25076# 0.197f
C7094 a_5082_26164# d4 6.91e-19
C7095 X1.X1.X1.X2.X1.X2.vout d1 0.033f
C7096 X2.X1.X2.X2.X1.X1.X3.vin2 X2.X1.X2.X2.X1.X1.X1.vin1 2.23e-19
C7097 X2.X1.X2.X2.X1.X2.vrefh a_39966_21264# 0.3f
C7098 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X3.vin1 0.0131f
C7099 X2.X1.X2.X2.X1.X1.X2.vin1 a_40352_19358# 1.78e-19
C7100 a_52792_20264# d1 0.521f
C7101 X2.X1.X1.X1.X2.X2.X3.vin1 d0 4.36e-19
C7102 X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin1 0.00437f
C7103 a_54606_6016# X2.X2.X2.X1.X1.X1.X3.vin2 0.567f
C7104 X2.X2.X2.X2.X2.X1.X2.vin1 vdd 0.576f
C7105 a_8872_31700# d1 0.515f
C7106 a_13696_892# vdd 1.05f
C7107 X1.X1.X2.X1.X2.X2.X3.vin1 vdd 0.962f
C7108 X1.X2.X1.X1.X1.X2.X2.vin1 a_16836_27070# 0.197f
C7109 a_46502_25164# X2.X2.X1.X1.X2.X1.X3.vin1 0.52f
C7110 d2 X1.X1.X2.X2.X2.X2.X1.vin2 7.2e-20
C7111 X2.X1.X1.X1.X1.X1.X3.vin2 d0 4.34e-19
C7112 d0 a_54606_4110# 0.0675f
C7113 a_54992_17452# vdd 1.05f
C7114 d4 X2.X1.X1.X1.X3.vin1 0.0378f
C7115 X2.X1.X2.X1.X1.X2.X2.vin1 a_40352_7922# 1.78e-19
C7116 X2.X1.X2.vrefh a_40352_4110# 9.79e-19
C7117 a_31862_15634# X2.X1.X1.X2.X1.X2.X1.vin1 8.22e-20
C7118 X2.X1.X2.X1.X1.X2.X3.vin2 X2.X1.X2.X1.X1.X2.X1.vin1 2.23e-19
C7119 X1.X2.X3.vin2 X3.vin1 0.00523f
C7120 a_6032_892# X1.X3.vin1 0.461f
C7121 X1.X2.X1.X2.X1.X2.vrefh a_16836_15634# 0.118f
C7122 d2 a_46502_15634# 0.0059f
C7123 a_38152_20264# d1 0.521f
C7124 a_48616_18540# X2.X2.X1.X2.X1.X1.X3.vin1 0.00232f
C7125 a_23512_27888# a_23212_29834# 6.1e-19
C7126 X2.X2.X1.X1.X2.X2.vrefh d2 0.168f
C7127 X2.X1.X2.X1.X2.X2.X3.vin2 vdd 0.761f
C7128 d2 a_19722_7064# 0.254f
C7129 d3 a_11072_32700# 2.56e-19
C7130 a_52792_20264# a_54606_19358# 1.06e-19
C7131 X2.X2.X2.X2.X1.X2.vrefh X2.X2.X2.X2.X1.X1.X1.vin2 0.076f
C7132 X2.X2.X2.X2.X1.X2.vout a_52492_22210# 0.0929f
C7133 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X2.vrefh 0.1f
C7134 a_25326_7922# X1.X2.X2.X1.X1.X2.vrefh 8.22e-20
C7135 d3 a_4782_20446# 4.67e-19
C7136 X1.X1.X1.X2.X2.X2.vout a_4396_5198# 0.36f
C7137 d4 a_4782_31882# 2.4e-19
C7138 a_5082_7064# a_4782_5198# 5.55e-20
C7139 a_5082_22312# X1.X1.X1.X1.X2.X2.vout 0.263f
C7140 a_10686_6016# X1.X1.X2.X1.X1.X2.X1.vin1 8.22e-20
C7141 a_19336_29936# a_19422_31882# 3.14e-19
C7142 a_19722_29936# a_19036_31882# 2.86e-19
C7143 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.X1.vin2 3.94e-19
C7144 a_34062_9010# X2.X1.X1.X2.X2.X1.vout 0.422f
C7145 X1.X1.X1.X1.X2.X2.X2.vin1 a_2582_19446# 0.402f
C7146 a_34362_26164# X2.X1.X1.X1.X2.X1.X3.vin2 3.49e-19
C7147 d2 a_25326_11734# 0.00328f
C7148 a_22826_22210# vdd 0.477f
C7149 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X2.vrefh 0.076f
C7150 X2.X1.X1.X1.X3.vin2 a_34062_24258# 0.00101f
C7151 a_31476_23258# d2 0.00464f
C7152 a_19036_28070# vdd 1.05f
C7153 d1 X2.X2.X1.X2.X2.X1.X2.vin1 1.03e-19
C7154 a_25326_21264# a_23512_20264# 1.15e-20
C7155 d1 X2.X2.X2.X1.X1.X1.X3.vin2 0.154f
C7156 a_23512_20264# d1 0.521f
C7157 a_39966_26982# d3 0.00112f
C7158 X1.X1.X1.X1.X2.X1.X1.vin1 a_2196_27070# 1.64e-19
C7159 X1.X1.X1.X3.vin1 X1.X1.X3.vin2 7.53e-21
C7160 a_40352_30794# X2.X1.X2.X2.X2.X2.vrefh 1.64e-19
C7161 X2.X2.X1.X1.X2.X1.X3.vin1 d1 0.151f
C7162 X1.X2.X2.X1.X1.X2.X2.vin1 a_25712_9828# 0.197f
C7163 X1.X1.X2.X2.X3.vin2 X1.X1.X2.X2.X2.X2.vout 0.0866f
C7164 X1.X2.X2.X1.X1.X1.X1.vin2 a_25326_4110# 0.273f
C7165 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X3.vin1 0.00836f
C7166 a_17222_21352# X1.X2.X1.X1.X2.X2.X2.vin1 8.88e-20
C7167 d0 a_25326_4110# 0.0675f
C7168 a_5082_26164# a_4396_24258# 2.97e-19
C7169 a_19722_29936# vdd 0.477f
C7170 X1.X1.X2.X2.X2.X2.X3.vin1 vdd 0.993f
C7171 X2.X2.X1.X2.X2.X2.X3.vin1 a_46502_4198# 0.00207f
C7172 a_4696_26164# a_4782_24258# 3.21e-19
C7173 X1.X1.X2.X1.X2.X2.vrefh d1 0.0124f
C7174 a_17222_9916# X1.X2.X1.X2.X2.X1.X3.vin1 0.52f
C7175 d3 X1.X2.X2.X3.vin2 0.481f
C7176 X2.X1.X1.X1.X2.vrefh a_31476_25164# 1.64e-19
C7177 d3 a_23212_10734# 0.621f
C7178 X2.X2.X2.X1.X1.X1.X3.vin2 X2.X2.X2.X1.X1.X1.X3.vin1 0.581f
C7179 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X1.vin2 0.216f
C7180 X2.X1.X1.X2.X1.X1.vout X2.X1.X1.X2.X1.X2.vout 0.507f
C7181 X1.X1.X1.X2.X1.X2.X1.vin2 X1.X1.X1.X2.X1.X2.X2.vin1 0.242f
C7182 X1.X2.X2.X1.X2.X1.vout a_23512_12640# 0.359f
C7183 X2.X1.X1.X2.X2.X1.X1.vin2 d1 4.01e-19
C7184 X2.X2.X1.X2.X1.X1.X3.vin2 a_46116_15634# 0.354f
C7185 X2.X1.X1.X2.X3.vin2 a_34062_9010# 0.00101f
C7186 a_37766_12640# vdd 0.561f
C7187 a_48616_18540# X2.X2.X3.vin1 0.354f
C7188 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X2.X1.X1.X1.X2.X2.vin1 0.00232f
C7189 d2 a_46502_30882# 4.64e-19
C7190 X2.X1.X1.X2.vrefh a_31476_19446# 0.118f
C7191 X1.X2.X1.X2.X2.X1.X3.vin1 d1 0.151f
C7192 a_4696_7064# X1.X1.X1.X2.X2.X2.vout 0.0929f
C7193 X1.X1.X1.X3.vin2 a_5082_14688# 0.00292f
C7194 X1.X2.X1.X1.X1.X1.X1.vin2 d4 8.21e-20
C7195 d0 a_16836_11822# 0.515f
C7196 X1.X2.X1.X1.X2.X2.vout X1.X2.X1.X1.X2.X2.X3.vin2 0.08f
C7197 d2 X2.X1.X1.X2.X2.X1.X1.vin1 0.0105f
C7198 a_40352_21264# d1 2.92e-22
C7199 a_31476_21352# X2.X1.X1.X1.X2.X2.X1.vin2 0.12f
C7200 d2 X1.X2.X2.X1.X1.X2.X1.vin2 0.226f
C7201 d0 X2.X2.X1.X2.X2.X1.X3.vin2 4.34e-19
C7202 X1.X1.X2.X3.vin1 vdd 1.26f
C7203 X2.X2.X2.X1.X2.X1.X2.vin1 a_54606_11734# 8.88e-20
C7204 a_54606_25076# X2.X2.X2.X2.X1.X2.X1.vin2 8.88e-20
C7205 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 0.049f
C7206 X2.X1.X1.X1.X3.vin2 d1 0.00807f
C7207 a_25712_28888# X1.X2.X2.X2.X2.X2.vrefh 0.118f
C7208 X2.X2.X2.X1.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X1.vin2 8.93e-19
C7209 a_25326_21264# X1.X2.X2.X2.X1.X1.X3.vin2 0.567f
C7210 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X3.vin1 0.00789f
C7211 X1.X2.X2.X2.X1.X1.X3.vin2 d1 0.15f
C7212 X2.X2.X2.X2.X3.vin1 a_52106_22210# 0.436f
C7213 a_2582_28976# X1.X1.X1.X1.X1.X2.X3.vin2 7.84e-19
C7214 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X1.X3.vin2 0.0523f
C7215 X1.X1.X1.X2.X2.X1.X1.vin2 a_2196_8010# 1.78e-19
C7216 X1.X1.X2.X1.X1.X1.X1.vin2 X1.X1.X2.X1.X1.X1.X1.vin1 0.668f
C7217 X1.X1.X1.X1.X1.X2.X3.vin1 a_4396_28070# 0.199f
C7218 X2.X1.X2.X2.X1.X1.X2.vin1 d2 0.031f
C7219 X1.X1.X2.X1.X1.X2.vout a_8186_6962# 0.254f
C7220 X1.X2.X2.X1.X3.vin1 a_23126_8828# 9.54e-19
C7221 a_34362_10916# X2.X1.X1.X2.X3.vin2 0.263f
C7222 a_4696_10916# X1.X1.X1.X2.X2.X1.X3.vin1 0.00251f
C7223 d0 a_46502_6104# 0.0675f
C7224 X2.X1.X2.X3.vin1 a_37766_16452# 5.31e-19
C7225 X1.X2.X3.vin1 X1.X2.X1.X3.vin2 1.04f
C7226 d0 X1.X2.X2.X1.X2.X2.X1.vin2 0.276f
C7227 X2.X1.X2.X1.X1.X2.X3.vin1 a_37466_6962# 0.00874f
C7228 X2.X1.X2.X2.X1.X2.X2.vin1 d0 0.262f
C7229 a_22826_25982# X1.X2.X2.X2.X2.X1.X3.vin2 3.49e-19
C7230 X1.X2.X1.X2.X2.vrefh a_16836_11822# 0.118f
C7231 a_40352_11734# a_40352_9828# 0.00396f
C7232 X1.X1.X2.X2.X2.X1.X1.vin1 a_10686_25076# 8.22e-20
C7233 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X1.X2.X3.vin2 3.94e-19
C7234 d3 X2.X2.X1.X3.vin2 0.483f
C7235 X1.X2.X2.X1.X1.X1.X2.vin1 a_25712_4110# 1.78e-19
C7236 X1.X2.vrefh X1.X1.X2.X2.X2.X2.X3.vin1 0.00118f
C7237 X1.X2.X2.X1.X1.X1.X3.vin2 X1.X2.X2.X1.X1.X1.X1.vin1 2.23e-19
C7238 d3 X1.X1.X1.X1.X3.vin1 0.088f
C7239 X1.X1.X2.X2.X2.X2.vrefh d1 0.0124f
C7240 a_54606_15546# a_54606_13640# 0.00198f
C7241 a_39966_17452# X2.X1.X2.X1.X2.X2.X2.vin1 0.402f
C7242 X1.X2.X2.X2.X3.vin1 d4 8.41e-19
C7243 a_2582_32788# X1.X1.X1.X1.X1.X1.X3.vin2 7.84e-19
C7244 d2 X2.X2.X1.X2.X3.vin1 0.0014f
C7245 X2.X2.X1.X2.X2.X2.X3.vin2 a_46502_4198# 0.567f
C7246 X1.X1.X2.X2.X1.X1.X3.vin1 vdd 0.997f
C7247 d4 X2.X2.X1.X2.X1.X1.X3.vin1 0.0205f
C7248 a_54992_19358# d1 2.25e-20
C7249 a_17222_27070# a_17222_28976# 0.00198f
C7250 X1.X2.X1.X2.vrefh a_16836_19446# 0.118f
C7251 a_2582_32788# vdd 0.554f
C7252 X1.X2.X2.X2.X3.vin1 a_23212_22210# 0.363f
C7253 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X1.vout 0.0524f
C7254 d2 a_5082_10916# 7.13e-19
C7255 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X3.vin1 0.00118f
C7256 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.X1.X3.vin2 0.581f
C7257 a_48616_22312# d2 0.526f
C7258 a_2582_17540# a_2582_15634# 0.00198f
C7259 X1.X2.X1.X1.X1.X2.vrefh a_16836_30882# 0.118f
C7260 X1.X1.X1.X2.X1.X1.X3.vin2 a_4696_14688# 0.00546f
C7261 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X1.vout 0.0215f
C7262 d0 X1.X1.X2.X1.X1.X2.X2.vin1 0.262f
C7263 a_39966_13640# a_38152_12640# 1.15e-20
C7264 a_25712_13640# vdd 1.05f
C7265 a_40352_21264# X2.X1.X2.X2.X1.X1.X1.vin2 1.78e-19
C7266 a_33976_29936# a_33676_31882# 6.1e-19
C7267 X2.X2.X1.X2.X1.X2.vout a_48316_12822# 0.36f
C7268 X1.X2.X1.X3.vin1 X1.X2.X2.X2.X3.vin2 7.46e-20
C7269 a_31862_13728# X2.X1.X1.X2.X1.X2.X2.vin1 8.88e-20
C7270 X1.X2.X2.X1.X2.X1.vout a_23212_14586# 0.169f
C7271 a_31862_25164# a_34062_24258# 4.2e-20
C7272 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X2.vin1 0.00117f
C7273 X1.X1.X2.X1.X2.X1.X3.vin2 vdd 0.903f
C7274 X2.X1.X2.X2.X1.X1.X1.vin1 d1 0.011f
C7275 d3 X2.X1.X1.X1.X1.X1.X1.vin1 0.00492f
C7276 a_46116_6104# a_46502_6104# 0.419f
C7277 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X2.X1.X2.X2.X2.X1.vin2 0.00232f
C7278 d2 X2.X2.X1.X2.X1.X2.X2.vin1 0.0329f
C7279 a_17222_21352# d0 0.0675f
C7280 X2.X1.X1.X1.X1.X2.X1.vin2 vdd 0.361f
C7281 a_54606_19358# a_54992_19358# 0.419f
C7282 X2.X2.X2.X2.X1.X2.X1.vin1 d2 0.0114f
C7283 d0 vrefl 0.0261f
C7284 a_39966_25076# X2.X1.X2.X2.X1.X2.X2.vin1 0.402f
C7285 a_40352_9828# X2.X1.X2.X1.X1.X2.X1.vin2 1.78e-19
C7286 X1.X2.X1.X1.X1.X2.X3.vin1 vdd 0.96f
C7287 a_23212_29834# X1.X2.X2.X2.X2.X2.vout 0.0929f
C7288 X1.X2.X2.X2.X2.X2.X1.vin2 d0 0.253f
C7289 d1 X1.X3.vin1 0.0299f
C7290 X2.X1.X1.X2.X2.X2.X3.vin2 a_31862_4198# 0.567f
C7291 a_8186_25982# vdd 0.487f
C7292 X2.X2.X1.X2.X1.X1.X3.vin2 a_49002_14688# 0.00815f
C7293 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 0.242f
C7294 a_39966_32700# a_39966_30794# 0.00198f
C7295 a_25326_17452# vdd 0.541f
C7296 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.X1.X3.vin1 1.22e-19
C7297 X1.X2.X2.X2.X1.X1.X2.vin1 a_25326_19358# 8.88e-20
C7298 X1.X2.X2.X2.X1.X1.X1.vin1 d1 0.011f
C7299 X1.X2.X2.X2.X1.X1.X3.vin2 X1.X2.X2.X2.X1.X1.X1.vin2 8.93e-19
C7300 X1.X2.X2.X2.vrefh a_25712_17452# 0.118f
C7301 d4 X2.X2.X3.vin1 0.286f
C7302 d2 a_48316_16634# 3.82e-19
C7303 X1.X2.X2.X2.vrefh d4 6.65e-20
C7304 X1.X2.X2.X1.X2.X1.X3.vin1 d1 0.151f
C7305 X2.X2.X1.X1.X1.X1.X3.vin2 a_46116_30882# 0.354f
C7306 a_2582_9916# a_4782_9010# 4.2e-20
C7307 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X2.vin1 0.00117f
C7308 X1.X2.X3.vin1 a_19722_10916# 6.09e-19
C7309 X2.X1.X2.X2.X2.X1.vout vdd 0.775f
C7310 X1.X2.X3.vin2 X1.X2.X2.X1.X2.X2.X3.vin2 0.0011f
C7311 a_54992_28888# a_54992_30794# 0.00396f
C7312 a_8572_25982# X1.X1.X2.X2.X1.X2.vout 7.93e-20
C7313 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X3.vin1 1.22e-19
C7314 a_52406_20264# a_52492_18358# 3.21e-19
C7315 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 0.0565f
C7316 a_4696_14688# vdd 1.05f
C7317 d0 a_40352_11734# 0.518f
C7318 d1 X1.X2.X2.X1.X1.X2.vrefh 0.0738f
C7319 d2 X1.X2.X1.X2.X1.X2.X3.vin2 0.121f
C7320 a_8572_29834# a_8486_31700# 3.38e-19
C7321 a_46502_23258# d0 0.0489f
C7322 X2.X2.X1.X1.X2.X2.X3.vin2 vdd 0.761f
C7323 d3 X2.X2.X1.X2.X3.vin2 0.156f
C7324 d1 a_39966_6016# 0.00148f
C7325 X1.X1.X2.X2.X1.X1.X1.vin1 d1 0.011f
C7326 a_33676_24258# d2 3.82e-19
C7327 X1.X2.X1.X2.X1.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X1.vin2 3.94e-19
C7328 a_31862_25164# d1 3.95e-19
C7329 X1.X1.X2.X2.vrefh d4 6.65e-20
C7330 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X1.X2.X2.X1.X1.X1.vin1 0.668f
C7331 d2 X2.X2.X1.X2.X2.X2.X1.vin2 7.2e-20
C7332 a_54606_6016# a_52792_5016# 1.15e-20
C7333 X2.X1.X1.X1.X1.X2.X3.vin2 d3 0.0251f
C7334 X1.X2.X2.X1.X3.vin2 a_23126_12640# 0.00101f
C7335 d2 a_4396_9010# 0.00167f
C7336 a_39966_32700# a_40352_32700# 0.419f
C7337 a_46116_25164# d2 0.00272f
C7338 X1.X2.X2.X1.X1.X1.vout a_23126_5016# 0.422f
C7339 X1.X1.X2.X2.X1.X1.vout a_8572_18358# 1.64e-19
C7340 a_10686_9828# X1.X1.X2.X1.X1.X2.X2.vin1 0.402f
C7341 a_52106_18358# a_52406_16452# 4.41e-20
C7342 d3 X2.X1.X2.X1.X3.vin2 0.387f
C7343 d6 a_28482_892# 0.00114f
C7344 a_46502_6104# X2.X2.X1.X2.X2.X2.X2.vin1 8.88e-20
C7345 d2 X2.X1.X1.X2.X2.X2.X3.vin1 0.0577f
C7346 X1.X2.X2.X1.X2.X1.X2.vin1 a_25712_13640# 0.197f
C7347 X1.X2.X1.X2.X2.X2.X1.vin1 d0 0.267f
C7348 X1.X1.X1.X2.X1.X1.X3.vin2 a_2582_15634# 0.567f
C7349 d5 a_42976_892# 9.9e-19
C7350 a_8572_18358# X1.X1.X2.X1.X2.X2.X3.vin2 0.00517f
C7351 a_34362_18540# vdd 0.478f
C7352 X2.X1.X1.X1.X2.X2.X3.vin2 vdd 0.761f
C7353 a_54606_26982# d2 0.00328f
C7354 X2.X2.X1.X2.X1.X1.X2.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 0.234f
C7355 a_17222_13728# X1.X2.X1.X2.X1.X2.X3.vin1 0.52f
C7356 X2.X2.X2.vrefh a_49566_892# 7.23e-19
C7357 vrefh vdd 9.92e-19
C7358 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X2.X1.X2.vin1 0.242f
C7359 a_39966_26982# a_39966_28888# 0.00198f
C7360 a_2582_9916# d1 3.95e-19
C7361 X1.X1.X1.X2.X1.X1.vout d1 0.0238f
C7362 a_48702_31882# X2.X2.X1.X1.X1.X1.X1.vin2 0.00743f
C7363 d2 a_48316_31882# 0.0017f
C7364 a_52492_29834# X2.X2.X2.X2.X2.X2.X3.vin1 0.00329f
C7365 d2 a_16836_9916# 0.00272f
C7366 X2.X1.X1.X1.X1.X2.X1.vin1 X2.X1.X1.X1.X1.X2.X1.vin2 0.668f
C7367 a_39966_32700# vdd 0.541f
C7368 d0 X2.X1.X2.X1.X1.X2.X1.vin2 0.276f
C7369 X1.X1.X2.X2.X2.X2.X3.vin2 a_10686_30794# 7.84e-19
C7370 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X1.X2.X2.X2.X2.X1.vin1 0.0689f
C7371 X1.X2.X1.X1.X2.X2.X3.vin2 vdd 0.761f
C7372 X1.X1.X2.X2.X1.X1.X2.vin1 X1.X2.X1.X1.X2.X2.X1.vin2 0.00232f
C7373 a_16836_21352# a_17222_21352# 0.419f
C7374 a_38152_24076# a_39966_23170# 1.06e-19
C7375 a_10686_21264# d1 0.00148f
C7376 X2.X1.X1.X1.X2.X2.vrefh a_31862_23258# 0.3f
C7377 X1.X1.X1.X1.X2.X1.X3.vin2 a_2582_23258# 0.567f
C7378 a_49002_26164# d4 3.47e-19
C7379 X2.X2.X1.X2.X1.X2.vout d1 0.033f
C7380 X1.X2.X2.X2.X1.X1.X1.vin2 X1.X2.X2.X2.X1.X1.X1.vin1 0.668f
C7381 X2.X2.X1.X1.X1.X1.X1.vin2 d1 0.00147f
C7382 d2 X1.X1.X1.X1.X1.X1.X2.vin1 6e-20
C7383 X1.X2.X1.X1.X2.X2.X1.vin2 d2 0.231f
C7384 d1 a_52792_5016# 0.522f
C7385 X1.X1.X1.X3.vin1 d1 0.00955f
C7386 a_17222_19446# a_19336_18540# 4.72e-20
C7387 a_19336_26164# X1.X2.X1.X1.X3.vin2 0.0927f
C7388 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X2.vrefh 0.00118f
C7389 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X1.vin2 0.216f
C7390 a_37766_16452# a_39966_15546# 4.2e-20
C7391 a_25712_6016# X1.X2.X2.X1.X1.X1.X1.vin2 1.78e-19
C7392 a_54992_32700# vrefl 0.118f
C7393 X1.X2.X1.X2.X1.X2.vrefh vdd 0.414f
C7394 X2.X2.X1.X2.X2.X1.X1.vin1 vdd 0.592f
C7395 d0 a_25712_6016# 0.515f
C7396 d0 X1.X1.X1.X2.X1.X2.X2.vin1 0.262f
C7397 X1.X2.X1.X1.X2.X1.X1.vin2 d0 0.276f
C7398 a_31862_11822# X2.X1.X1.X2.X2.X1.X1.vin1 8.22e-20
C7399 a_46116_27070# d0 0.515f
C7400 X1.X1.X1.X1.X2.X2.X3.vin1 d2 0.153f
C7401 d3 a_19036_24258# 0.00178f
C7402 a_2582_27070# X1.X1.X1.X1.X1.X2.X2.vin1 0.402f
C7403 a_25712_26982# d2 0.00272f
C7404 d2 X2.X2.X1.X1.X1.X1.X1.vin1 0.00798f
C7405 X2.X2.X1.X1.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X1.X1.vin2 0.23f
C7406 X2.X2.X2.X1.X1.X1.X3.vin1 a_52792_5016# 0.199f
C7407 X1.X1.X2.X2.X2.X1.X3.vin1 d0 4.36e-19
C7408 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X3.vin1 2.33e-19
C7409 X1.X1.X1.X1.X2.X1.X3.vin1 d0 4.36e-19
C7410 X1.X2.X2.X2.X2.X1.X3.vin2 X1.X2.X2.X2.X2.X2.X3.vin1 1.22e-19
C7411 d2 a_52406_5016# 0.00123f
C7412 a_17222_25164# X1.X2.X1.X1.X2.X1.X3.vin2 7.84e-19
C7413 X2.X1.X1.X1.X2.X1.X2.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 0.234f
C7414 X2.X3.vin1 vdd 1.78f
C7415 X1.X2.X1.X1.X2.X2.vout X1.X2.X1.X1.X2.X2.X3.vin1 0.335f
C7416 a_23512_27888# a_25326_28888# 1.15e-20
C7417 X2.X2.X2.X2.X1.X1.X2.vin1 vdd 0.576f
C7418 d3 X1.X2.X3.vin1 0.834f
C7419 d4 a_31862_17540# 0.00112f
C7420 a_2582_15634# vdd 0.541f
C7421 X2.X1.X2.X2.X1.X2.X3.vin2 a_37766_24076# 0.277f
C7422 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X3.vin1 0.00117f
C7423 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X3.vin1 0.0174f
C7424 a_16836_17540# d1 2.25e-20
C7425 X2.X2.X2.X2.X1.X1.X1.vin2 d2 0.231f
C7426 X1.X2.X1.X1.X1.X2.X2.vin1 a_17222_28976# 8.88e-20
C7427 d3 X1.X1.X1.X1.X2.X1.X3.vin2 2.81e-19
C7428 a_8186_22210# X1.X1.X2.X2.X1.X1.X3.vin2 0.00815f
C7429 a_54606_11734# a_54992_11734# 0.419f
C7430 a_16836_6104# a_16836_8010# 0.00396f
C7431 X2.X2.X1.X2.vrefh a_46116_17540# 1.64e-19
C7432 X1.X2.X2.X2.X2.vrefh d0 0.848f
C7433 X1.X1.X2.X2.X1.X1.vout d2 0.00169f
C7434 a_34362_22312# d4 3.79e-19
C7435 X1.X1.X1.X2.X2.X1.X2.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 0.234f
C7436 d3 X2.X2.X2.X2.X1.X2.X2.vin1 8.68e-20
C7437 a_31476_21352# a_31476_19446# 0.00396f
C7438 X2.X1.X1.X2.X2.X2.vrefh a_31476_8010# 0.118f
C7439 X1.X1.X1.X1.X1.X1.vout d1 0.0238f
C7440 a_52106_18358# X2.X2.X2.X1.X2.X2.X3.vin2 0.00846f
C7441 X2.X2.X1.X1.X3.vin1 X2.X2.X1.X1.X1.X2.vout 0.398f
C7442 X2.X2.X1.X2.X1.X1.X1.vin2 a_46502_15634# 8.88e-20
C7443 a_23212_25982# a_23512_24076# 6.48e-19
C7444 a_33976_26164# vdd 1.05f
C7445 X1.X1.X2.X1.X2.X2.X3.vin2 d2 0.113f
C7446 a_54992_4110# vdd 1.05f
C7447 a_19336_29936# a_17222_28976# 2.68e-20
C7448 X2.X2.X1.X3.vin2 X2.X2.X2.X1.X3.vin2 7.46e-20
C7449 X1.X1.X2.X2.X1.X1.X1.vin2 X1.X1.X2.X2.X1.X1.X1.vin1 0.668f
C7450 X2.X2.X2.X3.vin1 a_52106_14586# 7.98e-19
C7451 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X1.X3.vin2 1.22e-19
C7452 a_2582_8010# vdd 0.541f
C7453 d2 a_8186_29834# 0.273f
C7454 a_31476_9916# a_31476_8010# 0.00396f
C7455 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.vout 0.118f
C7456 a_2582_28976# X1.X1.X1.X1.X1.X1.X3.vin2 8.07e-19
C7457 X1.X1.X2.X1.X2.X1.vout X1.X1.X2.X1.X3.vin2 0.399f
C7458 X1.X1.X2.X1.X1.X1.X2.vin1 d1 0.0144f
C7459 X1.X2.X1.X1.X1.X2.vrefh vdd 0.43f
C7460 X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X2.X1.X3.vin1 0.0321f
C7461 X1.X1.X2.X2.X1.X2.X1.vin2 X1.X1.X2.X2.X1.X1.X3.vin2 3.94e-19
C7462 X1.X1.X2.X2.X1.X2.X1.vin1 a_10686_21264# 8.22e-20
C7463 d2 X1.X2.X2.X1.X1.X1.X3.vin1 3e-19
C7464 a_2582_28976# vdd 0.553f
C7465 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X3.vin1 0.00117f
C7466 X1.X1.X2.X1.X1.X2.X3.vin2 a_8486_8828# 0.277f
C7467 X1.X1.X3.vin1 a_4782_16634# 2.92e-19
C7468 d3 X1.X2.X2.X1.X1.X2.X2.vin1 8.68e-20
C7469 a_22826_14586# vdd 0.567f
C7470 X2.X1.X1.X1.X2.X2.X3.vin2 X2.X1.X1.X2.X1.X1.X1.vin2 3.94e-19
C7471 a_10686_23170# d2 0.00479f
C7472 a_46116_11822# vdd 1.05f
C7473 a_22826_29834# a_23212_29834# 0.419f
C7474 X1.X1.X1.X1.X2.X2.vrefh X1.X1.X1.X1.X2.X2.X1.vin1 0.267f
C7475 X2.X2.X2.X2.X2.X1.X3.vin1 a_54606_26982# 0.52f
C7476 X1.X2.X1.X1.X2.X1.X3.vin2 a_19722_22312# 0.00815f
C7477 X1.X1.X1.X1.X1.X1.X3.vin2 a_2582_30882# 0.567f
C7478 X2.X1.X2.X1.X2.X1.X1.vin1 a_40352_11734# 0.195f
C7479 a_2582_30882# vdd 0.541f
C7480 X2.X2.X2.X1.X2.X2.X1.vin2 X2.X2.X2.X1.X2.X2.X1.vin1 0.668f
C7481 a_46116_23258# a_46502_23258# 0.419f
C7482 a_52106_6962# a_52406_5016# 4.19e-20
C7483 X2.X2.X3.vin1 a_48702_12822# 2.12e-19
C7484 X2.X2.X1.X1.X1.X1.X2.vin1 X2.X2.X1.X1.X1.X1.X3.vin2 0.234f
C7485 a_4696_18540# d2 0.0111f
C7486 X2.X2.X1.X1.X1.X2.X1.vin1 a_46502_30882# 8.22e-20
C7487 X1.X1.X1.X3.vin1 a_5082_18540# 0.389f
C7488 X1.X1.X1.X3.vin2 a_4696_10916# 0.355f
C7489 a_25326_32700# d1 0.00148f
C7490 a_25712_4110# vdd 1.05f
C7491 X1.X1.X1.X1.X2.X1.vout d4 3.29e-19
C7492 X2.X1.X3.vin1 a_37766_5016# 8.66e-20
C7493 X2.X2.X2.X3.vin1 vdd 1.26f
C7494 a_52792_27888# a_52106_25982# 2.97e-19
C7495 X1.X2.X2.X1.X2.vrefh vdd 0.426f
C7496 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X3.vin2 0.161f
C7497 X2.X2.X2.X2.X3.vin1 a_52492_25982# 0.17f
C7498 a_2582_23258# a_4696_22312# 2.95e-20
C7499 a_52792_24076# vdd 1.05f
C7500 X2.vrefh X1.X2.X2.X2.X2.X2.X1.vin2 0.0763f
C7501 a_8572_6962# vdd 1.05f
C7502 a_31476_17540# X2.X1.X1.X2.X1.X1.X2.vin1 1.78e-19
C7503 d3 a_19722_26164# 0.284f
C7504 a_10686_21264# X1.X1.X2.X2.X1.X1.X1.vin2 8.88e-20
C7505 X1.X2.X2.X1.X1.X2.X3.vin1 a_25712_7922# 0.354f
C7506 X2.X1.X3.vin2 d0 0.034f
C7507 d4 a_33676_16634# 0.00176f
C7508 X2.X2.X2.X1.X2.X1.X3.vin2 d1 0.15f
C7509 a_11072_25076# d1 2.92e-22
C7510 X1.X2.X1.X1.X1.X1.X3.vin1 d2 0.00317f
C7511 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.X1.X1.X3.vin1 1.22e-19
C7512 a_19036_9010# a_17222_8010# 1.15e-20
C7513 a_52406_27888# d1 0.0749f
C7514 X2.X2.X3.vin1 X2.X2.X1.X2.X1.X1.vout 2.91e-19
C7515 a_2196_23258# d0 0.515f
C7516 X1.X2.X3.vin2 a_19722_7064# 5.84e-19
C7517 a_54606_11734# X2.X2.X2.X1.X1.X2.X3.vin2 8.07e-19
C7518 X1.X1.X1.X1.X1.X2.X2.vin1 d1 1.03e-19
C7519 a_2196_6104# d0 0.518f
C7520 X2.X2.X2.X2.X2.X2.X3.vin1 vrefl 0.00118f
C7521 X1.X2.X1.X2.X2.X2.X2.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 0.234f
C7522 a_19036_5198# a_19422_5198# 0.419f
C7523 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.X1.vin2 0.22f
C7524 a_8572_25982# a_10686_25076# 4.72e-20
C7525 a_37766_31700# a_39966_30794# 4.2e-20
C7526 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X2.vrefh 0.00118f
C7527 a_16836_6104# X1.X2.X1.X2.X2.X2.X3.vin1 0.354f
C7528 a_17222_6104# X1.X2.X1.X2.X2.X2.X1.vin1 0.417f
C7529 a_17222_6104# a_19422_5198# 4.2e-20
C7530 d3 X2.X2.X1.X1.X3.vin1 0.153f
C7531 X1.X1.X2.X2.X1.X2.X2.vin1 d2 0.0329f
C7532 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.X2.vin1 0.00117f
C7533 a_4396_16634# X1.X1.X1.X2.X1.X1.vout 0.359f
C7534 X2.X1.X2.X2.X2.X1.X3.vin1 a_40352_26982# 0.354f
C7535 a_23212_10734# a_23512_8828# 6.48e-19
C7536 X2.X2.X1.X1.X1.X1.X3.vin2 a_46502_32788# 7.84e-19
C7537 a_10686_13640# X1.X1.X2.X1.X2.X1.X2.vin1 0.402f
C7538 a_48702_28070# d2 0.00202f
C7539 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X2.X1.X2.X1.X1.X2.vin1 0.00232f
C7540 a_48616_7064# X2.X2.X1.X2.X2.X2.X3.vin1 0.00329f
C7541 d3 X1.X1.X2.X1.X2.X1.vout 0.00226f
C7542 a_37766_16452# vdd 0.471f
C7543 X2.X2.X1.X3.vin1 a_49002_22312# 7.98e-19
C7544 X2.X2.X1.X2.X2.X2.X3.vin1 vdd 0.993f
C7545 X1.X2.X2.X1.X2.X2.X1.vin1 vdd 0.592f
C7546 X2.X1.X1.X2.X2.X2.vrefh vdd 0.415f
C7547 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 0.581f
C7548 X1.X1.X1.X2.X2.X1.vout X1.X1.X1.X2.X2.X2.vout 0.514f
C7549 a_25326_28888# a_25712_28888# 0.419f
C7550 d2 X1.X1.X1.X2.X1.X1.X2.vin1 0.031f
C7551 a_52492_29834# a_54606_28888# 2.95e-20
C7552 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.X3.vin1 0.0131f
C7553 a_48316_28070# a_48616_29936# 6.71e-19
C7554 a_10686_32700# a_8872_31700# 1.15e-20
C7555 a_17222_28976# X1.X2.X1.X1.X1.X2.X1.vin1 0.417f
C7556 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.vrefh 0.00118f
C7557 a_16836_28976# X1.X2.X1.X1.X1.X2.X3.vin1 0.354f
C7558 a_23126_20264# X1.X2.X3.vin2 7.93e-20
C7559 X1.X1.X1.X2.X2.X2.X3.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 1.22e-19
C7560 d1 X2.X1.X2.X1.X1.X1.X1.vin1 0.013f
C7561 X2.X1.X2.X1.X1.X2.X1.vin1 X2.X2.X1.X2.X2.X2.vrefh 0.00437f
C7562 a_4396_24258# X1.X1.X1.X1.X2.X1.vout 0.359f
C7563 d0 a_46502_13728# 0.0675f
C7564 a_31476_9916# vdd 1.05f
C7565 X3.vin2 a_42976_892# 0.37f
C7566 a_25326_6016# a_23126_5016# 4.77e-21
C7567 a_17222_8010# vdd 0.541f
C7568 X1.X2.X2.X1.X3.vin2 X1.X2.X2.X1.X3.vin1 0.546f
C7569 X1.X2.X2.X1.X2.X1.vout a_23212_10734# 1.64e-19
C7570 X1.X2.X1.X2.X3.vin1 d1 0.00179f
C7571 a_8572_22210# d1 0.00613f
C7572 a_4696_26164# X1.X1.X1.X3.vin1 0.356f
C7573 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X2.vout 0.0866f
C7574 a_19422_28070# a_19722_26164# 4.41e-20
C7575 X1.X2.X1.X1.X1.X2.X3.vin2 a_19336_26164# 0.00535f
C7576 a_52106_25982# vdd 0.487f
C7577 X2.X2.X2.X2.X2.X1.X2.vin1 d0 0.262f
C7578 X1.X2.X2.X2.X1.X2.X1.vin2 X2.X1.X1.X1.X2.X1.X2.vin1 0.00232f
C7579 d0 a_13696_892# 2.73e-19
C7580 d0 X1.X1.X2.X1.X2.X2.X3.vin1 4.36e-19
C7581 X1.X2.X1.X3.vin2 a_19422_16634# 5.21e-19
C7582 a_19722_18540# X1.X2.X1.X2.X1.X1.X3.vin2 3.49e-19
C7583 X2.X1.X1.X1.X2.X2.X1.vin2 vdd 0.36f
C7584 X2.X2.X2.X1.X3.vin1 vdd 0.805f
C7585 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X3.vin2 0.102f
C7586 X1.X1.X2.X2.X2.X1.X3.vin2 a_10686_30794# 8.07e-19
C7587 a_31476_11822# d1 2.92e-22
C7588 d2 a_33976_29936# 0.606f
C7589 d0 a_54992_17452# 0.515f
C7590 X1.X2.X1.X1.X2.X2.X3.vin1 vdd 0.962f
C7591 a_37766_31700# vdd 0.471f
C7592 a_19722_26164# X1.X2.X1.X1.X3.vin1 0.385f
C7593 X1.X1.X2.X1.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin1 0.00437f
C7594 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X1.X3.vin2 5.19e-19
C7595 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X2.X3.vin1 0.0174f
C7596 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X2.vrefh 2.33e-19
C7597 a_25326_13640# X1.X2.X2.X1.X2.X1.X1.vin2 8.88e-20
C7598 X1.X2.X2.X2.X1.X2.X2.vin1 a_25326_23170# 8.88e-20
C7599 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X1.vin2 8.93e-19
C7600 d3 X1.X1.X1.X2.X2.vrefh 6.65e-20
C7601 a_49002_7064# a_48702_5198# 5.55e-20
C7602 a_54606_9828# X2.X2.X2.X1.X1.X2.X3.vin2 0.567f
C7603 d0 X2.X1.X2.X1.X2.X2.X3.vin2 4.34e-19
C7604 d3 X2.X1.X1.X1.X2.X1.X1.vin2 3.99e-21
C7605 X2.X2.X2.X2.X2.X2.X1.vin2 X2.X2.X2.X2.X2.X2.X1.vin1 0.668f
C7606 X1.X2.X2.X2.X2.X2.X1.vin1 vdd 0.592f
C7607 a_48616_14688# vdd 1.05f
C7608 d1 a_11072_4110# 5.03e-20
C7609 d3 X1.X2.X1.X1.X2.X1.X3.vin1 0.0195f
C7610 a_31862_15634# d1 0.00148f
C7611 X2.X2.X1.X2.X2.X2.X3.vin2 vdd 0.725f
C7612 X1.X1.X2.X1.X2.X1.X1.vin1 a_11072_9828# 1.64e-19
C7613 a_5082_29936# X1.X1.X1.X1.X1.X2.X3.vin1 0.00874f
C7614 X1.X2.X1.X3.vin2 a_19422_9010# 7.93e-20
C7615 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X1.X2.vout 0.398f
C7616 X2.X1.X1.X1.X2.X2.vrefh d1 0.0124f
C7617 a_11072_15546# X1.X1.X2.X1.X2.X2.vrefh 1.64e-19
C7618 X2.X1.X3.vin1 X2.X1.X2.X1.X3.vin2 6.26e-19
C7619 X2.X1.X3.vin2 X2.X1.X1.X2.X3.vin1 4.41e-19
C7620 a_25326_15546# X1.X2.X2.X1.X2.X1.X3.vin2 8.07e-19
C7621 X1.X1.X1.X2.X2.X2.vrefh d1 0.0124f
C7622 a_31862_9916# X2.X1.X1.X2.X2.X1.X2.vin1 8.88e-20
C7623 a_22826_18358# d2 0.00146f
C7624 a_48616_26164# X2.X2.X1.X1.X2.X1.X3.vin1 0.00251f
C7625 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X1.X2.X2.vrefh 0.267f
C7626 X2.X2.X1.X1.X2.vrefh a_46116_27070# 0.118f
C7627 X1.X2.X2.X1.X2.X1.X3.vin1 a_22826_10734# 0.00837f
C7628 X1.X1.X2.X2.X1.X2.X3.vin2 a_11072_25076# 0.354f
C7629 X2.X3.vin2 a_49566_892# 0.51f
C7630 d3 X1.X1.X1.X2.X2.X1.X1.vin2 3.99e-21
C7631 X1.X1.X1.X2.X1.X1.X1.vin1 X1.X1.X1.X2.X1.X1.X1.vin2 0.668f
C7632 X2.X2.X1.X1.X2.X2.X2.vin1 X2.X2.X1.X1.X2.X2.X3.vin2 0.234f
C7633 a_48316_20446# a_48702_20446# 0.419f
C7634 X1.X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X1.X2.X1.vin1 0.00437f
C7635 X1.X1.X2.X1.X2.X1.X1.vin2 d1 4.01e-19
C7636 d3 X2.X1.X2.X2.X3.vin1 0.376f
C7637 a_17222_23258# d1 0.00148f
C7638 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X2.X3.vin2 0.049f
C7639 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X1.X2.X3.vin2 3.94e-19
C7640 X2.X1.X1.X2.X2.X2.vout vdd 0.698f
C7641 X1.X1.X2.X2.X2.X2.X3.vin1 d0 4.36e-19
C7642 a_8486_27888# X1.X1.X2.X2.X2.X1.X3.vin1 0.428f
C7643 X1.X1.X1.X1.X1.X2.X2.vin1 X1.X1.X1.X1.X2.vrefh 0.564f
C7644 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X3.vin1 0.206f
C7645 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X3.vin1 0.00118f
C7646 X2.X2.X2.X2.X1.X2.X1.vin2 vdd 0.361f
C7647 X2.X2.X1.X2.X3.vin2 X2.X2.X1.X2.X2.X1.X3.vin1 0.0321f
C7648 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.X1.vin1 0.206f
C7649 a_8186_29834# X1.X1.X2.X2.X3.vin2 0.422f
C7650 X2.X1.X2.X1.X3.vin1 X2.X1.X2.X1.X1.X2.vout 0.398f
C7651 a_4396_31882# X1.X1.X1.X1.X1.X1.vout 0.359f
C7652 a_37466_10734# X2.X1.X2.X1.X1.X2.X3.vin2 0.00846f
C7653 X2.X1.X2.X2.X2.X2.X1.vin2 X2.X2.X1.X1.X1.X1.X2.vin1 0.00232f
C7654 X1.X1.X2.X1.X1.X1.vout a_8572_6962# 0.169f
C7655 X2.X1.X1.X1.X2.X1.vout a_34362_22312# 0.383f
C7656 X1.X1.X2.X2.X2.X2.X3.vin2 d1 0.0135f
C7657 X2.X2.X2.X2.X1.X2.vout a_52792_24076# 0.36f
C7658 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X2.vrefh 0.00118f
C7659 X2.X2.X1.X1.X2.X1.X2.vin1 a_46502_23258# 0.402f
C7660 d1 a_42976_892# 4.67e-19
C7661 X2.X2.X2.X2.X2.X2.vrefh a_54992_30794# 1.64e-19
C7662 a_52406_16452# X2.X2.X2.X1.X2.X2.vout 0.418f
C7663 a_39966_13640# d1 0.00148f
C7664 d3 a_34362_14688# 0.0469f
C7665 X1.X2.X3.vin2 a_20286_892# 0.0912f
C7666 X2.X2.X1.X3.vin1 d1 0.00955f
C7667 d2 X2.X2.X1.X2.X1.X2.X1.vin2 0.226f
C7668 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X3.vin2 0.449f
C7669 a_39966_6016# X2.X1.X2.X1.X1.X1.X1.vin2 8.88e-20
C7670 a_25326_17452# a_23512_16452# 1.15e-20
C7671 a_31862_30882# d1 0.00148f
C7672 a_46502_28976# d1 3.41e-19
C7673 a_38152_27888# a_39966_26982# 1.06e-19
C7674 a_2196_28976# a_2196_27070# 0.00396f
C7675 X2.X1.X1.X1.X2.vrefh a_31862_27070# 0.3f
C7676 a_52406_8828# vdd 0.47f
C7677 a_25326_19358# X1.X2.X2.X2.vrefh 8.22e-20
C7678 d2 X2.X1.X1.X2.X1.X2.X3.vin1 0.155f
C7679 a_33676_20446# a_33976_18540# 6.48e-19
C7680 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.X1.X1.vin1 5.19e-19
C7681 a_19036_12822# vdd 1.05f
C7682 X2.X1.X1.X1.X2.X2.X2.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 0.234f
C7683 a_33676_20446# a_34062_20446# 0.419f
C7684 X2.X1.X2.X1.X1.X2.X1.vin1 vdd 0.592f
C7685 X1.X1.X3.vin1 X1.X1.X1.X2.X2.X2.vout 0.0857f
C7686 a_34062_28070# X2.X1.X1.X3.vin1 1.64e-19
C7687 X2.X1.X1.X1.X1.X2.X3.vin2 a_34362_26164# 0.00846f
C7688 X2.X2.X2.X1.X1.X2.X3.vin1 a_54606_7922# 0.52f
C7689 d3 a_39966_11734# 0.00112f
C7690 a_19722_10916# a_19422_9010# 5.25e-20
C7691 a_19336_10916# X1.X2.X1.X2.X2.X1.vout 1.64e-19
C7692 a_34062_9010# a_34362_7064# 4.19e-20
C7693 X2.X2.X1.X2.X2.X1.X2.vin1 a_46116_8010# 0.197f
C7694 X2.X1.X1.X2.X1.X1.X1.vin1 d1 0.011f
C7695 X2.X1.X1.X2.X2.X1.vout a_33976_7064# 0.169f
C7696 a_31862_6104# vdd 0.553f
C7697 a_4782_12822# vdd 0.47f
C7698 X1.X2.X2.X2.X1.X2.X2.vin1 vdd 0.576f
C7699 d2 a_46502_17540# 0.00309f
C7700 a_37766_24076# X2.X1.X2.X2.X1.X2.vout 0.418f
C7701 a_25326_25076# a_23512_24076# 1.15e-20
C7702 X1.X1.X2.X2.X1.X1.X3.vin1 d0 4.36e-19
C7703 d3 a_52406_16452# 4.67e-19
C7704 X2.X1.X1.X1.X3.vin2 a_33976_22312# 0.363f
C7705 a_23512_27888# d1 0.521f
C7706 X2.X1.X1.X1.X2.X2.vout d1 0.033f
C7707 X1.X1.X2.X1.X2.X2.vout a_8186_14586# 0.263f
C7708 a_2582_32788# d0 0.0394f
C7709 d2 a_4396_5198# 0.00393f
C7710 a_16836_28976# X1.X2.X1.X1.X1.X2.vrefh 1.64e-19
C7711 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X2.vrefh 2.33e-19
C7712 a_8486_8828# X1.X1.X2.X1.X1.X2.vout 0.418f
C7713 X2.X2.X1.X3.vin1 X2.X2.X3.vin2 7.53e-21
C7714 d1 X2.X1.X1.X2.X2.X2.X3.vin2 0.214f
C7715 d2 a_52106_29834# 0.273f
C7716 a_37766_27888# a_37466_29834# 4.19e-20
C7717 X2.X2.X1.X1.X2.X2.vrefh X2.X2.X1.X1.X2.X2.X1.vin1 0.267f
C7718 d0 a_25712_13640# 0.515f
C7719 a_23126_27888# d2 0.00123f
C7720 a_33976_14688# X2.X1.X1.X2.X1.X2.vout 0.0929f
C7721 a_10686_19358# X1.X1.X2.X2.vrefh 8.22e-20
C7722 d6 a_34926_892# 0.00105f
C7723 a_54992_15546# d1 2.25e-20
C7724 d3 a_37766_24076# 0.00122f
C7725 d2 a_8572_14586# 0.526f
C7726 a_19036_20446# a_19422_20446# 0.419f
C7727 X1.X2.X1.X1.X2.X2.X2.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 0.234f
C7728 X3.vin1 X1.X3.vin2 0.246f
C7729 d0 X1.X1.X2.X1.X2.X1.X3.vin2 4.34e-19
C7730 a_23126_8828# a_22826_6962# 5.55e-20
C7731 a_11072_30794# X1.X1.X2.X2.X2.X2.vrefh 1.64e-19
C7732 a_2582_25164# a_2582_23258# 0.00198f
C7733 X2.X1.X1.X1.X1.X2.X1.vin2 d0 0.276f
C7734 X2.X1.X1.X2.X3.vin2 a_33976_7064# 0.363f
C7735 d3 a_8486_8828# 7.51e-19
C7736 a_10686_26982# X1.X1.X2.X2.X2.vrefh 8.22e-20
C7737 X1.X1.X2.X2.X2.X1.X1.vin2 a_10686_28888# 8.88e-20
C7738 a_52406_24076# d1 0.0749f
C7739 X1.X2.X1.X1.X3.vin2 vdd 1.32f
C7740 d3 a_25712_32700# 2.56e-19
C7741 X2.X2.X2.X1.X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.vout 0.08f
C7742 X1.X2.X1.X1.X1.X2.X3.vin1 d0 4.36e-19
C7743 X2.X1.X1.X1.X2.X2.X3.vin1 a_34062_20446# 0.42f
C7744 X1.X2.X1.X2.X3.vin2 vdd 1.29f
C7745 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X3.vin2 2.23e-19
C7746 a_25326_26982# vdd 0.553f
C7747 X2.X2.X1.X3.vin2 a_49002_14688# 0.00292f
C7748 X2.X1.X1.X2.X1.X2.vrefh a_31476_13728# 1.64e-19
C7749 a_2582_21352# vdd 0.553f
C7750 X2.X2.X2.X1.X2.X2.vout X2.X2.X2.X1.X2.X1.vout 0.514f
C7751 X2.X1.X2.X2.X1.X2.X1.vin1 d1 0.0118f
C7752 X2.X1.X2.X2.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin1 0.00437f
C7753 a_46116_32788# vdd 1.05f
C7754 a_48616_18540# d2 0.0111f
C7755 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X2.X1.X2.X2.X1.X1.vin2 0.00232f
C7756 a_46116_9916# a_46502_9916# 0.419f
C7757 X1.X2.X1.X2.X1.X1.X3.vin2 a_16836_15634# 0.354f
C7758 d2 a_52792_16452# 6.04e-19
C7759 d0 a_25326_17452# 0.0489f
C7760 d2 a_4696_7064# 0.608f
C7761 X1.X2.X1.X2.X1.X2.X1.vin2 X1.X2.X1.X2.X1.X2.X3.vin2 8.93e-19
C7762 X2.X1.X2.X3.vin2 a_37766_24076# 6.03e-19
C7763 a_39966_9828# a_37766_8828# 4.77e-21
C7764 d3 a_19422_16634# 4.67e-19
C7765 d3 a_2582_25164# 0.00112f
C7766 a_46502_19446# vdd 0.541f
C7767 a_2196_11822# X1.X1.X1.X2.X2.X1.X1.vin1 1.64e-19
C7768 a_2582_11822# a_2582_9916# 0.00198f
C7769 a_54606_13640# X2.X2.X2.X1.X2.X1.X3.vin2 0.567f
C7770 a_34062_16634# d1 0.0749f
C7771 a_52406_31700# X2.X2.X2.X2.X2.X2.vout 0.418f
C7772 X2.X1.X1.X1.X1.X1.X1.vin2 X2.X1.X1.X1.X1.X1.X3.vin2 8.93e-19
C7773 a_38152_24076# d2 6.04e-19
C7774 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.vrefh 2.33e-19
C7775 a_25712_19358# a_25712_17452# 0.00396f
C7776 X2.X2.X1.X1.X2.X2.X3.vin2 d0 4.34e-19
C7777 a_10686_17452# vdd 0.541f
C7778 d4 a_8572_18358# 0.63f
C7779 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X3.vin2 1.42e-20
C7780 a_2196_25164# X1.X1.X1.X1.X2.X1.X1.vin2 0.12f
C7781 d2 a_8872_8828# 0.00287f
C7782 a_8186_10734# a_8872_8828# 3.08e-19
C7783 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 0.139f
C7784 a_34926_892# a_35312_892# 0.419f
C7785 d3 a_19422_9010# 0.00148f
C7786 a_54992_30794# d1 2.25e-20
C7787 a_46502_27070# X2.X2.X1.X1.X1.X2.X1.vin2 8.88e-20
C7788 X2.X1.X2.X1.X2.X1.X3.vin1 a_39966_11734# 0.52f
C7789 a_37852_10734# a_37766_8828# 3.3e-19
C7790 X1.X2.X2.X1.X2.X2.vout d1 0.033f
C7791 d2 a_2196_11822# 0.00533f
C7792 a_31476_19446# vdd 1.05f
C7793 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X3.vin2 0.102f
C7794 d3 X2.X2.X2.X1.X2.X1.vout 0.00226f
C7795 X1.X2.X1.X2.X1.X2.vout a_19036_12822# 0.36f
C7796 X2.X2.X1.X1.X2.X1.vout vdd 0.805f
C7797 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X3.vin1 0.00118f
C7798 X2.X2.X1.X1.X1.X2.X3.vin2 a_46502_28976# 7.84e-19
C7799 X1.X1.X1.X1.X2.X2.X2.vin1 d1 1.03e-19
C7800 a_48316_28070# X2.X2.X1.X1.X1.X2.X3.vin1 0.199f
C7801 X2.X1.X1.X1.X2.X2.X3.vin2 d0 4.34e-19
C7802 a_37466_18358# a_37852_18358# 0.416f
C7803 d3 X2.X2.vrefh 0.00665f
C7804 X1.X1.X2.X2.vrefh a_11072_17452# 0.118f
C7805 a_2582_21352# X1.X1.X1.X1.X2.X2.X3.vin2 7.84e-19
C7806 d2 a_52792_31700# 0.00293f
C7807 a_54992_7922# X2.X2.X2.X1.X1.X2.vrefh 1.64e-19
C7808 X1.X1.X1.X2.X2.X2.X1.vin1 vdd 0.592f
C7809 a_52792_31700# a_54606_32700# 1.15e-20
C7810 X1.X1.X1.X1.X2.X2.X3.vin1 a_4396_20446# 0.199f
C7811 d0 vrefh 1.42e-19
C7812 X1.X2.X3.vin2 X1.X2.X2.X1.X1.X1.X3.vin1 0.00836f
C7813 d3 a_19422_31882# 3.23e-19
C7814 a_17222_32788# a_19036_31882# 1.06e-19
C7815 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X2.vin1 0.0689f
C7816 a_16836_19446# vdd 1.05f
C7817 d2 X1.X1.X2.X1.X2.X2.X1.vin1 0.0106f
C7818 a_23512_16452# a_22826_14586# 3.31e-19
C7819 a_8572_14586# a_8872_12640# 6.1e-19
C7820 d2 X1.X2.X1.X2.X2.X2.vrefh 0.168f
C7821 X1.X2.X2.X1.X1.X2.vout d1 0.033f
C7822 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X1.vin2 8.93e-19
C7823 a_39966_32700# d0 0.0489f
C7824 X2.X2.X1.X2.X2.vrefh a_46116_9916# 1.64e-19
C7825 X1.X1.X2.X1.X1.X1.X2.vin1 a_10686_4110# 8.88e-20
C7826 X1.X1.X1.X2.X1.X2.X1.vin1 d1 0.0118f
C7827 X1.X2.X1.X1.X2.X2.X3.vin2 d0 4.34e-19
C7828 a_25712_28888# d1 2.92e-22
C7829 X2.X2.X2.X2.X1.X2.X3.vin2 a_52792_24076# 0.101f
C7830 a_37852_25982# d2 0.0057f
C7831 a_34062_31882# d1 0.0394f
C7832 X2.X2.X1.X2.X2.X2.vrefh X2.X1.X2.X1.X1.X2.vrefh 0.117f
C7833 X2.X1.X1.X1.X1.X2.X2.vin1 X2.X1.X1.X1.X2.vrefh 0.564f
C7834 a_52406_27888# X2.X2.X2.X2.X2.X1.vout 0.422f
C7835 a_37766_27888# X2.X1.X2.X2.X2.X1.X3.vin1 0.428f
C7836 d2 a_17222_13728# 0.00479f
C7837 X2.X2.X2.X1.X1.X1.X1.vin2 a_54992_4110# 0.12f
C7838 a_54606_4110# X2.X2.X2.X1.X1.X1.X1.vin1 0.417f
C7839 a_33976_14688# a_31862_13728# 2.68e-20
C7840 X2.X2.X1.X2.X3.vin1 a_49002_10916# 0.372f
C7841 d2 a_23126_8828# 0.00138f
C7842 X1.X1.X2.X2.X2.X1.X3.vin2 d1 0.15f
C7843 X2.X2.X2.vrefh d5 0.00132f
C7844 d3 a_23512_24076# 0.00108f
C7845 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X2.vrefh 0.1f
C7846 d0 X1.X2.X1.X2.X1.X2.vrefh 0.848f
C7847 d0 X2.X2.X1.X2.X2.X1.X1.vin1 0.267f
C7848 a_17222_32788# vdd 0.554f
C7849 a_2196_19446# vdd 1.05f
C7850 d2 X1.X2.X2.X2.X2.X1.X2.vin1 0.0318f
C7851 d2 X1.X1.X2.X1.X1.X2.X1.vin1 0.0114f
C7852 d3 X2.X1.X1.X2.X1.X2.X3.vin2 0.0247f
C7853 X1.X2.X2.X2.X2.X2.vout d1 0.033f
C7854 X1.X2.X2.X1.X2.vrefh X1.X2.X2.X1.X1.X2.X3.vin2 0.161f
C7855 X2.X1.X3.vin2 X2.X1.X1.X2.X2.X1.vout 4.93e-20
C7856 d0 X2.X3.vin1 0.0254f
C7857 a_8872_27888# vdd 1.05f
C7858 X2.X2.X1.X2.X1.X2.X3.vin1 vdd 0.96f
C7859 X1.X1.X1.X1.X2.X1.X1.vin2 vdd 0.36f
C7860 X2.X1.X1.X2.X1.X2.X3.vin1 a_31862_11822# 0.00207f
C7861 a_10686_28888# X1.X1.X2.X2.X2.X2.vrefh 0.3f
C7862 X2.X1.X1.X1.X2.X1.X3.vin1 a_31862_23258# 0.00207f
C7863 X2.X2.X2.X2.X1.X1.X2.vin1 d0 0.262f
C7864 d2 a_25712_17452# 0.00441f
C7865 X1.X1.X2.X2.X2.X1.X1.vin1 d1 0.0118f
C7866 d4 d2 3.4f
C7867 d0 a_2582_15634# 0.0489f
C7868 a_48316_12822# a_48616_10916# 6.48e-19
C7869 d2 a_54606_11734# 0.00328f
C7870 X2.X2.X1.X1.X1.X2.X2.vin1 vdd 0.576f
C7871 d2 a_23126_31700# 0.00157f
C7872 a_23212_22210# d2 0.526f
C7873 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X3.vin2 0.161f
C7874 X2.X2.X1.X2.vrefh d1 0.00964f
C7875 X3.vin1 vdd 1.51f
C7876 X1.X1.X1.X1.X1.X2.vrefh X1.X1.X1.X1.X1.X1.X2.vin1 0.564f
C7877 X1.X2.X1.X1.X1.X1.X3.vin2 a_16836_30882# 0.354f
C7878 a_19036_28070# a_17222_27070# 1.15e-20
C7879 X3.vin1 a_28096_892# 0.196f
C7880 a_46502_9916# X2.X2.X1.X2.X2.X1.X3.vin2 7.84e-19
C7881 a_25326_11734# a_25326_9828# 0.00198f
C7882 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X2.vrefh 0.161f
C7883 d2 X1.X1.X2.X2.X2.X2.X1.vin1 9.24e-20
C7884 X2.X1.X2.X1.X1.X1.X1.vin2 X2.X1.X2.X1.X1.X1.X1.vin1 0.668f
C7885 d0 a_54992_4110# 0.518f
C7886 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.X2.vrefh 0.076f
C7887 d2 X1.X2.X1.X1.X1.X2.vout 0.109f
C7888 X1.X2.X2.vrefh d5 0.00132f
C7889 a_4696_29936# d1 0.00613f
C7890 X2.X2.X2.X2.X1.X1.vout a_52406_20264# 0.422f
C7891 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X2.vrefh 0.00118f
C7892 d0 a_2582_8010# 0.0489f
C7893 a_19336_14688# X1.X2.X1.X2.X3.vin1 0.363f
C7894 d4 a_17222_17540# 0.00112f
C7895 a_4396_20446# a_4696_18540# 6.48e-19
C7896 d2 X2.X2.X2.X1.X2.X2.X1.vin2 0.231f
C7897 X2.X1.X1.X1.X2.X2.X1.vin2 X2.X1.X1.X1.X2.X2.X2.vin1 0.242f
C7898 X2.X1.X2.X3.vin1 a_37466_10734# 0.509f
C7899 X2.X1.X3.vin2 X2.X1.X1.X2.X3.vin2 0.00254f
C7900 a_31476_23258# a_31476_21352# 0.00396f
C7901 X1.X2.X2.X1.X2.X2.vrefh a_25326_13640# 0.3f
C7902 X1.X1.X2.X2.X2.X1.vout X1.X1.X2.X2.X2.X1.X3.vin2 0.326f
C7903 a_52406_16452# X2.X2.X2.X1.X3.vin2 9.7e-20
C7904 a_2582_28976# d0 0.0675f
C7905 d3 a_34062_9010# 0.00148f
C7906 a_25712_7922# X1.X2.X2.X1.X1.X2.vrefh 1.64e-19
C7907 X1.X1.X1.X2.X2.X2.vout X1.X1.X1.X2.X2.X2.X3.vin2 0.08f
C7908 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X2.X1.X1.X1.X1.X1.vin2 0.00232f
C7909 X1.X2.X1.X1.X1.X2.vrefh d0 0.848f
C7910 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.vrefh 0.267f
C7911 X2.X1.X1.X2.X1.X2.vout vdd 0.697f
C7912 a_19722_29936# X1.X2.X1.X1.X1.X1.vout 0.386f
C7913 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X2.X1.vin1 5.19e-19
C7914 X1.X2.X1.X1.X3.vin1 a_19422_31882# 1.52e-19
C7915 X1.X2.X2.X2.X1.X2.vout d4 3.47e-19
C7916 a_52106_25982# X2.X2.X2.X2.X1.X2.X3.vin2 0.00846f
C7917 X1.X1.X1.X1.X2.X2.X3.vin2 a_2196_19446# 0.354f
C7918 a_4782_20446# a_2582_19446# 4.77e-21
C7919 d0 a_46116_11822# 0.515f
C7920 X1.X2.X1.X1.X1.X2.X3.vin2 vdd 0.787f
C7921 X1.X2.X2.X2.X1.X2.vout a_23212_22210# 0.0929f
C7922 X2.X1.X1.X2.X1.X2.vout a_34062_12822# 0.418f
C7923 d2 a_25712_11734# 0.00272f
C7924 d1 a_48702_9010# 0.0749f
C7925 X2.X1.X3.vin1 a_34362_14688# 3.28e-19
C7926 a_19036_16634# X1.X2.X1.X2.X1.X1.X3.vin2 0.1f
C7927 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X2.vrefh 0.076f
C7928 X1.X2.X2.X2.X1.X1.X3.vin2 a_23512_20264# 0.1f
C7929 X1.X1.X2.X3.vin2 a_8572_18358# 0.0927f
C7930 d3 X1.X2.X2.X1.X2.X1.X3.vin2 2.81e-19
C7931 a_31476_32788# d1 2.25e-20
C7932 a_2582_30882# d0 0.0489f
C7933 X1.X2.X1.X2.X2.X2.vrefh X1.X2.X1.X2.X2.X2.X1.vin2 0.1f
C7934 X1.X1.X2.X3.vin1 a_8572_10734# 0.356f
C7935 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X2.X1.X2.vrefh 0.0128f
C7936 X1.X1.X3.vin2 X1.X1.X2.X1.X3.vin1 0.0361f
C7937 a_25326_9828# X1.X2.X2.X1.X1.X2.X1.vin2 8.88e-20
C7938 X1.X2.X2.X1.X1.X1.X1.vin2 a_25712_4110# 0.12f
C7939 a_46116_13728# a_46502_13728# 0.419f
C7940 a_25326_4110# X1.X2.X2.X1.X1.X1.X1.vin1 0.417f
C7941 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X2.X1.X2.X1.X2.X1.vin2 0.00232f
C7942 X1.X2.X1.X1.X2.X2.X3.vin1 X1.X2.X1.X1.X2.X2.X2.vin1 0.00117f
C7943 d0 a_25712_4110# 0.518f
C7944 a_17222_21352# a_19422_20446# 4.2e-20
C7945 a_4396_24258# d2 3.82e-19
C7946 X1.X1.X1.X3.vin1 a_4782_24258# 5.28e-19
C7947 d4 a_38152_16452# 0.00119f
C7948 d0 X1.X2.X2.X1.X2.vrefh 0.848f
C7949 d3 X2.X1.X1.X1.X1.X2.X3.vin1 2.1e-19
C7950 X2.X2.X2.X2.X2.vrefh d1 0.00745f
C7951 a_17222_19446# X1.X2.X1.X2.X1.X1.X1.vin1 8.22e-20
C7952 d1 X2.X1.X2.X1.X1.X2.vout 0.033f
C7953 X2.X1.X1.X1.X2.vrefh X2.X1.X1.X1.X2.X1.X1.vin1 0.267f
C7954 a_52492_18358# a_52792_16452# 6.48e-19
C7955 d3 a_34362_10916# 0.29f
C7956 X2.X1.X2.X1.X1.X2.X2.vin1 d1 1.03e-19
C7957 d2 a_54606_9828# 0.00792f
C7958 d2 X2.X2.X2.X2.X2.X2.X1.vin2 7.2e-20
C7959 X2.X2.X2.X2.X2.X2.X1.vin2 a_54606_32700# 8.88e-20
C7960 d2 a_37766_8828# 0.00138f
C7961 a_54606_28888# X2.X2.X2.X2.X2.X1.X2.vin1 0.402f
C7962 a_19036_24258# X1.X2.X1.X1.X2.X1.X3.vin2 0.1f
C7963 X2.X1.X2.X1.X1.X2.vrefh vdd 0.43f
C7964 X1.X2.X2.X2.X2.X2.X2.vin1 a_23126_31700# 0.00351f
C7965 X1.X1.X1.X2.X1.X1.X2.vin1 X1.X1.X1.X2.X1.X2.vrefh 0.564f
C7966 a_39966_28888# X2.X1.X2.X2.X2.X2.X1.vin1 8.22e-20
C7967 a_8486_16452# X1.X1.X2.X1.X2.X2.X3.vin1 0.42f
C7968 a_25326_32700# X1.X2.X2.X2.X2.X2.X3.vin1 0.00207f
C7969 X2.X1.X2.X2.X2.X1.X3.vin2 X2.X1.X2.X2.X2.X2.X1.vin2 3.94e-19
C7970 a_46502_21352# d1 3.41e-19
C7971 X2.X1.X1.X1.X2.X2.X1.vin1 X2.X1.X1.X1.X2.X2.X1.vin2 0.668f
C7972 d2 X1.X2.X2.X1.X1.X2.X1.vin1 0.0114f
C7973 X2.X1.X2.X2.X1.X1.X3.vin1 a_37466_18358# 0.00837f
C7974 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X1.vin2 8.93e-19
C7975 X2.X2.X2.X2.X1.X2.X2.vin1 a_54606_23170# 8.88e-20
C7976 X2.X2.X2.X1.X2.X1.X2.vin1 a_54992_11734# 1.78e-19
C7977 X2.X2.X2.X1.X2.X1.X3.vin2 X2.X2.X2.X1.X2.X1.X1.vin1 2.23e-19
C7978 a_8186_25982# a_8486_27888# 5.25e-20
C7979 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X2.X3.vin2 0.587f
C7980 a_48616_10916# d1 0.0126f
C7981 a_10686_4110# a_11072_4110# 0.419f
C7982 a_19036_9010# X1.X2.X1.X2.X2.X1.X3.vin2 0.1f
C7983 X2.X2.X2.X2.X2.X1.X3.vin1 d4 0.00851f
C7984 a_22826_18358# X1.X2.X3.vin2 0.451f
C7985 d0 X2.X2.X1.X2.X2.X2.X3.vin1 4.36e-19
C7986 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X3.vin1 0.0321f
C7987 a_16836_11822# a_17222_11822# 0.419f
C7988 a_33676_28070# d1 0.521f
C7989 d0 X1.X2.X2.X1.X2.X2.X1.vin1 0.267f
C7990 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X2.X3.vin1 0.0131f
C7991 d0 X2.X1.X1.X2.X2.X2.vrefh 0.848f
C7992 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X1.X2.X3.vin2 5.19e-19
C7993 X2.X1.X1.X1.X2.vrefh d2 0.158f
C7994 X2.X2.X2.X1.X2.X1.vout X2.X2.X2.X1.X3.vin2 0.399f
C7995 a_46502_17540# X2.X2.X1.X2.X1.X1.X1.vin2 0.273f
C7996 X2.X1.X1.X1.X2.X1.X3.vin2 a_31862_23258# 0.567f
C7997 a_54606_15546# X2.X2.X2.X1.X2.X1.X3.vin2 8.07e-19
C7998 a_8486_24076# X1.X1.X2.X2.X1.X2.X3.vin1 0.42f
C7999 X1.X1.X1.X1.X2.X1.X2.vin1 X1.X1.X1.X1.X2.X2.vrefh 0.564f
C8000 d2 a_52492_14586# 0.526f
C8001 X1.X2.X3.vin1 a_19422_12822# 2.12e-19
C8002 a_17222_27070# X1.X2.X1.X1.X1.X2.X3.vin1 0.00207f
C8003 X2.X1.X1.X2.X1.X2.vout a_33976_10916# 7.93e-20
C8004 X2.X1.X2.X1.X2.X2.X2.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 0.234f
C8005 a_19722_14688# X1.X2.X1.X2.X1.X2.X3.vin1 0.00874f
C8006 X1.X1.X2.X3.vin2 d2 4.4e-19
C8007 X1.X1.X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.X3.vin2 0.581f
C8008 X1.X2.X1.X2.X1.X1.X3.vin2 vdd 0.905f
C8009 d0 a_31476_9916# 0.518f
C8010 X1.X1.X1.X1.X1.X1.X3.vin1 vdd 1.06f
C8011 d0 a_17222_8010# 0.0489f
C8012 X2.X1.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X1.X2.X1.vin1 0.00437f
C8013 d2 X1.X1.X1.X1.X1.X2.X1.vin2 0.226f
C8014 a_23512_27888# a_22826_25982# 2.97e-19
C8015 X1.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X3.vin1 0.0604f
C8016 X1.X1.X1.X2.X1.X1.X3.vin1 a_2582_15634# 0.00207f
C8017 X1.X1.X2.X2.X2.vrefh d2 0.158f
C8018 X2.X2.X1.X1.X2.X2.vout d2 0.00117f
C8019 X1.X1.X1.X2.X1.X1.vout X1.X1.X1.X2.X1.X2.vout 0.507f
C8020 a_52406_12640# d1 0.0749f
C8021 X2.X2.X1.X2.X2.X1.X3.vin2 X2.X2.X1.X2.X2.X2.X1.vin1 5.19e-19
C8022 X2.X1.X2.X1.X2.X1.X3.vin2 a_38152_12640# 0.1f
C8023 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X2.vrefh 0.076f
C8024 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.vout 0.2f
C8025 a_31862_13728# vdd 0.553f
C8026 a_54606_6016# a_54992_6016# 0.419f
C8027 a_34362_29936# a_34062_31882# 4.19e-20
C8028 a_22826_29834# d1 0.0422f
C8029 X1.X1.X2.X1.X2.X2.vout vdd 0.865f
C8030 X2.X1.X1.X1.X2.X2.X1.vin2 d0 0.276f
C8031 a_33976_29936# X2.X1.X1.X1.X1.X1.vout 0.169f
C8032 a_23212_25982# X1.X2.X2.X2.X3.vin2 0.0927f
C8033 X2.X2.X1.X3.vin1 a_49002_18540# 0.389f
C8034 d4 X2.X1.X2.X2.X2.X2.X3.vin2 1.57e-19
C8035 X2.X1.X1.X1.X2.X1.X3.vin1 a_34062_24258# 0.428f
C8036 X2.X1.X1.X2.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X2.vin1 0.00117f
C8037 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X3.vin2 0.0903f
C8038 X2.X2.X1.X2.X1.X2.vout X2.X2.X1.X2.X1.X2.X3.vin2 0.075f
C8039 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X1.vout 0.399f
C8040 a_46502_25164# X2.X2.X1.X1.X2.X1.X1.vin2 0.273f
C8041 a_31862_13728# a_34062_12822# 4.2e-20
C8042 X2.X1.X2.X2.X1.X2.vrefh d1 0.0071f
C8043 X1.X2.X2.X2.X2.X1.X3.vin1 a_23512_27888# 0.199f
C8044 X2.X1.X2.X2.X2.X1.X2.vin1 vdd 0.576f
C8045 d1 X1.X2.X2.X1.X1.X1.vout 0.0239f
C8046 X1.X2.X2.X1.X2.X2.X1.vin2 a_25326_15546# 0.273f
C8047 X2.X1.X2.X2.X1.X1.X3.vin2 a_37466_18358# 3.49e-19
C8048 X1.X2.X1.X2.X2.X1.X3.vin2 vdd 0.903f
C8049 X1.X2.X1.X1.X2.X2.X3.vin1 d0 4.36e-19
C8050 a_46116_6104# X2.X2.X1.X2.X2.X2.X3.vin1 0.354f
C8051 a_46502_6104# X2.X2.X1.X2.X2.X2.X1.vin1 0.417f
C8052 X2.X2.X2.X2.X1.X1.X1.vin2 X2.X2.X2.X2.vrefh 0.1f
C8053 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X3.vin2 0.234f
C8054 a_19036_31882# X1.X2.X1.X1.X1.X1.X3.vin2 0.1f
C8055 X2.X1.X1.X2.X2.X1.X3.vin2 a_31476_8010# 0.354f
C8056 a_54606_26982# a_54606_25076# 0.00198f
C8057 X1.X2.X2.X2.X2.X2.X1.vin1 d0 0.267f
C8058 a_40352_17452# vdd 1.05f
C8059 a_19722_26164# X1.X2.X1.X1.X2.X1.X3.vin2 3.49e-19
C8060 X1.X2.X1.X1.X3.vin2 a_19422_24258# 0.00101f
C8061 d0 X2.X2.X1.X2.X2.X2.X3.vin2 4.34e-19
C8062 d4 a_52492_18358# 0.63f
C8063 X1.X2.X2.X1.X2.X2.X3.vin2 vdd 0.761f
C8064 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X1.X2.X2.X2.X2.X1.vin1 0.0689f
C8065 d4 X1.X1.X2.X2.X3.vin2 0.0175f
C8066 X1.X1.X2.X3.vin1 a_8486_16452# 5.31e-19
C8067 X1.X2.X2.X2.X1.X1.X2.vin1 a_25712_19358# 1.78e-19
C8068 X1.X2.X2.X2.X1.X1.X3.vin2 X1.X2.X2.X2.X1.X1.X1.vin1 2.23e-19
C8069 d2 X2.X2.X1.X2.X1.X1.vout 0.00169f
C8070 a_19036_28070# a_19336_29936# 6.71e-19
C8071 X2.X1.X1.X3.vin2 d2 4.4e-19
C8072 a_19336_18540# d1 0.00616f
C8073 X2.X2.X1.X1.X2.X2.X2.vin1 a_46502_19446# 0.402f
C8074 X1.X1.X1.X2.X2.X1.X3.vin1 a_4782_9010# 0.428f
C8075 a_10686_32700# X1.X1.X2.X2.X2.X2.X3.vin2 0.567f
C8076 a_31476_4198# vdd 1.05f
C8077 X1.X2.X1.X1.X1.X1.X3.vin2 vdd 0.939f
C8078 a_25326_7922# a_25326_6016# 0.00198f
C8079 X2.X1.X2.vrefh vdd 0.704f
C8080 X2.X2.X3.vin2 a_52406_12640# 2.33e-19
C8081 a_11072_13640# a_11072_11734# 0.00396f
C8082 d1 a_54992_6016# 2.92e-22
C8083 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X1.vin1 5.19e-19
C8084 X2.X2.X1.X1.X2.X1.X1.vin2 d1 4.01e-19
C8085 X1.X1.X1.X2.X3.vin1 vdd 0.804f
C8086 a_19336_29936# a_19722_29936# 0.419f
C8087 X2.X2.X2.X2.X1.X2.X1.vin2 d0 0.276f
C8088 a_8486_31700# X1.X1.X2.X2.X2.X2.X3.vin1 0.42f
C8089 d1 X2.X1.X2.X1.X1.X1.X3.vin2 0.154f
C8090 X2.X1.X1.X1.X2.X1.vout d2 0.00174f
C8091 X2.X1.X1.X1.X2.X1.X3.vin1 d1 0.151f
C8092 X1.X1.X2.X2.X2.X2.vout vdd 0.698f
C8093 a_17222_9916# X1.X2.X1.X2.X2.X1.X1.vin2 0.273f
C8094 X2.X1.X2.X2.X1.X2.vout X2.X1.X2.X2.X1.X1.vout 0.507f
C8095 X2.X2.X1.X2.X2.X2.X1.vin2 a_46502_4198# 8.88e-20
C8096 d2 X2.X2.X2.X1.X1.X1.X2.vin1 6e-20
C8097 X2.X1.X2.X2.X1.X2.vrefh X2.X1.X2.X2.X1.X1.X1.vin2 0.076f
C8098 a_39966_19358# a_40352_19358# 0.419f
C8099 X2.X2.X2.X1.X1.X1.X3.vin2 a_52792_5016# 0.1f
C8100 d2 X1.X1.X1.X2.X2.X1.vout 0.0909f
C8101 X2.X2.X1.X1.X2.X1.X1.vin1 d2 0.0105f
C8102 X2.X1.X2.X2.X2.X2.X2.vin1 X2.X2.vrefh 0.597f
C8103 X1.X1.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X3.vin2 0.0533f
C8104 a_46116_28976# X2.X2.X1.X1.X1.X2.vrefh 1.64e-19
C8105 X2.X1.X2.X1.X1.X2.vrefh X2.X1.X2.X1.X1.X1.X3.vin1 0.00118f
C8106 a_4696_29936# a_4396_31882# 6.1e-19
C8107 X1.X1.X2.X1.X1.X2.X2.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 0.234f
C8108 X2.X1.X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X1.X3.vin1 0.00118f
C8109 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X3.vin1 0.0131f
C8110 X1.X2.X2.vrefh a_20672_892# 7.3e-19
C8111 d5 X2.X3.vin2 0.0456f
C8112 a_46502_6104# a_48702_5198# 4.2e-20
C8113 X2.X2.X1.X2.X2.X2.X3.vin1 X2.X2.X1.X2.X2.X2.X2.vin1 0.00117f
C8114 a_54992_26982# d2 0.00272f
C8115 X1.X2.X1.X2.X2.X1.X1.vin2 d1 4.01e-19
C8116 a_48616_26164# X2.X2.X1.X3.vin1 0.356f
C8117 d3 X2.X1.X2.X2.X1.X1.vout 0.00883f
C8118 X2.X1.X3.vin2 d6 0.013f
C8119 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.X1.X2.vin1 0.0689f
C8120 a_39966_26982# X2.X1.X2.X2.X2.X1.X3.vin2 7.84e-19
C8121 a_48702_16634# X2.X2.X1.X2.X1.X1.X3.vin2 0.267f
C8122 a_2582_4198# vdd 0.541f
C8123 X2.X1.X1.X1.X2.X2.X2.vin1 a_31476_19446# 0.197f
C8124 X1.X1.X1.X2.X2.X1.X3.vin1 d1 0.151f
C8125 d2 X2.X2.X1.X1.X1.X1.vout 0.0904f
C8126 a_54992_13640# X2.X2.X2.X1.X2.X1.X1.vin2 1.78e-19
C8127 a_52492_22210# a_54606_21264# 2.95e-20
C8128 a_25326_21264# a_25712_21264# 0.419f
C8129 X1.X2.X3.vin1 a_23126_5016# 8.66e-20
C8130 X1.X2.X1.X2.X1.X1.X3.vin1 X1.X2.X1.X2.X1.X1.X3.vin2 0.581f
C8131 d2 X1.X2.X1.X2.X2.X1.X1.vin1 0.0105f
C8132 a_25712_21264# d1 2.92e-22
C8133 d0 X2.X1.X2.X1.X1.X2.X1.vin1 0.267f
C8134 X1.X1.X2.X1.X1.X2.X3.vin1 a_8572_6962# 0.00329f
C8135 a_16836_21352# X1.X2.X1.X1.X2.X2.X3.vin1 0.354f
C8136 a_17222_21352# X1.X2.X1.X1.X2.X2.X1.vin1 0.417f
C8137 X2.X1.X2.X1.X1.X2.vout a_37466_6962# 0.254f
C8138 d1 a_46116_4198# 2.81e-20
C8139 X1.X1.X2.X2.X1.X1.X3.vin2 d1 0.15f
C8140 a_48616_29936# a_48702_31882# 3.14e-19
C8141 a_8572_25982# d1 0.0126f
C8142 a_49002_29936# a_48316_31882# 2.86e-19
C8143 a_25326_19358# a_25712_19358# 0.419f
C8144 d1 X2.X2.X2.vrefh 0.258f
C8145 X1.X2.X2.X2.X1.X1.X2.vin1 d2 0.031f
C8146 X1.X1.X2.X1.X3.vin1 d1 0.00179f
C8147 X2.X2.X2.X2.X2.X2.X2.vin1 d1 7.58e-19
C8148 d0 a_31862_6104# 0.0675f
C8149 X2.X1.X2.X2.X3.vin1 a_37852_22210# 0.363f
C8150 X2.X1.X2.X3.vin2 X2.X1.X2.X2.X1.X1.vout 0.0524f
C8151 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.X1.vin1 0.206f
C8152 X1.X2.X1.X3.vin1 X1.X2.X1.X1.X3.vin2 0.418f
C8153 a_52106_22210# d1 0.0422f
C8154 X2.X2.X1.X1.X2.X2.X1.vin2 a_46116_19446# 1.78e-19
C8155 X1.X2.X2.X2.X1.X2.X2.vin1 d0 0.262f
C8156 X2.X1.X1.X2.X2.X1.X3.vin2 vdd 0.903f
C8157 a_2582_27070# a_4782_28070# 4.77e-21
C8158 X1.X2.X1.X2.X1.X2.X2.vin1 a_16836_11822# 0.197f
C8159 X1.X1.X1.X3.vin2 X1.X1.X3.vin2 3.82e-19
C8160 a_8186_18358# X1.X1.X2.X3.vin1 0.374f
C8161 d3 X1.X2.X1.X1.X2.X1.vout 0.00226f
C8162 a_8872_20264# vdd 1.05f
C8163 X1.X2.X2.X2.X2.X2.X1.vin2 a_25326_30794# 0.273f
C8164 X2.X1.X1.X2.X1.X1.X2.vin1 a_31862_15634# 0.402f
C8165 d4 X2.X2.X1.X2.X1.X1.X1.vin2 3.99e-21
C8166 a_23512_27888# X1.X2.X2.X2.X2.X1.X3.vin2 0.1f
C8167 X1.X2.X1.X1.X2.X1.X3.vin1 X1.X2.X1.X1.X2.X1.X3.vin2 0.581f
C8168 a_34062_24258# X2.X1.X1.X1.X2.X1.X3.vin2 0.267f
C8169 d3 a_23212_18358# 7.7e-20
C8170 a_48616_29936# d1 0.00613f
C8171 a_52406_12640# a_52492_10734# 3.21e-19
C8172 X1.X2.X1.X1.X2.vrefh X1.X2.X1.X1.X1.X2.X1.vin2 0.076f
C8173 X2.X1.X3.vin1 a_34062_9010# 2.12e-19
C8174 X1.X1.X2.X1.X2.X2.X1.vin2 vdd 0.36f
C8175 a_31476_17540# X2.X1.X1.X2.X1.X1.X1.vin1 0.195f
C8176 X1.X2.X1.X1.X2.X2.X2.vin1 a_16836_19446# 0.197f
C8177 d4 X2.X1.X1.X2.X1.X1.X3.vin1 0.0205f
C8178 a_19422_28070# a_17222_28976# 4.2e-20
C8179 X1.X2.X3.vin2 a_23126_16452# 3.98e-19
C8180 a_48316_5198# a_48702_5198# 0.419f
C8181 a_54606_9828# a_52792_8828# 1.15e-20
C8182 X2.X1.X3.vin2 a_35312_892# 0.268f
C8183 a_10686_19358# a_8572_18358# 5.36e-21
C8184 X1.X2.X1.X1.X1.X2.X2.vin1 X1.X2.X1.X1.X1.X2.X3.vin1 0.00117f
C8185 X2.X2.X1.X2.X2.X2.X2.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 0.234f
C8186 d2 X1.X2.X2.X1.X3.vin2 0.00194f
C8187 X2.X2.X2.X2.X1.X1.X1.vin1 d2 0.0116f
C8188 a_33676_28070# a_34362_29936# 3.31e-19
C8189 a_34062_28070# a_33976_29936# 3.38e-19
C8190 X1.X2.X1.X2.X2.X2.X1.vin1 a_16836_8010# 1.64e-19
C8191 X2.X2.X2.X1.X2.X1.X1.vin2 X2.X2.X2.X1.X2.vrefh 0.1f
C8192 a_4782_9010# X1.X1.X1.X2.X2.X1.X3.vin2 0.267f
C8193 a_17222_6104# a_17222_8010# 0.00198f
C8194 X2.X1.X2.X1.X3.vin1 a_37852_6962# 0.363f
C8195 X2.X2.X1.X2.vrefh X2.X2.X1.X2.X1.X1.X1.vin1 0.267f
C8196 a_40352_7922# a_40352_6016# 0.00396f
C8197 a_52106_29834# X2.X2.X2.X2.X3.vin2 0.422f
C8198 a_33976_22312# X2.X1.X1.X1.X2.X2.vout 0.0929f
C8199 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X1.X2.vin1 0.242f
C8200 a_11072_13640# vdd 1.05f
C8201 a_31862_21352# a_31862_19446# 0.00198f
C8202 d1 a_16836_4198# 2.81e-20
C8203 X2.X1.X1.X3.vin1 vdd 1.27f
C8204 X1.X1.X2.X2.X1.X1.X3.vin1 a_8186_18358# 0.00837f
C8205 a_19336_29936# X1.X2.X1.X1.X1.X2.X3.vin1 0.00329f
C8206 a_19036_9010# a_19722_7064# 2.86e-19
C8207 a_19422_9010# a_19336_7064# 3.14e-19
C8208 d6 a_13696_892# 0.507f
C8209 a_37466_10734# vdd 0.489f
C8210 d1 X1.X2.X2.vrefh 0.258f
C8211 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X3.vin2 0.17f
C8212 a_10686_19358# a_11072_19358# 0.419f
C8213 X1.X2.X1.X1.X1.X2.X1.vin2 vdd 0.361f
C8214 a_8572_25982# X1.X1.X2.X2.X2.X1.vout 1.64e-19
C8215 X2.X2.X1.X2.X1.X1.X3.vin2 d1 0.15f
C8216 a_25326_26982# d0 0.0675f
C8217 X2.X2.X3.vin2 X2.X2.X2.vrefh 0.15f
C8218 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.vrefh 0.161f
C8219 a_37466_18358# d1 0.0424f
C8220 X1.X1.X2.X1.X1.X2.X1.vin2 vdd 0.361f
C8221 a_2582_21352# d0 0.0675f
C8222 a_39966_19358# d2 0.00309f
C8223 d0 a_46116_32788# 0.511f
C8224 X2.X1.X3.vin1 a_34362_10916# 6.09e-19
C8225 X1.X2.X2.X2.X1.X2.X3.vin1 d2 0.155f
C8226 X1.X2.X3.vin2 a_23126_8828# 2.33e-19
C8227 X1.X1.X1.X1.X1.X2.X3.vin1 X1.X1.X1.X1.X1.X1.X3.vin2 1.22e-19
C8228 a_31476_25164# X2.X1.X1.X1.X2.X1.X1.vin1 0.195f
C8229 a_31862_9916# a_31862_8010# 0.00198f
C8230 X1.X1.X1.X1.X1.X2.X3.vin1 vdd 0.96f
C8231 a_25712_21264# X1.X2.X2.X2.X1.X1.X1.vin2 1.78e-19
C8232 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X2.X1.X1.vin2 3.94e-19
C8233 X1.X1.X2.X2.X1.X2.X1.vin1 X1.X1.X2.X2.X1.X1.X3.vin2 5.19e-19
C8234 X1.X1.X1.X1.X2.X2.vrefh d1 0.0124f
C8235 a_33676_9010# X2.X1.X1.X2.X2.X1.X3.vin2 0.1f
C8236 X2.X2.X1.X2.vrefh X2.X1.X2.X2.vrefh 0.117f
C8237 a_11072_23170# d2 0.00351f
C8238 X1.X1.X2.X1.X2.X2.X3.vin2 a_8186_14586# 3.85e-19
C8239 X2.X2.X2.X1.X1.X1.vout d1 0.0239f
C8240 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.vout 0.335f
C8241 a_23512_12640# d1 0.521f
C8242 X2.X1.X1.X1.X2.X1.X3.vin2 d1 0.15f
C8243 X1.X1.X1.X1.X2.X2.X2.vin1 X1.X1.X1.X2.vrefh 0.564f
C8244 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X1.X2.vin1 0.242f
C8245 a_8486_20264# X1.X1.X2.X2.X1.X1.X3.vin1 0.428f
C8246 a_17222_11822# a_19336_10916# 4.72e-20
C8247 a_46502_19446# d0 0.0489f
C8248 a_33676_5198# X2.X1.X1.X2.X2.X2.X3.vin2 0.101f
C8249 X2.X2.X2.X2.X2.X1.X3.vin1 a_54992_26982# 0.354f
C8250 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X2.X1.X2.X1.X2.X2.vin1 0.00232f
C8251 a_2196_6104# a_2196_8010# 0.00396f
C8252 a_25326_19358# d2 0.00309f
C8253 X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X3.vin1 0.00836f
C8254 X1.X1.X2.X2.X2.X2.X1.vin2 vdd 0.387f
C8255 X1.X1.X1.X2.X1.X2.X3.vin2 X1.X1.X1.X2.X2.X1.X1.vin2 3.94e-19
C8256 X2.X2.X2.X1.X1.X1.vout X2.X2.X2.X1.X1.X1.X3.vin1 0.118f
C8257 a_2196_32788# a_2582_32788# 0.419f
C8258 d4 X1.X2.X3.vin2 0.297f
C8259 X1.X1.X1.X2.X2.X1.X3.vin2 d1 0.15f
C8260 a_54606_15546# a_54992_15546# 0.419f
C8261 a_10686_17452# d0 0.0489f
C8262 a_33976_7064# a_34362_7064# 0.419f
C8263 X1.X1.X3.vin1 a_8186_10734# 3.93e-19
C8264 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X3.vin2 0.17f
C8265 X1.X2.X2.X2.X1.X1.vout a_23212_18358# 1.64e-19
C8266 a_52406_20264# vdd 0.561f
C8267 X1.X2.X2.X2.X2.X2.X3.vin2 d1 0.0135f
C8268 X1.X1.X3.vin1 d2 0.1f
C8269 a_48702_31882# X2.X2.X1.X1.X1.X1.X3.vin2 0.267f
C8270 a_37766_24076# a_37852_22210# 3.38e-19
C8271 a_46502_15634# vdd 0.541f
C8272 a_37766_27888# d3 0.00195f
C8273 a_31476_19446# d0 0.515f
C8274 X1.X1.X2.X2.X1.X1.X2.vin1 a_10686_19358# 8.88e-20
C8275 a_31862_17540# a_33676_16634# 1.06e-19
C8276 X2.X2.X1.X1.X2.X2.vrefh vdd 0.415f
C8277 a_25712_32700# a_25712_30794# 0.00396f
C8278 a_19722_7064# vdd 0.477f
C8279 X1.X1.X2.X2.X1.X1.X3.vin2 X1.X1.X2.X2.X1.X1.X1.vin2 8.93e-19
C8280 X2.X1.X1.X2.X1.X1.X1.vin1 X2.X1.X1.X2.X1.X1.X2.vin1 0.0689f
C8281 a_39966_28888# X2.X1.X2.X2.X2.X2.vrefh 0.3f
C8282 d4 X2.X1.X1.X2.X1.X1.vout 0.00145f
C8283 a_22826_6962# a_23512_5016# 2.86e-19
C8284 d1 a_25326_6016# 0.00148f
C8285 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.vout 0.326f
C8286 a_17222_25164# d1 3.95e-19
C8287 d2 X2.X1.X1.X2.X2.X2.X1.vin2 7.2e-20
C8288 a_10686_19358# d2 0.00309f
C8289 d2 X1.X1.X2.X1.X2.X1.X3.vin1 0.104f
C8290 X1.X1.X2.X1.X2.X1.X3.vin1 a_8186_10734# 0.00837f
C8291 X1.X3.vin2 a_20286_892# 0.51f
C8292 X2.X2.X1.X1.X1.X1.X3.vin2 d1 0.152f
C8293 a_31476_25164# d2 0.00272f
C8294 a_2196_9916# X1.X1.X1.X2.X2.X1.X1.vin1 0.195f
C8295 a_37766_20264# vdd 0.561f
C8296 a_4782_28070# d1 0.0749f
C8297 a_8572_25982# X1.X1.X2.X2.X1.X2.X3.vin2 0.00535f
C8298 X1.X1.X1.X2.X2.X2.X1.vin1 d0 0.267f
C8299 a_25326_11734# vdd 0.553f
C8300 a_19422_5198# X1.X2.X1.X2.X2.X2.X3.vin2 0.277f
C8301 a_17222_13728# X1.X2.X1.X2.X1.X2.X1.vin2 0.273f
C8302 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X3.vin2 2.23e-19
C8303 X1.X2.X1.X2.X2.X2.X3.vin1 a_19422_5198# 0.42f
C8304 a_31476_23258# vdd 1.05f
C8305 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.X1.vin1 0.206f
C8306 X2.X2.X3.vin2 X2.X2.X2.X1.X1.X1.vout 0.033f
C8307 X1.X2.X1.X2.X2.X2.X1.vin1 X1.X2.X1.X2.X2.X2.X3.vin1 0.206f
C8308 a_16836_19446# d0 0.515f
C8309 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.vout 0.326f
C8310 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X1.X3.vin1 0.581f
C8311 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X1.X2.X2.X1.X2.X1.vin1 0.668f
C8312 a_52492_29834# X2.X2.X2.X2.X2.X2.vout 0.0929f
C8313 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X3.vin2 0.234f
C8314 X2.X1.X1.X1.X1.X1.X2.vin1 a_31862_30882# 0.402f
C8315 X2.X2.X2.X3.vin2 d2 4.4e-19
C8316 a_37766_27888# X2.X1.X2.X3.vin2 7.93e-20
C8317 a_4396_20446# d4 0.00107f
C8318 d3 X1.X1.X1.X1.X2.X2.vout 8.47e-19
C8319 a_11072_19358# a_11072_17452# 0.00396f
C8320 a_37466_6962# X2.X1.X2.X1.X1.X1.X3.vin2 0.00815f
C8321 d2 a_2196_9916# 0.00272f
C8322 a_23126_20264# vdd 0.561f
C8323 X1.X2.vrefh X1.X1.X2.X2.X2.X2.X1.vin2 0.0763f
C8324 a_46116_13728# a_46116_11822# 0.00396f
C8325 X1.X2.X2.X2.X2.X1.X3.vin2 a_25712_28888# 0.354f
C8326 a_52492_29834# X2.X2.X2.X2.X2.X1.X3.vin2 0.00546f
C8327 a_54606_13640# a_52406_12640# 4.77e-21
C8328 a_48702_28070# a_49002_29936# 5.55e-20
C8329 X2.X1.X1.X2.X1.X2.vrefh X1.X2.X2.X1.X2.X2.vrefh 0.117f
C8330 a_17222_32788# d0 0.0394f
C8331 X2.X2.X2.X1.X1.X1.vout X2.X2.X2.X1.X1.X2.vout 0.507f
C8332 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X2.vrefh 0.076f
C8333 a_2196_19446# d0 0.515f
C8334 X1.X2.X2.X1.X2.X1.vout X1.X2.X2.X1.X2.X1.X3.vin2 0.326f
C8335 X1.X1.X2.X2.X2.X2.X3.vin2 a_8872_31700# 0.101f
C8336 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X2.X3.vin1 0.206f
C8337 a_46502_30882# vdd 0.541f
C8338 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X2.vrefh 0.00118f
C8339 a_23212_14586# d1 0.00613f
C8340 X1.X1.X1.X1.X2.X2.X1.vin2 d2 0.231f
C8341 d4 X2.X1.X1.X1.X1.X1.vout 0.0336f
C8342 X2.X1.X1.X2.X2.X1.X1.vin1 vdd 0.592f
C8343 X1.X2.X2.X1.X1.X1.X2.vin1 X1.X2.X2.X1.X1.X1.X3.vin1 0.00117f
C8344 X2.X2.X1.X2.X2.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin2 0.1f
C8345 X3.vin2 X2.X3.vin2 0.215f
C8346 X1.X1.X1.X1.X2.X1.X1.vin2 d0 0.276f
C8347 d0 X2.X2.X1.X2.X1.X2.X3.vin1 4.36e-19
C8348 X1.X2.X2.X1.X1.X1.X3.vin2 a_23126_5016# 0.267f
C8349 X1.X2.X2.X1.X1.X2.X1.vin2 vdd 0.361f
C8350 a_5082_26164# d2 7.13e-19
C8351 a_54606_9828# X2.X2.X2.X1.X1.X2.X1.vin2 8.88e-20
C8352 a_19722_22312# d1 0.0422f
C8353 X2.X1.X1.X2.X1.X2.X3.vin2 a_31862_9916# 8.07e-19
C8354 X2.X2.X1.X1.X1.X2.X2.vin1 d0 0.262f
C8355 X1.X1.X1.X3.vin2 a_4782_9010# 7.93e-20
C8356 d0 X3.vin1 0.0184f
C8357 X2.X1.X2.X1.X3.vin1 a_37766_5016# 1.52e-19
C8358 d3 a_8486_24076# 0.00122f
C8359 d3 X2.X2.X1.X2.X2.X1.X3.vin2 7.71e-19
C8360 X2.X1.X2.X1.X1.X2.X1.vin2 a_39966_7922# 0.273f
C8361 d4 X2.X2.X2.X2.X3.vin2 0.0939f
C8362 X2.X1.X2.X2.X1.X1.X2.vin1 vdd 0.576f
C8363 X2.X2.X1.X1.X2.X1.X3.vin2 a_46502_21352# 8.07e-19
C8364 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.vout 0.335f
C8365 d2 X2.X1.X1.X1.X3.vin1 0.0594f
C8366 a_2196_17540# d1 2.25e-20
C8367 a_11072_17452# d2 0.00441f
C8368 X1.X2.X1.X1.X2.X2.vrefh a_17222_21352# 8.22e-20
C8369 X1.X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.X1.X1.vin2 0.076f
C8370 a_31862_8010# X2.X1.X1.X2.X2.X2.X1.vin1 8.22e-20
C8371 d2 X2.X1.X2.X1.X1.X1.vout 0.115f
C8372 X1.X2.X2.X1.X2.X1.X2.vin1 a_25326_11734# 8.88e-20
C8373 X1.X2.X2.X2.X1.X2.X3.vin2 X1.X2.X2.X2.X1.X2.X1.vin1 2.23e-19
C8374 d3 X2.X1.X2.X2.X1.X2.X2.vin1 8.68e-20
C8375 X1.X2.X2.X1.X3.vin1 a_22826_6962# 0.436f
C8376 X1.X2.X2.X1.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X1.vin2 8.93e-19
C8377 X1.X2.X2.X2.X1.X2.X2.vin1 a_25712_23170# 1.78e-19
C8378 a_54606_30794# a_54992_30794# 0.419f
C8379 X2.X2.X1.X2.X3.vin1 vdd 0.804f
C8380 X1.X1.X2.X1.X2.X1.X3.vin1 a_8872_12640# 0.199f
C8381 d2 a_4782_31882# 7.51e-19
C8382 a_37466_29834# X2.X1.X2.X2.X2.X1.vout 0.383f
C8383 a_23126_27888# X1.X2.X2.X2.X2.X1.vout 0.422f
C8384 a_52492_6962# X2.X2.X2.X1.X3.vin1 0.363f
C8385 a_5082_10916# vdd 0.487f
C8386 X2.X1.X2.X1.X2.X2.X1.vin2 d1 2.18e-19
C8387 d2 a_23512_5016# 0.00251f
C8388 a_48616_22312# vdd 1.05f
C8389 X1.X2.X1.X1.X1.X2.X3.vin2 d0 4.34e-19
C8390 d4 a_5082_29936# 0.00116f
C8391 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X1.X3.vin1 0.0425f
C8392 a_46116_27070# a_46502_27070# 0.419f
C8393 X1.X1.X1.X3.vin2 d1 0.0129f
C8394 X1.X2.X1.X3.vin2 a_19336_10916# 0.355f
C8395 a_10686_6016# d2 4.64e-19
C8396 a_31862_9916# a_34062_9010# 4.2e-20
C8397 a_16836_21352# a_16836_19446# 0.00396f
C8398 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X2.vin1 0.00117f
C8399 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X3.vin1 0.0131f
C8400 a_52792_27888# a_54606_26982# 1.06e-19
C8401 X2.X1.X1.X2.vrefh d4 6.65e-20
C8402 d3 X1.X1.X2.X1.X1.X2.X2.vin1 8.68e-20
C8403 a_8872_24076# d2 6.04e-19
C8404 a_48702_20446# X2.X2.X1.X1.X2.X2.X3.vin2 0.277f
C8405 X1.X1.X2.X1.X2.X1.X1.vin1 d1 0.0118f
C8406 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X1.X3.vin1 0.0425f
C8407 X1.X2.X2.X2.X1.X2.X1.vin2 d1 0.00406f
C8408 X2.X2.X1.X2.X1.X2.X2.vin1 vdd 0.576f
C8409 a_39966_17452# X2.X1.X2.X1.X2.X2.X3.vin1 0.00207f
C8410 X2.X2.X2.X2.X1.X2.X1.vin1 vdd 0.592f
C8411 X1.X2.X2.X2.X2.vrefh a_25326_25076# 0.3f
C8412 X1.X1.X2.X2.X1.X2.vrefh a_11072_21264# 0.118f
C8413 a_48702_24258# a_46502_23258# 4.77e-21
C8414 X2.X1.X3.vin2 a_34362_7064# 5.84e-19
C8415 a_20286_892# vdd 1.05f
C8416 a_54992_13640# d1 2.92e-22
C8417 X1.X2.X1.X2.vrefh d4 6.65e-20
C8418 a_31862_32788# d4 8.99e-20
C8419 X1.X2.X1.X2.X1.X1.X2.vin1 d1 1.03e-19
C8420 d1 X2.X3.vin2 0.00146f
C8421 X1.X2.X1.X1.X2.X2.X3.vin2 X1.X2.X1.X2.X1.X1.X1.vin2 3.94e-19
C8422 X1.X2.X1.X1.X1.X1.X1.vin2 d2 1.68e-19
C8423 a_48316_16634# vdd 1.05f
C8424 X2.X1.X2.X1.X2.X1.X3.vin2 d1 0.15f
C8425 a_52492_25982# d1 0.0126f
C8426 d0 X2.X1.X2.X1.X1.X2.vrefh 0.848f
C8427 a_17222_9916# X1.X2.X1.X2.X2.X1.X2.vin1 8.88e-20
C8428 X2.X1.X2.X1.X1.X1.X2.vin1 a_39966_4110# 8.88e-20
C8429 X2.X1.X2.X1.X1.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X1.vin2 8.93e-19
C8430 d2 X2.X2.X2.X1.X2.X1.X2.vin1 0.0318f
C8431 X2.X1.X1.X1.X1.X2.vrefh X1.X2.X2.X2.X2.X2.vrefh 0.117f
C8432 X1.X2.X2.X1.X2.X2.X3.vin2 a_23512_16452# 0.101f
C8433 X2.X1.X2.X2.X2.X2.X1.vin2 d1 0.0985f
C8434 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X2.vrefh 0.076f
C8435 a_10686_7922# X1.X1.X2.X1.X1.X2.vrefh 8.22e-20
C8436 a_25712_19358# X1.X2.X2.X2.vrefh 1.64e-19
C8437 X2.X2.X1.X1.X1.X2.X3.vin1 d1 0.146f
C8438 a_4696_18540# a_2582_17540# 5.36e-21
C8439 a_33976_18540# a_34362_18540# 0.413f
C8440 X1.X2.X1.X2.X1.X2.X3.vin2 vdd 0.787f
C8441 X1.X1.X3.vin2 a_8186_6962# 0.00111f
C8442 a_34062_20446# a_34362_18540# 4.41e-20
C8443 a_34062_20446# X2.X1.X1.X1.X2.X2.X3.vin2 0.277f
C8444 X2.X1.X2.X1.X2.X2.X3.vin1 X2.X1.X2.X1.X2.X2.vrefh 2.33e-19
C8445 X2.X1.X1.X1.X2.X2.X3.vin2 a_33976_18540# 0.00504f
C8446 a_5082_26164# a_4396_28070# 3.08e-19
C8447 a_4696_26164# a_4782_28070# 3.3e-19
C8448 a_10686_6016# X1.X1.X2.X1.X1.X1.X3.vin2 0.567f
C8449 a_37766_27888# a_39966_28888# 4.77e-21
C8450 X1.X2.X1.X2.X2.X1.X2.vin1 d1 1.03e-19
C8451 d3 X1.X2.X2.X2.X3.vin2 0.157f
C8452 a_33676_24258# vdd 1.05f
C8453 a_54606_17452# d1 0.00148f
C8454 X2.X2.X2.X1.X1.X2.X3.vin1 a_54992_7922# 0.354f
C8455 X2.X2.X1.X2.X2.X2.X1.vin2 vdd 0.387f
C8456 a_2196_13728# X1.X1.X1.X2.X1.X2.X1.vin1 0.195f
C8457 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X2.vrefh 0.1f
C8458 a_4396_9010# vdd 1.05f
C8459 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X1.vout 0.399f
C8460 a_46116_25164# vdd 1.05f
C8461 a_2582_19446# X1.X1.X1.X2.X1.X1.X1.vin1 8.22e-20
C8462 X2.X2.X1.X1.X2.X1.X1.vin2 X2.X2.X1.X1.X2.X1.X3.vin2 8.93e-19
C8463 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X1.vout 0.0524f
C8464 d1 X1.X1.X2.X1.X1.X1.X3.vin1 0.16f
C8465 X2.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 8.36e-19
C8466 a_48316_9010# a_46502_8010# 1.15e-20
C8467 X2.X1.X1.X2.X2.X1.vout X2.X1.X1.X2.X2.X2.vout 0.514f
C8468 X2.X1.X1.X2.X2.X2.X3.vin1 vdd 0.993f
C8469 a_52492_6962# a_52406_8828# 3.38e-19
C8470 X2.X1.X2.X1.X2.X1.vout a_37852_10734# 1.64e-19
C8471 X1.X2.X2.X2.X3.vin1 d2 0.0014f
C8472 X2.X1.X2.X1.X3.vin2 X2.X1.X2.X1.X3.vin1 0.546f
C8473 d2 X2.X2.X1.X2.X1.X1.X3.vin1 0.104f
C8474 a_16836_28976# X1.X2.X1.X1.X1.X2.X1.vin2 0.12f
C8475 X2.X2.X2.X1.X2.vrefh d1 0.00745f
C8476 a_54606_7922# a_54606_6016# 0.00198f
C8477 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X2.vout 0.0866f
C8478 X1.X2.X2.X2.X1.X2.X3.vin2 a_23512_24076# 0.101f
C8479 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X2.vrefh 0.076f
C8480 a_19336_10916# a_19722_10916# 0.414f
C8481 a_54606_26982# vdd 0.553f
C8482 d0 X1.X2.X1.X2.X1.X1.X3.vin2 4.34e-19
C8483 d2 X1.X2.X2.X1.X3.vin1 0.0619f
C8484 X1.X1.X1.X2.X2.X2.X1.vin2 X1.X1.X1.X2.X2.X1.X3.vin2 3.94e-19
C8485 X2.X2.X3.vin2 X2.X3.vin2 0.147f
C8486 d2 X1.X1.X1.X2.X2.X2.X3.vin2 8.42e-19
C8487 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X2.X3.vin1 1.42e-20
C8488 X1.X1.X1.X1.X1.X1.X3.vin1 d0 4.36e-19
C8489 a_49952_892# vdd 0.477f
C8490 a_5082_18540# X1.X1.X1.X3.vin2 0.233f
C8491 a_34062_28070# d4 2.4e-19
C8492 a_10686_28888# X1.X1.X2.X2.X2.X1.X3.vin2 0.567f
C8493 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X2.vrefh 0.267f
C8494 X1.X2.X1.X1.X1.X1.X2.vin1 d1 0.0144f
C8495 X2.X2.X2.X3.vin2 a_52492_18358# 0.0927f
C8496 a_48316_31882# vdd 1.05f
C8497 a_54606_19358# a_54606_17452# 0.00198f
C8498 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X1.vout 0.118f
C8499 a_52106_29834# X2.X2.X2.X2.X2.X2.X3.vin2 3.85e-19
C8500 X2.X1.X1.X1.X1.X2.vout d1 0.033f
C8501 d0 a_31862_13728# 0.0675f
C8502 a_16836_9916# vdd 1.05f
C8503 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.vout 0.398f
C8504 X2.X1.X2.X1.X1.X1.X1.vin2 X2.X2.X2.vrefh 0.0128f
C8505 a_11072_19358# X1.X1.X2.X2.vrefh 1.64e-19
C8506 a_8572_22210# a_10686_21264# 2.95e-20
C8507 d1 a_37852_6962# 0.00613f
C8508 d6 X2.X3.vin1 0.0293f
C8509 d2 a_19722_14688# 0.0191f
C8510 X2.X1.X3.vin1 a_34926_892# 0.17f
C8511 a_2582_17540# X1.X1.X1.X2.X1.X1.X2.vin1 8.88e-20
C8512 a_19422_20446# X1.X2.X1.X1.X2.X2.X3.vin2 0.277f
C8513 a_22826_29834# X1.X2.X2.X2.X2.X1.X3.vin2 0.00815f
C8514 X1.X1.X1.X1.X2.X1.X3.vin1 a_2582_23258# 0.00207f
C8515 X2.X1.X2.X2.X2.X1.X2.vin1 d0 0.262f
C8516 X2.X2.X2.X2.vrefh d4 6.65e-20
C8517 a_10686_26982# X1.X1.X2.X2.X2.X1.X2.vin1 8.88e-20
C8518 d0 X1.X2.X1.X2.X2.X1.X3.vin2 4.34e-19
C8519 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X2.vout 0.0866f
C8520 X1.X1.X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X1.X1.X2.vin1 0.234f
C8521 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.X1.X3.vin2 8.93e-19
C8522 a_11072_26982# X1.X1.X2.X2.X2.vrefh 1.64e-19
C8523 X1.X1.X1.X1.X1.X1.X2.vin1 vdd 0.578f
C8524 X2.X1.X2.X2.X1.X2.X1.vin1 a_40352_21264# 1.64e-19
C8525 X1.X1.X2.X1.X2.X1.X3.vin1 a_10686_11734# 0.52f
C8526 X1.X2.X1.X1.X2.X2.X1.vin2 vdd 0.36f
C8527 X1.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X1.X2.vout 0.398f
C8528 d0 a_40352_17452# 0.515f
C8529 X2.X2.X2.X1.X2.X1.X3.vin1 a_54606_11734# 0.52f
C8530 a_54606_9828# a_54992_9828# 0.419f
C8531 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.vrefh 0.1f
C8532 a_25712_25076# X1.X2.X2.X2.X1.X2.X1.vin2 1.78e-19
C8533 a_33676_12822# d1 0.521f
C8534 X2.X1.X1.X2.X1.X2.vrefh X2.X1.X1.X2.X1.X2.X1.vin1 0.267f
C8535 X1.X2.X2.X2.X1.X2.vrefh X2.X1.X1.X1.X2.X2.X1.vin2 0.0128f
C8536 d4 X1.X2.X2.X2.X2.X1.vout 0.0233f
C8537 X1.X1.X1.X1.X2.X2.X3.vin1 vdd 0.962f
C8538 a_25712_26982# vdd 1.05f
C8539 d2 X2.X2.X1.X2.X1.X2.vrefh 0.177f
C8540 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.vout 0.326f
C8541 d1 a_54606_7922# 3.41e-19
C8542 d3 X1.X2.X1.X1.X2.X1.X1.vin2 3.99e-21
C8543 a_46116_9916# X2.X2.X1.X2.X2.X1.X3.vin1 0.354f
C8544 d0 X1.X2.X2.X1.X2.X2.X3.vin2 4.34e-19
C8545 X2.X2.X1.X2.X1.X1.X1.vin1 X2.X2.X1.X2.X1.X1.X3.vin2 2.23e-19
C8546 a_46502_9916# X2.X2.X1.X2.X2.X1.X1.vin1 0.417f
C8547 a_22826_29834# X1.X2.X2.X2.X2.X2.X3.vin1 0.00874f
C8548 a_52406_5016# vdd 0.562f
C8549 d3 X1.X1.X1.X2.X1.X2.X2.vin1 8.68e-20
C8550 d2 X2.X1.X1.X2.X2.vrefh 0.158f
C8551 X2.X2.X1.X1.X1.X1.X1.vin1 vdd 0.596f
C8552 X2.X2.X3.vin1 d2 0.1f
C8553 a_8186_14586# a_8572_14586# 0.419f
C8554 d2 X1.X1.X1.X2.X2.X2.vout 0.11f
C8555 X1.X2.X2.X2.vrefh d2 0.173f
C8556 X2.X2.X2.X2.vrefh X2.X2.X2.X1.X2.X2.X1.vin2 0.076f
C8557 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.X1.X1.vin1 0.668f
C8558 a_37852_14586# a_37766_12640# 3.14e-19
C8559 X2.X1.X2.X1.X1.X2.X2.vin1 X2.X1.X2.X1.X1.X2.X3.vin1 0.00117f
C8560 X1.X2.X3.vin1 d5 0.0539f
C8561 X2.X1.X2.X1.X1.X2.X3.vin2 a_37766_8828# 0.277f
C8562 d3 X1.X1.X2.X2.X2.X1.X3.vin1 0.0332f
C8563 d0 a_31476_4198# 0.515f
C8564 X1.X2.X1.X1.X1.X1.X3.vin2 d0 4.34e-19
C8565 d3 X1.X1.X1.X1.X2.X1.X3.vin1 0.0195f
C8566 X1.X2.X2.X1.X1.X1.X1.vin2 X2.X1.X2.vrefh 0.0128f
C8567 a_40352_26982# a_40352_25076# 0.00396f
C8568 d0 X2.X1.X2.vrefh 4.78f
C8569 X2.X2.X2.X2.X1.X1.X1.vin2 vdd 0.36f
C8570 a_2196_23258# a_2196_21352# 0.00396f
C8571 d2 a_31476_15634# 0.00414f
C8572 X1.X2.X1.X1.X3.vin1 X1.X2.X2.X2.X3.vin2 0.0604f
C8573 a_37466_22210# a_37766_20264# 4.19e-20
C8574 d2 X1.X1.X2.X1.X2.vrefh 0.158f
C8575 X1.X1.X2.X2.X1.X1.vout vdd 0.78f
C8576 a_23512_12640# a_22826_10734# 2.97e-19
C8577 X1.X1.X2.X2.X3.vin1 a_8486_24076# 9.54e-19
C8578 X1.X2.X3.vin2 X1.X2.X2.X1.X3.vin2 0.039f
C8579 a_8486_27888# a_8872_27888# 0.419f
C8580 X1.X1.X2.X1.X2.X2.X3.vin2 vdd 0.761f
C8581 X1.X1.X2.X2.vrefh d2 0.173f
C8582 X1.X1.X1.X1.X2.X1.X1.vin1 X1.X1.X1.X1.X2.X1.X1.vin2 0.668f
C8583 X1.X2.X2.X2.X2.vrefh d3 6.65e-20
C8584 X1.X1.X3.vin1 a_8486_5016# 8.66e-20
C8585 a_35312_892# X2.X3.vin1 0.461f
C8586 a_31476_32788# X2.X1.X1.X1.X1.X1.X2.vin1 1.78e-19
C8587 d4 a_19722_18540# 0.256f
C8588 X2.X2.X1.X1.X1.X2.X2.vin1 X2.X2.X1.X1.X2.vrefh 0.564f
C8589 X2.X1.X2.X1.X2.X1.X3.vin1 a_40352_11734# 0.354f
C8590 a_54606_21264# X2.X2.X2.X2.X1.X1.X2.vin1 0.402f
C8591 a_8186_29834# vdd 0.477f
C8592 a_2196_15634# a_2582_15634# 0.419f
C8593 a_11072_32700# d1 2.92e-22
C8594 X2.X1.X2.X2.X2.X2.X3.vin1 X2.X1.X2.X2.X2.X2.vrefh 2.33e-19
C8595 a_16836_23258# d2 0.00464f
C8596 d1 X2.X1.X1.X2.X2.X1.X2.vin1 1.03e-19
C8597 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X1.X2.X3.vin1 0.587f
C8598 a_4782_20446# d1 0.0749f
C8599 X1.X2.X2.X1.X1.X1.X3.vin1 vdd 1.03f
C8600 X1.X2.X1.X2.X1.X2.vout X1.X2.X1.X2.X1.X2.X3.vin2 0.075f
C8601 d3 a_19336_10916# 0.621f
C8602 a_25326_17452# a_25326_15546# 0.00198f
C8603 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 0.242f
C8604 a_25326_9828# a_23126_8828# 4.77e-21
C8605 d3 a_52492_22210# 7.7e-20
C8606 X2.X1.X2.X2.X1.X2.X1.vin2 X2.X1.X2.X2.X1.X2.vrefh 0.1f
C8607 X2.X2.X1.X3.vin2 a_48702_16634# 5.21e-19
C8608 a_49002_18540# X2.X2.X1.X2.X1.X1.X3.vin2 3.49e-19
C8609 a_10686_23170# vdd 0.553f
C8610 X1.X1.X1.X1.X2.X2.X3.vin1 X1.X1.X1.X1.X2.X2.X3.vin2 0.587f
C8611 a_52792_31700# X2.X2.X2.X2.X2.X2.X3.vin2 0.101f
C8612 d0 a_2582_4198# 0.049f
C8613 a_48316_24258# a_48702_24258# 0.419f
C8614 d2 X2.X2.X1.X1.X1.X2.vrefh 6.65e-20
C8615 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X2.vout 0.0857f
C8616 a_25326_13640# d1 0.00148f
C8617 a_39966_26982# d1 3.95e-19
C8618 X1.X1.X1.X2.X1.X1.X2.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 0.234f
C8619 X1.X2.X1.X1.X1.X1.X3.vin1 a_19036_31882# 0.199f
C8620 X2.X2.X3.vin1 a_52106_6962# 6.45e-19
C8621 d2 X2.X1.X1.X2.X1.X2.X1.vin2 0.226f
C8622 X1.X1.X2.X1.X1.X1.X2.vin1 a_11072_4110# 1.78e-19
C8623 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.X1.vin1 2.23e-19
C8624 X2.X2.X1.X2.X2.vrefh X2.X2.X1.X2.X2.X1.X1.vin1 0.267f
C8625 a_4696_18540# vdd 1.05f
C8626 X2.X1.X1.X1.X1.X2.X2.vin1 a_31862_27070# 0.402f
C8627 X1.X2.X2.X3.vin2 d1 0.0129f
C8628 a_49002_22312# X2.X2.X1.X1.X2.X2.X3.vin1 0.00874f
C8629 a_31862_28976# d1 3.41e-19
C8630 a_49002_26164# d2 7.13e-19
C8631 a_2196_23258# a_2582_23258# 0.419f
C8632 a_23212_10734# d1 0.0126f
C8633 d2 X1.X2.X1.X2.X1.X2.X3.vin1 0.155f
C8634 X2.X2.X1.X1.X3.vin2 a_48616_22312# 0.363f
C8635 d2 a_46116_28976# 0.00351f
C8636 X2.X2.X2.X1.X1.X1.X1.vin1 a_54992_4110# 0.195f
C8637 a_33976_14688# X2.X1.X1.X2.X1.X2.X3.vin1 0.00329f
C8638 a_2196_6104# a_2582_6104# 0.419f
C8639 X1.X2.X3.vin2 a_23126_12640# 2.33e-19
C8640 X1.X1.X1.X2.X2.X1.X3.vin2 a_5082_7064# 0.00815f
C8641 X1.X2.X1.X1.X1.X1.X3.vin1 vdd 1.06f
C8642 d0 X2.X1.X1.X2.X2.X1.X3.vin2 4.34e-19
C8643 d3 X2.X1.X3.vin2 0.77f
C8644 a_2196_8010# a_2582_8010# 0.419f
C8645 X1.X2.X1.X2.X1.X1.X1.vin1 d1 0.011f
C8646 d3 a_48316_24258# 0.00178f
C8647 X1.X1.X1.X1.X2.X1.X2.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 0.234f
C8648 X1.X1.X2.X1.X2.X2.X3.vin1 X1.X1.X2.X1.X3.vin2 1.42e-20
C8649 d2 a_31862_17540# 0.00309f
C8650 d2 X2.X1.X2.X1.X2.X1.vout 0.00174f
C8651 X1.X1.X2.X2.X1.X2.X2.vin1 vdd 0.576f
C8652 d0 X1.X1.X2.X1.X2.X2.X1.vin2 0.276f
C8653 X1.X1.X2.X2.X2.X1.X3.vin2 X1.X1.X2.X2.X2.X2.vrefh 0.161f
C8654 d4 X2.X2.X2.X2.X2.X2.X3.vin2 0.0533f
C8655 a_37466_29834# a_37766_31700# 5.55e-20
C8656 d2 a_54992_11734# 0.00272f
C8657 a_48702_28070# vdd 0.47f
C8658 a_48702_12822# a_49002_10916# 4.41e-20
C8659 X2.X2.X2.X2.X1.X1.vout d4 0.00164f
C8660 a_10686_17452# a_8486_16452# 4.77e-21
C8661 X2.X2.X1.X2.X1.X2.X3.vin2 a_48616_10916# 0.00535f
C8662 d1 a_37766_5016# 0.0752f
C8663 a_2196_28976# a_2582_28976# 0.419f
C8664 a_34362_22312# d2 0.0191f
C8665 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X3.vin1 0.0131f
C8666 X2.X1.X2.X2.X1.X1.vout a_37852_22210# 0.169f
C8667 X3.vin1 vout 0.104f
C8668 X1.X2.X1.X1.X1.X2.X3.vin2 a_17222_27070# 0.567f
C8669 X2.X2.X1.X2.X2.X1.X3.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 0.581f
C8670 d0 a_11072_13640# 0.515f
C8671 a_25326_11734# X1.X2.X2.X1.X1.X2.X3.vin2 8.07e-19
C8672 a_39966_4110# a_40352_4110# 0.419f
C8673 d4 a_49002_29936# 5.68e-19
C8674 X1.X1.X1.X2.X1.X1.X2.vin1 vdd 0.576f
C8675 a_19336_26164# X1.X2.X1.X1.X1.X2.vout 7.93e-20
C8676 X2.X1.X2.X3.vin2 X2.X1.X3.vin2 0.171f
C8677 d2 a_34062_5198# 0.00202f
C8678 X2.X2.X1.X3.vin2 d1 0.0129f
C8679 X1.X1.X1.X1.X3.vin1 d1 0.00179f
C8680 d1 a_8186_6962# 0.0422f
C8681 a_4782_20446# a_5082_18540# 4.41e-20
C8682 X1.X2.X2.X3.vin2 a_23126_24076# 6.03e-19
C8683 d2 X2.X2.X2.X1.X2.X2.X1.vin1 0.0106f
C8684 X1.X2.X1.X1.X1.X2.X1.vin2 d0 0.276f
C8685 X1.X1.X1.X1.X2.X2.X3.vin2 a_4696_18540# 0.00504f
C8686 d0 X1.X1.X2.X1.X1.X2.X1.vin2 0.276f
C8687 X2.X2.X1.X2.X2.vrefh a_46116_11822# 0.118f
C8688 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X1.X3.vin2 1.22e-19
C8689 X1.X2.X2.X1.X2.X2.vrefh X1.X2.X2.X1.X2.X1.X3.vin2 0.161f
C8690 a_31476_23258# X2.X1.X1.X1.X2.X2.X1.vin1 1.64e-19
C8691 a_31862_23258# a_31862_21352# 0.00198f
C8692 a_17222_6104# X1.X2.X1.X2.X2.X1.X3.vin2 8.07e-19
C8693 X1.X1.X1.X1.X1.X2.X3.vin1 d0 4.36e-19
C8694 a_16836_25164# a_16836_23258# 0.00396f
C8695 a_34362_29936# X2.X1.X1.X1.X1.X2.vout 0.254f
C8696 a_37466_25982# a_38152_24076# 3.08e-19
C8697 X2.X2.X1.X2.X2.X2.vout X2.X2.X1.X2.X3.vin2 0.0866f
C8698 a_40352_17452# a_40352_15546# 0.00396f
C8699 a_2196_30882# a_2582_30882# 0.419f
C8700 d2 a_46502_8010# 0.00665f
C8701 X1.X2.X1.X2.X1.X1.vout X1.X2.X1.X2.X1.X1.X3.vin2 0.342f
C8702 a_10686_6016# a_8486_5016# 4.77e-21
C8703 a_39966_23170# d2 0.00479f
C8704 d4 X2.X1.X2.X3.vin1 0.0865f
C8705 a_54606_13640# a_54992_13640# 0.419f
C8706 X1.X1.X2.X2.X2.X2.X1.vin2 d0 0.253f
C8707 a_37466_6962# a_37852_6962# 0.419f
C8708 X2.X1.X2.X2.X1.X1.X1.vin1 X2.X2.X1.X2.vrefh 0.00437f
C8709 X2.X1.X1.X1.X1.X1.X1.vin1 d1 1.51e-19
C8710 X1.X2.X2.X1.X1.X1.X1.vin1 a_25712_4110# 0.195f
C8711 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X1.vin2 8.93e-19
C8712 X1.X2.X2.X1.X1.X2.X2.vin1 a_25326_7922# 8.88e-20
C8713 a_33976_29936# vdd 1.05f
C8714 a_46116_13728# X2.X2.X1.X2.X1.X2.X3.vin1 0.354f
C8715 X1.X2.X1.X1.X2.X2.X3.vin1 a_19422_20446# 0.42f
C8716 a_31862_27070# X2.X1.X1.X1.X2.X1.X1.vin1 8.22e-20
C8717 a_46502_13728# X2.X2.X1.X2.X1.X2.X1.vin1 0.417f
C8718 X1.X1.X1.X1.X2.X1.vout d2 0.00174f
C8719 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X3.vin2 2.23e-19
C8720 d0 a_46502_15634# 0.0489f
C8721 X2.X1.X2.X1.X2.X2.vout X2.X1.X2.X1.X3.vin2 0.0866f
C8722 d2 a_33676_16634# 3.82e-19
C8723 a_37466_10734# a_38152_8828# 3.08e-19
C8724 X2.X2.X1.X1.X2.X2.vrefh d0 0.848f
C8725 X2.X1.X1.X2.X2.vrefh a_31862_11822# 0.3f
C8726 a_38152_12640# a_39966_11734# 1.06e-19
C8727 X2.X2.X1.X3.vin2 X2.X2.X3.vin2 3.82e-19
C8728 a_52106_18358# X2.X2.X2.X3.vin1 0.374f
C8729 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X1.vin2 0.076f
C8730 a_37852_10734# a_39966_9828# 4.72e-20
C8731 X2.X1.X1.X1.X2.X1.X3.vin2 a_33976_22312# 0.00546f
C8732 d2 X2.X2.X2.X1.X1.X2.X3.vin2 0.121f
C8733 X1.X1.X2.X3.vin1 X1.X1.X2.X1.X3.vin2 0.418f
C8734 X1.X1.X3.vin2 X1.X1.X2.X1.X2.X1.vout 3.2e-19
C8735 a_54606_30794# X2.X2.X2.X2.X2.X2.X2.vin1 8.88e-20
C8736 X2.X2.X2.X2.X2.X2.X1.vin2 X2.X2.X2.X2.X2.X2.X3.vin2 8.93e-19
C8737 X2.X2.X2.X2.X2.X1.X2.vin1 X2.X2.X2.X2.X2.X1.X3.vin2 0.234f
C8738 d2 X2.X2.X2.X2.X2.X2.X1.vin1 9.24e-20
C8739 X1.X2.X1.X1.X2.X1.vout X1.X2.X1.X1.X2.X1.X3.vin2 0.326f
C8740 d0 a_25326_11734# 0.0675f
C8741 a_13696_892# a_14082_892# 0.419f
C8742 d1 X1.X1.X2.X1.X1.X2.vrefh 0.0738f
C8743 X2.X1.X2.X2.X2.X1.X3.vin2 X2.X1.X2.X2.X2.X2.X1.vin1 5.19e-19
C8744 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.X3.vin1 0.587f
C8745 X2.X2.X1.X1.X2.X2.X3.vin1 d1 0.146f
C8746 a_31476_23258# d0 0.515f
C8747 a_37466_25982# a_37852_25982# 0.414f
C8748 X2.X1.X2.X2.X2.vrefh d2 0.158f
C8749 a_22826_18358# vdd 0.476f
C8750 d3 a_22826_22210# 0.0474f
C8751 X1.X2.X3.vin1 a_20672_892# 0.386f
C8752 a_19036_28070# d3 0.00108f
C8753 X2.X2.X2.X2.X1.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X1.vin1 2.23e-19
C8754 X1.X2.X2.X1.X2.X2.X3.vin1 a_23212_14586# 0.00329f
C8755 X2.X2.X2.X2.X1.X2.X2.vin1 a_54992_23170# 1.78e-19
C8756 a_10686_9828# X1.X1.X2.X1.X1.X2.X1.vin2 8.88e-20
C8757 X2.X2.X1.X2.X3.vin2 d1 0.00807f
C8758 a_11072_6016# X1.X1.X2.X1.X1.X1.X1.vin2 1.78e-19
C8759 X1.X2.X1.X2.X2.X1.vout X1.X2.X1.X2.X2.X1.X3.vin2 0.326f
C8760 a_52792_27888# a_52106_29834# 2.86e-19
C8761 d4 X1.X1.X1.X1.X1.X2.X3.vin2 0.0533f
C8762 a_52492_25982# X2.X2.X2.X2.X2.X1.vout 1.64e-19
C8763 a_31862_27070# d2 0.00792f
C8764 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X3.vin2 0.17f
C8765 X2.X1.X1.X1.X1.X2.X3.vin2 d1 0.171f
C8766 a_37766_27888# a_38152_27888# 0.419f
C8767 d3 a_19722_29936# 0.00177f
C8768 a_4696_14688# a_4396_12822# 6.71e-19
C8769 d3 X1.X1.X2.X2.X2.X2.X3.vin1 0.0137f
C8770 X2.X2.X1.X2.X1.X1.X3.vin1 X2.X2.X1.X2.X1.X1.X1.vin2 0.216f
C8771 a_11072_28888# d1 2.92e-22
C8772 X2.X1.X2.X1.X3.vin2 d1 0.00807f
C8773 X1.X1.X1.X2.vrefh a_2196_17540# 1.64e-19
C8774 d2 a_2582_13728# 0.00479f
C8775 d2 a_33676_31882# 0.0017f
C8776 a_37466_25982# d4 3.58e-19
C8777 a_46502_30882# d0 0.0489f
C8778 d3 a_37766_12640# 0.00195f
C8779 d0 X2.X1.X1.X2.X2.X1.X1.vin1 0.267f
C8780 d2 X1.X1.X2.X2.X2.X1.X2.vin1 0.0318f
C8781 X2.X2.X1.X2.X1.X2.X1.vin2 vdd 0.361f
C8782 d0 X1.X2.X2.X1.X1.X2.X1.vin2 0.276f
C8783 X2.X1.X2.X3.vin1 a_37766_8828# 1.64e-19
C8784 a_10686_11734# X1.X1.X2.X1.X2.vrefh 8.22e-20
C8785 X1.X2.X2.X1.X2.vrefh a_25712_9828# 0.118f
C8786 X2.X1.X1.X1.X2.X1.X1.vin2 a_31862_23258# 8.88e-20
C8787 X2.X1.X1.X2.X1.X2.X1.vin2 a_31862_11822# 8.88e-20
C8788 X1.X1.X2.X1.X3.vin2 X1.X1.X2.X1.X2.X1.X3.vin2 0.0533f
C8789 X2.X1.X1.X2.X1.X2.X3.vin1 vdd 0.96f
C8790 X2.X1.X2.X2.X1.X2.vrefh a_40352_21264# 0.118f
C8791 a_52106_6962# X2.X2.X2.X1.X1.X2.X3.vin2 3.85e-19
C8792 X2.X2.X2.X1.X1.X1.X3.vin2 a_54992_6016# 0.354f
C8793 d3 X1.X1.X2.X3.vin1 0.676f
C8794 X2.X1.X2.X2.X1.X1.X2.vin1 d0 0.262f
C8795 X2.X1.X1.X1.X3.vin1 X2.X1.X1.X1.X1.X1.vout 0.13f
C8796 X2.X2.X1.X1.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X1.X1.vin2 0.216f
C8797 X2.X1.X1.X2.X1.X2.X3.vin1 a_34062_12822# 0.42f
C8798 X2.X1.X1.X2.X1.X2.X1.vin1 X2.X1.X1.X2.X1.X2.X3.vin2 2.23e-19
C8799 X2.X2.X2.X3.vin1 a_52106_10734# 0.509f
C8800 X2.X2.X3.vin2 X2.X2.X1.X2.X3.vin2 0.00254f
C8801 X1.X2.X2.X1.X2.X2.X1.vin2 a_25712_15546# 0.12f
C8802 a_25326_15546# X1.X2.X2.X1.X2.X2.X1.vin1 0.417f
C8803 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X3.vin1 0.206f
C8804 a_10686_26982# d2 0.00328f
C8805 X2.X2.X2.X2.X1.X1.X1.vin1 X2.X2.X2.X2.vrefh 0.267f
C8806 X1.X2.X1.X1.X2.X2.vout d4 6.02e-19
C8807 X2.X2.X2.X2.X1.X2.vrefh d2 0.177f
C8808 a_54606_26982# X2.X2.X2.X2.X1.X2.X3.vin2 8.07e-19
C8809 a_22826_22210# X1.X2.X2.X2.X1.X1.vout 0.387f
C8810 a_52106_22210# a_52792_20264# 2.86e-19
C8811 X1.X2.X1.X1.X1.X1.vout X1.X2.X1.X1.X1.X1.X3.vin2 0.342f
C8812 X2.X2.X1.X2.X1.X1.X1.vin2 X2.X2.X1.X2.X1.X2.vrefh 0.076f
C8813 a_19036_28070# a_19422_28070# 0.419f
C8814 X1.X2.X1.X1.X1.X2.X2.vin1 X1.X2.X1.X1.X1.X2.X3.vin2 0.234f
C8815 a_46502_17540# vdd 0.553f
C8816 a_19036_24258# d1 0.521f
C8817 a_52792_16452# a_52106_14586# 3.31e-19
C8818 d4 a_2582_17540# 0.00112f
C8819 a_4396_5198# vdd 1.05f
C8820 a_4696_26164# X1.X1.X1.X1.X3.vin1 0.169f
C8821 X1.X2.X3.vin1 d1 0.0876f
C8822 a_11072_6016# X1.X1.X2.X1.X1.X2.X1.vin1 1.64e-19
C8823 X1.X2.X2.X3.vin2 X1.X2.X2.X3.vin1 0.559f
C8824 a_19422_28070# a_19722_29936# 5.55e-20
C8825 X1.X2.X3.vin2 X1.X2.X2.X1.X3.vin1 0.0361f
C8826 a_48702_20446# a_46502_19446# 4.77e-21
C8827 X2.X2.X1.X1.X2.X2.X3.vin2 a_46116_19446# 0.354f
C8828 X1.X2.X2.X3.vin1 a_23212_10734# 0.356f
C8829 a_52106_29834# vdd 0.477f
C8830 X1.X1.X1.X1.X2.X1.X3.vin2 d1 0.15f
C8831 a_23126_27888# vdd 0.561f
C8832 X1.X1.X2.X1.X1.X1.X3.vin1 a_10686_4110# 0.52f
C8833 a_37466_6962# a_37766_5016# 4.19e-20
C8834 a_25326_7922# X1.X2.X2.X1.X1.X1.X3.vin2 8.07e-19
C8835 a_8572_14586# vdd 1.05f
C8836 X2.X2.X2.X2.X1.X2.X2.vin1 d1 1.03e-19
C8837 d0 X2.X2.X1.X2.X1.X2.X2.vin1 0.262f
C8838 a_19722_29936# X1.X2.X1.X1.X3.vin1 0.434f
C8839 X2.X2.X2.X2.X1.X2.X1.vin1 d0 0.267f
C8840 X1.X2.X1.X1.X2.X2.X1.vin2 X1.X2.X1.X1.X2.X2.X2.vin1 0.242f
C8841 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X1.X3.vin1 0.0321f
C8842 d2 a_48316_9010# 0.00167f
C8843 a_8486_8828# a_10686_7922# 4.2e-20
C8844 d3 X1.X1.X2.X1.X2.X1.X3.vin2 2.81e-19
C8845 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.X1.vin2 0.216f
C8846 a_16836_8010# a_17222_8010# 0.419f
C8847 a_37766_16452# a_37852_14586# 3.38e-19
C8848 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.X1.vin2 0.216f
C8849 X1.X2.X3.vin2 a_19722_14688# 2.04e-19
C8850 X2.X2.X1.X1.X2.X2.vrefh a_46116_23258# 0.118f
C8851 X1.X2.X1.X1.X3.vin2 a_19422_20446# 9.7e-20
C8852 X2.X2.X1.X1.X1.X2.X1.vin1 X2.X2.X1.X1.X1.X2.vrefh 0.267f
C8853 a_4696_29936# X1.X1.X1.X1.X1.X1.vout 0.169f
C8854 a_5082_29936# a_4782_31882# 4.19e-20
C8855 d0 a_20286_892# 2.73e-19
C8856 d3 X1.X2.X1.X1.X1.X2.X3.vin1 0.0105f
C8857 a_52792_16452# vdd 1.05f
C8858 a_48616_18540# vdd 1.05f
C8859 X2.X2.X1.X2.X2.X2.X3.vin1 a_48702_5198# 0.42f
C8860 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X3.vin2 2.23e-19
C8861 d3 a_8186_25982# 0.292f
C8862 a_4696_7064# vdd 1.05f
C8863 a_19336_7064# a_19422_5198# 3.38e-19
C8864 a_19722_7064# a_19036_5198# 3.31e-19
C8865 X1.X2.X2.X1.X1.X2.X2.vin1 d1 1.03e-19
C8866 a_37766_12640# X2.X1.X2.X1.X2.X1.X3.vin1 0.428f
C8867 a_25326_23170# a_23212_22210# 2.68e-20
C8868 X2.X1.X1.X2.X1.X2.X2.vin1 X2.X1.X1.X2.X2.vrefh 0.564f
C8869 a_8486_16452# X1.X1.X2.X1.X2.X2.vout 0.418f
C8870 d2 a_39966_9828# 0.00792f
C8871 X2.X1.X1.X3.vin2 X2.X1.X2.X3.vin1 1.22e-19
C8872 a_33676_20446# a_31862_19446# 1.15e-20
C8873 X1.X1.X2.X1.X1.X1.X1.vin2 vdd 0.387f
C8874 X2.X1.X3.vin1 X2.X1.X3.vin2 3.25f
C8875 a_38152_20264# a_37466_18358# 2.97e-19
C8876 a_46116_28976# X2.X2.X1.X1.X1.X2.X1.vin1 0.195f
C8877 X1.X1.X2.X2.X2.vrefh X1.X2.X1.X1.X2.X1.X1.vin1 0.00437f
C8878 a_52106_10734# X2.X2.X2.X1.X3.vin1 0.385f
C8879 a_38152_24076# vdd 1.05f
C8880 d0 X1.X2.X1.X2.X1.X2.X3.vin2 4.34e-19
C8881 a_31862_21352# d1 3.41e-19
C8882 a_54992_25076# X2.X2.X2.X2.X1.X2.X1.vin2 1.78e-19
C8883 a_52492_22210# X2.X2.X2.X2.X1.X1.X3.vin2 0.00546f
C8884 X1.X2.X2.X2.X1.X1.X3.vin2 a_25712_21264# 0.354f
C8885 d3 X2.X1.X2.X2.X2.X1.vout 0.0421f
C8886 d4 a_19036_16634# 0.00176f
C8887 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X2.X3.vin2 8.93e-19
C8888 a_8872_8828# vdd 1.05f
C8889 a_37466_14586# X2.X1.X2.X1.X2.X1.X3.vin2 0.00815f
C8890 a_46116_21352# d2 0.00274f
C8891 d3 a_4696_14688# 7.7e-20
C8892 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X3.vin1 0.206f
C8893 d0 X2.X2.X1.X2.X2.X2.X1.vin2 0.276f
C8894 a_46116_25164# d0 0.518f
C8895 a_22826_25982# X1.X2.X2.X3.vin2 0.452f
C8896 a_2196_6104# a_2196_4198# 0.00396f
C8897 a_19722_26164# d1 0.0318f
C8898 X2.X2.X1.X1.X3.vin1 a_48702_31882# 1.52e-19
C8899 X1.X1.X2.X2.X2.X1.X1.vin1 a_11072_25076# 1.64e-19
C8900 X2.X2.X1.X2.X1.X2.vout a_48616_10916# 7.93e-20
C8901 a_2196_11822# vdd 1.05f
C8902 a_49002_29936# X2.X2.X1.X1.X1.X1.vout 0.386f
C8903 d2 a_37852_10734# 0.0057f
C8904 d0 X2.X1.X1.X2.X2.X2.X3.vin1 4.36e-19
C8905 a_22826_10734# a_23212_10734# 0.414f
C8906 a_25326_26982# a_23212_25982# 5.36e-21
C8907 d4 X1.X1.X1.X2.X1.X1.X3.vin2 4.77e-19
C8908 a_8486_24076# X1.X1.X2.X2.X1.X2.vout 0.418f
C8909 a_54606_26982# d0 0.0675f
C8910 a_19036_12822# a_17222_11822# 1.15e-20
C8911 X2.X1.X1.X1.X1.X2.X2.vin1 d2 0.0329f
C8912 a_34062_16634# a_31862_15634# 4.77e-21
C8913 X2.X1.X2.X1.X2.X2.X2.vin1 a_40352_17452# 0.197f
C8914 X1.X2.X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.vrefh 0.161f
C8915 d0 a_49952_892# 3.19e-19
C8916 X1.X1.X1.X1.X1.X1.X1.vin2 X1.X1.X1.X1.X1.X1.X3.vin2 8.93e-19
C8917 a_17222_27070# X1.X2.X1.X1.X1.X2.X1.vin2 8.88e-20
C8918 a_25326_30794# X1.X2.X2.X2.X2.X2.X1.vin1 0.417f
C8919 X1.X2.X2.X2.X2.X2.X1.vin2 a_25712_30794# 0.12f
C8920 a_23126_16452# vdd 0.471f
C8921 X1.X1.X1.X1.X1.X1.X1.vin2 vdd 0.399f
C8922 a_52792_31700# vdd 1.05f
C8923 X2.X1.X2.X2.X3.vin1 X2.X1.X2.X2.X3.vin2 0.552f
C8924 d4 X2.X2.X2.X1.X2.X2.X2.vin1 8.68e-20
C8925 X2.X2.X2.X1.X1.X1.vout X2.X2.X2.X1.X1.X1.X3.vin2 0.342f
C8926 X2.X2.X1.X1.X3.vin1 d1 0.00179f
C8927 X1.X1.X1.X2.X1.X1.X1.vin2 a_2582_15634# 8.88e-20
C8928 d3 a_34362_18540# 0.0469f
C8929 X1.X1.X3.vin2 a_8486_8828# 2.33e-19
C8930 a_31862_17540# X2.X1.X1.X2.X1.X1.X3.vin1 0.52f
C8931 X1.X1.X2.X1.X2.X2.X1.vin1 vdd 0.592f
C8932 a_19036_20446# a_17222_19446# 1.15e-20
C8933 X2.X2.X2.X1.X1.X2.X3.vin2 a_52792_8828# 0.101f
C8934 d0 a_16836_9916# 0.518f
C8935 a_48702_5198# X2.X2.X1.X2.X2.X2.X3.vin2 0.277f
C8936 X1.X1.X2.X1.X2.X1.vout d1 0.0238f
C8937 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X1.X2.X1.vin1 2.23e-19
C8938 a_19422_28070# X1.X2.X1.X1.X1.X2.X3.vin1 0.42f
C8939 a_4696_22312# d1 0.00613f
C8940 X1.X1.X1.X1.X3.vin2 d4 0.0401f
C8941 X1.X2.X1.X2.X2.X2.vrefh vdd 0.415f
C8942 d4 a_40352_32700# 1.8e-19
C8943 X2.X2.X2.X1.X2.X1.X1.vin1 X2.X2.X2.X1.X2.vrefh 0.267f
C8944 a_34062_28070# X2.X1.X1.X1.X3.vin1 9.54e-19
C8945 X2.X1.X1.X1.X1.X2.X3.vin2 a_34362_29936# 3.85e-19
C8946 X2.X2.X2.X2.X1.X1.X3.vin1 X2.X2.X2.X1.X2.X2.X3.vin2 1.22e-19
C8947 a_37852_25982# vdd 1.05f
C8948 a_17222_13728# vdd 0.553f
C8949 X2.X1.X1.X2.X1.X2.X1.vin2 X2.X1.X1.X2.X1.X2.X2.vin1 0.242f
C8950 d3 a_39966_32700# 1.28e-19
C8951 a_5082_22312# X1.X1.X1.X1.X2.X2.X3.vin1 0.00874f
C8952 X2.X1.X1.X1.X2.X2.X3.vin1 a_31862_19446# 0.00207f
C8953 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 0.242f
C8954 a_54606_17452# a_54606_15546# 0.00198f
C8955 a_46116_6104# X2.X2.X1.X2.X2.X2.X1.vin2 0.12f
C8956 a_23126_8828# vdd 0.47f
C8957 X1.X2.X1.X1.X2.X2.X1.vin2 d0 0.276f
C8958 d6 X3.vin1 2.49f
C8959 d0 X1.X1.X1.X1.X1.X1.X2.vin1 0.262f
C8960 d5 a_28482_892# 4.95e-19
C8961 X1.X2.X1.X2.X2.X1.vout a_19722_7064# 0.383f
C8962 X2.X1.X2.X2.X1.X2.X2.vin1 a_40352_25076# 0.197f
C8963 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X2.X3.vin1 0.0174f
C8964 X1.X2.X2.X2.X2.X1.X2.vin1 vdd 0.576f
C8965 a_39966_6016# X2.X1.X2.X1.X1.X1.X3.vin2 0.567f
C8966 X1.X1.X2.X1.X1.X2.X1.vin1 vdd 0.592f
C8967 X1.X1.X1.X1.X2.X2.X3.vin1 d0 4.36e-19
C8968 X1.X2.X1.X2.X2.vrefh a_16836_9916# 1.64e-19
C8969 a_25712_26982# d0 0.518f
C8970 X1.X2.X1.X1.X2.X1.X3.vin2 a_17222_21352# 8.07e-19
C8971 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin1 0.52f
C8972 X2.X1.X1.X2.X2.X1.X3.vin1 a_31862_8010# 0.00207f
C8973 a_2582_25164# X1.X1.X1.X1.X2.X1.X2.vin1 8.88e-20
C8974 d2 a_22826_6962# 0.272f
C8975 X2.X1.X1.X2.X2.X2.vrefh a_31476_6104# 1.64e-19
C8976 a_40352_19358# d2 0.00256f
C8977 d0 X2.X2.X1.X1.X1.X1.X1.vin1 0.0488f
C8978 d3 X2.X2.X1.X2.X2.X1.X1.vin1 6.34e-20
C8979 a_37852_18358# a_39966_17452# 4.72e-20
C8980 a_25712_17452# vdd 1.05f
C8981 d4 X1.X1.X1.X1.X1.X1.X3.vin2 0.0533f
C8982 a_19336_29936# X1.X2.X1.X1.X1.X1.X3.vin2 0.00546f
C8983 X2.X1.X1.X2.X2.X1.vout X2.X1.X1.X2.X2.X1.X3.vin2 0.326f
C8984 a_52106_10734# a_52406_8828# 4.41e-20
C8985 d4 vdd 4.64f
C8986 a_54606_11734# vdd 0.553f
C8987 a_23212_22210# vdd 1.05f
C8988 X2.X1.X1.X2.X1.X2.vrefh d1 0.0071f
C8989 a_23126_31700# vdd 0.471f
C8990 a_10686_32700# a_11072_32700# 0.419f
C8991 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X1.X3.vin2 0.0533f
C8992 X2.X2.X2.X2.X1.X1.X1.vin2 d0 0.276f
C8993 X1.X1.X1.X2.X2.X2.X1.vin1 a_2196_8010# 1.64e-19
C8994 a_2582_6104# a_2582_8010# 0.00198f
C8995 a_25712_19358# d2 0.00256f
C8996 X1.X1.X2.X2.X2.X2.X1.vin1 vdd 0.592f
C8997 a_2582_32788# X1.X1.X1.X1.X1.X1.X1.vin1 0.42f
C8998 a_2196_32788# X1.X1.X1.X1.X1.X1.X3.vin1 0.354f
C8999 X2.X2.X2.X1.X2.X2.X1.vin2 X2.X2.X2.X1.X2.X2.vrefh 0.1f
C9000 a_8572_18358# d2 0.0113f
C9001 X1.X1.X2.X1.X2.X2.X3.vin2 d0 4.34e-19
C9002 a_34362_7064# X2.X1.X1.X2.X2.X2.vout 0.263f
C9003 X2.X1.X1.X2.X2.X2.X2.vin1 vdd 0.578f
C9004 a_8486_31700# X1.X1.X2.X2.X2.X2.vout 0.418f
C9005 a_17222_15634# d1 0.00148f
C9006 X1.X2.X1.X1.X1.X2.vout vdd 0.696f
C9007 d1 a_40352_6016# 2.92e-22
C9008 X1.X1.X1.X2.X2.vrefh d1 0.00745f
C9009 X2.X2.X2.X1.X2.X2.X1.vin2 vdd 0.36f
C9010 X2.X1.X1.X1.X2.X1.X1.vin2 d1 4.01e-19
C9011 d3 a_33976_26164# 0.621f
C9012 X2.X1.X1.X2.X1.X1.X3.vin1 a_33676_16634# 0.199f
C9013 X1.X1.X2.X2.X1.X1.X3.vin2 X1.X1.X2.X2.X1.X1.X1.vin1 2.23e-19
C9014 X2.X1.X2.X2.X2.X1.X3.vin2 X2.X1.X2.X2.X2.X2.vrefh 0.161f
C9015 X1.X1.X2.X2.X1.X1.X2.vin1 a_11072_19358# 1.78e-19
C9016 X2.X1.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X3.vin2 0.0533f
C9017 a_23126_5016# a_25326_4110# 4.2e-20
C9018 X1.X2.X2.X1.X1.X1.X3.vin1 X1.X2.X2.X1.X1.X1.X1.vin2 0.22f
C9019 d1 X1.X2.X2.X1.X1.X1.X3.vin2 0.154f
C9020 X1.X2.X1.X1.X2.X1.X3.vin1 d1 0.151f
C9021 d0 X1.X2.X2.X1.X1.X1.X3.vin1 4.36e-19
C9022 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.vout 0.2f
C9023 a_49002_18540# X2.X2.X1.X3.vin2 0.233f
C9024 X1.X1.X2.X1.X1.X2.X2.vin1 a_11072_9828# 0.197f
C9025 d2 X2.X1.X2.X1.X1.X1.X2.vin1 6e-20
C9026 a_11072_19358# d2 0.00256f
C9027 X2.X2.X1.X2.X2.X2.X1.vin2 X2.X2.X1.X2.X2.X2.X2.vin1 0.242f
C9028 X2.X2.X1.X1.X2.X1.X2.vin1 X2.X2.X1.X1.X2.X2.vrefh 0.564f
C9029 X2.X1.X1.X1.X2.X1.X1.vin1 d2 0.0105f
C9030 a_8486_24076# a_8186_22210# 5.55e-20
C9031 a_10686_23170# d0 0.0675f
C9032 X2.X2.X2.X1.X2.vrefh X2.X2.X2.X1.X1.X2.X2.vin1 0.564f
C9033 X1.X2.X2.vrefh X1.X3.vin1 0.00136f
C9034 X1.X1.X3.vin1 a_8186_14586# 2.24e-19
C9035 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.vout 0.197f
C9036 a_25712_11734# vdd 1.05f
C9037 X2.X1.X1.X2.vrefh X1.X2.X2.X2.vrefh 0.117f
C9038 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin1 0.52f
C9039 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X1.X2.X1.vin2 0.216f
C9040 X2.X1.X3.vin1 a_37766_12640# 8.66e-20
C9041 d3 a_22826_14586# 9.23e-19
C9042 X1.X1.X1.X2.X2.X1.X1.vin2 d1 4.01e-19
C9043 X1.X2.vrefh d4 0.00449f
C9044 a_31476_28976# a_31476_30882# 0.00396f
C9045 X1.X2.X1.X2.X1.X1.X1.vin2 X1.X2.X1.X2.X1.X1.X3.vin2 8.93e-19
C9046 a_34062_31882# a_31862_30882# 4.77e-21
C9047 X2.X1.X2.X2.X3.vin1 d1 0.00179f
C9048 a_39966_23170# a_40352_23170# 0.419f
C9049 X2.X1.X1.X1.X1.X2.vrefh d1 0.0738f
C9050 X1.X1.X1.X1.X2.X2.X3.vin2 d4 0.0265f
C9051 a_4396_24258# vdd 1.05f
C9052 X2.X1.X2.X1.X2.vrefh a_39966_9828# 0.3f
C9053 X1.X1.X2.X1.X2.X1.vout a_8486_12640# 0.422f
C9054 X2.X2.X2.X2.X3.vin1 a_52492_22210# 0.363f
C9055 X2.X2.X3.vin1 X2.X2.X1.X2.X2.X1.vout 0.0215f
C9056 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X1.vout 0.0524f
C9057 d2 X1.X1.X1.X2.X2.X1.X1.vin1 0.0105f
C9058 X1.X1.X2.X1.X1.X2.vout a_8572_6962# 0.0929f
C9059 X1.X2.X3.vin1 X1.X2.X2.X3.vin1 3.45e-19
C9060 a_11072_32700# a_11072_30794# 0.00396f
C9061 a_46116_25164# a_46116_23258# 0.00396f
C9062 a_11072_21264# d1 2.92e-22
C9063 a_46502_13728# a_46502_11822# 0.00198f
C9064 a_16836_21352# X1.X2.X1.X1.X2.X2.X1.vin2 0.12f
C9065 X2.X1.X2.X1.X1.X2.X3.vin1 a_37852_6962# 0.00329f
C9066 X2.X2.X2.X1.X2.X1.X3.vin2 a_52406_12640# 0.267f
C9067 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X3.vin1 0.0565f
C9068 X2.X2.X1.X2.X1.X2.X3.vin1 X2.X2.X1.X2.X2.vrefh 0.00118f
C9069 X2.X2.X2.X1.X2.X1.X2.vin1 X2.X2.X2.X1.X2.X1.X3.vin1 0.00117f
C9070 d3 X1.X2.X2.X1.X2.vrefh 6.65e-20
C9071 X1.X2.X1.X1.X1.X1.X3.vin1 d0 4.36e-19
C9072 a_52106_14586# a_52492_14586# 0.419f
C9073 a_54606_9828# vdd 0.542f
C9074 d3 X2.X2.X2.X3.vin1 0.676f
C9075 a_17222_30882# d1 0.00148f
C9076 a_10686_21264# X1.X1.X2.X2.X1.X1.X3.vin2 0.567f
C9077 d3 a_52792_24076# 0.00108f
C9078 X2.X2.X2.X2.X2.X2.X1.vin2 vdd 0.387f
C9079 a_37766_8828# vdd 0.47f
C9080 a_2582_27070# a_2582_25164# 0.00198f
C9081 X1.X1.X2.X2.X1.X1.X2.vin1 d2 0.031f
C9082 a_34362_14688# d1 0.0422f
C9083 X1.X2.X2.X1.X2.X1.X3.vin1 a_23512_12640# 0.199f
C9084 X1.X1.X2.X2.X1.X2.X2.vin1 d0 0.262f
C9085 X1.X1.X1.X1.X3.vin2 X1.X1.X2.X3.vin2 7.46e-20
C9086 X1.X2.X1.X1.X2.X1.X1.vin2 X1.X2.X1.X1.X2.X1.X3.vin2 8.93e-19
C9087 d2 a_8186_10734# 7.13e-19
C9088 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X1.vin2 8.93e-19
C9089 a_8186_25982# X1.X1.X2.X2.X3.vin1 0.372f
C9090 X2.X2.X2.X1.X1.X2.X2.vin1 a_54606_7922# 8.88e-20
C9091 X1.X2.X2.X1.X1.X2.X1.vin1 vdd 0.592f
C9092 X1.X2.X1.X2.vrefh X1.X1.X2.X2.vrefh 0.117f
C9093 X1.X2.X2.X1.X2.X2.X1.vin2 X1.X2.X2.X1.X2.X2.vrefh 0.1f
C9094 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X3.vin1 1.22e-19
C9095 a_33676_16634# X2.X1.X1.X2.X1.X1.vout 0.359f
C9096 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 5.19e-19
C9097 d4 X2.X1.X1.X2.X1.X1.X1.vin2 3.99e-21
C9098 X1.X2.X1.X1.X1.X2.X2.vin1 X1.X2.X1.X1.X1.X2.X1.vin2 0.242f
C9099 a_22826_18358# a_23512_16452# 3.08e-19
C9100 a_25326_17452# X1.X2.X2.X1.X2.X2.X2.vin1 0.402f
C9101 X1.X2.X1.X1.X2.vrefh X1.X1.X2.X2.X2.vrefh 0.117f
C9102 X2.X1.X2.X1.X1.X2.X1.vin2 a_40352_7922# 0.12f
C9103 a_39966_7922# X2.X1.X2.X1.X1.X2.X1.vin1 0.417f
C9104 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X3.vin1 1.22e-19
C9105 d2 a_37852_29834# 0.627f
C9106 d4 X1.X2.X1.X2.X1.X1.X3.vin1 0.0205f
C9107 d3 a_37766_16452# 4.67e-19
C9108 a_39966_11734# d1 3.95e-19
C9109 X1.X1.X1.X2.X1.X1.X1.vin1 d1 0.011f
C9110 d0 X1.X1.X1.X2.X1.X1.X2.vin1 0.262f
C9111 a_31862_25164# X2.X1.X1.X1.X2.X1.X3.vin2 7.84e-19
C9112 X1.X1.X1.X1.X1.X1.X1.vin1 vrefh 0.103f
C9113 a_8872_20264# a_8186_18358# 2.97e-19
C9114 X2.X1.X1.X1.X2.vrefh vdd 0.426f
C9115 a_17222_17540# d2 0.00309f
C9116 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X3.vin1 2.33e-19
C9117 X2.X2.X3.vin1 a_49002_10916# 6.09e-19
C9118 a_10686_25076# a_8486_24076# 4.77e-21
C9119 X1.X2.X2.X1.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X1.vin1 2.23e-19
C9120 a_52492_14586# vdd 1.05f
C9121 X1.X2.X2.X1.X2.X1.X2.vin1 a_25712_11734# 1.78e-19
C9122 a_54606_23170# a_52492_22210# 2.68e-20
C9123 a_52406_16452# d1 0.0749f
C9124 X1.X1.X2.X3.vin2 vdd 0.716f
C9125 X1.X1.X1.X1.X1.X2.X1.vin2 X1.X1.X1.X1.X1.X1.X3.vin2 3.94e-19
C9126 d1 X1.X2.X1.X2.X2.X2.X2.vin1 0.0144f
C9127 X1.X2.X2.X1.X1.X2.vrefh a_25326_6016# 0.3f
C9128 a_16836_6104# d1 2.25e-20
C9129 X1.X2.X2.X2.X1.X2.vout d2 0.00124f
C9130 X1.X1.X1.X1.X1.X2.X1.vin2 vdd 0.361f
C9131 X1.X2.X2.X1.X1.X1.X2.vin1 X2.X1.X1.X2.X2.X2.X1.vin2 0.00232f
C9132 a_31476_6104# a_31862_6104# 0.419f
C9133 X2.X1.X1.X2.X1.X1.X3.vin2 X2.X1.X1.X2.X1.X2.X1.vin1 5.19e-19
C9134 X2.X1.X2.X1.X2.X2.X1.vin1 d1 0.0118f
C9135 X2.X2.X1.X1.X2.X2.vout vdd 0.865f
C9136 X1.X1.X1.X2.X1.X2.X2.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 0.234f
C9137 X2.X2.X1.X1.X2.vrefh a_46116_25164# 1.64e-19
C9138 X1.X1.X2.X2.X2.vrefh vdd 0.426f
C9139 X1.X1.X2.X2.X1.X2.X1.vin1 a_11072_21264# 1.64e-19
C9140 a_4396_12822# a_4782_12822# 0.419f
C9141 a_25326_25076# X1.X2.X2.X2.X1.X2.X2.vin1 0.402f
C9142 X2.X2.X2.X2.X1.X2.vout d4 3.47e-19
C9143 X2.X1.X1.X2.X2.X1.X3.vin1 a_34062_9010# 0.428f
C9144 X2.X1.X2.X2.X1.X1.vout a_37852_18358# 1.64e-19
C9145 X2.X1.X1.X2.vrefh a_31862_17540# 8.22e-20
C9146 a_4696_14688# a_5082_14688# 0.419f
C9147 a_2582_9916# X1.X1.X1.X2.X2.X1.X3.vin2 7.84e-19
C9148 a_17222_21352# a_17222_19446# 0.00198f
C9149 a_8486_20264# a_8872_20264# 0.419f
C9150 X1.X1.X2.X1.X1.X1.X3.vin2 d2 0.0682f
C9151 a_37766_24076# d1 0.0749f
C9152 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X3.vin2 0.17f
C9153 X1.X2.X3.vin1 a_22826_10734# 3.93e-19
C9154 a_8572_29834# a_10686_30794# 2.68e-20
C9155 d3 a_52106_25982# 0.29f
C9156 a_8486_8828# d1 0.0749f
C9157 a_48702_12822# vdd 0.47f
C9158 X1.X2.X2.X2.X1.X2.X1.vin2 X1.X2.X2.X2.X1.X1.X3.vin2 3.94e-19
C9159 X1.X2.X2.X2.X1.X2.X1.vin1 d1 0.0118f
C9160 a_52106_6962# d2 0.272f
C9161 X1.X2.X2.X2.X1.X2.X1.vin1 a_25326_21264# 8.22e-20
C9162 X2.X2.X2.X1.X1.X1.vout a_52792_5016# 0.359f
C9163 d3 X2.X2.X2.X1.X3.vin1 0.0869f
C9164 d1 a_31862_8010# 0.00148f
C9165 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.X3.vin1 0.587f
C9166 d2 a_38152_16452# 6.04e-19
C9167 X2.X2.X2.X2.X1.X2.X3.vin1 X2.X2.X2.X2.X1.X2.vrefh 2.33e-19
C9168 a_19422_12822# a_19336_10916# 3.3e-19
C9169 X2.X1.X2.vrefh d6 4.63e-19
C9170 a_19036_12822# a_19722_10916# 3.08e-19
C9171 X1.X1.X1.X2.X1.X2.X1.vin2 a_2196_11822# 1.78e-19
C9172 a_25712_32700# d1 2.92e-22
C9173 d3 a_37766_31700# 4.75e-19
C9174 a_38152_24076# a_37466_22210# 3.31e-19
C9175 X1.X2.X2.X2.X2.vrefh X1.X2.X2.X2.X1.X2.X3.vin2 0.161f
C9176 X2.X1.X2.X2.X2.X1.X1.vin2 X2.X1.X2.X2.X2.vrefh 0.1f
C9177 a_28482_892# X3.vin2 0.263f
C9178 a_11072_21264# X1.X1.X2.X2.X1.X1.X1.vin2 1.78e-19
C9179 d7 vdd 0.445f
C9180 d7 a_28096_892# 0.502f
C9181 X2.X2.X3.vin2 a_52406_16452# 3.98e-19
C9182 X2.X1.X1.X1.X1.X1.X3.vin1 d4 0.00851f
C9183 d3 a_48616_14688# 7.7e-20
C9184 a_52106_25982# X2.X2.X2.X2.X2.X1.X3.vin2 3.49e-19
C9185 d2 a_8872_12640# 3.82e-19
C9186 a_19422_16634# d1 0.0749f
C9187 X2.X2.X1.X2.X1.X1.vout vdd 0.78f
C9188 a_8872_12640# a_8186_10734# 2.97e-19
C9189 a_34362_10916# X2.X1.X1.X2.X2.X1.X3.vin1 0.00837f
C9190 a_52406_31700# d1 0.0489f
C9191 X2.X1.X1.X3.vin2 vdd 0.716f
C9192 a_10686_15546# a_10686_13640# 0.00198f
C9193 X2.X2.X1.X2.X2.X2.vout a_49002_7064# 0.263f
C9194 a_25326_26982# a_25326_25076# 0.00198f
C9195 a_2582_25164# d1 3.95e-19
C9196 a_54992_11734# a_54992_9828# 0.00396f
C9197 a_17222_9916# a_19422_9010# 4.2e-20
C9198 X2.X1.X2.X1.X1.X1.X3.vin2 X2.X1.X2.X1.X1.X1.X1.vin1 2.23e-19
C9199 X1.X2.X1.X2.X2.X1.X3.vin1 X1.X2.X1.X2.X2.X1.X2.vin1 0.00117f
C9200 d2 X1.X2.X1.X2.X2.X2.X1.vin2 7.2e-20
C9201 X2.X1.X2.X1.X1.X1.X2.vin1 a_40352_4110# 1.78e-19
C9202 X2.X1.X2.X2.X2.X2.X1.vin1 d1 0.0118f
C9203 a_11072_7922# X1.X1.X2.X1.X1.X2.vrefh 1.64e-19
C9204 X2.X1.X1.X3.vin2 a_34062_12822# 6.03e-19
C9205 a_16836_25164# d2 0.00272f
C9206 X1.X1.X1.X2.X1.X2.vrefh a_2582_13728# 8.22e-20
C9207 a_4696_18540# X1.X1.X1.X2.X1.X1.X3.vin1 0.00232f
C9208 X2.X2.X1.X1.X1.X1.X3.vin2 X2.X2.X1.X1.X1.X1.X1.vin2 8.93e-19
C9209 a_34362_18540# X2.X1.X3.vin1 0.47f
C9210 X2.X2.X2.X2.X2.X1.X3.vin1 d2 0.104f
C9211 d2 a_4396_28070# 0.00393f
C9212 X1.X1.X2.X1.X2.X1.X2.vin1 a_11072_13640# 0.197f
C9213 X1.X1.X1.X3.vin1 a_4782_28070# 1.64e-19
C9214 X2.X1.X1.X1.X2.X1.vout vdd 0.805f
C9215 a_5082_26164# X1.X1.X1.X1.X1.X2.X3.vin2 0.00846f
C9216 a_19422_9010# d1 0.0749f
C9217 X2.X1.X2.X2.X2.X1.X3.vin1 X2.X1.X2.X2.X2.X1.X2.vin1 0.00117f
C9218 a_37766_27888# X2.X1.X2.X2.X2.X1.X3.vin2 0.267f
C9219 X2.X2.X2.X1.X2.X2.X3.vin2 d1 0.151f
C9220 X1.X2.X2.X2.X2.X2.X1.vin2 X1.X2.X2.X2.X2.X2.vrefh 0.1f
C9221 X1.X1.X1.X2.X2.X1.vout vdd 0.775f
C9222 X2.X2.X2.X1.X1.X1.X2.vin1 vdd 0.578f
C9223 a_2582_13728# X1.X1.X1.X2.X1.X2.X3.vin1 0.52f
C9224 X2.X2.X1.X1.X2.X1.X1.vin1 vdd 0.592f
C9225 X2.X2.X2.X1.X2.X1.vout d1 0.0238f
C9226 X1.X2.X2.X2.X2.X1.X1.vin1 X1.X2.X2.X2.X2.vrefh 0.267f
C9227 d2 a_38152_31700# 0.00293f
C9228 a_33676_31882# X2.X1.X1.X1.X1.X1.vout 0.359f
C9229 X2.X2.X1.X1.X3.vin2 d4 0.00419f
C9230 X1.X2.X2.X2.X1.X2.X3.vin1 a_25326_23170# 0.52f
C9231 X2.X1.X2.vrefh a_35312_892# 7.3e-19
C9232 X1.X2.X1.X1.X1.X2.X1.vin1 X1.X2.X1.X1.X1.X2.X1.vin2 0.668f
C9233 a_16836_27070# d1 2.92e-22
C9234 a_54606_7922# X2.X2.X2.X1.X1.X1.X3.vin2 8.07e-19
C9235 X1.X2.X1.X1.X2.X1.X2.vin1 a_16836_23258# 0.197f
C9236 X2.X2.vrefh d1 7.29e-21
C9237 a_46116_13728# X2.X2.X1.X2.X1.X2.X2.vin1 1.78e-19
C9238 a_46116_25164# X2.X2.X1.X1.X2.X1.X2.vin1 1.78e-19
C9239 a_54992_26982# vdd 1.05f
C9240 a_19722_10916# X1.X2.X1.X2.X3.vin2 0.263f
C9241 a_2196_21352# a_2582_21352# 0.419f
C9242 d0 X2.X2.X1.X2.X1.X2.X1.vin2 0.276f
C9243 a_37852_29834# a_38152_31700# 6.71e-19
C9244 X2.X1.X2.X1.X1.X2.vrefh X2.X2.X1.X2.X2.X2.X1.vin1 0.00437f
C9245 X1.X2.X2.X2.X2.X1.X1.vin2 a_25326_26982# 0.273f
C9246 a_19422_31882# d1 0.0394f
C9247 a_8186_29834# a_8486_27888# 4.19e-20
C9248 a_54606_19358# X2.X2.X2.X1.X2.X2.X3.vin2 8.07e-19
C9249 a_37466_14586# X2.X1.X2.X1.X3.vin2 0.423f
C9250 X2.X2.X1.X1.X1.X1.vout vdd 0.781f
C9251 X1.X2.X1.X2.X2.X1.X1.vin1 vdd 0.592f
C9252 a_39966_32700# X2.X1.X2.X2.X2.X2.X2.vin1 0.402f
C9253 d0 X2.X1.X1.X2.X1.X2.X3.vin1 4.36e-19
C9254 d2 X2.X1.X2.X2.X2.X2.X3.vin2 0.00427f
C9255 X2.X1.X2.X1.X1.X1.X1.vin1 X2.X2.X2.vrefh 0.00437f
C9256 a_8572_22210# X1.X1.X2.X2.X1.X1.X3.vin2 0.00546f
C9257 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X2.vrefh 0.00118f
C9258 d2 X2.X1.X2.X1.X2.vrefh 0.158f
C9259 d3 a_52406_8828# 7.51e-19
C9260 d1 a_49002_7064# 0.0422f
C9261 X1.X1.X1.X2.X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X2.vin1 0.00117f
C9262 X2.X1.X3.vin1 X2.X3.vin1 0.273f
C9263 a_2582_17540# a_4782_16634# 4.2e-20
C9264 a_37466_22210# d4 1.54e-19
C9265 a_19336_22312# d2 0.526f
C9266 d3 a_19036_12822# 0.00108f
C9267 a_11072_28888# a_11072_30794# 0.00396f
C9268 a_11072_26982# X1.X1.X2.X2.X2.X1.X2.vin1 1.78e-19
C9269 X1.X1.X2.X2.X2.X1.X1.vin1 X1.X1.X2.X2.X2.X1.X3.vin2 2.23e-19
C9270 X1.X2.X2.X2.X1.X1.X2.vin1 vdd 0.576f
C9271 a_23512_24076# d1 0.521f
C9272 X1.X1.X2.X1.X2.X1.X3.vin1 a_11072_11734# 0.354f
C9273 d1 a_28482_892# 2.34e-19
C9274 X2.X2.X3.vin2 X2.X2.X2.X1.X2.X2.X3.vin2 0.0011f
C9275 a_25712_13640# X1.X2.X2.X1.X2.X1.X1.vin2 1.78e-19
C9276 X2.X2.X2.X1.X1.X2.X3.vin2 a_54992_9828# 0.354f
C9277 X2.X2.X2.X3.vin1 X2.X2.X2.X1.X3.vin2 0.418f
C9278 X2.X2.X3.vin2 X2.X2.X2.X1.X2.X1.vout 3.2e-19
C9279 d0 a_46502_17540# 0.0675f
C9280 a_25326_32700# X1.X2.X2.X2.X2.X2.X3.vin2 0.567f
C9281 X2.X2.X2.X1.X2.X1.X3.vin1 a_54992_11734# 0.354f
C9282 d2 a_31862_11822# 0.00792f
C9283 X2.X1.X1.X2.X1.X2.X3.vin2 d1 0.171f
C9284 a_52492_18358# d2 0.0113f
C9285 a_46116_19446# a_46502_19446# 0.419f
C9286 d2 X1.X1.X2.X2.X3.vin2 0.0685f
C9287 X2.X1.X1.X3.vin1 a_33976_18540# 0.17f
C9288 d1 a_54992_7922# 2.25e-20
C9289 d3 a_4782_12822# 0.00122f
C9290 a_23512_27888# a_22826_29834# 2.86e-19
C9291 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X3.vin1 0.206f
C9292 X2.X1.X1.X3.vin2 a_33976_10916# 0.355f
C9293 X2.X2.X1.X1.X2.X2.X2.vin1 d4 8.68e-20
C9294 X2.X1.X1.X3.vin1 a_34062_20446# 5.31e-19
C9295 d3 X1.X2.X2.X2.X1.X2.X2.vin1 8.68e-20
C9296 a_10686_26982# a_11072_26982# 0.419f
C9297 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X2.vrefh 0.00118f
C9298 a_23126_16452# a_23512_16452# 0.419f
C9299 X1.X1.X3.vin1 X1.X1.X1.X2.X1.X1.X3.vin2 8.36e-19
C9300 X1.X2.X2.X1.X3.vin2 vdd 1.32f
C9301 X1.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X1.vout 0.0524f
C9302 X1.X2.X2.X2.X3.vin2 a_23212_29834# 0.363f
C9303 X2.X1.X1.X2.X2.X1.X1.vin2 X2.X1.X1.X2.X2.X1.X2.vin1 0.242f
C9304 a_25712_15546# a_25712_13640# 0.00396f
C9305 X2.X2.X2.X2.X1.X1.X1.vin1 vdd 0.592f
C9306 X1.X2.X2.X1.X1.X1.X1.vin1 X2.X1.X2.vrefh 0.00437f
C9307 a_2582_23258# a_2582_21352# 0.00198f
C9308 a_2196_23258# X1.X1.X1.X1.X2.X2.X1.vin1 1.64e-19
C9309 X2.X1.X2.X2.X1.X1.vout X2.X1.X2.X2.X1.X1.X3.vin1 0.118f
C9310 d2 a_52792_8828# 0.00287f
C9311 X2.X2.X3.vin2 a_49002_7064# 5.84e-19
C9312 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X2.X3.vin2 0.102f
C9313 a_52492_6962# a_52406_5016# 3.14e-19
C9314 X2.X1.X1.X1.X2.X2.X2.vin1 d4 8.68e-20
C9315 X2.X2.X1.X1.X1.X2.X2.vin1 a_46502_27070# 0.402f
C9316 a_2582_25164# X1.X1.X1.X1.X2.vrefh 8.22e-20
C9317 a_54606_26982# a_54606_28888# 0.00198f
C9318 a_31862_32788# a_33676_31882# 1.06e-19
C9319 X2.X2.X2.X2.X2.X1.X1.vin2 X2.X2.X2.X2.X2.X1.X2.vin1 0.242f
C9320 X2.X1.X1.X1.X1.X1.X1.vin1 X2.X1.X1.X1.X1.X1.X2.vin1 0.0689f
C9321 X1.X1.X1.X3.vin1 X1.X1.X1.X3.vin2 0.552f
C9322 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X3.vin2 0.234f
C9323 a_39966_19358# vdd 0.553f
C9324 d2 a_10686_11734# 0.00328f
C9325 d3 X1.X2.X1.X1.X3.vin2 0.433f
C9326 X1.X2.X2.X2.X1.X2.X3.vin1 vdd 0.96f
C9327 d3 X1.X2.X1.X2.X3.vin2 0.156f
C9328 a_23126_24076# a_23512_24076# 0.419f
C9329 d1 a_34062_9010# 0.0749f
C9330 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X1.vin1 0.0689f
C9331 a_25326_26982# d3 0.00112f
C9332 X1.X2.X2.X1.X1.X2.X2.vin1 X1.X2.X2.X1.X1.X2.X3.vin1 0.00117f
C9333 X1.X2.X2.X1.X2.X2.X3.vin2 a_25326_15546# 7.84e-19
C9334 X1.X2.X2.X1.X1.X2.X3.vin2 a_23126_8828# 0.277f
C9335 X1.X2.X1.X2.X2.X1.X3.vin2 a_16836_8010# 0.354f
C9336 a_2196_21352# a_2196_19446# 0.00396f
C9337 X1.X2.X1.X1.X2.X2.X2.vin1 d4 8.68e-20
C9338 X2.X1.X2.X2.X1.X2.X1.vin1 X2.X1.X2.X2.X1.X2.vrefh 0.267f
C9339 X1.X2.X1.X1.X1.X1.X1.vin2 a_16836_30882# 1.78e-19
C9340 d5 a_34926_892# 0.508f
C9341 d3 a_46116_32788# 2.56e-19
C9342 a_40352_13640# d1 2.92e-22
C9343 a_11072_23170# vdd 1.05f
C9344 X1.X2.X3.vin2 a_22826_6962# 0.00111f
C9345 a_48702_24258# X2.X2.X1.X1.X2.X1.vout 0.422f
C9346 d0 X1.X1.X2.X1.X1.X1.X1.vin2 0.276f
C9347 a_40352_6016# X2.X1.X2.X1.X1.X1.X1.vin2 1.78e-19
C9348 X1.X2.X2.X1.X2.X1.X3.vin2 d1 0.15f
C9349 a_40352_26982# d1 2.25e-20
C9350 a_17222_15634# a_19336_14688# 2.95e-20
C9351 d4 a_23512_16452# 0.00119f
C9352 a_4782_16634# X1.X1.X1.X2.X1.X1.X3.vin2 0.267f
C9353 a_25326_19358# vdd 0.553f
C9354 a_46502_11822# X2.X2.X1.X2.X2.X1.X1.vin1 8.22e-20
C9355 X2.X2.X1.X1.X1.X2.X1.vin2 d1 0.00406f
C9356 X1.X2.X1.X1.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X1.vout 0.118f
C9357 d2 X2.X1.X2.X1.X2.X1.X2.vin1 0.0318f
C9358 X1.X2.X2.X2.X1.X2.X3.vin2 a_22826_22210# 3.85e-19
C9359 X1.X1.X3.vin1 vdd 0.855f
C9360 a_23126_12640# vdd 0.561f
C9361 X2.X2.X2.X1.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.X3.vin2 1.22e-19
C9362 X2.X1.X1.X1.X1.X2.X3.vin2 a_31476_27070# 0.354f
C9363 a_10686_6016# a_11072_6016# 0.419f
C9364 a_34062_28070# a_31862_27070# 4.77e-21
C9365 a_4696_26164# a_2582_25164# 5.36e-21
C9366 a_33976_26164# a_34362_26164# 0.414f
C9367 X2.X1.X1.X1.X1.X2.X3.vin1 d1 0.146f
C9368 X2.X2.X2.X1.X3.vin2 X2.X2.X2.X1.X3.vin1 0.546f
C9369 X2.X2.X2.X1.X2.X1.vout a_52492_10734# 1.64e-19
C9370 X1.X2.X2.X3.vin2 X1.X2.X2.X2.X1.X1.X3.vin2 0.0943f
C9371 X2.X1.X1.X2.X3.vin1 X2.X1.X1.X2.X1.X2.X3.vin1 0.0174f
C9372 a_37852_6962# a_39966_6016# 2.95e-20
C9373 a_34362_10916# d1 0.0316f
C9374 d0 a_2196_11822# 0.515f
C9375 X2.X2.X1.X1.X3.vin2 X2.X2.X1.X1.X2.X2.vout 0.0866f
C9376 d2 X2.X2.X1.X1.X1.X2.X1.vin1 0.0114f
C9377 a_2582_6104# X1.X1.X1.X2.X2.X2.X1.vin1 0.417f
C9378 a_2196_6104# X1.X1.X1.X2.X2.X2.X3.vin1 0.354f
C9379 X2.X1.X2.X2.X1.X1.vout X2.X1.X2.X2.X1.X1.X3.vin2 0.342f
C9380 X2.X1.X3.vin1 a_37766_16452# 8.66e-20
C9381 a_2582_27070# a_2196_27070# 0.419f
C9382 X2.X1.X1.X1.X1.X2.X2.vin1 a_31476_28976# 1.78e-19
C9383 d1 a_8872_5016# 0.522f
C9384 a_39966_17452# d1 0.00148f
C9385 a_10686_19358# vdd 0.553f
C9386 X1.X1.X2.X1.X2.X1.X3.vin1 vdd 0.997f
C9387 a_52106_6962# a_52792_8828# 3.31e-19
C9388 a_16836_17540# X1.X2.X1.X2.X1.X1.X2.vin1 1.78e-19
C9389 X2.X1.X1.X2.X2.X2.X1.vin2 vdd 0.387f
C9390 X1.X2.X2.X2.X1.X1.X3.vin1 a_23212_18358# 0.00255f
C9391 a_31476_25164# vdd 1.05f
C9392 a_48616_26164# X2.X2.X1.X1.X3.vin1 0.169f
C9393 d2 X2.X2.X1.X2.X1.X1.X1.vin2 0.231f
C9394 X2.X1.X1.X1.X2.X1.X3.vin2 X2.X1.X1.X1.X2.X2.vrefh 0.161f
C9395 a_38152_31700# X2.X1.X2.X2.X2.X2.X3.vin2 0.101f
C9396 a_33976_22312# a_31862_21352# 2.68e-20
C9397 d3 X2.X2.X1.X1.X2.X1.vout 0.00226f
C9398 a_48616_29936# a_46502_28976# 2.68e-20
C9399 a_39966_7922# X2.X1.X2.X1.X1.X2.vrefh 8.22e-20
C9400 a_4782_24258# X1.X1.X1.X1.X2.X1.X3.vin2 0.267f
C9401 X1.X1.X1.X1.X1.X1.X1.vin2 d0 0.201f
C9402 d2 a_8486_5016# 0.00123f
C9403 a_54606_21264# a_52406_20264# 4.77e-21
C9404 a_10686_28888# a_11072_28888# 0.419f
C9405 a_48316_9010# X2.X2.X1.X2.X2.X1.vout 0.359f
C9406 d2 X2.X1.X1.X2.X1.X1.X3.vin1 0.104f
C9407 d0 X1.X1.X2.X1.X2.X2.X1.vin1 0.267f
C9408 X1.X2.X1.X3.vin1 d4 0.509f
C9409 a_5082_26164# X1.X1.X1.X1.X3.vin2 0.241f
C9410 a_38152_27888# X2.X1.X2.X2.X2.X1.vout 0.359f
C9411 X1.X1.X2.X1.X2.X2.X3.vin2 a_8486_16452# 0.277f
C9412 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X3.vin1 0.00117f
C9413 d0 X1.X2.X1.X2.X2.X2.vrefh 0.848f
C9414 X1.X1.X1.X2.X2.X1.X3.vin2 X1.X1.X1.X2.X2.X2.vrefh 0.161f
C9415 a_2582_28976# X1.X1.X1.X1.X1.X2.X1.vin1 0.417f
C9416 a_39966_25076# a_38152_24076# 1.15e-20
C9417 a_2196_28976# X1.X1.X1.X1.X1.X2.X3.vin1 0.354f
C9418 X2.X2.X2.X3.vin2 vdd 0.716f
C9419 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X1.X3.vin2 0.0943f
C9420 X1.X2.X2.X1.X1.X2.vout X1.X2.X2.X1.X1.X1.vout 0.507f
C9421 a_2196_9916# vdd 1.05f
C9422 d0 a_17222_13728# 0.0675f
C9423 X1.X1.X1.X1.X2.X1.X1.vin2 a_2582_23258# 8.88e-20
C9424 a_4782_16634# vdd 0.561f
C9425 X1.X1.X2.X2.X2.X1.X1.vin2 a_11072_28888# 1.78e-19
C9426 a_23126_31700# a_23512_31700# 0.419f
C9427 a_8572_29834# d1 0.00613f
C9428 a_22826_14586# X1.X2.X2.X1.X2.X1.vout 0.383f
C9429 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X3.vin1 0.546f
C9430 X2.X1.X2.X1.X2.X2.vrefh d1 0.0124f
C9431 a_8872_12640# a_10686_11734# 1.06e-19
C9432 X1.X1.X1.X2.X2.vrefh a_2582_11822# 0.3f
C9433 a_46116_11822# a_46502_11822# 0.419f
C9434 d0 X1.X1.X2.X1.X1.X2.X1.vin1 0.267f
C9435 X1.X1.X1.X1.X1.X2.X1.vin1 a_2582_30882# 8.22e-20
C9436 X1.X2.X2.X2.X2.X1.X2.vin1 d0 0.262f
C9437 a_52792_12640# a_54606_11734# 1.06e-19
C9438 a_5082_22312# d4 3.79e-19
C9439 X1.X1.X1.X1.X2.X2.X1.vin2 vdd 0.36f
C9440 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X1.X3.vin2 1.22e-19
C9441 d3 a_17222_32788# 1.28e-19
C9442 a_48616_22312# a_48702_20446# 3.38e-19
C9443 a_49002_22312# a_48316_20446# 3.31e-19
C9444 a_16836_32788# a_17222_32788# 0.419f
C9445 a_17222_25164# a_17222_23258# 0.00198f
C9446 a_22826_29834# X1.X2.X2.X2.X2.X2.vout 0.263f
C9447 d0 a_25712_17452# 0.515f
C9448 a_46116_9916# X2.X2.X1.X2.X2.X1.X1.vin2 0.12f
C9449 X2.X2.X2.X2.X1.X2.X3.vin1 d2 0.155f
C9450 a_16836_13728# a_16836_11822# 0.00396f
C9451 X1.X1.X1.X1.X1.X2.vout X1.X1.X1.X1.X1.X2.X3.vin1 0.326f
C9452 a_5082_26164# vdd 0.489f
C9453 d4 d0 5.4e-19
C9454 d0 a_54606_11734# 0.0675f
C9455 a_25326_13640# X1.X2.X2.X1.X2.X1.X3.vin1 0.00207f
C9456 a_10686_9828# a_8872_8828# 1.15e-20
C9457 a_52406_24076# a_52106_22210# 5.55e-20
C9458 d2 X2.X1.X1.X2.X1.X2.X2.vin1 0.0329f
C9459 d3 X2.X2.X1.X2.X1.X2.X3.vin1 2.1e-19
C9460 d3 a_8872_27888# 0.00178f
C9461 a_39966_9828# X2.X1.X2.X1.X1.X2.X3.vin2 0.567f
C9462 d3 X1.X1.X1.X1.X2.X1.X1.vin2 3.99e-21
C9463 a_40352_23170# d2 0.00351f
C9464 X2.X1.X2.X3.vin1 X2.X1.X2.X1.X2.X1.vout 0.038f
C9465 X1.X1.X2.X1.X1.X1.X3.vin2 a_8486_5016# 0.267f
C9466 a_49002_10916# a_48316_9010# 2.97e-19
C9467 a_48616_10916# a_48702_9010# 3.21e-19
C9468 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X1.X3.vin1 0.00117f
C9469 d2 X2.X2.X2.X1.X1.X2.X1.vin2 0.226f
C9470 X1.X2.X3.vin2 d2 0.1f
C9471 X2.X2.X2.X1.X2.X1.X3.vin2 a_54992_13640# 0.354f
C9472 X1.X1.X2.X2.X2.X2.X1.vin1 d0 0.267f
C9473 X2.X2.X1.X1.X1.X2.X2.vin1 d3 8.68e-20
C9474 a_39966_32700# X2.X1.X2.X2.X2.X2.X3.vin1 0.00207f
C9475 X1.X2.X2.X1.X2.X1.X3.vin1 a_23212_10734# 0.00251f
C9476 X2.X1.X2.X2.X2.X2.X2.vin1 a_37766_31700# 0.00351f
C9477 X1.X2.X2.X1.X1.X1.X1.vin2 X2.X1.X1.X2.X2.X2.X2.vin1 0.00232f
C9478 X2.X1.X1.X1.X3.vin1 vdd 0.805f
C9479 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X3.vin1 0.206f
C9480 a_37852_25982# a_39966_25076# 4.72e-20
C9481 X1.X2.X2.X1.X1.X2.X3.vin2 X1.X2.X2.X1.X1.X2.X1.vin1 2.23e-19
C9482 X1.X2.X2.X1.X1.X2.X2.vin1 a_25712_7922# 1.78e-19
C9483 a_17222_15634# X1.X2.X1.X2.X1.X2.X1.vin1 8.22e-20
C9484 d0 X2.X1.X1.X2.X2.X2.X2.vin1 0.262f
C9485 a_11072_17452# vdd 1.05f
C9486 a_52406_20264# a_52106_18358# 5.25e-20
C9487 d0 X2.X2.X2.X1.X2.X2.X1.vin2 0.276f
C9488 X2.X1.X2.X1.X1.X1.vout vdd 0.78f
C9489 X1.X1.X2.X2.X2.X1.vout a_8572_29834# 0.169f
C9490 a_8186_29834# a_8486_31700# 5.55e-20
C9491 d2 X2.X1.X1.X2.X1.X1.vout 0.00169f
C9492 X1.X2.X2.X1.X1.X2.X3.vin1 X1.X2.X2.X1.X1.X1.X3.vin2 1.22e-19
C9493 a_52406_27888# a_52492_25982# 3.21e-19
C9494 a_4782_31882# X1.X1.X1.X1.X1.X1.X3.vin2 0.267f
C9495 a_4782_31882# vdd 0.565f
C9496 X2.X1.X2.X2.X2.X2.vrefh d1 0.0124f
C9497 a_37852_10734# X2.X1.X2.X1.X1.X2.X3.vin2 0.00535f
C9498 a_46502_28976# X2.X2.X1.X1.X1.X1.X3.vin2 8.07e-19
C9499 X2.X2.X2.X2.X2.X2.X1.vin1 X2.X2.X2.X2.X2.X2.X3.vin2 2.23e-19
C9500 a_23512_5016# vdd 1.05f
C9501 a_2196_27070# d1 2.92e-22
C9502 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.vout 0.0857f
C9503 a_54992_30794# X2.X2.X2.X2.X2.X2.X2.vin1 1.78e-19
C9504 X2.X2.X1.X1.X1.X2.X3.vin2 X2.X2.X1.X1.X1.X2.X1.vin2 8.93e-19
C9505 a_46116_21352# X2.X2.X1.X1.X2.X2.X1.vin1 0.195f
C9506 X2.X2.X2.X1.X2.X2.X3.vin1 a_52792_16452# 0.199f
C9507 d0 a_25712_11734# 0.518f
C9508 a_2196_32788# X1.X1.X1.X1.X1.X1.X2.vin1 1.78e-19
C9509 a_14082_892# X3.vin1 0.472f
C9510 d6 a_20286_892# 0.00105f
C9511 d3 X2.X1.X1.X2.X1.X2.vout 0.0232f
C9512 X1.X1.X1.X1.X2.X2.X1.vin2 X1.X1.X1.X1.X2.X2.X3.vin2 8.93e-19
C9513 a_8186_18358# X1.X1.X2.X1.X2.X2.X3.vin2 0.00846f
C9514 a_4396_24258# a_5082_22312# 2.86e-19
C9515 X1.X2.X2.X1.X2.X1.X1.vin2 X1.X2.X2.X1.X2.vrefh 0.1f
C9516 a_4782_24258# a_4696_22312# 3.14e-19
C9517 a_10686_6016# vdd 0.541f
C9518 a_4396_20446# d2 6.04e-19
C9519 X1.X2.X1.X1.X1.X2.X3.vin2 d3 0.103f
C9520 X1.X2.X1.X1.X1.X1.X1.vin2 a_19036_31882# 0.00113f
C9521 a_8872_24076# vdd 1.05f
C9522 X1.X1.X1.X3.vin1 a_4782_20446# 5.31e-19
C9523 a_31476_6104# a_31476_4198# 0.00396f
C9524 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.X1.vin2 8.93e-19
C9525 X1.X1.X2.X1.X1.X2.X2.vin1 a_10686_7922# 8.88e-20
C9526 a_52106_29834# X2.X2.X2.X2.X2.X2.X3.vin1 0.00874f
C9527 a_39966_6016# a_37766_5016# 4.77e-21
C9528 a_10686_13640# d1 0.00148f
C9529 d2 X1.X1.X1.X2.X1.X2.vrefh 0.177f
C9530 X1.X1.X3.vin1 X1.X1.X2.X1.X1.X1.vout 5.53e-20
C9531 d2 X1.X2.X1.X2.X1.X2.X1.vin2 0.226f
C9532 a_19036_16634# a_19722_14688# 2.86e-19
C9533 a_19422_16634# a_19336_14688# 3.14e-19
C9534 X2.X1.X2.X2.X2.X1.X1.vin2 d2 0.231f
C9535 a_5082_14688# a_4782_12822# 5.55e-20
C9536 X1.X1.X2.X2.X1.X1.vout a_8486_20264# 0.422f
C9537 a_19722_10916# X1.X2.X1.X2.X2.X1.X3.vin2 3.49e-19
C9538 a_17222_28976# d1 3.41e-19
C9539 d0 a_54606_9828# 0.0489f
C9540 X2.X1.X1.X2.X2.X1.X3.vin2 a_34362_7064# 0.00815f
C9541 X2.X2.X2.X1.X2.X2.vrefh X2.X2.X2.X1.X2.X1.X2.vin1 0.564f
C9542 X2.X2.X2.X2.X2.X2.X1.vin2 d0 0.253f
C9543 X1.X1.X1.X2.vrefh X1.X1.X1.X2.X1.X1.X1.vin1 0.267f
C9544 X1.X2.X1.X1.X1.X1.X1.vin2 vdd 0.399f
C9545 d2 X1.X1.X1.X2.X1.X2.X3.vin1 0.155f
C9546 d2 X2.X1.X1.X1.X1.X1.vout 0.0903f
C9547 d2 a_31476_28976# 0.00351f
C9548 X2.X1.X2.X2.X1.X1.vout d1 0.0238f
C9549 X2.X1.X2.X2.X1.X2.X3.vin1 a_38152_24076# 0.199f
C9550 X1.X1.X2.X1.X2.X2.vout X1.X1.X2.X1.X3.vin2 0.0866f
C9551 d0 X1.X2.X2.X1.X1.X2.X1.vin1 0.267f
C9552 a_11072_11734# X1.X1.X2.X1.X2.vrefh 1.64e-19
C9553 X2.X2.X2.X2.X1.X2.X1.vin2 X2.X2.X2.X2.X1.X1.X3.vin2 3.94e-19
C9554 X2.X2.X2.X2.X1.X2.X1.vin1 a_54606_21264# 8.22e-20
C9555 X2.X2.X2.X1.X2.X1.X2.vin1 vdd 0.576f
C9556 a_37766_16452# X2.X1.X2.X1.X2.X2.X3.vin1 0.42f
C9557 X2.X1.X1.X2.X1.X1.X2.vin1 X2.X1.X1.X2.X1.X2.vrefh 0.564f
C9558 a_11072_28888# X1.X1.X2.X2.X2.X2.vrefh 0.118f
C9559 X3.vin2 a_34926_892# 4.87e-19
C9560 X1.X2.X2.X2.X1.X2.X1.vin2 X2.X1.X1.X1.X2.X2.vrefh 0.0128f
C9561 a_17222_8010# a_19336_7064# 2.95e-20
C9562 X1.X1.X2.X1.X1.X2.X3.vin1 a_8872_8828# 0.199f
C9563 a_37766_27888# X2.X1.X2.X2.X3.vin2 0.00101f
C9564 d2 X2.X2.X2.X2.X3.vin2 0.0685f
C9565 a_34362_29936# X2.X1.X1.X1.X1.X2.X3.vin1 0.00874f
C9566 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X2.vout 0.197f
C9567 a_52492_14586# a_52792_12640# 6.1e-19
C9568 X2.X2.X1.X2.X2.X1.X1.vin2 X2.X2.X1.X2.X2.X1.X3.vin2 8.93e-19
C9569 X1.X1.X2.X1.X2.X1.X1.vin2 X1.X1.X2.X1.X2.X1.X1.vin1 0.668f
C9570 a_48316_20446# d1 0.521f
C9571 a_23126_8828# a_23212_6962# 3.38e-19
C9572 a_11072_26982# d2 0.00272f
C9573 X1.X2.X2.X1.X2.X2.X1.vin1 a_25712_15546# 0.195f
C9574 a_17222_6104# X1.X2.X1.X2.X2.X2.vrefh 8.22e-20
C9575 X2.X1.X1.X1.X2.vrefh d0 0.848f
C9576 X1.X2.X3.vin1 X1.X2.X1.X2.X2.X1.X3.vin1 0.00789f
C9577 d2 X1.X1.X1.X1.X1.X2.vrefh 6.65e-20
C9578 a_22826_25982# a_23512_24076# 3.08e-19
C9579 a_19422_28070# X1.X2.X1.X1.X1.X2.X3.vin2 0.277f
C9580 X1.X2.X2.X2.X3.vin1 vdd 0.804f
C9581 X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 0.0903f
C9582 X1.X2.X2.X1.X3.vin1 vdd 0.805f
C9583 X2.X2.X1.X2.X1.X1.X3.vin1 vdd 0.997f
C9584 X1.X2.X1.X1.X2.X1.vout d1 0.0238f
C9585 X1.X2.X2.X1.X2.X2.vrefh a_25712_13640# 0.118f
C9586 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X2.vout 0.197f
C9587 X2.X2.X3.vin1 a_52106_14586# 2.24e-19
C9588 a_16836_17540# X1.X2.X1.X2.X1.X1.X1.vin1 0.195f
C9589 X1.X1.X1.X2.X2.X2.X3.vin2 vdd 0.725f
C9590 d4 X1.X1.X1.X2.X1.X1.X3.vin1 0.0205f
C9591 a_23212_18358# d1 0.00638f
C9592 X1.X2.vrefh X1.X2.X1.X1.X1.X1.X1.vin2 0.109f
C9593 X1.X1.X1.X1.X1.X2.X1.vin2 d0 0.276f
C9594 a_37766_8828# a_38152_8828# 0.419f
C9595 d2 a_5082_29936# 0.254f
C9596 X1.X1.X2.X2.X2.vrefh d0 0.848f
C9597 a_33676_20446# d1 0.521f
C9598 X1.X1.X2.X2.X1.X2.vrefh X1.X1.X2.X2.X1.X1.X3.vin1 0.00118f
C9599 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X3.vin1 0.199f
C9600 X1.X2.X1.X1.X1.X2.X3.vin2 X1.X2.X1.X1.X3.vin1 0.0565f
C9601 X2.X2.X1.X2.X1.X2.X2.vin1 X2.X2.X1.X2.X2.vrefh 0.564f
C9602 X2.X1.X1.X2.vrefh d2 0.173f
C9603 a_39966_4110# vdd 0.553f
C9604 X1.X1.X2.X1.X1.X1.X3.vin1 a_11072_4110# 0.354f
C9605 d4 X2.X2.X2.X1.X2.X2.X3.vin1 2.52e-19
C9606 X2.X1.X2.X1.X1.X1.vout X2.X1.X2.X1.X1.X1.X3.vin1 0.118f
C9607 a_19722_14688# vdd 0.477f
C9608 X2.X1.X1.X2.X1.X1.X3.vin2 d1 0.15f
C9609 X1.X1.X1.X1.X2.vrefh a_2196_27070# 0.118f
C9610 a_31476_9916# a_31862_9916# 0.419f
C9611 X1.X2.X2.X1.X1.X2.X2.vin1 X2.X1.X1.X2.X2.X1.X1.vin2 0.00232f
C9612 X2.X2.X2.X2.X2.X2.X3.vin1 a_52792_31700# 0.199f
C9613 d3 X1.X1.X2.X1.X2.X2.vout 8.47e-19
C9614 a_42976_892# X2.X3.vin2 0.0927f
C9615 a_2196_6104# X1.X1.X1.X2.X2.X2.X2.vin1 1.78e-19
C9616 a_25712_9828# X1.X2.X2.X1.X1.X2.X1.vin2 1.78e-19
C9617 a_46116_13728# X2.X2.X1.X2.X1.X2.X1.vin2 0.12f
C9618 a_19036_20446# d1 0.521f
C9619 d2 X2.X2.X1.X2.X2.X1.vout 0.0909f
C9620 X1.X1.X2.X1.X1.X2.X3.vin1 X1.X1.X2.X1.X1.X2.X1.vin1 0.206f
C9621 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X1.vin2 0.242f
C9622 a_54606_6016# a_54606_4110# 0.00198f
C9623 X1.X2.X1.X2.vrefh d2 0.173f
C9624 a_52792_24076# a_54606_23170# 1.06e-19
C9625 d3 X1.X2.X1.X2.X2.X1.X3.vin2 7.71e-19
C9626 a_8572_10734# a_8872_8828# 6.48e-19
C9627 a_39966_13640# X2.X1.X2.X1.X2.X1.X3.vin2 0.567f
C9628 a_10686_13640# a_8486_12640# 4.77e-21
C9629 a_31862_32788# d2 1.95e-19
C9630 X1.X1.X1.X2.X2.X1.X2.vin1 a_2582_8010# 0.402f
C9631 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X1.vin2 0.216f
C9632 a_46116_9916# d1 2.25e-20
C9633 a_52406_16452# a_54606_15546# 4.2e-20
C9634 d0 d7 1.37e-19
C9635 X1.X1.X1.X1.X3.vin1 X1.X1.X1.X1.X1.X1.vout 0.13f
C9636 X2.X2.X3.vin1 vdd 0.852f
C9637 X2.X1.X1.X2.X2.vrefh vdd 0.426f
C9638 X2.X1.X1.X1.X1.X2.X3.vin2 a_31862_25164# 8.07e-19
C9639 X2.X2.X1.X2.X1.X2.vrefh vdd 0.414f
C9640 d2 a_54992_9828# 0.00533f
C9641 X2.X2.X1.X1.X3.vin2 X2.X2.X2.X3.vin2 7.46e-20
C9642 a_33676_16634# a_33976_14688# 6.1e-19
C9643 a_52106_25982# X2.X2.X2.X2.X3.vin1 0.372f
C9644 X1.X2.X2.X2.vrefh vdd 0.414f
C9645 X2.X1.X1.X2.X1.X2.X2.vin1 a_31862_11822# 0.402f
C9646 X2.X2.X2.X2.X2.X2.X1.vin2 a_54992_32700# 1.78e-19
C9647 X1.X1.X1.X2.X2.X2.vout vdd 0.698f
C9648 a_19722_7064# X1.X2.X1.X2.X2.X2.X3.vin2 3.85e-19
C9649 X1.X2.X1.X2.X2.X2.vout a_19422_5198# 0.418f
C9650 X2.X2.X2.X2.X2.X1.X2.vin1 a_54992_28888# 0.197f
C9651 X2.vrefh d4 0.00449f
C9652 X2.X1.X3.vin2 a_37852_18358# 0.355f
C9653 X1.X2.X1.X2.X2.X2.X3.vin1 a_19722_7064# 0.00874f
C9654 d2 X2.X1.X2.X1.X1.X2.X3.vin2 0.121f
C9655 a_40352_28888# X2.X1.X2.X2.X2.X2.X1.vin1 1.64e-19
C9656 X1.X2.X2.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X2.vout 0.08f
C9657 d1 a_34926_892# 4.67e-19
C9658 X2.X1.X1.X1.X2.X2.X3.vin2 a_31862_19446# 0.567f
C9659 X2.X2.X1.X1.X2.X2.X1.vin2 d1 2.18e-19
C9660 X1.X1.X2.X1.X1.X1.X1.vin1 vdd 0.592f
C9661 X1.X2.X1.X2.vrefh a_17222_17540# 8.22e-20
C9662 a_46502_28976# X2.X2.X1.X1.X1.X2.X3.vin1 0.52f
C9663 X1.X1.X2.X1.X2.vrefh vdd 0.426f
C9664 a_31476_15634# vdd 1.05f
C9665 d3 X1.X2.X1.X1.X1.X1.X3.vin2 0.0678f
C9666 X2.X1.X1.X1.X1.X2.X1.vin2 X1.X2.X2.X2.X2.X2.vrefh 0.0128f
C9667 X1.X2.X2.X1.X2.X2.vout a_23212_14586# 0.0929f
C9668 X2.X1.X1.X1.X2.X2.X3.vin1 d1 0.146f
C9669 X1.X1.X2.X2.vrefh vdd 0.414f
C9670 d4 X1.X2.X1.X2.X1.X1.vout 0.00145f
C9671 X1.X2.X2.X1.X2.X1.X3.vin2 a_22826_10734# 3.49e-19
C9672 d4 X2.X2.X2.X2.X2.X2.X3.vin1 0.00851f
C9673 X2.X2.X1.X1.X2.X2.X1.vin1 d2 0.0106f
C9674 d3 X1.X1.X1.X2.X3.vin1 0.375f
C9675 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X3.vin2 0.0321f
C9676 X2.X1.X1.X1.X1.X1.X3.vin2 d1 0.152f
C9677 a_37766_31700# X2.X1.X2.X2.X2.X2.X3.vin1 0.42f
C9678 X2.X1.X1.X1.X1.X1.X2.vin1 X2.X1.X1.X1.X1.X2.vrefh 0.564f
C9679 d0 X2.X2.X2.X1.X1.X1.X2.vin1 0.262f
C9680 d1 a_54606_4110# 0.00106f
C9681 X2.X2.X1.X1.X2.X1.X1.vin1 d0 0.267f
C9682 X2.X2.X1.X2.X2.X2.vrefh a_46502_8010# 0.3f
C9683 a_37766_27888# d1 0.0749f
C9684 a_2582_6104# a_2582_4198# 0.00198f
C9685 d3 X1.X1.X2.X2.X2.X2.vout 0.222f
C9686 a_16836_23258# vdd 1.05f
C9687 d2 a_49002_10916# 7.13e-19
C9688 a_54606_21264# X2.X2.X2.X2.X1.X1.X1.vin2 8.88e-20
C9689 X1.X2.X1.X2.X1.X2.X3.vin2 a_17222_11822# 0.567f
C9690 a_54992_15546# a_54992_13640# 0.00396f
C9691 a_54992_26982# d0 0.518f
C9692 a_34062_28070# d2 0.00202f
C9693 X2.X2.X2.X1.X1.X1.X3.vin1 a_54606_4110# 0.52f
C9694 X1.X2.X2.X2.X2.X2.X1.vin1 a_25712_30794# 0.195f
C9695 a_52492_29834# d1 0.00613f
C9696 a_48616_14688# a_49002_14688# 0.419f
C9697 X1.X1.X2.X2.X2.X2.X2.vin1 vdd 0.578f
C9698 X2.X2.X1.X1.X1.X2.vrefh vdd 0.43f
C9699 a_8486_16452# a_8572_14586# 3.38e-19
C9700 d0 X1.X2.X1.X2.X2.X1.X1.vin1 0.267f
C9701 X1.X2.X1.X1.X2.X2.X3.vin2 a_17222_19446# 0.567f
C9702 X2.X1.X1.X2.X1.X2.X1.vin2 vdd 0.361f
C9703 X2.X2.X2.X2.vrefh d2 0.173f
C9704 X1.X1.X1.X1.X2.X2.vout d1 0.033f
C9705 a_4696_29936# a_4782_28070# 3.38e-19
C9706 a_5082_29936# a_4396_28070# 3.31e-19
C9707 a_52492_25982# a_52406_24076# 3.3e-19
C9708 a_2196_30882# X1.X1.X1.X1.X1.X1.X2.vin1 0.197f
C9709 a_31476_30882# vdd 1.05f
C9710 a_49002_26164# vdd 0.489f
C9711 X1.X2.X1.X2.X1.X2.X3.vin1 vdd 0.96f
C9712 X2.X2.X2.X1.X2.X2.X2.vin1 X2.X2.X2.X1.X2.X2.X1.vin1 0.0689f
C9713 X2.X2.X1.X2.X2.X2.X1.vin1 X2.X2.X1.X2.X2.X2.X1.vin2 0.668f
C9714 X2.X1.X2.X2.vrefh a_39966_17452# 0.3f
C9715 d1 a_25326_4110# 0.00107f
C9716 d2 X2.X2.X2.X1.X2.X1.X3.vin1 0.104f
C9717 X1.X2.X2.X2.X1.X1.X2.vin1 d0 0.262f
C9718 a_46116_28976# vdd 1.05f
C9719 X2.X2.X2.X1.X2.X2.X3.vin2 a_54606_15546# 7.84e-19
C9720 X1.X1.X2.X1.X1.X1.X2.vin1 X1.X1.X2.X1.X1.X2.vrefh 0.564f
C9721 d4 X1.X2.X1.X1.X1.X1.vout 4.78e-20
C9722 d2 X1.X2.X2.X2.X2.X1.vout 0.115f
C9723 a_19722_14688# X1.X2.X1.X2.X1.X2.vout 0.254f
C9724 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X3.vin1 1.22e-19
C9725 X2.X1.X3.vin2 X2.X1.X2.X1.X3.vin1 0.0361f
C9726 X2.X1.X2.X3.vin1 a_37852_10734# 0.356f
C9727 X2.X1.X3.vin2 d5 0.0353f
C9728 X1.X2.X1.X2.X2.vrefh X1.X2.X1.X2.X2.X1.X1.vin1 0.267f
C9729 X2.X2.X2.X1.X2.X2.X3.vin1 a_52492_14586# 0.00329f
C9730 X2.X1.X1.X2.X2.X2.vrefh X2.X1.X1.X2.X2.X2.X1.vin1 0.267f
C9731 X1.X2.X1.X2.X3.vin2 a_19336_7064# 0.363f
C9732 X2.X1.X2.X1.X1.X1.X3.vin1 a_39966_4110# 0.52f
C9733 a_2582_25164# a_4782_24258# 4.2e-20
C9734 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X2.vin1 0.00117f
C9735 d3 X2.X1.X1.X2.X2.X1.X3.vin2 7.71e-19
C9736 a_37852_18358# X2.X1.X2.X1.X2.X2.X3.vin2 0.00517f
C9737 X2.X1.X2.X1.X2.X1.vout vdd 0.805f
C9738 a_31862_17540# vdd 0.553f
C9739 X1.X2.X1.X1.X1.X2.vout X1.X2.X1.X1.X1.X1.vout 0.507f
C9740 X2.X2.X2.X3.vin2 X2.X2.X2.X2.X1.X2.X3.vin2 0.102f
C9741 X1.X2.X2.X2.vrefh X2.X1.X1.X2.X1.X1.X1.vin2 0.0128f
C9742 X2.X2.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.X3.vin1 0.0174f
C9743 a_16836_11822# d1 2.92e-22
C9744 X1.X2.X1.X1.X2.X1.X2.vin1 d2 0.0318f
C9745 a_54992_11734# vdd 1.05f
C9746 a_34362_22312# vdd 0.567f
C9747 X2.X2.X2.X2.X1.X1.X1.vin1 d0 0.267f
C9748 X1.X1.X2.X2.X2.X2.X3.vin2 a_11072_32700# 0.354f
C9749 X1.X1.X2.X2.X2.X2.X2.vin1 X1.X2.vrefh 0.597f
C9750 X1.X1.X2.vrefh a_2582_4198# 0.301f
C9751 d1 X2.X2.X1.X2.X2.X1.X3.vin2 0.15f
C9752 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.X1.vin2 0.22f
C9753 a_8872_5016# a_10686_4110# 1.06e-19
C9754 a_52406_31700# a_54606_30794# 4.2e-20
C9755 a_8486_24076# d1 0.0749f
C9756 X2.X1.X3.vin1 X2.X1.X1.X2.X1.X2.vout 3.08e-19
C9757 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X3.vin1 0.449f
C9758 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X3.vin1 0.206f
C9759 X2.X1.X1.X2.X1.X1.X1.vin2 a_31476_15634# 1.78e-19
C9760 a_19722_18540# d2 0.00132f
C9761 X2.X2.X2.X1.X2.X2.X1.vin1 X2.X2.X2.X1.X2.X2.vrefh 0.267f
C9762 X2.X2.X2.X2.X1.X2.X1.vin2 a_54606_23170# 0.273f
C9763 a_34062_5198# vdd 0.47f
C9764 d1 a_46502_6104# 3.41e-19
C9765 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X1.X3.vin2 0.0903f
C9766 X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X2.X1.vout 0.399f
C9767 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X1.X3.vin2 1.22e-19
C9768 X1.X2.X2.X1.X2.X2.X1.vin2 d1 2.18e-19
C9769 X2.X2.X2.X1.X2.X2.X1.vin1 vdd 0.592f
C9770 X2.X1.X2.X2.X1.X2.X2.vin1 d1 1.03e-19
C9771 X2.X2.X1.X2.X2.X2.vout a_48316_5198# 0.36f
C9772 d3 X2.X1.X1.X3.vin1 0.675f
C9773 a_39966_19358# d0 0.0675f
C9774 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.vout 0.118f
C9775 d3 a_37466_10734# 0.284f
C9776 a_16836_9916# a_16836_8010# 0.00396f
C9777 a_54606_25076# d2 0.00792f
C9778 X1.X2.X2.X1.X1.X1.X3.vin1 X1.X2.X2.X1.X1.X1.X1.vin1 0.206f
C9779 X1.X2.X2.X2.X1.X2.X3.vin1 d0 4.36e-19
C9780 X1.X2.X2.X1.X2.X1.X2.vin1 X2.X1.X1.X2.X1.X2.X1.vin2 0.00232f
C9781 a_46502_8010# a_48616_7064# 2.95e-20
C9782 a_31476_13728# a_31862_13728# 0.419f
C9783 X1.X1.X2.X1.X2.X2.X3.vin1 a_10686_15546# 0.52f
C9784 a_37766_12640# a_38152_12640# 0.419f
C9785 a_11072_23170# d0 0.518f
C9786 d3 X1.X1.X1.X1.X1.X2.X3.vin1 2.1e-19
C9787 a_4396_12822# a_5082_10916# 3.08e-19
C9788 a_39966_23170# vdd 0.553f
C9789 X1.X1.X1.X2.X1.X1.X2.vin1 a_2196_15634# 0.197f
C9790 a_4782_12822# a_4696_10916# 3.3e-19
C9791 a_46502_8010# vdd 0.541f
C9792 a_46116_30882# a_46116_32788# 0.00396f
C9793 a_40352_26982# a_40352_28888# 0.00396f
C9794 X1.X1.X2.X1.X1.X2.X2.vin1 d1 1.03e-19
C9795 a_25326_19358# d0 0.0675f
C9796 d5 a_13696_892# 9.9e-19
C9797 X2.X1.X1.X3.vin1 X2.X1.X2.X3.vin2 1.22e-19
C9798 X2.X1.X1.X1.X1.X2.X1.vin1 a_31476_30882# 1.64e-19
C9799 X1.X1.X2.X3.vin2 a_8486_27888# 7.93e-20
C9800 d2 a_25326_9828# 0.00792f
C9801 a_31862_28976# a_31862_30882# 0.00198f
C9802 X1.X1.X3.vin1 d0 0.0427f
C9803 a_39966_28888# X2.X1.X2.X2.X2.X1.X2.vin1 0.402f
C9804 X1.X1.X1.X2.X1.X1.X3.vin2 a_2582_13728# 8.07e-19
C9805 X1.X1.X1.X1.X2.X1.vout vdd 0.805f
C9806 X2.X1.X2.X1.X2.vrefh X2.X1.X2.X1.X1.X2.X3.vin2 0.161f
C9807 X1.X2.X2.X3.vin1 a_23212_18358# 0.17f
C9808 a_46502_25164# a_46502_23258# 0.00198f
C9809 X2.X2.X1.X2.X1.X2.X3.vin1 a_46502_11822# 0.00207f
C9810 X1.X2.X2.X2.X2.X2.X3.vin2 a_22826_29834# 3.85e-19
C9811 a_33676_16634# vdd 1.05f
C9812 X1.X2.X1.X1.X2.X2.X1.vin1 X1.X2.X1.X1.X2.X2.X1.vin2 0.668f
C9813 d3 a_52406_20264# 4.67e-19
C9814 a_17222_21352# d1 3.41e-19
C9815 X1.X1.X2.X2.X1.X2.X3.vin1 a_10686_23170# 0.52f
C9816 vrefl d1 7.29e-21
C9817 a_31476_21352# d2 0.00274f
C9818 a_10686_19358# d0 0.0675f
C9819 a_34362_7064# X2.X1.X1.X2.X2.X2.X3.vin1 0.00874f
C9820 d0 X2.X1.X1.X2.X2.X2.X1.vin2 0.276f
C9821 X2.X2.X2.X1.X1.X2.X3.vin2 vdd 0.787f
C9822 X1.X2.X2.X2.X2.X2.X1.vin2 d1 0.0985f
C9823 d0 X1.X1.X2.X1.X2.X1.X3.vin1 4.36e-19
C9824 X2.X2.X2.X2.X2.X2.X1.vin1 vdd 0.592f
C9825 a_31476_25164# d0 0.518f
C9826 X1.X1.X1.X1.X2.X1.X2.vin1 a_2196_23258# 0.197f
C9827 d4 a_8486_16452# 8.66e-19
C9828 X1.X2.X1.X3.vin2 X1.X2.X1.X2.X1.X2.X3.vin2 0.102f
C9829 X2.X2.X2.vrefh a_46116_4198# 0.119f
C9830 d1 a_48316_5198# 0.522f
C9831 a_52406_8828# X2.X2.X2.X1.X1.X2.X3.vin1 0.42f
C9832 X1.X2.X1.X2.X1.X2.vout X1.X2.X1.X2.X1.X2.X3.vin1 0.326f
C9833 a_54606_32700# X2.X2.X2.X2.X2.X2.X3.vin2 0.567f
C9834 d2 X2.X2.X2.X2.X2.X2.X3.vin2 5.81e-19
C9835 a_19336_26164# d2 0.0057f
C9836 a_46502_15634# X2.X2.X1.X2.X1.X2.X1.vin1 8.22e-20
C9837 X2.X2.X2.X1.X1.X2.X3.vin2 X2.X2.X2.X1.X1.X2.X1.vin1 2.23e-19
C9838 X2.X2.X2.X1.X1.X2.X2.vin1 a_54992_7922# 1.78e-19
C9839 X2.X2.X2.X2.X1.X1.vout d2 0.00169f
C9840 d3 a_37766_20264# 4.67e-19
C9841 X2.X1.X2.X2.X2.vrefh vdd 0.426f
C9842 X2.X1.X2.X2.X2.X1.vout X2.X1.X2.X2.X2.X1.X3.vin2 0.326f
C9843 X1.X2.X1.X2.X1.X2.X2.vin1 X1.X2.X1.X2.X1.X2.X3.vin2 0.234f
C9844 a_31862_17540# X2.X1.X1.X2.X1.X1.X1.vin2 0.273f
C9845 X1.X2.X2.X1.X2.X2.X1.vin1 X1.X2.X2.X1.X2.X2.vrefh 0.267f
C9846 a_19036_12822# a_19422_12822# 0.419f
C9847 d3 a_25326_11734# 0.00112f
C9848 d4 X2.X1.X2.X1.X2.X2.X2.vin1 8.68e-20
C9849 a_16836_25164# X1.X2.X1.X1.X2.X1.X2.vin1 1.78e-19
C9850 X1.X2.X2.X2.X3.vin2 d1 0.00807f
C9851 X1.X2.X2.X1.X2.X2.X2.vin1 X1.X2.X2.X1.X2.X2.X3.vin2 0.234f
C9852 X2.X1.X2.X1.X1.X2.X1.vin1 a_40352_7922# 0.195f
C9853 a_34362_29936# X2.X1.X1.X1.X1.X1.X3.vin2 0.00815f
C9854 d2 a_49002_29936# 0.254f
C9855 d0 a_2196_9916# 0.518f
C9856 a_40352_11734# d1 2.25e-20
C9857 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X3.vin2 0.581f
C9858 X2.X2.X1.X3.vin1 X2.X2.X1.X3.vin2 0.552f
C9859 d1 a_33976_7064# 0.00613f
C9860 X2.X1.X1.X1.X2.X2.X1.vin2 a_31862_19446# 8.88e-20
C9861 a_31862_27070# vdd 0.542f
C9862 a_46502_23258# d1 0.00148f
C9863 d2 a_8186_14586# 0.0191f
C9864 d3 a_23126_20264# 4.67e-19
C9865 X1.X1.X2.X2.X1.X2.X3.vin2 a_8486_24076# 0.277f
C9866 X1.X1.X2.X2.X1.X2.X2.vin1 X1.X1.X2.X2.X1.X2.X3.vin1 0.00117f
C9867 a_2582_13728# vdd 0.553f
C9868 X1.X1.X1.X1.X2.X2.X1.vin2 d0 0.276f
C9869 a_33676_31882# vdd 1.05f
C9870 a_39966_6016# a_40352_6016# 0.419f
C9871 X2.X1.X2.X3.vin2 a_37766_20264# 5.21e-19
C9872 X2.X1.X2.X1.X2.X1.X3.vin1 a_37466_10734# 0.00837f
C9873 X1.X2.X1.X1.X3.vin2 X1.X2.X1.X1.X2.X1.X3.vin2 0.0533f
C9874 X1.X2.X2.X1.X1.X2.vrefh X1.X2.X2.X1.X1.X1.X3.vin2 0.165f
C9875 a_31862_25164# X2.X1.X1.X1.X2.X1.X1.vin2 0.273f
C9876 X2.X1.X1.X2.X2.X1.X1.vin2 a_31862_8010# 8.88e-20
C9877 d1 a_19422_5198# 0.0751f
C9878 X1.X2.X1.X2.X2.X2.X1.vin1 d1 0.0118f
C9879 a_31862_6104# X2.X1.X1.X2.X2.X2.X1.vin1 0.417f
C9880 a_31476_6104# X2.X1.X1.X2.X2.X2.X3.vin1 0.354f
C9881 a_4782_12822# X1.X1.X1.X2.X1.X2.X3.vin2 0.277f
C9882 X1.X1.X2.X2.X2.X1.X2.vin1 vdd 0.576f
C9883 X2.X2.X1.X1.X2.vrefh X2.X2.X1.X1.X2.X1.X1.vin1 0.267f
C9884 d3 X2.X1.X1.X2.X2.X1.X1.vin1 6.34e-20
C9885 X2.X1.X2.X3.vin1 d2 6.42e-19
C9886 X1.X2.X2.X2.X1.X2.X2.vin1 X1.X2.X2.X2.X1.X2.X3.vin2 0.234f
C9887 X2.X1.X2.X2.X1.X1.X3.vin1 X2.X1.X2.X1.X2.X2.X3.vin2 1.22e-19
C9888 X2.X1.X1.X2.vrefh X2.X1.X1.X2.X1.X1.X3.vin1 2.33e-19
C9889 a_5082_14688# X1.X1.X1.X2.X3.vin1 0.436f
C9890 X1.X1.X1.X2.X2.X1.X3.vin1 X1.X1.X1.X2.X2.X1.X3.vin2 0.581f
C9891 X1.X2.X1.X1.X2.X2.X3.vin1 a_17222_19446# 0.00207f
C9892 a_48316_24258# a_49002_22312# 2.86e-19
C9893 a_48702_24258# a_48616_22312# 3.14e-19
C9894 X1.X1.X2.X2.X2.X2.X3.vin1 a_10686_30794# 0.52f
C9895 a_2196_32788# X1.X1.X1.X1.X1.X1.X1.vin2 0.12f
C9896 X1.X1.X1.X2.X2.vrefh a_2582_9916# 8.22e-20
C9897 a_10686_26982# vdd 0.553f
C9898 a_11072_17452# d0 0.515f
C9899 d1 X2.X1.X2.X1.X1.X2.X1.vin2 0.00406f
C9900 X1.X2.X2.X2.X1.X2.X1.vin1 X1.X2.X2.X2.X1.X1.X3.vin2 5.19e-19
C9901 X2.X2.X2.X2.X1.X2.vrefh vdd 0.414f
C9902 X1.X2.X1.X2.X1.X2.X3.vin2 a_19722_10916# 0.00846f
C9903 a_19336_29936# X1.X2.X1.X1.X1.X2.vout 0.0929f
C9904 X2.X1.X3.vin1 X2.X1.X2.vrefh 0.178f
C9905 d4 a_8186_18358# 0.281f
C9906 X2.X1.X2.X2.X2.X1.X1.vin1 X2.X1.X2.X2.X2.vrefh 0.267f
C9907 a_48702_20446# a_48616_18540# 3.3e-19
C9908 a_40352_28888# X2.X1.X2.X2.X2.X2.vrefh 0.118f
C9909 a_48316_20446# a_49002_18540# 3.08e-19
C9910 d1 a_25712_6016# 2.92e-22
C9911 X1.X2.X3.vin1 X1.X2.X1.X2.X3.vin1 7.18e-19
C9912 X1.X2.X2.vrefh a_16836_4198# 0.119f
C9913 X1.X1.X1.X2.X1.X2.X2.vin1 d1 1.03e-19
C9914 a_46116_27070# d1 2.92e-22
C9915 X1.X2.X1.X1.X2.X1.X1.vin2 d1 4.01e-19
C9916 d3 X2.X2.X1.X2.X3.vin1 0.375f
C9917 X2.X1.X3.vin2 X3.vin2 0.00486f
C9918 d2 a_16836_15634# 0.00414f
C9919 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X2.X2.X3.vin1 0.0131f
C9920 X1.X1.X2.X2.X2.X1.X3.vin1 d1 0.151f
C9921 d3 a_5082_10916# 0.29f
C9922 a_49002_26164# X2.X2.X1.X1.X3.vin2 0.241f
C9923 a_10686_15546# X1.X1.X2.X1.X2.X1.X3.vin2 8.07e-19
C9924 X1.X2.X2.X2.X1.X1.vout a_23126_20264# 0.422f
C9925 a_25326_26982# X1.X2.X2.X2.X1.X2.X3.vin2 8.07e-19
C9926 X1.X1.X1.X1.X2.X1.X3.vin1 d1 0.151f
C9927 a_2582_9916# X1.X1.X1.X2.X2.X1.X1.vin2 0.273f
C9928 d2 X1.X2.X2.X1.X1.X1.X2.vin1 6e-20
C9929 a_10686_6016# d0 0.0489f
C9930 X1.X2.X1.X2.X2.X1.X3.vin1 a_19422_9010# 0.428f
C9931 X1.X2.X1.X1.X2.X1.X1.vin1 d2 0.0105f
C9932 X1.X2.X2.X1.X3.vin1 X1.X2.X2.X1.X1.X2.X3.vin2 0.0565f
C9933 a_49002_14688# X2.X2.X1.X2.X1.X2.X3.vin1 0.00874f
C9934 a_48316_9010# a_48616_7064# 6.1e-19
C9935 X1.X1.X1.X2.X1.X2.vrefh X1.X1.X1.X2.X1.X2.X3.vin1 2.33e-19
C9936 d2 X1.X1.X1.X1.X1.X2.X3.vin2 0.122f
C9937 a_8486_20264# d4 0.0013f
C9938 X1.X2.X2.X2.X2.vrefh d1 0.00745f
C9939 a_19336_10916# a_17222_9916# 5.36e-21
C9940 a_48316_9010# vdd 1.05f
C9941 a_8186_14586# a_8872_12640# 2.86e-19
C9942 X2.X2.X1.X1.X1.X1.X2.vin1 a_46116_32788# 1.78e-19
C9943 a_23212_10734# X1.X2.X2.X1.X1.X2.vout 7.93e-20
C9944 X1.X2.X2.X2.X2.X2.X1.vin1 X1.X2.X2.X2.X2.X2.vrefh 0.267f
C9945 d3 X2.X2.X1.X2.X1.X2.X2.vin1 8.68e-20
C9946 X2.X1.X3.vin2 X2.X1.X2.X1.X2.X2.vout 3.38e-19
C9947 X2.X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X2.X1.X2.vin1 0.564f
C9948 X1.X2.X2.X2.X1.X2.X3.vin1 a_25712_23170# 0.354f
C9949 X2.X1.X2.X1.X1.X2.vout a_37852_6962# 0.0929f
C9950 a_2196_4198# a_2582_4198# 0.419f
C9951 X2.X2.X1.X2.X1.X2.X1.vin2 X2.X2.X1.X2.X2.vrefh 0.076f
C9952 a_48616_29936# X2.X2.X1.X1.X1.X1.X3.vin2 0.00546f
C9953 a_37466_25982# d2 7.13e-19
C9954 X1.X2.X1.X1.X1.X1.X1.vin2 d0 0.201f
C9955 a_19336_10916# d1 0.0126f
C9956 a_10686_21264# a_11072_21264# 0.419f
C9957 a_52492_22210# d1 0.00613f
C9958 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X2.vin1 0.0689f
C9959 X2.X2.X1.X1.X2.X1.X1.vin1 X2.X2.X1.X1.X2.X1.X2.vin1 0.0689f
C9960 a_46502_13728# a_48316_12822# 1.06e-19
C9961 a_19036_24258# a_17222_23258# 1.15e-20
C9962 a_46502_25164# a_48316_24258# 1.06e-19
C9963 X1.X1.X2.X3.vin1 X1.X1.X3.vin2 1.16f
C9964 X1.X2.X1.X2.X2.X2.X1.vin2 a_17222_4198# 8.88e-20
C9965 a_39966_9828# vdd 0.542f
C9966 a_2196_21352# X1.X1.X1.X1.X2.X2.X3.vin1 0.354f
C9967 a_2582_21352# X1.X1.X1.X1.X2.X2.X1.vin1 0.417f
C9968 d0 X2.X2.X2.X1.X2.X1.X2.vin1 0.262f
C9969 X1.X2.X2.X2.X2.X1.X1.vin2 a_25712_26982# 0.12f
C9970 a_25326_26982# X1.X2.X2.X2.X2.X1.X1.vin1 0.417f
C9971 a_54992_9828# X2.X2.X2.X1.X1.X2.X1.vin2 1.78e-19
C9972 a_23126_27888# a_23212_25982# 3.21e-19
C9973 X1.X1.X2.X2.X2.X1.vout X1.X1.X2.X2.X2.X1.X3.vin1 0.118f
C9974 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X1.X3.vin2 0.049f
C9975 X2.X1.X1.X2.X1.X2.X3.vin2 X2.X1.X1.X2.X2.X1.X1.vin2 3.94e-19
C9976 a_46116_32788# a_46502_32788# 0.419f
C9977 d2 a_33976_14688# 0.526f
C9978 a_46116_21352# vdd 1.05f
C9979 d4 X1.X2.X1.X2.X1.X1.X1.vin2 3.99e-21
C9980 X1.X2.X1.X1.X2.X2.vout d2 0.00117f
C9981 a_33676_28070# X2.X1.X1.X1.X1.X2.vout 0.36f
C9982 X2.X2.X1.X1.X2.X1.X3.vin2 X2.X2.X1.X1.X2.X2.X1.vin2 3.94e-19
C9983 X1.X1.X1.X2.X1.X1.X3.vin1 a_4782_16634# 0.428f
C9984 d3 X1.X2.X1.X2.X1.X2.X3.vin2 0.0247f
C9985 X2.X2.X2.X2.X2.X1.vout a_52492_29834# 0.169f
C9986 d3 a_33676_24258# 0.00178f
C9987 X1.X2.X1.X1.X2.X2.vrefh X1.X2.X1.X1.X2.X2.X1.vin2 0.1f
C9988 a_37852_10734# vdd 1.05f
C9989 X1.X2.X1.X2.X2.X1.X3.vin2 a_19336_7064# 0.00546f
C9990 d3 a_4396_9010# 0.00178f
C9991 d4 a_37466_29834# 5.68e-19
C9992 d0 X2.X2.X1.X2.X1.X1.X3.vin1 4.36e-19
C9993 X2.X1.X3.vin2 d1 0.0804f
C9994 a_2582_17540# d2 0.00309f
C9995 d2 X2.X1.X2.X1.X2.X1.X1.vin2 0.231f
C9996 X2.X1.X1.X1.X1.X2.X2.vin1 vdd 0.576f
C9997 X2.X1.X1.X3.vin1 X2.X1.X3.vin1 0.188f
C9998 a_48316_24258# d1 0.521f
C9999 X2.X2.X2.X2.X1.X1.vout a_52492_18358# 1.64e-19
C10000 a_8572_29834# a_10686_28888# 2.95e-20
C10001 d0 X1.X1.X1.X2.X2.X2.X3.vin2 4.34e-19
C10002 X2.X1.X3.vin1 a_37466_10734# 3.93e-19
C10003 a_48702_20446# d4 7.27e-19
C10004 X2.X1.X1.X3.vin2 X2.X1.X1.X2.X3.vin2 0.17f
C10005 a_54606_26982# d3 0.00112f
C10006 a_2196_23258# d1 2.92e-22
C10007 X2.X1.X1.X1.X2.X2.vrefh a_31862_21352# 8.22e-20
C10008 a_2196_6104# d1 2.25e-20
C10009 d0 a_39966_4110# 0.0675f
C10010 d2 a_39966_15546# 0.00393f
C10011 a_16836_25164# X1.X2.X1.X1.X2.X1.X1.vin1 0.195f
C10012 a_10686_17452# X1.X1.X2.X1.X2.X2.X2.vin1 0.402f
C10013 d2 X2.X2.X1.X2.X2.X2.vrefh 0.168f
C10014 d4 a_33976_18540# 0.63f
C10015 a_34062_20446# d4 9.67e-19
C10016 X1.X1.X2.X3.vin2 a_8186_18358# 0.263f
C10017 X2.X1.X1.X1.X1.X1.X3.vin1 a_33676_31882# 0.199f
C10018 X2.X1.X2.X1.X2.X2.X3.vin2 X2.X1.X2.X1.X2.X2.vout 0.08f
C10019 a_8572_29834# a_8872_31700# 6.71e-19
C10020 X1.X1.X1.X1.X2.X1.X3.vin1 X1.X1.X1.X1.X2.vrefh 2.33e-19
C10021 X2.X2.X1.X1.X1.X2.X3.vin2 a_46116_27070# 0.354f
C10022 a_48702_28070# a_46502_27070# 4.77e-21
C10023 X1.X1.X2.X2.X1.X2.X3.vin2 X1.X1.X2.X2.X2.X1.X3.vin1 1.22e-19
C10024 X2.X2.X2.X2.X2.X1.X1.vin1 X2.X2.X2.X2.X2.X1.X2.vin1 0.0689f
C10025 a_33976_22312# a_33676_20446# 6.71e-19
C10026 a_54606_26982# X2.X2.X2.X2.X2.X1.X3.vin2 7.84e-19
C10027 X1.X1.X2.X3.vin1 X1.X1.X1.X2.X3.vin2 7.46e-20
C10028 X1.X2.X1.X2.X1.X2.vrefh a_16836_13728# 1.64e-19
C10029 X1.X2.X2.X2.X2.vrefh a_25712_25076# 0.118f
C10030 a_23212_14586# a_23512_12640# 6.1e-19
C10031 a_4396_28070# X1.X1.X1.X1.X1.X2.X3.vin2 0.101f
C10032 d2 a_11072_11734# 0.00272f
C10033 a_40352_19358# vdd 1.05f
C10034 a_22826_6962# vdd 0.477f
C10035 X2.X2.X3.vin1 d0 0.04f
C10036 d0 X2.X1.X1.X2.X2.vrefh 0.848f
C10037 d0 X2.X2.X1.X2.X1.X2.vrefh 0.848f
C10038 a_25326_23170# d2 0.00479f
C10039 d2 a_31476_8010# 0.00464f
C10040 a_23212_6962# a_23512_5016# 6.1e-19
C10041 X1.X2.X2.X2.vrefh d0 0.848f
C10042 X2.X1.X1.X1.X1.X1.X1.vin2 d4 8.21e-20
C10043 a_31476_19446# a_31862_19446# 0.419f
C10044 a_52106_18358# a_52792_16452# 3.08e-19
C10045 a_4696_29936# X1.X1.X1.X1.X3.vin1 0.363f
C10046 X1.X1.X2.X1.X2.X1.X3.vin1 a_8572_10734# 0.00251f
C10047 a_2582_21352# a_2582_19446# 0.00198f
C10048 a_19422_20446# d4 7.27e-19
C10049 d3 X2.X2.X1.X1.X1.X1.X1.vin1 0.00492f
C10050 a_46502_13728# d1 3.41e-19
C10051 d5 X2.X3.vin1 0.0932f
C10052 d0 X1.X1.X2.X1.X1.X1.X1.vin1 0.269f
C10053 X1.X2.X1.X2.X2.X1.X1.vin2 X1.X2.X1.X2.X2.X1.X2.vin1 0.242f
C10054 X1.X1.X2.X3.vin2 a_8486_20264# 5.21e-19
C10055 d0 X1.X1.X2.X1.X2.vrefh 0.848f
C10056 d0 a_31476_15634# 0.515f
C10057 X2.X2.X2.vrefh X2.X3.vin2 4.75e-20
C10058 d2 a_19036_16634# 3.82e-19
C10059 a_25712_19358# vdd 1.05f
C10060 X2.X2.X2.X2.X2.X1.X2.vin1 d1 1.03e-19
C10061 a_8572_18358# vdd 1.05f
C10062 X1.X1.X2.X1.X2.X2.X3.vin1 d1 0.146f
C10063 a_52792_27888# d2 0.00251f
C10064 X1.X1.X2.X2.vrefh d0 0.848f
C10065 d1 a_13696_892# 4.67e-19
C10066 X1.X1.X2.X1.X1.X1.X3.vin2 a_11072_6016# 0.354f
C10067 a_2196_25164# d2 0.00272f
C10068 d3 X1.X1.X2.X2.X1.X1.vout 0.00883f
C10069 X2.X1.X2.X2.X2.X1.X3.vin1 a_37852_25982# 0.00251f
C10070 X2.X2.X1.X3.vin2 a_48702_9010# 7.93e-20
C10071 a_4696_26164# X1.X1.X1.X1.X2.X1.X3.vin1 0.00251f
C10072 a_34362_26164# X2.X1.X1.X3.vin1 0.509f
C10073 d2 a_39966_30794# 6.36e-19
C10074 a_54992_17452# d1 2.92e-22
C10075 a_2582_13728# X1.X1.X1.X2.X1.X2.X1.vin2 0.273f
C10076 a_37852_6962# X2.X1.X2.X1.X1.X1.X3.vin2 0.00546f
C10077 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X3.vin1 0.206f
C10078 a_19722_18540# X1.X2.X3.vin2 6.58e-20
C10079 a_37852_18358# a_37766_16452# 3.3e-19
C10080 a_54606_25076# X2.X2.X2.X2.X1.X2.X3.vin1 0.00207f
C10081 d2 X1.X1.X1.X2.X1.X1.X3.vin2 0.169f
C10082 a_16836_23258# d0 0.515f
C10083 a_48702_28070# X2.X2.X1.X1.X1.X2.vout 0.418f
C10084 a_33676_28070# a_31862_28976# 1.06e-19
C10085 X2.X1.X1.X1.X1.X2.X2.vin1 X2.X1.X1.X1.X1.X2.X1.vin1 0.0689f
C10086 X2.X1.X2.X1.X2.X2.X3.vin2 d1 0.151f
C10087 X1.X2.X1.X2.X2.vrefh X1.X1.X2.X1.X2.vrefh 0.117f
C10088 a_11072_19358# vdd 1.05f
C10089 a_38152_16452# a_39966_15546# 1.06e-19
C10090 X1.X1.X1.X1.X1.X1.X1.vin2 a_2196_30882# 1.78e-19
C10091 X2.X1.X1.X2.X1.X2.vrefh a_31862_15634# 0.3f
C10092 d2 a_19036_9010# 0.00167f
C10093 X2.X1.X2.X1.X1.X1.X2.vin1 vdd 0.578f
C10094 a_17222_17540# a_19036_16634# 1.06e-19
C10095 d3 a_8186_29834# 0.00329f
C10096 a_37852_29834# a_39966_30794# 2.68e-20
C10097 X2.X1.X1.X1.X2.X1.X1.vin1 vdd 0.592f
C10098 d2 X2.X2.X2.X1.X2.X2.X2.vin1 0.0314f
C10099 X2.X2.X1.X3.vin1 X2.X2.X1.X1.X3.vin1 0.199f
C10100 a_40352_7922# X2.X1.X2.X1.X1.X2.vrefh 1.64e-19
C10101 a_33976_22312# X2.X1.X1.X1.X2.X2.X3.vin1 0.00329f
C10102 a_16836_19446# a_17222_19446# 0.419f
C10103 a_48616_29936# X2.X2.X1.X1.X1.X2.X3.vin1 0.00329f
C10104 X1.X1.X2.X2.X2.X2.X2.vin1 d0 0.199f
C10105 X2.X2.X1.X1.X1.X2.vrefh d0 0.848f
C10106 d2 a_52106_14586# 0.0191f
C10107 X2.X2.X2.X2.X1.X1.X3.vin2 a_52406_20264# 0.267f
C10108 X2.X2.X2.X2.X1.X1.X2.vin1 X2.X2.X2.X2.X1.X1.X3.vin1 0.00117f
C10109 X2.X2.X1.X1.X2.X2.X3.vin1 X2.X2.X1.X2.vrefh 0.00118f
C10110 X1.X1.X2.X2.X2.X1.X3.vin2 a_11072_28888# 0.354f
C10111 a_22826_22210# d1 0.0422f
C10112 X1.X1.X1.X1.X3.vin2 d2 0.00194f
C10113 a_19036_28070# d1 0.521f
C10114 X2.X2.vrefh X2.X2.X1.X1.X1.X1.X1.vin2 0.109f
C10115 d2 a_40352_32700# 3.9e-19
C10116 d0 X2.X1.X1.X2.X1.X2.X1.vin2 0.276f
C10117 X1.X1.X1.X1.X1.X2.X1.vin1 X1.X1.X1.X1.X1.X2.X3.vin1 0.206f
C10118 a_46116_9916# a_46116_8010# 0.00396f
C10119 X2.X1.X2.X2.X1.X2.X3.vin2 a_38152_24076# 0.101f
C10120 X2.X1.X1.X1.X2.X1.X1.vin2 X2.X1.X1.X1.X2.X2.vrefh 0.076f
C10121 X1.X2.X1.X1.X2.vrefh d2 0.158f
C10122 X2.X1.X1.X2.X1.X1.X2.vin1 X2.X1.X1.X2.X1.X1.X3.vin2 0.234f
C10123 X1.X1.X1.X2.X1.X1.X1.vin2 X1.X1.X1.X2.X1.X1.X2.vin1 0.242f
C10124 a_31476_32788# X2.X1.X1.X1.X1.X1.X1.vin1 0.195f
C10125 a_31476_30882# d0 0.515f
C10126 d2 a_19036_31882# 0.0017f
C10127 d0 X1.X2.X1.X2.X1.X2.X3.vin1 4.36e-19
C10128 X1.X1.X1.X2.X2.X1.X1.vin1 vdd 0.592f
C10129 a_19722_29936# d1 0.0422f
C10130 d3 a_4696_18540# 7.7e-20
C10131 a_46116_28976# d0 0.518f
C10132 a_22826_25982# X1.X2.X2.X2.X3.vin2 0.263f
C10133 X1.X1.X2.X2.X2.X2.X3.vin1 d1 0.147f
C10134 X2.X2.X1.X3.vin2 a_48616_10916# 0.355f
C10135 d2 a_48616_7064# 0.608f
C10136 d2 X2.X2.X2.X1.X2.X2.vrefh 0.168f
C10137 a_25326_32700# a_25712_32700# 0.419f
C10138 X1.X1.X1.X2.X3.vin1 a_4696_10916# 0.17f
C10139 X1.X2.X2.X1.X3.vin1 a_23212_6962# 0.363f
C10140 a_37766_12640# d1 0.0749f
C10141 X1.X1.X2.X2.X1.X1.X2.vin1 vdd 0.576f
C10142 X1.X1.X2.X1.X2.vrefh a_10686_9828# 0.3f
C10143 a_49002_22312# X2.X2.X1.X1.X2.X2.X3.vin2 3.85e-19
C10144 X2.X2.X1.X1.X2.X2.vout a_48702_20446# 0.418f
C10145 a_19336_22312# X1.X2.X1.X1.X2.X2.vout 0.0929f
C10146 X2.X1.X2.X2.X1.X1.X1.vin1 a_39966_17452# 8.22e-20
C10147 d2 X1.X1.X1.X1.X1.X1.X3.vin2 0.0661f
C10148 a_10686_7922# a_8572_6962# 2.68e-20
C10149 X2.X1.X2.X2.X1.X1.X1.vin2 X2.X1.X2.X1.X2.X2.X3.vin2 3.94e-19
C10150 d3 X1.X2.X1.X1.X1.X1.X3.vin1 0.0103f
C10151 a_54606_32700# vdd 0.541f
C10152 X1.X2.X1.X1.X2.X1.X3.vin1 a_17222_23258# 0.00207f
C10153 X1.X2.X2.X1.X2.X2.X3.vin1 X1.X2.X2.X1.X2.X2.X1.vin2 0.216f
C10154 X2.X1.X2.X2.X2.X1.vout X2.X1.X2.X2.X3.vin2 0.399f
C10155 a_17222_13728# a_17222_11822# 0.00198f
C10156 a_16836_32788# X1.X2.X1.X1.X1.X1.X3.vin1 0.354f
C10157 a_17222_32788# X1.X2.X1.X1.X1.X1.X1.vin1 0.42f
C10158 d2 vdd 63.9f
C10159 a_23126_16452# a_25326_15546# 4.2e-20
C10160 a_2196_19446# a_2582_19446# 0.419f
C10161 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X3.vin2 0.0321f
C10162 a_8186_10734# vdd 0.489f
C10163 d0 a_31862_17540# 0.0675f
C10164 X2.X2.X1.X2.X2.X1.X1.vin1 X2.X2.X1.X2.X2.X1.X1.vin2 0.668f
C10165 X1.X2.X1.X2.X1.X2.X3.vin1 X1.X2.X1.X2.X2.vrefh 0.00118f
C10166 X1.X2.X2.X1.X2.X1.X3.vin2 X1.X2.X2.X1.X2.X1.X3.vin1 0.581f
C10167 X1.X2.X3.vin1 X1.X2.X2.X1.X1.X2.vout 1.71e-19
C10168 d0 a_54992_11734# 0.518f
C10169 X1.X2.X2.X2.X1.X2.vrefh X1.X2.X2.X2.X1.X1.X2.vin1 0.564f
C10170 X1.X1.X1.X2.X2.X1.X1.vin2 X1.X1.X1.X2.X2.X2.vrefh 0.076f
C10171 X1.X1.X2.X1.X1.X2.X3.vin2 a_8872_8828# 0.101f
C10172 X1.X1.X3.vin1 a_8486_16452# 8.66e-20
C10173 d4 a_52106_18358# 0.281f
C10174 d4 X1.X1.X1.X1.X1.X2.vout 0.0921f
C10175 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X1.X2.X1.X2.vrefh 0.1f
C10176 d3 X1.X1.X2.X2.X1.X2.X2.vin1 8.68e-20
C10177 a_31862_9916# X2.X1.X1.X2.X2.X1.X3.vin2 7.84e-19
C10178 d2 X2.X2.X2.X1.X1.X2.X1.vin1 0.0114f
C10179 X1.X1.X2.X3.vin1 d1 0.00955f
C10180 X2.X2.X1.X2.X3.vin2 a_48702_9010# 0.00101f
C10181 a_37852_29834# vdd 1.05f
C10182 a_48702_28070# d3 0.00107f
C10183 a_23126_24076# a_22826_22210# 5.55e-20
C10184 X2.X1.X2.X2.X1.X1.vout a_38152_20264# 0.359f
C10185 a_37852_25982# X2.X1.X2.X2.X1.X2.X3.vin2 0.00535f
C10186 a_17222_17540# vdd 0.553f
C10187 d0 X2.X2.X2.X1.X2.X2.X1.vin1 0.267f
C10188 a_46116_15634# a_46502_15634# 0.419f
C10189 X2.X2.X2.X2.X2.X1.X3.vin1 a_52792_27888# 0.199f
C10190 X1.X1.X2.X1.X2.X2.vrefh a_10686_13640# 0.3f
C10191 X1.X2.X1.X2.X2.X2.vrefh a_16836_8010# 0.118f
C10192 a_16836_23258# a_16836_21352# 0.00396f
C10193 X2.X2.X2.X2.X1.X1.X2.vin1 a_54992_21264# 0.197f
C10194 X2.X1.X3.vin2 a_37466_6962# 0.00111f
C10195 a_19336_7064# a_19722_7064# 0.419f
C10196 X2.X2.X1.X1.X2.X1.X3.vin2 a_46502_23258# 0.567f
C10197 X1.X2.X2.X2.X1.X2.vout vdd 0.697f
C10198 X2.X2.X1.X1.X1.X2.X3.vin1 X2.X2.X1.X1.X1.X1.X3.vin2 1.22e-19
C10199 X1.X1.X2.X2.X1.X1.X3.vin1 d1 0.146f
C10200 a_46502_21352# X2.X2.X1.X1.X2.X2.X3.vin1 0.52f
C10201 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X2.vin1 0.0689f
C10202 a_2582_32788# d1 2.7e-19
C10203 a_39966_23170# d0 0.0675f
C10204 X1.X2.X2.X1.X2.X1.X1.vin1 X1.X2.X2.X1.X2.vrefh 0.267f
C10205 d6 d7 5.23e-19
C10206 X1.X1.X1.X1.X2.X1.vout a_5082_22312# 0.383f
C10207 X2.X2.X2.X1.X2.X1.vout X2.X2.X2.X1.X2.X1.X3.vin2 0.326f
C10208 X1.X2.vrefh d2 0.0108f
C10209 X1.X1.X2.X1.X1.X1.X3.vin2 vdd 0.937f
C10210 d0 a_46502_8010# 0.0489f
C10211 d2 a_33676_9010# 0.00167f
C10212 a_38152_31700# a_39966_30794# 1.06e-19
C10213 X2.X1.X1.X1.X1.X2.vrefh a_31862_30882# 0.3f
C10214 a_52492_29834# a_54606_30794# 2.68e-20
C10215 X1.X1.X1.X1.X2.X2.X3.vin2 d2 0.113f
C10216 a_25712_13640# d1 2.92e-22
C10217 X1.X2.X2.X2.X1.X2.X3.vin1 X1.X2.X2.X2.X1.X2.vrefh 2.33e-19
C10218 a_33976_18540# X2.X1.X1.X3.vin2 0.0927f
C10219 a_52106_6962# vdd 0.477f
C10220 a_31862_6104# a_31862_4198# 0.00198f
C10221 X1.X1.X2.X1.X1.X2.X3.vin2 X1.X1.X2.X1.X1.X2.X1.vin1 2.23e-19
C10222 X1.X1.X2.X1.X1.X2.X2.vin1 a_11072_7922# 1.78e-19
C10223 a_48616_10916# X2.X2.X1.X2.X3.vin2 0.0927f
C10224 X1.X2.X1.X1.X2.vrefh a_16836_25164# 1.64e-19
C10225 a_38152_16452# vdd 1.05f
C10226 X1.X2.X2.X1.X2.X1.X1.vin2 a_25326_11734# 0.273f
C10227 X2.X1.X1.X1.X1.X2.X1.vin2 d1 0.00406f
C10228 X2.X1.X2.X1.X1.X1.X2.vin1 X2.X1.X2.X1.X1.X1.X3.vin1 0.00117f
C10229 X1.X1.X2.X1.X2.X1.X3.vin2 d1 0.15f
C10230 X2.X1.X2.X1.X1.X1.X3.vin2 a_37766_5016# 0.267f
C10231 a_19422_16634# X1.X2.X1.X2.X3.vin1 1.52e-19
C10232 X1.X1.X1.X2.X3.vin1 X1.X1.X1.X2.X1.X2.X3.vin2 0.0565f
C10233 X2.X1.X2.X2.X2.X1.X1.vin1 d2 0.0105f
C10234 X1.X2.X1.X2.X1.X1.vout a_19722_14688# 0.387f
C10235 d2 X1.X2.X2.X1.X2.X1.X2.vin1 0.0318f
C10236 a_2196_6104# X1.X1.X1.X2.X2.X2.X1.vin2 0.12f
C10237 X1.X2.X1.X1.X1.X2.X3.vin1 d1 0.146f
C10238 X2.X1.X1.X1.X1.X1.X2.vin1 X2.X1.X1.X1.X1.X1.X3.vin2 0.234f
C10239 a_39966_30794# X2.X1.X2.X2.X2.X2.X3.vin2 7.84e-19
C10240 X2.X2.X1.X2.X2.X1.X3.vin2 a_46116_8010# 0.354f
C10241 d0 X2.X2.X2.X1.X1.X2.X3.vin2 4.34e-19
C10242 a_33676_28070# X2.X1.X1.X1.X1.X2.X3.vin2 0.101f
C10243 X1.X2.X2.X2.X2.X2.X2.vin1 vdd 0.578f
C10244 a_8186_25982# d1 0.0316f
C10245 X2.X2.X2.X2.X2.X2.X1.vin1 d0 0.267f
C10246 d2 X2.X1.X1.X1.X1.X2.X1.vin1 0.0114f
C10247 a_8872_12640# vdd 1.05f
C10248 d2 a_33976_10916# 0.0057f
C10249 a_23512_20264# a_23212_18358# 6.2e-19
C10250 a_25326_28888# X1.X2.X2.X2.X2.X2.X1.vin1 8.22e-20
C10251 X1.X2.X2.X2.X2.X1.X3.vin2 X1.X2.X2.X2.X2.X2.X1.vin2 3.94e-19
C10252 a_25326_17452# d1 0.00148f
C10253 X1.X1.X2.X1.X2.vrefh X1.X1.X2.X1.X1.X2.X3.vin1 0.00118f
C10254 X1.X2.X1.X2.X2.X2.X1.vin2 vdd 0.387f
C10255 X1.X2.X2.X2.X2.X1.X3.vin1 X1.X2.X2.X2.X2.vrefh 2.33e-19
C10256 X2.X1.X2.X2.X2.vrefh d0 0.848f
C10257 X1.X1.X3.vin1 a_8186_18358# 5.87e-20
C10258 X2.X2.X2.X2.X1.X2.X1.vin1 X2.X2.X2.X2.X1.X1.X3.vin2 5.19e-19
C10259 X2.X1.X2.X1.X2.X1.X2.vin1 X2.X1.X2.X1.X2.X1.X1.vin2 0.242f
C10260 X1.X2.X2.X2.X1.X2.X1.vin1 X2.X1.X1.X1.X2.X2.vrefh 0.00437f
C10261 X2.X2.X2.X2.X3.vin1 a_52406_20264# 1.52e-19
C10262 d2 X2.X1.X1.X2.X1.X1.X1.vin2 0.231f
C10263 X2.X1.X2.X2.X1.X2.X2.vin1 X2.X1.X2.X2.X1.X2.X1.vin2 0.242f
C10264 X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.X3.vin1 0.00789f
C10265 a_39966_13640# a_39966_11734# 0.00198f
C10266 a_39966_25076# a_39966_23170# 0.00198f
C10267 a_16836_25164# vdd 1.05f
C10268 X3.vin2 X2.X3.vin1 0.145f
C10269 X2.X1.X2.X2.X2.X1.vout X2.X1.X2.X2.X2.X2.vout 0.514f
C10270 X2.X2.X2.X2.X2.X1.X3.vin1 vdd 0.997f
C10271 d3 a_22826_18358# 0.0469f
C10272 X2.X1.X2.X2.X2.X1.vout d1 0.0238f
C10273 a_46116_21352# X2.X2.X1.X1.X2.X2.X2.vin1 1.78e-19
C10274 a_2196_28976# X1.X1.X1.X1.X1.X2.X1.vin2 0.12f
C10275 a_23126_31700# a_25326_30794# 4.2e-20
C10276 X1.X2.X2.X2.X2.X2.X3.vin1 X1.X2.X2.X2.X2.X2.X1.vin2 0.22f
C10277 d2 X1.X2.X1.X2.X1.X1.X3.vin1 0.104f
C10278 a_4396_28070# vdd 1.05f
C10279 a_4696_14688# d1 0.00613f
C10280 d2 X1.X2.X1.X2.X1.X2.vout 0.00124f
C10281 a_25712_11734# a_25712_9828# 0.00396f
C10282 a_10686_11734# a_11072_11734# 0.419f
C10283 X1.X1.X2.X3.vin1 a_8486_12640# 5.28e-19
C10284 a_31862_27070# d0 0.0489f
C10285 X2.X1.X2.X2.X2.X2.X3.vin2 a_40352_32700# 0.354f
C10286 X2.X2.X1.X1.X2.X2.X3.vin2 d1 0.151f
C10287 X1.X2.X2.X2.X3.vin2 X1.X2.X2.X2.X2.X1.X3.vin2 0.0533f
C10288 X1.X2.X2.X1.X2.X2.X1.vin2 X2.X1.X1.X2.X1.X1.X2.vin1 0.00232f
C10289 X1.X1.X2.X2.X3.vin1 X1.X1.X2.X2.X1.X1.vout 0.131f
C10290 X1.X2.X1.X2.X2.X2.X3.vin1 X1.X2.X1.X2.X2.X2.vrefh 2.33e-19
C10291 a_38152_31700# vdd 1.05f
C10292 X2.X1.X2.X1.X2.X2.X1.vin2 X2.X1.X2.X1.X2.X1.X3.vin2 3.94e-19
C10293 d2 X2.X1.X2.X1.X1.X1.X3.vin1 3e-19
C10294 X2.X1.X2.X1.X2.X2.X1.vin1 a_39966_13640# 8.22e-20
C10295 a_46116_9916# X2.X2.X1.X2.X2.X1.X2.vin1 1.78e-19
C10296 X2.X2.X2.X2.X2.vrefh X2.X2.X2.X2.X1.X2.X2.vin1 0.564f
C10297 d0 a_2582_13728# 0.0675f
C10298 a_2582_27070# a_2582_28976# 0.00198f
C10299 a_39966_21264# a_37766_20264# 4.77e-21
C10300 X1.X1.X1.X2.X1.X2.X2.vin1 a_2582_11822# 0.402f
C10301 a_17222_17540# X1.X2.X1.X2.X1.X1.X3.vin1 0.52f
C10302 X2.X2.X1.X2.X1.X2.X2.vin1 a_46502_11822# 0.402f
C10303 a_34362_18540# d1 0.0424f
C10304 X1.X1.X2.X1.X3.vin2 a_8572_14586# 0.363f
C10305 X1.X1.X2.X2.X2.X1.X2.vin1 d0 0.262f
C10306 X2.X1.X1.X2.X2.X1.X3.vin2 X2.X1.X1.X2.X2.X2.X1.vin1 5.19e-19
C10307 d2 X1.X1.X2.X1.X1.X1.vout 0.115f
C10308 X2.X1.X1.X1.X2.X2.X3.vin2 d1 0.151f
C10309 X2.X2.X2.X2.X1.X2.vout d2 0.00124f
C10310 X2.X1.X1.X2.X2.X1.X3.vin1 X2.X1.X1.X2.X2.X2.vrefh 0.00118f
C10311 a_46116_30882# a_46502_30882# 0.419f
C10312 a_25326_13640# a_23512_12640# 1.15e-20
C10313 X1.X1.X2.X1.X3.vin1 a_8186_6962# 0.436f
C10314 X2.X1.X2.X2.X2.vrefh a_39966_25076# 0.3f
C10315 a_8486_20264# a_10686_19358# 4.2e-20
C10316 X1.X1.X2.X2.X1.X1.X3.vin1 X1.X1.X2.X2.X1.X1.X1.vin2 0.216f
C10317 a_39966_9828# a_40352_9828# 0.419f
C10318 X2.X1.X2.X2.X2.X2.X3.vin2 vdd 0.738f
C10319 a_40352_4110# vdd 1.05f
C10320 a_17222_13728# X1.X2.X1.X2.X1.X2.X2.vin1 8.88e-20
C10321 X2.X1.X2.X1.X2.vrefh vdd 0.426f
C10322 a_34362_26164# a_33676_24258# 2.97e-19
C10323 a_31862_9916# X2.X1.X1.X2.X2.X1.X1.vin1 0.417f
C10324 a_19336_22312# vdd 1.05f
C10325 a_31476_9916# X2.X1.X1.X2.X2.X1.X3.vin1 0.354f
C10326 d3 X2.X1.X1.X2.X1.X2.X3.vin1 2.1e-19
C10327 a_23512_12640# a_23212_10734# 6.2e-19
C10328 a_33976_26164# a_34062_24258# 3.21e-19
C10329 a_39966_32700# d1 0.00148f
C10330 X1.X1.X1.X2.X2.X2.X1.vin1 X1.X1.X1.X2.X2.X2.X2.vin1 0.0689f
C10331 a_10686_26982# d0 0.0675f
C10332 a_2582_6104# a_4396_5198# 1.06e-19
C10333 a_37852_22210# a_37766_20264# 3.14e-19
C10334 X1.X1.X2.X3.vin2 X1.X1.X2.X2.X1.X2.X3.vin1 0.0131f
C10335 X2.X2.X2.X2.X1.X2.vrefh d0 0.844f
C10336 X2.X2.X1.X2.X1.X2.X1.vin1 X2.X2.X1.X2.X1.X2.X1.vin2 0.668f
C10337 a_33976_7064# a_33676_5198# 6.71e-19
C10338 X1.X2.X1.X1.X2.X2.X3.vin2 d1 0.151f
C10339 X2.X2.X2.X1.X1.X1.X2.vin1 X2.X2.X2.X1.X1.X1.X1.vin1 0.0689f
C10340 d4 X1.X2.X1.X3.vin2 0.12f
C10341 X2.X2.X2.X1.X1.X1.X3.vin2 a_54606_4110# 7.84e-19
C10342 X1.X1.X2.X2.X2.vrefh X1.X1.X2.X2.X1.X2.X3.vin1 0.00118f
C10343 X1.X1.X2.X1.X2.X1.X2.vin1 X1.X1.X2.X1.X2.X1.X3.vin1 0.00117f
C10344 X1.X1.X2.X1.X2.X1.X3.vin2 a_8486_12640# 0.267f
C10345 a_52492_18358# vdd 1.05f
C10346 a_31862_11822# vdd 0.542f
C10347 X2.X1.X1.X1.X1.X1.X3.vin1 d2 0.00317f
C10348 X1.X1.X2.X2.X3.vin2 vdd 1.29f
C10349 X1.X2.X1.X2.X1.X2.vrefh d1 0.0071f
C10350 X2.X2.X2.X1.X2.X2.X3.vin1 X2.X2.X2.X1.X2.X2.X1.vin1 0.206f
C10351 X2.X2.X1.X2.X2.X1.X1.vin1 d1 0.0118f
C10352 a_4782_9010# a_2582_8010# 4.77e-21
C10353 X2.X1.X1.X1.X1.X2.X3.vin2 X2.X1.X1.X1.X2.X1.X3.vin1 1.22e-19
C10354 a_34062_12822# a_31862_11822# 4.77e-21
C10355 a_34062_16634# a_34362_14688# 4.19e-20
C10356 X2.X1.X1.X2.X1.X1.vout a_33976_14688# 0.169f
C10357 X2.X1.X1.X2.X1.X2.X3.vin2 a_31476_11822# 0.354f
C10358 X2.X2.X2.X1.X2.X2.vout a_52792_16452# 0.36f
C10359 X2.X2.X1.X3.vin2 X2.X2.X1.X2.X1.X1.X3.vin2 0.0943f
C10360 X2.X2.X1.X2.X1.X1.X2.vin1 a_46502_15634# 0.402f
C10361 d1 X2.X3.vin1 0.0443f
C10362 a_48316_24258# X2.X2.X1.X1.X2.X1.X3.vin2 0.1f
C10363 a_39966_21264# X2.X1.X2.X2.X1.X1.X2.vin1 0.402f
C10364 X2.X2.X2.X2.X1.X1.X2.vin1 d1 1.03e-19
C10365 a_2582_15634# d1 0.00148f
C10366 X1.X1.X2.X1.X1.X1.X3.vin2 X1.X1.X2.X1.X1.X1.vout 0.342f
C10367 X1.X2.X3.vin1 X1.X2.X2.X1.X1.X1.vout 5.53e-20
C10368 d3 a_52106_29834# 2.73e-19
C10369 X1.X2.X3.vin2 X1.X3.vin2 0.147f
C10370 a_8186_25982# X1.X1.X2.X2.X1.X2.X3.vin2 0.00846f
C10371 X1.X2.X1.X1.X1.X1.X1.vin1 X1.X2.X1.X1.X1.X1.X3.vin2 2.23e-19
C10372 X2.X1.X1.X1.X3.vin2 X2.X1.X1.X1.X2.X2.X3.vin1 1.42e-20
C10373 a_23126_27888# d3 0.00148f
C10374 a_52792_8828# vdd 1.05f
C10375 a_11072_9828# X1.X1.X2.X1.X1.X2.X1.vin2 1.78e-19
C10376 a_2582_6104# a_4696_7064# 2.68e-20
C10377 a_52106_29834# X2.X2.X2.X2.X2.X2.vout 0.263f
C10378 a_33976_26164# d1 0.0126f
C10379 d1 a_54992_4110# 2.25e-20
C10380 X2.X2.X1.X1.X3.vin2 d2 0.00194f
C10381 X1.X1.X1.X2.X2.X2.X3.vin1 a_2582_4198# 0.00207f
C10382 a_8186_22210# a_8872_20264# 2.86e-19
C10383 a_10686_11734# vdd 0.553f
C10384 a_31476_6104# X2.X1.X1.X2.X2.X2.X2.vin1 1.78e-19
C10385 X2.X1.X2.X2.X1.X2.X3.vin1 a_39966_23170# 0.52f
C10386 a_2582_8010# d1 0.00148f
C10387 X2.X2.X2.X2.X1.X1.X3.vin2 X2.X2.X2.X2.X1.X1.X1.vin2 8.93e-19
C10388 X2.X2.X2.X2.X1.X1.X2.vin1 a_54606_19358# 8.88e-20
C10389 a_19336_18540# X1.X2.X3.vin1 0.354f
C10390 a_52106_29834# X2.X2.X2.X2.X2.X1.X3.vin2 0.00815f
C10391 d2 X1.X1.X1.X2.X1.X2.X1.vin2 0.226f
C10392 a_23212_14586# a_25326_13640# 2.95e-20
C10393 d3 a_48616_18540# 7.7e-20
C10394 X2.X1.X2.X2.X1.X2.vout a_38152_24076# 0.36f
C10395 X2.X2.X2.X1.X1.X1.X3.vin1 a_54992_4110# 0.354f
C10396 X2.X1.X1.X1.X2.X1.X2.vin1 a_31476_23258# 0.197f
C10397 a_2582_28976# d1 3.41e-19
C10398 X1.X2.X2.X2.X2.X2.X1.vin2 X2.X1.X1.X1.X1.X1.X2.vin1 0.00232f
C10399 X1.X2.X1.X1.X1.X2.vrefh d1 0.0738f
C10400 X1.X2.X2.X2.X2.X1.X1.vin2 X1.X2.X2.X2.X2.X1.X2.vin1 0.242f
C10401 a_25326_26982# a_25326_28888# 0.00198f
C10402 d0 a_39966_9828# 0.0489f
C10403 a_49002_14688# X2.X2.X1.X2.X3.vin1 0.436f
C10404 X1.X1.X2.X1.X2.X2.X2.vin1 X1.X1.X2.X1.X2.X2.X1.vin2 0.242f
C10405 a_10686_17452# a_10686_15546# 0.00198f
C10406 a_22826_14586# d1 0.0422f
C10407 d2 a_16836_28976# 0.00351f
C10408 X2.X2.X1.X2.X2.X1.X2.vin1 X2.X2.X1.X2.X2.X1.X3.vin2 0.234f
C10409 a_2582_32788# a_4396_31882# 1.06e-19
C10410 X1.X2.X2.X1.X1.X2.X3.vin2 a_22826_6962# 3.85e-19
C10411 a_37766_16452# X2.X1.X2.X1.X2.X2.vout 0.418f
C10412 a_46116_11822# d1 2.92e-22
C10413 a_43362_892# vdd 0.473f
C10414 X1.X1.X2.X1.X1.X2.vout a_8872_8828# 0.36f
C10415 X2.X2.X1.X2.X2.X2.vout X2.X2.X1.X2.X2.X2.X3.vin1 0.335f
C10416 a_4696_10916# a_5082_10916# 0.414f
C10417 X2.X2.X1.X2.X1.X2.vrefh a_46116_13728# 1.64e-19
C10418 X2.X1.X2.X2.X3.vin2 a_37766_31700# 9.7e-20
C10419 X2.X1.X2.X1.X2.X1.X2.vin1 vdd 0.576f
C10420 a_37466_22210# d2 0.0191f
C10421 a_5082_29936# X1.X1.X1.X1.X1.X2.X3.vin2 3.85e-19
C10422 a_4396_16634# a_4696_14688# 6.1e-19
C10423 X1.X1.X1.X1.X3.vin1 a_4782_28070# 9.54e-19
C10424 a_46116_21352# d0 0.518f
C10425 a_2582_30882# d1 0.00148f
C10426 d3 a_38152_24076# 0.00108f
C10427 d1 a_25712_4110# 5.03e-20
C10428 X2.X2.X1.X1.X1.X2.X1.vin1 vdd 0.592f
C10429 X2.X1.X2.X2.vrefh X2.X1.X2.X1.X2.X2.X3.vin2 0.161f
C10430 d4 X2.X2.X1.X1.X1.X2.vout 1.45e-19
C10431 d3 a_8872_8828# 0.00108f
C10432 a_48616_14688# a_48316_12822# 6.71e-19
C10433 a_31862_11822# a_33976_10916# 4.72e-20
C10434 X1.X2.X2.X1.X2.vrefh d1 0.00745f
C10435 a_17222_11822# X1.X2.X1.X2.X2.X1.X1.vin1 8.22e-20
C10436 X2.X2.X2.X3.vin1 d1 0.00955f
C10437 a_48616_26164# a_48316_24258# 6.2e-19
C10438 X2.X1.X2.X2.X2.vrefh X2.X1.X2.X2.X1.X2.X3.vin1 0.00118f
C10439 a_52792_24076# d1 0.521f
C10440 a_54992_26982# a_54992_25076# 0.00396f
C10441 d1 a_8572_6962# 0.00613f
C10442 X2.X1.X2.X1.X1.X2.X3.vin1 X2.X1.X2.X1.X1.X2.X1.vin2 0.216f
C10443 a_37766_8828# a_39966_7922# 4.2e-20
C10444 X2.X2.X1.X2.X1.X1.X1.vin2 vdd 0.36f
C10445 X2.X1.X1.X1.X1.X2.X2.vin1 d0 0.262f
C10446 X2.X2.X1.X1.X2.X2.X2.vin1 d2 0.0314f
C10447 X1.X2.X1.X2.X3.vin2 X1.X2.X1.X2.X2.X2.vout 0.0866f
C10448 X2.X1.X2.X1.X1.X1.X3.vin1 a_40352_4110# 0.354f
C10449 X1.X1.X1.X1.X2.X1.X3.vin1 a_4782_24258# 0.428f
C10450 a_8486_5016# vdd 0.562f
C10451 X2.X1.X1.X2.X1.X1.X3.vin1 vdd 0.997f
C10452 d4 X1.X1.X1.X2.X1.X1.X1.vin2 3.99e-21
C10453 a_37852_25982# X2.X1.X2.X2.X1.X2.vout 7.93e-20
C10454 a_39966_9828# a_38152_8828# 1.15e-20
C10455 d3 a_23126_16452# 4.67e-19
C10456 a_48702_16634# a_48616_14688# 3.14e-19
C10457 X2.X2.X2.X2.X2.X2.X3.vin1 X2.X2.X2.X2.X2.X2.X1.vin1 0.206f
C10458 a_48316_16634# a_49002_14688# 2.86e-19
C10459 X2.X1.X3.vin2 a_37466_14586# 3.67e-19
C10460 a_25712_7922# a_25712_6016# 0.00396f
C10461 d4 X2.X2.X2.X1.X2.X2.vout 6.95e-19
C10462 X1.X1.X2.vrefh X1.X1.X2.X1.X1.X1.X1.vin2 0.096f
C10463 X2.X1.X2.X1.X1.X1.vout a_38152_5016# 0.359f
C10464 X2.X1.X1.X1.X2.X2.X2.vin1 d2 0.0314f
C10465 a_37766_16452# d1 0.0749f
C10466 X2.X2.X2.X2.X1.X2.X1.vin2 a_54992_23170# 0.12f
C10467 X2.X2.X1.X1.X1.X1.X2.vin1 a_46502_30882# 0.402f
C10468 X2.X2.X2.X2.X2.X2.vout a_52792_31700# 0.36f
C10469 a_54606_23170# X2.X2.X2.X2.X1.X2.X1.vin1 0.417f
C10470 X2.X2.X1.X1.X2.vrefh X2.X1.X2.X2.X2.vrefh 0.117f
C10471 X1.X2.X2.X1.X2.X2.X1.vin1 d1 0.0118f
C10472 d1 X2.X2.X1.X2.X2.X2.X3.vin1 0.149f
C10473 d3 a_37852_25982# 0.621f
C10474 X2.X2.X1.X2.X2.X2.vout X2.X2.X1.X2.X2.X2.X3.vin2 0.08f
C10475 X1.X1.X1.X1.X1.X2.X2.vin1 a_2196_27070# 0.197f
C10476 d1 X2.X1.X1.X2.X2.X2.vrefh 0.0124f
C10477 d3 a_23126_8828# 7.51e-19
C10478 a_17222_9916# a_17222_8010# 0.00198f
C10479 a_40352_19358# d0 0.518f
C10480 a_39966_13640# a_40352_13640# 0.419f
C10481 a_37852_10734# a_38152_8828# 6.48e-19
C10482 X2.X2.X2.X2.X1.X2.X3.vin2 d2 0.121f
C10483 X2.X2.X2.X3.vin1 X2.X2.X3.vin2 1.16f
C10484 X1.X2.X1.X1.X2.X2.X2.vin1 d2 0.0314f
C10485 X1.X1.X2.X1.X2.X2.X3.vin1 a_11072_15546# 0.354f
C10486 X2.X2.X2.X2.X1.X2.X3.vin1 vdd 0.96f
C10487 a_4696_10916# a_4396_9010# 6.2e-19
C10488 a_2196_13728# X1.X1.X1.X2.X1.X2.X2.vin1 1.78e-19
C10489 a_31862_13728# X2.X1.X1.X2.X1.X2.X1.vin1 0.417f
C10490 a_31476_13728# X2.X1.X1.X2.X1.X2.X3.vin1 0.354f
C10491 a_31476_9916# d1 2.25e-20
C10492 d1 a_17222_8010# 0.00148f
C10493 X2.X1.X1.X2.X1.X2.X2.vin1 vdd 0.576f
C10494 X2.X2.X2.X1.X1.X2.X1.vin2 vdd 0.361f
C10495 d2 a_40352_9828# 0.00533f
C10496 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.vrefh 0.161f
C10497 d2 a_23512_16452# 6.04e-19
C10498 a_40352_23170# vdd 1.05f
C10499 a_4396_16634# a_2582_15634# 1.15e-20
C10500 X1.X1.X1.X2.X1.X2.X3.vin2 a_5082_10916# 0.00846f
C10501 d3 d4 18.5f
C10502 X1.X2.X3.vin2 vdd 0.834f
C10503 a_46502_30882# a_46502_32788# 0.00198f
C10504 X2.X1.X2.X3.vin2 a_37852_25982# 0.355f
C10505 a_52106_25982# d1 0.0316f
C10506 d3 a_54606_11734# 0.00112f
C10507 a_16836_32788# d4 1.8e-19
C10508 a_46502_28976# X2.X2.X1.X1.X1.X2.X1.vin2 0.273f
C10509 a_25712_19358# d0 0.518f
C10510 d3 a_23212_22210# 7.7e-20
C10511 d5 X3.vin1 0.0663f
C10512 d2 X1.X2.X2.X1.X1.X2.X3.vin2 0.121f
C10513 X1.X2.X3.vin1 X1.X2.X2.vrefh 0.178f
C10514 X2.X2.X2.X1.X1.X2.X1.vin2 X2.X2.X2.X1.X1.X2.X1.vin1 0.668f
C10515 X2.X1.X1.X1.X2.X2.X1.vin2 d1 2.18e-19
C10516 X2.X2.X2.X1.X3.vin1 d1 0.00179f
C10517 X1.X1.X1.X2.X1.X1.X3.vin2 X1.X1.X1.X2.X1.X2.X3.vin1 1.22e-19
C10518 X2.X1.X2.X2.X2.X1.X2.vin1 X2.X1.X2.X2.X2.X1.X3.vin2 0.234f
C10519 a_10686_28888# X1.X1.X2.X2.X2.X1.X3.vin1 0.00207f
C10520 d4 X2.X2.X2.X2.X2.X2.vout 0.0955f
C10521 a_37766_31700# X2.X1.X2.X2.X2.X2.vout 0.418f
C10522 X2.X2.X1.X1.X2.X1.X3.vin1 a_46502_23258# 0.00207f
C10523 X1.X2.X1.X2.X1.X1.X1.vin1 X1.X2.X1.X2.X1.X1.X2.vin1 0.0689f
C10524 X2.X1.X1.X2.X1.X1.vout vdd 0.78f
C10525 a_37766_31700# d1 0.0489f
C10526 a_2196_9916# a_2196_8010# 0.00396f
C10527 X1.X2.X1.X1.X2.X2.X3.vin1 d1 0.146f
C10528 X1.X1.X2.X2.X1.X2.X3.vin1 a_11072_23170# 0.354f
C10529 d3 X1.X2.X1.X1.X1.X2.vout 0.125f
C10530 X2.X1.X1.X1.X2.X2.X1.vin1 d2 0.0106f
C10531 a_11072_19358# d0 0.518f
C10532 d4 X2.X2.X2.X2.X2.X1.X3.vin2 0.0533f
C10533 d0 X2.X1.X2.X1.X1.X1.X2.vin1 0.262f
C10534 a_48616_14688# d1 0.00613f
C10535 X1.X2.X2.X2.X2.X2.X1.vin1 d1 0.0118f
C10536 X1.X2.X2.X2.X2.X1.X1.vin2 X2.X1.X1.X1.X2.vrefh 0.0128f
C10537 a_4396_24258# a_2582_23258# 1.15e-20
C10538 X2.X1.X2.X1.X2.X1.X1.vin1 a_39966_9828# 8.22e-20
C10539 X2.X1.X1.X1.X2.X1.X1.vin1 d0 0.267f
C10540 X1.X1.X1.X1.X2.X1.X3.vin2 X1.X1.X1.X1.X2.X2.vrefh 0.161f
C10541 X2.X1.X2.X3.vin2 d4 0.535f
C10542 X2.X1.X2.X1.X2.X1.X1.vin2 X2.X1.X2.X1.X1.X2.X3.vin2 3.94e-19
C10543 a_10686_26982# a_8486_27888# 4.2e-20
C10544 X1.X2.X2.X1.X1.X1.vout X1.X2.X2.X1.X1.X1.X3.vin2 0.342f
C10545 d1 X2.X2.X1.X2.X2.X2.X3.vin2 0.214f
C10546 X1.X1.X2.X2.X2.X1.X1.vin2 X1.X1.X2.X2.X2.X1.X3.vin1 0.216f
C10547 X1.X1.X2.X2.X2.X2.X2.vin1 a_8486_31700# 0.00351f
C10548 a_10686_32700# X1.X1.X2.X2.X2.X2.X3.vin1 0.00207f
C10549 a_52792_5016# a_54606_4110# 1.06e-19
C10550 X1.X2.X1.X3.vin1 d2 6.42e-19
C10551 X2.X1.X3.vin2 X2.X1.X2.X1.X1.X2.X3.vin1 0.00836f
C10552 a_19422_12822# X1.X2.X1.X2.X1.X2.X3.vin2 0.277f
C10553 X2.X1.X2.X1.X2.X2.X3.vin2 a_37466_14586# 3.85e-19
C10554 a_4396_20446# vdd 1.05f
C10555 X2.X1.X1.X2.X1.X1.X3.vin1 X2.X1.X1.X2.X1.X1.X1.vin2 0.216f
C10556 a_17222_25164# a_19036_24258# 1.06e-19
C10557 a_46116_23258# a_46116_21352# 0.00396f
C10558 X1.X2.X1.X1.X2.X1.X1.vin1 X1.X2.X1.X1.X2.X1.X2.vin1 0.0689f
C10559 X2.X1.X2.X1.X2.X2.vrefh a_39966_13640# 0.3f
C10560 d2 a_23512_31700# 0.00293f
C10561 X2.X2.X2.X3.vin2 a_52106_18358# 0.263f
C10562 X2.X1.X2.X1.X1.X2.X1.vin2 X2.X2.X1.X2.X2.X1.X2.vin1 0.00232f
C10563 X1.X1.X1.X2.X1.X2.vrefh vdd 0.414f
C10564 d0 X1.X1.X1.X2.X2.X1.X1.vin1 0.267f
C10565 X2.X1.X2.X2.X2.X1.X1.vin2 vdd 0.36f
C10566 X2.X1.X1.X2.X3.vin2 a_34062_5198# 9.7e-20
C10567 X2.X2.X3.vin2 X2.X2.X2.X1.X3.vin1 0.0361f
C10568 d3 a_4396_24258# 0.00178f
C10569 X2.X2.X2.X2.X1.X2.X1.vin2 d1 0.00406f
C10570 d1 X2.X1.X1.X2.X2.X2.vout 0.0331f
C10571 X2.X2.X2.X3.vin1 a_52492_10734# 0.356f
C10572 X1.X2.X1.X2.X1.X2.X1.vin2 vdd 0.361f
C10573 d2 a_52792_12640# 3.82e-19
C10574 X1.X2.X2.X2.X1.X1.vout d4 0.00164f
C10575 X2.X2.X1.X1.X2.X2.X3.vin2 X2.X2.X1.X2.X1.X1.X1.vin1 5.19e-19
C10576 a_5082_22312# d2 0.0191f
C10577 X1.X1.X1.X3.vin1 X1.X1.X1.X1.X2.X2.vout 0.2f
C10578 X1.X2.X2.X2.X1.X1.vout a_23212_22210# 0.169f
C10579 X1.X1.X1.X2.X1.X2.X3.vin1 vdd 0.96f
C10580 a_31476_28976# vdd 1.05f
C10581 a_52492_22210# a_52792_20264# 6.1e-19
C10582 X1.X1.X2.X2.X1.X1.X2.vin1 d0 0.262f
C10583 a_31476_4198# a_31862_4198# 0.419f
C10584 a_48616_29936# X2.X2.X1.X1.X3.vin1 0.363f
C10585 X2.X1.X1.X1.X1.X1.vout vdd 0.781f
C10586 X1.X2.X1.X1.X2.X1.X3.vin2 X1.X2.X1.X1.X2.X2.X1.vin2 3.94e-19
C10587 X2.X1.X2.X1.X1.X1.X3.vin2 a_40352_6016# 0.354f
C10588 d3 a_54606_9828# 1.89e-19
C10589 X2.X1.X2.vrefh a_31862_4198# 0.301f
C10590 X2.X1.X1.X1.X2.X1.X3.vin1 X2.X1.X1.X1.X2.X1.X1.vin2 0.216f
C10591 a_38152_5016# a_39966_4110# 1.06e-19
C10592 X2.X2.X2.X1.X2.X2.vout a_52492_14586# 0.0929f
C10593 d2 d0 0.0111f
C10594 d0 a_54606_32700# 0.0489f
C10595 X1.X1.X1.X1.X2.X1.X1.vin2 X1.X1.X1.X1.X2.X1.X2.vin1 0.242f
C10596 a_46502_27070# X2.X2.X1.X1.X2.X1.X1.vin1 8.22e-20
C10597 d3 a_37766_8828# 7.51e-19
C10598 X1.X1.X2.X1.X1.X1.vout a_8486_5016# 0.422f
C10599 d4 X1.X2.X1.X1.X3.vin1 0.00246f
C10600 X2.X1.X1.X2.X2.X2.X1.vin1 X2.X1.X1.X2.X2.X2.X3.vin1 0.206f
C10601 X2.X2.X2.X2.X2.X1.X3.vin1 X2.X2.X2.X2.X1.X2.X3.vin2 1.22e-19
C10602 a_19422_28070# X1.X2.X1.X1.X1.X2.vout 0.418f
C10603 X2.X2.X2.X1.X3.vin1 X2.X2.X2.X1.X1.X2.vout 0.398f
C10604 X2.X2.X2.X2.X3.vin2 vdd 1.29f
C10605 X2.X2.X2.X2.X2.X1.X1.vin2 a_54606_26982# 0.273f
C10606 a_37466_14586# a_37766_12640# 4.19e-20
C10607 X2.X2.X1.X1.X2.X1.vout a_49002_22312# 0.383f
C10608 X2.X1.X1.X1.X2.X1.X3.vin2 a_31862_21352# 8.07e-19
C10609 d1 a_52406_8828# 0.0749f
C10610 X1.X1.X2.X2.X2.X2.X3.vin1 a_11072_30794# 0.354f
C10611 a_37852_6962# a_37766_5016# 3.14e-19
C10612 a_19036_12822# d1 0.521f
C10613 X1.X1.X1.X1.X1.X1.X1.vin1 X1.X1.X1.X1.X1.X1.X1.vin2 0.696f
C10614 a_49566_892# a_49952_892# 0.406f
C10615 X1.X1.X2.X1.X2.X1.X3.vin1 X1.X1.X2.X1.X1.X2.X3.vin2 1.22e-19
C10616 a_11072_26982# vdd 1.05f
C10617 X1.X1.X1.X2.X2.vrefh X1.X1.X1.X2.X2.X1.X3.vin1 2.33e-19
C10618 a_4396_20446# X1.X1.X1.X1.X2.X2.X3.vin2 0.101f
C10619 d1 X2.X1.X2.X1.X1.X2.X1.vin1 0.0118f
C10620 X1.X2.X1.X1.X3.vin1 X1.X2.X1.X1.X1.X2.vout 0.398f
C10621 a_17222_17540# d0 0.0675f
C10622 X1.X1.X1.X2.X2.X2.X2.vin1 a_2582_4198# 0.402f
C10623 a_10686_13640# X1.X1.X2.X1.X2.X1.X1.vin2 8.88e-20
C10624 a_4396_31882# a_2582_30882# 1.15e-20
C10625 X2.X2.X2.X2.X2.X1.X3.vin2 X2.X2.X2.X2.X2.X2.X1.vin2 3.94e-19
C10626 d2 X1.X2.X1.X2.X2.vrefh 0.158f
C10627 a_54606_28888# X2.X2.X2.X2.X2.X2.X1.vin1 8.22e-20
C10628 a_19422_24258# a_19336_22312# 3.14e-19
C10629 a_19036_24258# a_19722_22312# 2.86e-19
C10630 X1.X1.X1.X1.X1.X1.X3.vin2 X1.X1.X1.X1.X1.X2.vrefh 0.165f
C10631 a_49952_892# vss 0.973f
C10632 a_49566_892# vss 1.67f
C10633 X2.X3.vin2 vss 3.86f
C10634 a_43362_892# vss 0.997f
C10635 a_42976_892# vss 1.67f
C10636 X2.X3.vin1 vss 2.94f
C10637 a_35312_892# vss 1.01f
C10638 a_34926_892# vss 1.67f
C10639 X3.vin2 vss 6.29f
C10640 vout vss 0.355f
C10641 a_28482_892# vss 1.03f
C10642 a_28096_892# vss 1.67f
C10643 d7 vss 0.864f
C10644 a_20672_892# vss 0.97f
C10645 a_20286_892# vss 1.67f
C10646 X1.X3.vin2 vss 3.74f
C10647 X3.vin1 vss 5.65f
C10648 a_14082_892# vss 0.996f
C10649 a_13696_892# vss 1.67f
C10650 d6 vss 15.3f
C10651 X1.X3.vin1 vss 2.98f
C10652 a_6032_892# vss 1.01f
C10653 a_5646_892# vss 1.67f
C10654 d5 vss 11.4f
C10655 a_54992_4110# vss 1.66f
C10656 X2.X2.X2.X1.X1.X1.X1.vin1 vss 2.17f
C10657 a_54606_4110# vss 0.858f
C10658 X2.X2.X2.X1.X1.X1.X1.vin2 vss 2.21f
C10659 a_46502_4198# vss 0.888f
C10660 a_46116_4198# vss 1.67f
C10661 X2.X2.X2.vrefh vss 12.4f
C10662 a_52792_5016# vss 1.67f
C10663 X2.X2.X2.X1.X1.X1.X3.vin1 vss 0.982f
C10664 a_52406_5016# vss 0.854f
C10665 X2.X2.X1.X2.X2.X2.X3.vin2 vss 1.69f
C10666 a_48702_5198# vss 0.947f
C10667 a_48316_5198# vss 1.67f
C10668 X2.X2.X1.X2.X2.X2.X2.vin1 vss 1.8f
C10669 a_40352_4110# vss 1.66f
C10670 X2.X1.X2.X1.X1.X1.X1.vin1 vss 2.16f
C10671 a_39966_4110# vss 0.858f
C10672 X2.X1.X2.X1.X1.X1.X1.vin2 vss 2.19f
C10673 a_31862_4198# vss 0.888f
C10674 a_31476_4198# vss 1.67f
C10675 X2.X1.X2.vrefh vss 12.3f
C10676 a_38152_5016# vss 1.67f
C10677 X2.X1.X2.X1.X1.X1.X3.vin1 vss 0.982f
C10678 a_37766_5016# vss 0.854f
C10679 X2.X1.X1.X2.X2.X2.X3.vin2 vss 1.69f
C10680 a_34062_5198# vss 0.947f
C10681 a_33676_5198# vss 1.67f
C10682 X2.X1.X1.X2.X2.X2.X2.vin1 vss 1.8f
C10683 a_25712_4110# vss 1.66f
C10684 X1.X2.X2.X1.X1.X1.X1.vin1 vss 2.16f
C10685 a_25326_4110# vss 0.858f
C10686 X1.X2.X2.X1.X1.X1.X1.vin2 vss 2.19f
C10687 a_17222_4198# vss 0.888f
C10688 a_16836_4198# vss 1.67f
C10689 X1.X2.X2.vrefh vss 12.3f
C10690 a_23512_5016# vss 1.67f
C10691 X1.X2.X2.X1.X1.X1.X3.vin1 vss 0.982f
C10692 a_23126_5016# vss 0.854f
C10693 X1.X2.X1.X2.X2.X2.X3.vin2 vss 1.69f
C10694 a_19422_5198# vss 0.947f
C10695 a_19036_5198# vss 1.67f
C10696 X1.X2.X1.X2.X2.X2.X2.vin1 vss 1.8f
C10697 a_11072_4110# vss 1.66f
C10698 X1.X1.X2.X1.X1.X1.X1.vin1 vss 2.16f
C10699 a_10686_4110# vss 0.858f
C10700 X1.X1.X2.X1.X1.X1.X1.vin2 vss 2.19f
C10701 a_2582_4198# vss 0.888f
C10702 a_2196_4198# vss 1.67f
C10703 X1.X1.X2.vrefh vss 12.5f
C10704 a_8872_5016# vss 1.67f
C10705 X1.X1.X2.X1.X1.X1.X3.vin1 vss 0.982f
C10706 a_8486_5016# vss 0.854f
C10707 X1.X1.X1.X2.X2.X2.X3.vin2 vss 1.69f
C10708 a_4782_5198# vss 0.947f
C10709 a_4396_5198# vss 1.67f
C10710 X1.X1.X1.X2.X2.X2.X2.vin1 vss 1.8f
C10711 a_54992_6016# vss 1.66f
C10712 X2.X2.X2.X1.X1.X1.X3.vin2 vss 1.34f
C10713 X2.X2.X2.X1.X1.X1.X2.vin1 vss 1.8f
C10714 a_54606_6016# vss 0.883f
C10715 X2.X2.X1.X2.X2.X2.X1.vin2 vss 2.19f
C10716 X2.X2.X1.X2.X2.X2.X3.vin1 vss 0.896f
C10717 X2.X2.X1.X2.X2.X2.X1.vin1 vss 2.05f
C10718 a_46502_6104# vss 0.856f
C10719 a_46116_6104# vss 1.66f
C10720 a_40352_6016# vss 1.66f
C10721 X2.X1.X2.X1.X1.X1.X3.vin2 vss 1.34f
C10722 X2.X1.X2.X1.X1.X1.X2.vin1 vss 1.8f
C10723 a_39966_6016# vss 0.883f
C10724 X2.X1.X1.X2.X2.X2.X1.vin2 vss 2.19f
C10725 X2.X1.X1.X2.X2.X2.X3.vin1 vss 0.896f
C10726 X2.X1.X1.X2.X2.X2.X1.vin1 vss 2.05f
C10727 a_31862_6104# vss 0.856f
C10728 a_31476_6104# vss 1.66f
C10729 a_25712_6016# vss 1.66f
C10730 X1.X2.X2.X1.X1.X1.X3.vin2 vss 1.34f
C10731 X1.X2.X2.X1.X1.X1.X2.vin1 vss 1.8f
C10732 a_25326_6016# vss 0.883f
C10733 X1.X2.X1.X2.X2.X2.X1.vin2 vss 2.19f
C10734 X1.X2.X1.X2.X2.X2.X3.vin1 vss 0.896f
C10735 X1.X2.X1.X2.X2.X2.X1.vin1 vss 2.05f
C10736 a_17222_6104# vss 0.856f
C10737 a_16836_6104# vss 1.66f
C10738 a_11072_6016# vss 1.66f
C10739 X1.X1.X2.X1.X1.X1.X3.vin2 vss 1.34f
C10740 X1.X1.X2.X1.X1.X1.X2.vin1 vss 1.8f
C10741 a_10686_6016# vss 0.883f
C10742 X1.X1.X1.X2.X2.X2.X1.vin2 vss 2.21f
C10743 X1.X1.X1.X2.X2.X2.X3.vin1 vss 0.896f
C10744 X1.X1.X1.X2.X2.X2.X1.vin1 vss 2.05f
C10745 a_2582_6104# vss 0.856f
C10746 a_2196_6104# vss 1.66f
C10747 a_52492_6962# vss 1.66f
C10748 X2.X2.X2.X1.X1.X1.vout vss 0.861f
C10749 a_52106_6962# vss 0.96f
C10750 X2.X2.X1.X2.X2.X2.vout vss 1.18f
C10751 a_49002_7064# vss 0.962f
C10752 a_48616_7064# vss 1.66f
C10753 a_37852_6962# vss 1.66f
C10754 X2.X1.X2.X1.X1.X1.vout vss 0.861f
C10755 a_37466_6962# vss 0.96f
C10756 X2.X1.X1.X2.X2.X2.vout vss 1.18f
C10757 a_34362_7064# vss 0.962f
C10758 a_33976_7064# vss 1.66f
C10759 a_23212_6962# vss 1.66f
C10760 X1.X2.X2.X1.X1.X1.vout vss 0.861f
C10761 a_22826_6962# vss 0.96f
C10762 X1.X2.X1.X2.X2.X2.vout vss 1.18f
C10763 a_19722_7064# vss 0.962f
C10764 a_19336_7064# vss 1.66f
C10765 a_8572_6962# vss 1.66f
C10766 X1.X1.X2.X1.X1.X1.vout vss 0.861f
C10767 a_8186_6962# vss 0.96f
C10768 X1.X1.X1.X2.X2.X2.vout vss 1.18f
C10769 a_5082_7064# vss 0.962f
C10770 a_4696_7064# vss 1.66f
C10771 X2.X2.X2.X1.X1.X2.vrefh vss 4.22f
C10772 a_54992_7922# vss 1.66f
C10773 X2.X2.X2.X1.X1.X2.X1.vin1 vss 2.05f
C10774 a_54606_7922# vss 0.856f
C10775 X2.X2.X2.X1.X1.X2.X1.vin2 vss 2.19f
C10776 a_46502_8010# vss 0.883f
C10777 a_46116_8010# vss 1.66f
C10778 X2.X1.X2.X1.X1.X2.vrefh vss 4.07f
C10779 X2.X2.X1.X2.X2.X2.vrefh vss 4.05f
C10780 a_52792_8828# vss 1.67f
C10781 X2.X2.X2.X1.X1.X2.vout vss 1.11f
C10782 X2.X2.X2.X1.X1.X2.X3.vin1 vss 0.892f
C10783 a_52406_8828# vss 0.945f
C10784 X2.X2.X1.X2.X2.X1.X3.vin2 vss 1.32f
C10785 X2.X2.X1.X2.X2.X1.vout vss 0.816f
C10786 a_48702_9010# vss 0.854f
C10787 a_48316_9010# vss 1.67f
C10788 X2.X2.X1.X2.X2.X1.X2.vin1 vss 1.79f
C10789 a_40352_7922# vss 1.66f
C10790 X2.X1.X2.X1.X1.X2.X1.vin1 vss 2.05f
C10791 a_39966_7922# vss 0.856f
C10792 X2.X1.X2.X1.X1.X2.X1.vin2 vss 2.17f
C10793 a_31862_8010# vss 0.883f
C10794 a_31476_8010# vss 1.66f
C10795 X1.X2.X2.X1.X1.X2.vrefh vss 4.07f
C10796 X2.X1.X1.X2.X2.X2.vrefh vss 4.05f
C10797 a_38152_8828# vss 1.67f
C10798 X2.X1.X2.X1.X1.X2.vout vss 1.11f
C10799 X2.X1.X2.X1.X1.X2.X3.vin1 vss 0.892f
C10800 a_37766_8828# vss 0.945f
C10801 X2.X1.X1.X2.X2.X1.X3.vin2 vss 1.32f
C10802 X2.X1.X1.X2.X2.X1.vout vss 0.816f
C10803 a_34062_9010# vss 0.854f
C10804 a_33676_9010# vss 1.67f
C10805 X2.X1.X1.X2.X2.X1.X2.vin1 vss 1.79f
C10806 a_25712_7922# vss 1.66f
C10807 X1.X2.X2.X1.X1.X2.X1.vin1 vss 2.05f
C10808 a_25326_7922# vss 0.856f
C10809 X1.X2.X2.X1.X1.X2.X1.vin2 vss 2.17f
C10810 a_17222_8010# vss 0.883f
C10811 a_16836_8010# vss 1.66f
C10812 X1.X1.X2.X1.X1.X2.vrefh vss 4.07f
C10813 X1.X2.X1.X2.X2.X2.vrefh vss 4.05f
C10814 a_23512_8828# vss 1.67f
C10815 X1.X2.X2.X1.X1.X2.vout vss 1.11f
C10816 X1.X2.X2.X1.X1.X2.X3.vin1 vss 0.892f
C10817 a_23126_8828# vss 0.945f
C10818 X1.X2.X1.X2.X2.X1.X3.vin2 vss 1.32f
C10819 X1.X2.X1.X2.X2.X1.vout vss 0.816f
C10820 a_19422_9010# vss 0.854f
C10821 a_19036_9010# vss 1.67f
C10822 X1.X2.X1.X2.X2.X1.X2.vin1 vss 1.79f
C10823 a_11072_7922# vss 1.66f
C10824 X1.X1.X2.X1.X1.X2.X1.vin1 vss 2.05f
C10825 a_10686_7922# vss 0.856f
C10826 X1.X1.X2.X1.X1.X2.X1.vin2 vss 2.17f
C10827 a_2582_8010# vss 0.883f
C10828 a_2196_8010# vss 1.66f
C10829 X1.X1.X1.X2.X2.X2.vrefh vss 4.21f
C10830 a_8872_8828# vss 1.67f
C10831 X1.X1.X2.X1.X1.X2.vout vss 1.11f
C10832 X1.X1.X2.X1.X1.X2.X3.vin1 vss 0.892f
C10833 a_8486_8828# vss 0.945f
C10834 X1.X1.X1.X2.X2.X1.X3.vin2 vss 1.32f
C10835 X1.X1.X1.X2.X2.X1.vout vss 0.816f
C10836 a_4782_9010# vss 0.854f
C10837 a_4396_9010# vss 1.67f
C10838 X1.X1.X1.X2.X2.X1.X2.vin1 vss 1.8f
C10839 a_54992_9828# vss 1.66f
C10840 X2.X2.X2.X1.X1.X2.X3.vin2 vss 1.55f
C10841 X2.X2.X2.X1.X1.X2.X2.vin1 vss 1.8f
C10842 a_54606_9828# vss 0.884f
C10843 X2.X2.X1.X2.X2.X1.X1.vin2 vss 2.17f
C10844 X2.X2.X1.X2.X2.X1.X3.vin1 vss 0.91f
C10845 X2.X2.X1.X2.X2.X1.X1.vin1 vss 2.05f
C10846 a_46502_9916# vss 0.855f
C10847 a_46116_9916# vss 1.66f
C10848 a_40352_9828# vss 1.66f
C10849 X2.X1.X2.X1.X1.X2.X3.vin2 vss 1.55f
C10850 X2.X1.X2.X1.X1.X2.X2.vin1 vss 1.79f
C10851 a_39966_9828# vss 0.884f
C10852 X2.X1.X1.X2.X2.X1.X1.vin2 vss 2.17f
C10853 X2.X1.X1.X2.X2.X1.X3.vin1 vss 0.91f
C10854 X2.X1.X1.X2.X2.X1.X1.vin1 vss 2.05f
C10855 a_31862_9916# vss 0.855f
C10856 a_31476_9916# vss 1.66f
C10857 a_25712_9828# vss 1.66f
C10858 X1.X2.X2.X1.X1.X2.X3.vin2 vss 1.55f
C10859 X1.X2.X2.X1.X1.X2.X2.vin1 vss 1.79f
C10860 a_25326_9828# vss 0.884f
C10861 X1.X2.X1.X2.X2.X1.X1.vin2 vss 2.17f
C10862 X1.X2.X1.X2.X2.X1.X3.vin1 vss 0.91f
C10863 X1.X2.X1.X2.X2.X1.X1.vin1 vss 2.05f
C10864 a_17222_9916# vss 0.855f
C10865 a_16836_9916# vss 1.66f
C10866 a_11072_9828# vss 1.66f
C10867 X1.X1.X2.X1.X1.X2.X3.vin2 vss 1.55f
C10868 X1.X1.X2.X1.X1.X2.X2.vin1 vss 1.79f
C10869 a_10686_9828# vss 0.884f
C10870 X1.X1.X1.X2.X2.X1.X1.vin2 vss 2.18f
C10871 X1.X1.X1.X2.X2.X1.X3.vin1 vss 0.91f
C10872 X1.X1.X1.X2.X2.X1.X1.vin1 vss 2.05f
C10873 a_2582_9916# vss 0.855f
C10874 a_2196_9916# vss 1.66f
C10875 a_52492_10734# vss 1.67f
C10876 X2.X2.X2.X1.X3.vin1 vss 2.32f
C10877 a_52106_10734# vss 0.926f
C10878 X2.X2.X1.X2.X3.vin2 vss 1.96f
C10879 a_49002_10916# vss 0.93f
C10880 a_48616_10916# vss 1.67f
C10881 a_37852_10734# vss 1.67f
C10882 X2.X1.X2.X1.X3.vin1 vss 2.32f
C10883 a_37466_10734# vss 0.926f
C10884 X2.X1.X1.X2.X3.vin2 vss 1.96f
C10885 a_34362_10916# vss 0.93f
C10886 a_33976_10916# vss 1.67f
C10887 a_23212_10734# vss 1.67f
C10888 X1.X2.X2.X1.X3.vin1 vss 2.32f
C10889 a_22826_10734# vss 0.926f
C10890 X1.X2.X1.X2.X3.vin2 vss 1.96f
C10891 a_19722_10916# vss 0.93f
C10892 a_19336_10916# vss 1.67f
C10893 a_8572_10734# vss 1.67f
C10894 X1.X1.X2.X1.X3.vin1 vss 2.32f
C10895 a_8186_10734# vss 0.926f
C10896 X1.X1.X1.X2.X3.vin2 vss 1.96f
C10897 a_5082_10916# vss 0.93f
C10898 a_4696_10916# vss 1.67f
C10899 X2.X2.X2.X1.X2.vrefh vss 4.21f
C10900 a_54992_11734# vss 1.66f
C10901 X2.X2.X2.X1.X2.X1.X1.vin1 vss 2.05f
C10902 a_54606_11734# vss 0.855f
C10903 X2.X2.X2.X1.X2.X1.X1.vin2 vss 2.18f
C10904 a_46502_11822# vss 0.884f
C10905 a_46116_11822# vss 1.66f
C10906 X2.X1.X2.X1.X2.vrefh vss 4.06f
C10907 X2.X2.X1.X2.X2.vrefh vss 4.06f
C10908 a_52792_12640# vss 1.67f
C10909 X2.X2.X2.X1.X2.X1.X3.vin1 vss 0.905f
C10910 a_52406_12640# vss 0.854f
C10911 X2.X2.X1.X2.X1.X2.X3.vin2 vss 1.5f
C10912 a_48702_12822# vss 0.945f
C10913 a_48316_12822# vss 1.67f
C10914 X2.X2.X1.X2.X1.X2.X2.vin1 vss 1.79f
C10915 a_40352_11734# vss 1.66f
C10916 X2.X1.X2.X1.X2.X1.X1.vin1 vss 2.05f
C10917 a_39966_11734# vss 0.855f
C10918 X2.X1.X2.X1.X2.X1.X1.vin2 vss 2.17f
C10919 a_31862_11822# vss 0.884f
C10920 a_31476_11822# vss 1.66f
C10921 X1.X2.X2.X1.X2.vrefh vss 4.06f
C10922 X2.X1.X1.X2.X2.vrefh vss 4.06f
C10923 a_38152_12640# vss 1.67f
C10924 X2.X1.X2.X1.X2.X1.X3.vin1 vss 0.905f
C10925 a_37766_12640# vss 0.854f
C10926 X2.X1.X1.X2.X1.X2.X3.vin2 vss 1.5f
C10927 a_34062_12822# vss 0.945f
C10928 a_33676_12822# vss 1.67f
C10929 X2.X1.X1.X2.X1.X2.X2.vin1 vss 1.79f
C10930 a_25712_11734# vss 1.66f
C10931 X1.X2.X2.X1.X2.X1.X1.vin1 vss 2.05f
C10932 a_25326_11734# vss 0.855f
C10933 X1.X2.X2.X1.X2.X1.X1.vin2 vss 2.17f
C10934 a_17222_11822# vss 0.884f
C10935 a_16836_11822# vss 1.66f
C10936 X1.X1.X2.X1.X2.vrefh vss 4.06f
C10937 X1.X2.X1.X2.X2.vrefh vss 4.06f
C10938 a_23512_12640# vss 1.67f
C10939 X1.X2.X2.X1.X2.X1.X3.vin1 vss 0.905f
C10940 a_23126_12640# vss 0.854f
C10941 X1.X2.X1.X2.X1.X2.X3.vin2 vss 1.5f
C10942 a_19422_12822# vss 0.945f
C10943 a_19036_12822# vss 1.67f
C10944 X1.X2.X1.X2.X1.X2.X2.vin1 vss 1.79f
C10945 a_11072_11734# vss 1.66f
C10946 X1.X1.X2.X1.X2.X1.X1.vin1 vss 2.05f
C10947 a_10686_11734# vss 0.855f
C10948 X1.X1.X2.X1.X2.X1.X1.vin2 vss 2.17f
C10949 a_2582_11822# vss 0.884f
C10950 a_2196_11822# vss 1.66f
C10951 X1.X1.X1.X2.X2.vrefh vss 4.21f
C10952 a_8872_12640# vss 1.67f
C10953 X1.X1.X2.X1.X2.X1.X3.vin1 vss 0.905f
C10954 a_8486_12640# vss 0.854f
C10955 X1.X1.X1.X2.X1.X2.X3.vin2 vss 1.5f
C10956 a_4782_12822# vss 0.945f
C10957 a_4396_12822# vss 1.67f
C10958 X1.X1.X1.X2.X1.X2.X2.vin1 vss 1.8f
C10959 a_54992_13640# vss 1.66f
C10960 X2.X2.X2.X1.X2.X1.X3.vin2 vss 1.28f
C10961 X2.X2.X2.X1.X2.X1.X2.vin1 vss 1.8f
C10962 a_54606_13640# vss 0.883f
C10963 X2.X2.X1.X2.X1.X2.X1.vin2 vss 2.17f
C10964 X2.X2.X1.X2.X1.X2.X3.vin1 vss 0.887f
C10965 X2.X2.X1.X2.X1.X2.X1.vin1 vss 2.05f
C10966 a_46502_13728# vss 0.856f
C10967 a_46116_13728# vss 1.66f
C10968 a_40352_13640# vss 1.66f
C10969 X2.X1.X2.X1.X2.X1.X3.vin2 vss 1.28f
C10970 X2.X1.X2.X1.X2.X1.X2.vin1 vss 1.79f
C10971 a_39966_13640# vss 0.883f
C10972 X2.X1.X1.X2.X1.X2.X1.vin2 vss 2.17f
C10973 X2.X1.X1.X2.X1.X2.X3.vin1 vss 0.887f
C10974 X2.X1.X1.X2.X1.X2.X1.vin1 vss 2.05f
C10975 a_31862_13728# vss 0.856f
C10976 a_31476_13728# vss 1.66f
C10977 a_25712_13640# vss 1.66f
C10978 X1.X2.X2.X1.X2.X1.X3.vin2 vss 1.28f
C10979 X1.X2.X2.X1.X2.X1.X2.vin1 vss 1.79f
C10980 a_25326_13640# vss 0.883f
C10981 X1.X2.X1.X2.X1.X2.X1.vin2 vss 2.17f
C10982 X1.X2.X1.X2.X1.X2.X3.vin1 vss 0.887f
C10983 X1.X2.X1.X2.X1.X2.X1.vin1 vss 2.05f
C10984 a_17222_13728# vss 0.856f
C10985 a_16836_13728# vss 1.66f
C10986 a_11072_13640# vss 1.66f
C10987 X1.X1.X2.X1.X2.X1.X3.vin2 vss 1.28f
C10988 X1.X1.X2.X1.X2.X1.X2.vin1 vss 1.79f
C10989 a_10686_13640# vss 0.883f
C10990 X1.X1.X1.X2.X1.X2.X1.vin2 vss 2.19f
C10991 X1.X1.X1.X2.X1.X2.X3.vin1 vss 0.887f
C10992 X1.X1.X1.X2.X1.X2.X1.vin1 vss 2.05f
C10993 a_2582_13728# vss 0.856f
C10994 a_2196_13728# vss 1.66f
C10995 a_52492_14586# vss 1.66f
C10996 X2.X2.X2.X1.X3.vin2 vss 1.74f
C10997 X2.X2.X2.X1.X2.X1.vout vss 0.788f
C10998 a_52106_14586# vss 0.876f
C10999 X2.X2.X1.X2.X1.X2.vout vss 1.04f
C11000 X2.X2.X1.X2.X3.vin1 vss 2.11f
C11001 a_49002_14688# vss 0.909f
C11002 a_48616_14688# vss 1.66f
C11003 a_37852_14586# vss 1.66f
C11004 X2.X1.X2.X1.X3.vin2 vss 1.74f
C11005 X2.X1.X2.X1.X2.X1.vout vss 0.788f
C11006 a_37466_14586# vss 0.876f
C11007 X2.X1.X1.X2.X1.X2.vout vss 1.04f
C11008 X2.X1.X1.X2.X3.vin1 vss 2.11f
C11009 a_34362_14688# vss 0.909f
C11010 a_33976_14688# vss 1.66f
C11011 a_23212_14586# vss 1.66f
C11012 X1.X2.X2.X1.X3.vin2 vss 1.74f
C11013 X1.X2.X2.X1.X2.X1.vout vss 0.788f
C11014 a_22826_14586# vss 0.876f
C11015 X1.X2.X1.X2.X1.X2.vout vss 1.04f
C11016 X1.X2.X1.X2.X3.vin1 vss 2.11f
C11017 a_19722_14688# vss 0.909f
C11018 a_19336_14688# vss 1.66f
C11019 a_8572_14586# vss 1.66f
C11020 X1.X1.X2.X1.X3.vin2 vss 1.74f
C11021 X1.X1.X2.X1.X2.X1.vout vss 0.788f
C11022 a_8186_14586# vss 0.876f
C11023 X1.X1.X1.X2.X1.X2.vout vss 1.04f
C11024 X1.X1.X1.X2.X3.vin1 vss 2.11f
C11025 a_5082_14688# vss 0.909f
C11026 a_4696_14688# vss 1.66f
C11027 X2.X2.X2.X1.X2.X2.vrefh vss 4.21f
C11028 a_54992_15546# vss 1.66f
C11029 X2.X2.X2.X1.X2.X2.X1.vin1 vss 2.05f
C11030 a_54606_15546# vss 0.856f
C11031 X2.X2.X2.X1.X2.X2.X1.vin2 vss 2.18f
C11032 a_46502_15634# vss 0.883f
C11033 a_46116_15634# vss 1.66f
C11034 X2.X1.X2.X1.X2.X2.vrefh vss 4.05f
C11035 X2.X2.X1.X2.X1.X2.vrefh vss 4.05f
C11036 a_52792_16452# vss 1.67f
C11037 X2.X2.X2.X1.X2.X2.vout vss 1.04f
C11038 X2.X2.X2.X1.X2.X2.X3.vin1 vss 0.888f
C11039 a_52406_16452# vss 0.945f
C11040 X2.X2.X1.X2.X1.X1.X3.vin2 vss 1.3f
C11041 X2.X2.X1.X2.X1.X1.vout vss 0.842f
C11042 a_48702_16634# vss 0.854f
C11043 a_48316_16634# vss 1.67f
C11044 X2.X2.X1.X2.X1.X1.X2.vin1 vss 1.79f
C11045 a_40352_15546# vss 1.66f
C11046 X2.X1.X2.X1.X2.X2.X1.vin1 vss 2.05f
C11047 a_39966_15546# vss 0.856f
C11048 X2.X1.X2.X1.X2.X2.X1.vin2 vss 2.17f
C11049 a_31862_15634# vss 0.883f
C11050 a_31476_15634# vss 1.66f
C11051 X1.X2.X2.X1.X2.X2.vrefh vss 4.05f
C11052 X2.X1.X1.X2.X1.X2.vrefh vss 4.05f
C11053 a_38152_16452# vss 1.67f
C11054 X2.X1.X2.X1.X2.X2.vout vss 1.04f
C11055 X2.X1.X2.X1.X2.X2.X3.vin1 vss 0.888f
C11056 a_37766_16452# vss 0.945f
C11057 X2.X1.X1.X2.X1.X1.X3.vin2 vss 1.3f
C11058 X2.X1.X1.X2.X1.X1.vout vss 0.842f
C11059 a_34062_16634# vss 0.854f
C11060 a_33676_16634# vss 1.67f
C11061 X2.X1.X1.X2.X1.X1.X2.vin1 vss 1.79f
C11062 a_25712_15546# vss 1.66f
C11063 X1.X2.X2.X1.X2.X2.X1.vin1 vss 2.05f
C11064 a_25326_15546# vss 0.856f
C11065 X1.X2.X2.X1.X2.X2.X1.vin2 vss 2.17f
C11066 a_17222_15634# vss 0.883f
C11067 a_16836_15634# vss 1.66f
C11068 X1.X1.X2.X1.X2.X2.vrefh vss 4.05f
C11069 X1.X2.X1.X2.X1.X2.vrefh vss 4.05f
C11070 a_23512_16452# vss 1.67f
C11071 X1.X2.X2.X1.X2.X2.vout vss 1.04f
C11072 X1.X2.X2.X1.X2.X2.X3.vin1 vss 0.888f
C11073 a_23126_16452# vss 0.945f
C11074 X1.X2.X1.X2.X1.X1.X3.vin2 vss 1.3f
C11075 X1.X2.X1.X2.X1.X1.vout vss 0.842f
C11076 a_19422_16634# vss 0.854f
C11077 a_19036_16634# vss 1.67f
C11078 X1.X2.X1.X2.X1.X1.X2.vin1 vss 1.79f
C11079 a_11072_15546# vss 1.66f
C11080 X1.X1.X2.X1.X2.X2.X1.vin1 vss 2.05f
C11081 a_10686_15546# vss 0.856f
C11082 X1.X1.X2.X1.X2.X2.X1.vin2 vss 2.17f
C11083 a_2582_15634# vss 0.883f
C11084 a_2196_15634# vss 1.66f
C11085 X1.X1.X1.X2.X1.X2.vrefh vss 4.21f
C11086 a_8872_16452# vss 1.67f
C11087 X1.X1.X2.X1.X2.X2.vout vss 1.04f
C11088 X1.X1.X2.X1.X2.X2.X3.vin1 vss 0.888f
C11089 a_8486_16452# vss 0.945f
C11090 X1.X1.X1.X2.X1.X1.X3.vin2 vss 1.3f
C11091 X1.X1.X1.X2.X1.X1.vout vss 0.842f
C11092 a_4782_16634# vss 0.854f
C11093 a_4396_16634# vss 1.67f
C11094 X1.X1.X1.X2.X1.X1.X2.vin1 vss 1.8f
C11095 a_54992_17452# vss 1.66f
C11096 X2.X2.X2.X1.X2.X2.X3.vin2 vss 1.52f
C11097 X2.X2.X2.X1.X2.X2.X2.vin1 vss 1.8f
C11098 a_54606_17452# vss 0.884f
C11099 X2.X2.X1.X2.X1.X1.X1.vin2 vss 2.17f
C11100 X2.X2.X1.X2.X1.X1.X3.vin1 vss 0.912f
C11101 X2.X2.X1.X2.X1.X1.X1.vin1 vss 2.05f
C11102 a_46502_17540# vss 0.855f
C11103 a_46116_17540# vss 1.66f
C11104 a_40352_17452# vss 1.66f
C11105 X2.X1.X2.X1.X2.X2.X3.vin2 vss 1.52f
C11106 X2.X1.X2.X1.X2.X2.X2.vin1 vss 1.79f
C11107 a_39966_17452# vss 0.884f
C11108 X2.X1.X1.X2.X1.X1.X1.vin2 vss 2.17f
C11109 X2.X1.X1.X2.X1.X1.X3.vin1 vss 0.912f
C11110 X2.X1.X1.X2.X1.X1.X1.vin1 vss 2.05f
C11111 a_31862_17540# vss 0.855f
C11112 a_31476_17540# vss 1.66f
C11113 a_25712_17452# vss 1.66f
C11114 X1.X2.X2.X1.X2.X2.X3.vin2 vss 1.52f
C11115 X1.X2.X2.X1.X2.X2.X2.vin1 vss 1.79f
C11116 a_25326_17452# vss 0.884f
C11117 X1.X2.X1.X2.X1.X1.X1.vin2 vss 2.17f
C11118 X1.X2.X1.X2.X1.X1.X3.vin1 vss 0.912f
C11119 X1.X2.X1.X2.X1.X1.X1.vin1 vss 2.05f
C11120 a_17222_17540# vss 0.855f
C11121 a_16836_17540# vss 1.66f
C11122 a_11072_17452# vss 1.66f
C11123 X1.X1.X2.X1.X2.X2.X3.vin2 vss 1.52f
C11124 X1.X1.X2.X1.X2.X2.X2.vin1 vss 1.79f
C11125 a_10686_17452# vss 0.884f
C11126 X1.X1.X1.X2.X1.X1.X1.vin2 vss 2.18f
C11127 X1.X1.X1.X2.X1.X1.X3.vin1 vss 0.912f
C11128 X1.X1.X1.X2.X1.X1.X1.vin1 vss 2.05f
C11129 a_2582_17540# vss 0.855f
C11130 a_2196_17540# vss 1.66f
C11131 a_52492_18358# vss 1.67f
C11132 X2.X2.X3.vin2 vss 3.99f
C11133 X2.X2.X2.X3.vin1 vss 1.68f
C11134 a_52106_18358# vss 0.909f
C11135 X2.X2.X1.X3.vin2 vss 2.13f
C11136 X2.X2.X3.vin1 vss 3.21f
C11137 a_49002_18540# vss 0.91f
C11138 a_48616_18540# vss 1.67f
C11139 a_37852_18358# vss 1.67f
C11140 X2.X1.X3.vin2 vss 3.97f
C11141 X2.X1.X2.X3.vin1 vss 1.68f
C11142 a_37466_18358# vss 0.909f
C11143 X2.X1.X1.X3.vin2 vss 2.12f
C11144 X2.X1.X3.vin1 vss 3.19f
C11145 a_34362_18540# vss 0.91f
C11146 a_33976_18540# vss 1.67f
C11147 a_23212_18358# vss 1.67f
C11148 X1.X2.X3.vin2 vss 3.94f
C11149 X1.X2.X2.X3.vin1 vss 1.68f
C11150 a_22826_18358# vss 0.909f
C11151 X1.X2.X1.X3.vin2 vss 2.13f
C11152 X1.X2.X3.vin1 vss 3.19f
C11153 a_19722_18540# vss 0.91f
C11154 a_19336_18540# vss 1.67f
C11155 a_8572_18358# vss 1.67f
C11156 X1.X1.X3.vin2 vss 4f
C11157 X1.X1.X2.X3.vin1 vss 1.68f
C11158 a_8186_18358# vss 0.909f
C11159 X1.X1.X1.X3.vin2 vss 2.12f
C11160 X1.X1.X3.vin1 vss 3.21f
C11161 a_5082_18540# vss 0.91f
C11162 a_4696_18540# vss 1.67f
C11163 d4 vss 34.8f
C11164 X2.X2.X2.X2.vrefh vss 4.21f
C11165 a_54992_19358# vss 1.66f
C11166 X2.X2.X2.X2.X1.X1.X1.vin1 vss 2.05f
C11167 a_54606_19358# vss 0.855f
C11168 X2.X2.X2.X2.X1.X1.X1.vin2 vss 2.18f
C11169 a_46502_19446# vss 0.884f
C11170 a_46116_19446# vss 1.66f
C11171 X2.X1.X2.X2.vrefh vss 4.05f
C11172 X2.X2.X1.X2.vrefh vss 4.05f
C11173 a_52792_20264# vss 1.67f
C11174 X2.X2.X2.X2.X1.X1.X3.vin1 vss 0.912f
C11175 a_52406_20264# vss 0.854f
C11176 X2.X2.X1.X1.X2.X2.X3.vin2 vss 1.52f
C11177 a_48702_20446# vss 0.945f
C11178 a_48316_20446# vss 1.67f
C11179 X2.X2.X1.X1.X2.X2.X2.vin1 vss 1.79f
C11180 a_40352_19358# vss 1.66f
C11181 X2.X1.X2.X2.X1.X1.X1.vin1 vss 2.05f
C11182 a_39966_19358# vss 0.855f
C11183 X2.X1.X2.X2.X1.X1.X1.vin2 vss 2.17f
C11184 a_31862_19446# vss 0.884f
C11185 a_31476_19446# vss 1.66f
C11186 X1.X2.X2.X2.vrefh vss 4.05f
C11187 X2.X1.X1.X2.vrefh vss 4.05f
C11188 a_38152_20264# vss 1.67f
C11189 X2.X1.X2.X2.X1.X1.X3.vin1 vss 0.912f
C11190 a_37766_20264# vss 0.854f
C11191 X2.X1.X1.X1.X2.X2.X3.vin2 vss 1.52f
C11192 a_34062_20446# vss 0.945f
C11193 a_33676_20446# vss 1.67f
C11194 X2.X1.X1.X1.X2.X2.X2.vin1 vss 1.79f
C11195 a_25712_19358# vss 1.66f
C11196 X1.X2.X2.X2.X1.X1.X1.vin1 vss 2.05f
C11197 a_25326_19358# vss 0.855f
C11198 X1.X2.X2.X2.X1.X1.X1.vin2 vss 2.17f
C11199 a_17222_19446# vss 0.884f
C11200 a_16836_19446# vss 1.66f
C11201 X1.X1.X2.X2.vrefh vss 4.05f
C11202 X1.X2.X1.X2.vrefh vss 4.05f
C11203 a_23512_20264# vss 1.67f
C11204 X1.X2.X2.X2.X1.X1.X3.vin1 vss 0.912f
C11205 a_23126_20264# vss 0.854f
C11206 X1.X2.X1.X1.X2.X2.X3.vin2 vss 1.52f
C11207 a_19422_20446# vss 0.945f
C11208 a_19036_20446# vss 1.67f
C11209 X1.X2.X1.X1.X2.X2.X2.vin1 vss 1.79f
C11210 a_11072_19358# vss 1.66f
C11211 X1.X1.X2.X2.X1.X1.X1.vin1 vss 2.05f
C11212 a_10686_19358# vss 0.855f
C11213 X1.X1.X2.X2.X1.X1.X1.vin2 vss 2.17f
C11214 a_2582_19446# vss 0.884f
C11215 a_2196_19446# vss 1.66f
C11216 X1.X1.X1.X2.vrefh vss 4.21f
C11217 a_8872_20264# vss 1.67f
C11218 X1.X1.X2.X2.X1.X1.X3.vin1 vss 0.912f
C11219 a_8486_20264# vss 0.854f
C11220 X1.X1.X1.X1.X2.X2.X3.vin2 vss 1.52f
C11221 a_4782_20446# vss 0.945f
C11222 a_4396_20446# vss 1.67f
C11223 X1.X1.X1.X1.X2.X2.X2.vin1 vss 1.8f
C11224 a_54992_21264# vss 1.66f
C11225 X2.X2.X2.X2.X1.X1.X3.vin2 vss 1.3f
C11226 X2.X2.X2.X2.X1.X1.X2.vin1 vss 1.8f
C11227 a_54606_21264# vss 0.883f
C11228 X2.X2.X1.X1.X2.X2.X1.vin2 vss 2.17f
C11229 X2.X2.X1.X1.X2.X2.X3.vin1 vss 0.888f
C11230 X2.X2.X1.X1.X2.X2.X1.vin1 vss 2.05f
C11231 a_46502_21352# vss 0.856f
C11232 a_46116_21352# vss 1.66f
C11233 a_40352_21264# vss 1.66f
C11234 X2.X1.X2.X2.X1.X1.X3.vin2 vss 1.3f
C11235 X2.X1.X2.X2.X1.X1.X2.vin1 vss 1.79f
C11236 a_39966_21264# vss 0.883f
C11237 X2.X1.X1.X1.X2.X2.X1.vin2 vss 2.17f
C11238 X2.X1.X1.X1.X2.X2.X3.vin1 vss 0.888f
C11239 X2.X1.X1.X1.X2.X2.X1.vin1 vss 2.05f
C11240 a_31862_21352# vss 0.856f
C11241 a_31476_21352# vss 1.66f
C11242 a_25712_21264# vss 1.66f
C11243 X1.X2.X2.X2.X1.X1.X3.vin2 vss 1.3f
C11244 X1.X2.X2.X2.X1.X1.X2.vin1 vss 1.79f
C11245 a_25326_21264# vss 0.883f
C11246 X1.X2.X1.X1.X2.X2.X1.vin2 vss 2.17f
C11247 X1.X2.X1.X1.X2.X2.X3.vin1 vss 0.888f
C11248 X1.X2.X1.X1.X2.X2.X1.vin1 vss 2.05f
C11249 a_17222_21352# vss 0.856f
C11250 a_16836_21352# vss 1.66f
C11251 a_11072_21264# vss 1.66f
C11252 X1.X1.X2.X2.X1.X1.X3.vin2 vss 1.3f
C11253 X1.X1.X2.X2.X1.X1.X2.vin1 vss 1.79f
C11254 a_10686_21264# vss 0.883f
C11255 X1.X1.X1.X1.X2.X2.X1.vin2 vss 2.18f
C11256 X1.X1.X1.X1.X2.X2.X3.vin1 vss 0.888f
C11257 X1.X1.X1.X1.X2.X2.X1.vin1 vss 2.05f
C11258 a_2582_21352# vss 0.856f
C11259 a_2196_21352# vss 1.66f
C11260 a_52492_22210# vss 1.66f
C11261 X2.X2.X2.X2.X1.X1.vout vss 0.841f
C11262 a_52106_22210# vss 0.909f
C11263 X2.X2.X1.X1.X2.X2.vout vss 1.04f
C11264 a_49002_22312# vss 0.876f
C11265 a_48616_22312# vss 1.66f
C11266 a_37852_22210# vss 1.66f
C11267 X2.X1.X2.X2.X1.X1.vout vss 0.842f
C11268 a_37466_22210# vss 0.909f
C11269 X2.X1.X1.X1.X2.X2.vout vss 1.04f
C11270 a_34362_22312# vss 0.876f
C11271 a_33976_22312# vss 1.66f
C11272 a_23212_22210# vss 1.66f
C11273 X1.X2.X2.X2.X1.X1.vout vss 0.841f
C11274 a_22826_22210# vss 0.909f
C11275 X1.X2.X1.X1.X2.X2.vout vss 1.04f
C11276 a_19722_22312# vss 0.876f
C11277 a_19336_22312# vss 1.66f
C11278 a_8572_22210# vss 1.66f
C11279 X1.X1.X2.X2.X1.X1.vout vss 0.842f
C11280 a_8186_22210# vss 0.909f
C11281 X1.X1.X1.X1.X2.X2.vout vss 1.04f
C11282 a_5082_22312# vss 0.876f
C11283 a_4696_22312# vss 1.66f
C11284 X2.X2.X2.X2.X1.X2.vrefh vss 4.21f
C11285 a_54992_23170# vss 1.66f
C11286 X2.X2.X2.X2.X1.X2.X1.vin1 vss 2.05f
C11287 a_54606_23170# vss 0.856f
C11288 X2.X2.X2.X2.X1.X2.X1.vin2 vss 2.19f
C11289 a_46502_23258# vss 0.883f
C11290 a_46116_23258# vss 1.66f
C11291 X2.X1.X2.X2.X1.X2.vrefh vss 4.05f
C11292 X2.X2.X1.X1.X2.X2.vrefh vss 4.05f
C11293 a_52792_24076# vss 1.67f
C11294 X2.X2.X2.X2.X1.X2.vout vss 1.04f
C11295 X2.X2.X2.X2.X1.X2.X3.vin1 vss 0.887f
C11296 a_52406_24076# vss 0.945f
C11297 X2.X2.X1.X1.X2.X1.X3.vin2 vss 1.28f
C11298 X2.X2.X1.X1.X2.X1.vout vss 0.789f
C11299 a_48702_24258# vss 0.854f
C11300 a_48316_24258# vss 1.67f
C11301 X2.X2.X1.X1.X2.X1.X2.vin1 vss 1.79f
C11302 a_40352_23170# vss 1.66f
C11303 X2.X1.X2.X2.X1.X2.X1.vin1 vss 2.05f
C11304 a_39966_23170# vss 0.856f
C11305 X2.X1.X2.X2.X1.X2.X1.vin2 vss 2.17f
C11306 a_31862_23258# vss 0.883f
C11307 a_31476_23258# vss 1.66f
C11308 X1.X2.X2.X2.X1.X2.vrefh vss 4.05f
C11309 X2.X1.X1.X1.X2.X2.vrefh vss 4.05f
C11310 a_38152_24076# vss 1.67f
C11311 X2.X1.X2.X2.X1.X2.vout vss 1.04f
C11312 X2.X1.X2.X2.X1.X2.X3.vin1 vss 0.887f
C11313 a_37766_24076# vss 0.945f
C11314 X2.X1.X1.X1.X2.X1.X3.vin2 vss 1.28f
C11315 X2.X1.X1.X1.X2.X1.vout vss 0.788f
C11316 a_34062_24258# vss 0.854f
C11317 a_33676_24258# vss 1.67f
C11318 X2.X1.X1.X1.X2.X1.X2.vin1 vss 1.79f
C11319 a_25712_23170# vss 1.66f
C11320 X1.X2.X2.X2.X1.X2.X1.vin1 vss 2.05f
C11321 a_25326_23170# vss 0.856f
C11322 X1.X2.X2.X2.X1.X2.X1.vin2 vss 2.17f
C11323 a_17222_23258# vss 0.883f
C11324 a_16836_23258# vss 1.66f
C11325 X1.X1.X2.X2.X1.X2.vrefh vss 4.05f
C11326 X1.X2.X1.X1.X2.X2.vrefh vss 4.05f
C11327 a_23512_24076# vss 1.67f
C11328 X1.X2.X2.X2.X1.X2.vout vss 1.04f
C11329 X1.X2.X2.X2.X1.X2.X3.vin1 vss 0.887f
C11330 a_23126_24076# vss 0.945f
C11331 X1.X2.X1.X1.X2.X1.X3.vin2 vss 1.28f
C11332 X1.X2.X1.X1.X2.X1.vout vss 0.789f
C11333 a_19422_24258# vss 0.854f
C11334 a_19036_24258# vss 1.67f
C11335 X1.X2.X1.X1.X2.X1.X2.vin1 vss 1.79f
C11336 a_11072_23170# vss 1.66f
C11337 X1.X1.X2.X2.X1.X2.X1.vin1 vss 2.05f
C11338 a_10686_23170# vss 0.856f
C11339 X1.X1.X2.X2.X1.X2.X1.vin2 vss 2.17f
C11340 a_2582_23258# vss 0.883f
C11341 a_2196_23258# vss 1.66f
C11342 X1.X1.X1.X1.X2.X2.vrefh vss 4.21f
C11343 a_8872_24076# vss 1.67f
C11344 X1.X1.X2.X2.X1.X2.vout vss 1.04f
C11345 X1.X1.X2.X2.X1.X2.X3.vin1 vss 0.887f
C11346 a_8486_24076# vss 0.945f
C11347 X1.X1.X1.X1.X2.X1.X3.vin2 vss 1.28f
C11348 X1.X1.X1.X1.X2.X1.vout vss 0.788f
C11349 a_4782_24258# vss 0.854f
C11350 a_4396_24258# vss 1.67f
C11351 X1.X1.X1.X1.X2.X1.X2.vin1 vss 1.8f
C11352 a_54992_25076# vss 1.66f
C11353 X2.X2.X2.X2.X1.X2.X3.vin2 vss 1.5f
C11354 X2.X2.X2.X2.X1.X2.X2.vin1 vss 1.8f
C11355 a_54606_25076# vss 0.884f
C11356 X2.X2.X1.X1.X2.X1.X1.vin2 vss 2.17f
C11357 X2.X2.X1.X1.X2.X1.X3.vin1 vss 0.905f
C11358 X2.X2.X1.X1.X2.X1.X1.vin1 vss 2.05f
C11359 a_46502_25164# vss 0.855f
C11360 a_46116_25164# vss 1.66f
C11361 a_40352_25076# vss 1.66f
C11362 X2.X1.X2.X2.X1.X2.X3.vin2 vss 1.5f
C11363 X2.X1.X2.X2.X1.X2.X2.vin1 vss 1.79f
C11364 a_39966_25076# vss 0.884f
C11365 X2.X1.X1.X1.X2.X1.X1.vin2 vss 2.17f
C11366 X2.X1.X1.X1.X2.X1.X3.vin1 vss 0.905f
C11367 X2.X1.X1.X1.X2.X1.X1.vin1 vss 2.05f
C11368 a_31862_25164# vss 0.855f
C11369 a_31476_25164# vss 1.66f
C11370 a_25712_25076# vss 1.66f
C11371 X1.X2.X2.X2.X1.X2.X3.vin2 vss 1.5f
C11372 X1.X2.X2.X2.X1.X2.X2.vin1 vss 1.79f
C11373 a_25326_25076# vss 0.884f
C11374 X1.X2.X1.X1.X2.X1.X1.vin2 vss 2.17f
C11375 X1.X2.X1.X1.X2.X1.X3.vin1 vss 0.905f
C11376 X1.X2.X1.X1.X2.X1.X1.vin1 vss 2.05f
C11377 a_17222_25164# vss 0.855f
C11378 a_16836_25164# vss 1.66f
C11379 a_11072_25076# vss 1.66f
C11380 X1.X1.X2.X2.X1.X2.X3.vin2 vss 1.5f
C11381 X1.X1.X2.X2.X1.X2.X2.vin1 vss 1.79f
C11382 a_10686_25076# vss 0.884f
C11383 X1.X1.X1.X1.X2.X1.X1.vin2 vss 2.18f
C11384 X1.X1.X1.X1.X2.X1.X3.vin1 vss 0.905f
C11385 X1.X1.X1.X1.X2.X1.X1.vin1 vss 2.05f
C11386 a_2582_25164# vss 0.855f
C11387 a_2196_25164# vss 1.66f
C11388 a_52492_25982# vss 1.67f
C11389 X2.X2.X2.X3.vin2 vss 2.05f
C11390 X2.X2.X2.X2.X3.vin1 vss 2.11f
C11391 a_52106_25982# vss 0.93f
C11392 X2.X2.X1.X1.X3.vin2 vss 1.73f
C11393 X2.X2.X1.X3.vin1 vss 1.91f
C11394 a_49002_26164# vss 0.926f
C11395 a_48616_26164# vss 1.67f
C11396 a_37852_25982# vss 1.67f
C11397 X2.X1.X2.X3.vin2 vss 2.29f
C11398 X2.X1.X2.X2.X3.vin1 vss 2.11f
C11399 a_37466_25982# vss 0.93f
C11400 X2.X1.X1.X1.X3.vin2 vss 1.74f
C11401 X2.X1.X1.X3.vin1 vss 1.67f
C11402 a_34362_26164# vss 0.926f
C11403 a_33976_26164# vss 1.67f
C11404 a_23212_25982# vss 1.67f
C11405 X1.X2.X2.X3.vin2 vss 2.05f
C11406 X1.X2.X2.X2.X3.vin1 vss 2.11f
C11407 a_22826_25982# vss 0.93f
C11408 X1.X2.X1.X1.X3.vin2 vss 1.73f
C11409 X1.X2.X1.X3.vin1 vss 1.91f
C11410 a_19722_26164# vss 0.926f
C11411 a_19336_26164# vss 1.67f
C11412 a_8572_25982# vss 1.67f
C11413 X1.X1.X2.X3.vin2 vss 2.29f
C11414 X1.X1.X2.X2.X3.vin1 vss 2.11f
C11415 a_8186_25982# vss 0.93f
C11416 X1.X1.X1.X1.X3.vin2 vss 1.74f
C11417 X1.X1.X1.X3.vin1 vss 1.67f
C11418 a_5082_26164# vss 0.926f
C11419 a_4696_26164# vss 1.67f
C11420 d3 vss 83.5f
C11421 X2.X2.X2.X2.X2.vrefh vss 4.21f
C11422 a_54992_26982# vss 1.66f
C11423 X2.X2.X2.X2.X2.X1.X1.vin1 vss 2.05f
C11424 a_54606_26982# vss 0.855f
C11425 X2.X2.X2.X2.X2.X1.X1.vin2 vss 2.18f
C11426 a_46502_27070# vss 0.884f
C11427 a_46116_27070# vss 1.66f
C11428 X2.X1.X2.X2.X2.vrefh vss 4.06f
C11429 X2.X2.X1.X1.X2.vrefh vss 4.06f
C11430 a_52792_27888# vss 1.67f
C11431 X2.X2.X2.X2.X2.X1.X3.vin1 vss 0.91f
C11432 a_52406_27888# vss 0.854f
C11433 X2.X2.X1.X1.X1.X2.X3.vin2 vss 1.52f
C11434 a_48702_28070# vss 0.945f
C11435 a_48316_28070# vss 1.67f
C11436 X2.X2.X1.X1.X1.X2.X2.vin1 vss 1.79f
C11437 a_40352_26982# vss 1.66f
C11438 X2.X1.X2.X2.X2.X1.X1.vin1 vss 2.05f
C11439 a_39966_26982# vss 0.855f
C11440 X2.X1.X2.X2.X2.X1.X1.vin2 vss 2.17f
C11441 a_31862_27070# vss 0.884f
C11442 a_31476_27070# vss 1.66f
C11443 X1.X2.X2.X2.X2.vrefh vss 4.06f
C11444 X2.X1.X1.X1.X2.vrefh vss 4.06f
C11445 a_38152_27888# vss 1.67f
C11446 X2.X1.X2.X2.X2.X1.X3.vin1 vss 0.905f
C11447 a_37766_27888# vss 0.854f
C11448 X2.X1.X1.X1.X1.X2.X3.vin2 vss 1.54f
C11449 a_34062_28070# vss 0.945f
C11450 a_33676_28070# vss 1.67f
C11451 X2.X1.X1.X1.X1.X2.X2.vin1 vss 1.79f
C11452 a_25712_26982# vss 1.66f
C11453 X1.X2.X2.X2.X2.X1.X1.vin1 vss 2.05f
C11454 a_25326_26982# vss 0.855f
C11455 X1.X2.X2.X2.X2.X1.X1.vin2 vss 2.17f
C11456 a_17222_27070# vss 0.884f
C11457 a_16836_27070# vss 1.66f
C11458 X1.X1.X2.X2.X2.vrefh vss 4.06f
C11459 X1.X2.X1.X1.X2.vrefh vss 4.06f
C11460 a_23512_27888# vss 1.67f
C11461 X1.X2.X2.X2.X2.X1.X3.vin1 vss 0.91f
C11462 a_23126_27888# vss 0.854f
C11463 X1.X2.X1.X1.X1.X2.X3.vin2 vss 1.52f
C11464 a_19422_28070# vss 0.945f
C11465 a_19036_28070# vss 1.67f
C11466 X1.X2.X1.X1.X1.X2.X2.vin1 vss 1.79f
C11467 a_11072_26982# vss 1.66f
C11468 X1.X1.X2.X2.X2.X1.X1.vin1 vss 2.05f
C11469 a_10686_26982# vss 0.855f
C11470 X1.X1.X2.X2.X2.X1.X1.vin2 vss 2.17f
C11471 a_2582_27070# vss 0.884f
C11472 a_2196_27070# vss 1.66f
C11473 X1.X1.X1.X1.X2.vrefh vss 4.21f
C11474 a_8872_27888# vss 1.67f
C11475 X1.X1.X2.X2.X2.X1.X3.vin1 vss 0.905f
C11476 a_8486_27888# vss 0.854f
C11477 X1.X1.X1.X1.X1.X2.X3.vin2 vss 1.54f
C11478 a_4782_28070# vss 0.945f
C11479 a_4396_28070# vss 1.67f
C11480 X1.X1.X1.X1.X1.X2.X2.vin1 vss 1.8f
C11481 a_54992_28888# vss 1.66f
C11482 X2.X2.X2.X2.X2.X1.X3.vin2 vss 1.31f
C11483 X2.X2.X2.X2.X2.X1.X2.vin1 vss 1.8f
C11484 a_54606_28888# vss 0.883f
C11485 X2.X2.X1.X1.X1.X2.X1.vin2 vss 2.17f
C11486 X2.X2.X1.X1.X1.X2.X3.vin1 vss 0.89f
C11487 X2.X2.X1.X1.X1.X2.X1.vin1 vss 2.05f
C11488 a_46502_28976# vss 0.856f
C11489 a_46116_28976# vss 1.66f
C11490 a_40352_28888# vss 1.66f
C11491 X2.X1.X2.X2.X2.X1.X3.vin2 vss 1.28f
C11492 X2.X1.X2.X2.X2.X1.X2.vin1 vss 1.79f
C11493 a_39966_28888# vss 0.883f
C11494 X2.X1.X1.X1.X1.X2.X1.vin2 vss 2.17f
C11495 X2.X1.X1.X1.X1.X2.X3.vin1 vss 0.892f
C11496 X2.X1.X1.X1.X1.X2.X1.vin1 vss 2.05f
C11497 a_31862_28976# vss 0.856f
C11498 a_31476_28976# vss 1.66f
C11499 a_25712_28888# vss 1.66f
C11500 X1.X2.X2.X2.X2.X1.X3.vin2 vss 1.31f
C11501 X1.X2.X2.X2.X2.X1.X2.vin1 vss 1.79f
C11502 a_25326_28888# vss 0.883f
C11503 X1.X2.X1.X1.X1.X2.X1.vin2 vss 2.17f
C11504 X1.X2.X1.X1.X1.X2.X3.vin1 vss 0.89f
C11505 X1.X2.X1.X1.X1.X2.X1.vin1 vss 2.05f
C11506 a_17222_28976# vss 0.856f
C11507 a_16836_28976# vss 1.66f
C11508 a_11072_28888# vss 1.66f
C11509 X1.X1.X2.X2.X2.X1.X3.vin2 vss 1.28f
C11510 X1.X1.X2.X2.X2.X1.X2.vin1 vss 1.79f
C11511 a_10686_28888# vss 0.883f
C11512 X1.X1.X1.X1.X1.X2.X1.vin2 vss 2.19f
C11513 X1.X1.X1.X1.X1.X2.X3.vin1 vss 0.892f
C11514 X1.X1.X1.X1.X1.X2.X1.vin1 vss 2.05f
C11515 a_2582_28976# vss 0.856f
C11516 a_2196_28976# vss 1.66f
C11517 a_52492_29834# vss 1.66f
C11518 X2.X2.X2.X2.X3.vin2 vss 1.95f
C11519 X2.X2.X2.X2.X2.X1.vout vss 0.814f
C11520 a_52106_29834# vss 0.962f
C11521 X2.X2.X1.X1.X1.X2.vout vss 1.08f
C11522 X2.X2.X1.X1.X3.vin1 vss 2.31f
C11523 a_49002_29936# vss 0.96f
C11524 a_48616_29936# vss 1.66f
C11525 a_37852_29834# vss 1.66f
C11526 X2.X1.X2.X2.X3.vin2 vss 1.92f
C11527 X2.X1.X2.X2.X2.X1.vout vss 0.8f
C11528 a_37466_29834# vss 0.962f
C11529 X2.X1.X1.X1.X1.X2.vout vss 1.11f
C11530 X2.X1.X1.X1.X3.vin1 vss 2.32f
C11531 a_34362_29936# vss 0.96f
C11532 a_33976_29936# vss 1.66f
C11533 a_23212_29834# vss 1.66f
C11534 X1.X2.X2.X2.X3.vin2 vss 1.95f
C11535 X1.X2.X2.X2.X2.X1.vout vss 0.814f
C11536 a_22826_29834# vss 0.962f
C11537 X1.X2.X1.X1.X1.X2.vout vss 1.08f
C11538 X1.X2.X1.X1.X3.vin1 vss 2.31f
C11539 a_19722_29936# vss 0.96f
C11540 a_19336_29936# vss 1.66f
C11541 a_8572_29834# vss 1.66f
C11542 X1.X1.X2.X2.X3.vin2 vss 1.92f
C11543 X1.X1.X2.X2.X2.X1.vout vss 0.8f
C11544 a_8186_29834# vss 0.962f
C11545 X1.X1.X1.X1.X1.X2.vout vss 1.11f
C11546 X1.X1.X1.X1.X3.vin1 vss 2.32f
C11547 a_5082_29936# vss 0.96f
C11548 a_4696_29936# vss 1.66f
C11549 d2 vss 88.9f
C11550 X2.X2.X2.X2.X2.X2.vrefh vss 4.21f
C11551 a_54992_30794# vss 1.66f
C11552 X2.X2.X2.X2.X2.X2.X1.vin1 vss 2.05f
C11553 a_54606_30794# vss 0.856f
C11554 X2.X2.X2.X2.X2.X2.X1.vin2 vss 2.24f
C11555 a_46502_30882# vss 0.883f
C11556 a_46116_30882# vss 1.66f
C11557 X2.X1.X2.X2.X2.X2.vrefh vss 4.05f
C11558 X2.X2.X1.X1.X1.X2.vrefh vss 4.07f
C11559 a_52792_31700# vss 1.67f
C11560 X2.X2.X2.X2.X2.X2.vout vss 1.17f
C11561 X2.X2.X2.X2.X2.X2.X3.vin1 vss 0.899f
C11562 a_52406_31700# vss 0.967f
C11563 X2.X2.X1.X1.X1.X1.X3.vin2 vss 1.32f
C11564 X2.X2.X1.X1.X1.X1.vout vss 0.853f
C11565 a_48702_31882# vss 0.879f
C11566 a_48316_31882# vss 1.67f
C11567 X2.X2.X1.X1.X1.X1.X2.vin1 vss 1.8f
C11568 a_40352_30794# vss 1.66f
C11569 X2.X1.X2.X2.X2.X2.X1.vin1 vss 2.05f
C11570 a_39966_30794# vss 0.856f
C11571 X2.X1.X2.X2.X2.X2.X1.vin2 vss 2.22f
C11572 a_31862_30882# vss 0.883f
C11573 a_31476_30882# vss 1.66f
C11574 X1.X2.X2.X2.X2.X2.vrefh vss 4.05f
C11575 X2.X1.X1.X1.X1.X2.vrefh vss 4.07f
C11576 a_38152_31700# vss 1.67f
C11577 X2.X1.X2.X2.X2.X2.vout vss 1.11f
C11578 X2.X1.X2.X2.X2.X2.X3.vin1 vss 0.894f
C11579 a_37766_31700# vss 0.967f
C11580 X2.X1.X1.X1.X1.X1.X3.vin2 vss 1.34f
C11581 X2.X1.X1.X1.X1.X1.vout vss 0.861f
C11582 a_34062_31882# vss 0.879f
C11583 a_33676_31882# vss 1.67f
C11584 X2.X1.X1.X1.X1.X1.X2.vin1 vss 1.8f
C11585 a_25712_30794# vss 1.66f
C11586 X1.X2.X2.X2.X2.X2.X1.vin1 vss 2.05f
C11587 a_25326_30794# vss 0.856f
C11588 X1.X2.X2.X2.X2.X2.X1.vin2 vss 2.22f
C11589 a_17222_30882# vss 0.883f
C11590 a_16836_30882# vss 1.66f
C11591 X1.X1.X2.X2.X2.X2.vrefh vss 4.05f
C11592 X1.X2.X1.X1.X1.X2.vrefh vss 4.07f
C11593 a_23512_31700# vss 1.67f
C11594 X1.X2.X2.X2.X2.X2.vout vss 1.17f
C11595 X1.X2.X2.X2.X2.X2.X3.vin1 vss 0.899f
C11596 a_23126_31700# vss 0.967f
C11597 X1.X2.X1.X1.X1.X1.X3.vin2 vss 1.32f
C11598 X1.X2.X1.X1.X1.X1.vout vss 0.853f
C11599 a_19422_31882# vss 0.879f
C11600 a_19036_31882# vss 1.67f
C11601 X1.X2.X1.X1.X1.X1.X2.vin1 vss 1.8f
C11602 a_11072_30794# vss 1.66f
C11603 X1.X1.X2.X2.X2.X2.X1.vin1 vss 2.05f
C11604 a_10686_30794# vss 0.856f
C11605 X1.X1.X2.X2.X2.X2.X1.vin2 vss 2.22f
C11606 a_2582_30882# vss 0.883f
C11607 a_2196_30882# vss 1.66f
C11608 X1.X1.X1.X1.X1.X2.vrefh vss 4.22f
C11609 a_8872_31700# vss 1.67f
C11610 X1.X1.X2.X2.X2.X2.vout vss 1.11f
C11611 X1.X1.X2.X2.X2.X2.X3.vin1 vss 0.894f
C11612 a_8486_31700# vss 0.967f
C11613 X1.X1.X1.X1.X1.X1.X3.vin2 vss 1.34f
C11614 X1.X1.X1.X1.X1.X1.vout vss 0.861f
C11615 a_4782_31882# vss 0.879f
C11616 a_4396_31882# vss 1.67f
C11617 d1 vss 0.112p
C11618 X1.X1.X1.X1.X1.X1.X2.vin1 vss 1.8f
C11619 vrefh vss 1.34f
C11620 vrefl vss 3.21f
C11621 a_54992_32700# vss 1.66f
C11622 X2.X2.X2.X2.X2.X2.X3.vin2 vss 1.76f
C11623 X2.X2.X2.X2.X2.X2.X2.vin1 vss 1.83f
C11624 a_54606_32700# vss 0.887f
C11625 X2.X2.X1.X1.X1.X1.X1.vin2 vss 2.31f
C11626 X2.X2.X1.X1.X1.X1.X3.vin1 vss 0.999f
C11627 X2.X2.X1.X1.X1.X1.X1.vin1 vss 2.3f
C11628 a_46502_32788# vss 0.884f
C11629 a_46116_32788# vss 1.67f
C11630 X2.X2.vrefh vss 4.97f
C11631 a_40352_32700# vss 1.67f
C11632 X2.X1.X2.X2.X2.X2.X3.vin2 vss 1.69f
C11633 X2.X1.X2.X2.X2.X2.X2.vin1 vss 1.82f
C11634 a_39966_32700# vss 0.888f
C11635 X2.X1.X1.X1.X1.X1.X1.vin2 vss 2.31f
C11636 X2.X1.X1.X1.X1.X1.X3.vin1 vss 1f
C11637 X2.X1.X1.X1.X1.X1.X1.vin1 vss 2.3f
C11638 a_31862_32788# vss 0.884f
C11639 a_31476_32788# vss 1.67f
C11640 X2.vrefh vss 4.97f
C11641 a_25712_32700# vss 1.67f
C11642 X1.X2.X2.X2.X2.X2.X3.vin2 vss 1.74f
C11643 X1.X2.X2.X2.X2.X2.X2.vin1 vss 1.82f
C11644 a_25326_32700# vss 0.888f
C11645 X1.X2.X1.X1.X1.X1.X1.vin2 vss 2.31f
C11646 X1.X2.X1.X1.X1.X1.X3.vin1 vss 0.999f
C11647 X1.X2.X1.X1.X1.X1.X1.vin1 vss 2.3f
C11648 a_17222_32788# vss 0.884f
C11649 a_16836_32788# vss 1.67f
C11650 X1.X2.vrefh vss 4.97f
C11651 a_11072_32700# vss 1.67f
C11652 X1.X1.X2.X2.X2.X2.X3.vin2 vss 1.69f
C11653 X1.X1.X2.X2.X2.X2.X2.vin1 vss 1.82f
C11654 a_10686_32700# vss 0.888f
C11655 X1.X1.X1.X1.X1.X1.X1.vin2 vss 2.33f
C11656 X1.X1.X1.X1.X1.X1.X3.vin1 vss 1.01f
C11657 X1.X1.X1.X1.X1.X1.X1.vin1 vss 2.34f
C11658 a_2582_32788# vss 0.884f
C11659 a_2196_32788# vss 1.67f
C11660 d0 vss 0.206p
C11661 vdd vss 1.43p
.ends

