* NGSPICE file created from sw.ext - technology: sky130B

.subckt sky130_fd_pr__pfet_01v8_XPYSY6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFH27D a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt sw vdd vss din vin1 vin2 vout
XM1 vdd din m1_994_178# vdd sky130_fd_pr__pfet_01v8_XPYSY6
XM2 vdd m1_994_178# m1_688_n494# vdd sky130_fd_pr__pfet_01v8_XPYSY6
XM3 vdd m1_994_178# vout vin1 sky130_fd_pr__pfet_01v8_XPYSY6
XM4 vdd m1_688_n494# vin2 vout sky130_fd_pr__pfet_01v8_XPYSY6
XM5 m1_994_178# vss vss din sky130_fd_pr__nfet_01v8_ZFH27D
XM6 m1_688_n494# vss vss m1_994_178# sky130_fd_pr__nfet_01v8_ZFH27D
XM7 vout vss vin2 m1_994_178# sky130_fd_pr__nfet_01v8_ZFH27D
XM8 vin1 vss vout m1_688_n494# sky130_fd_pr__nfet_01v8_ZFH27D
.ends

