magic
tech sky130B
timestamp 1687755428
<< nwell >>
rect 141 0 244 200
rect 343 0 447 200
rect 554 0 630 200
<< metal1 >>
rect -6 50 44 150
rect 100 50 150 150
rect 200 50 250 150
rect 306 50 356 150
rect 406 50 456 150
rect 512 50 562 150
rect 612 50 662 150
rect 718 50 768 150
rect -200 0 -160 40
rect -200 -200 -160 -160
rect -200 -400 -160 -360
rect -200 -600 -160 -560
rect -200 -800 -160 -760
rect -200 -1000 -160 -960
use sky130_fd_pr__pfet_01v8_XPG7Y6  XM1
timestamp 1687754106
transform 1 0 72 0 1 100
box -72 -100 72 100
use sky130_fd_pr__pfet_01v8_XPG7Y6  XM2
timestamp 1687754106
transform 1 0 278 0 1 100
box -72 -100 72 100
use sky130_fd_pr__pfet_01v8_XPG7Y6  XM3
timestamp 1687754106
transform 1 0 484 0 1 100
box -72 -100 72 100
use sky130_fd_pr__pfet_01v8_XPG7Y6  XM4
timestamp 1687754106
transform 1 0 690 0 1 100
box -72 -100 72 100
use sky130_fd_pr__nfet_01v8_J3M27M  XM5
timestamp 1687754370
transform 1 0 72 0 1 -165
box -54 -65 54 65
use sky130_fd_pr__nfet_01v8_J3M27M  XM6
timestamp 1687754370
transform 1 0 278 0 1 -165
box -54 -65 54 65
use sky130_fd_pr__nfet_01v8_J3M27M  XM7
timestamp 1687754370
transform 1 0 484 0 1 -165
box -54 -65 54 65
use sky130_fd_pr__nfet_01v8_J3M27M  XM8
timestamp 1687754370
transform 1 0 690 0 1 -165
box -54 -65 54 65
<< labels >>
flabel metal1 -200 0 -160 40 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 -200 -200 -160 -160 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 -200 -400 -160 -360 0 FreeSans 128 0 0 0 din
port 2 nsew
flabel metal1 -200 -600 -160 -560 0 FreeSans 128 0 0 0 vin1
port 3 nsew
flabel metal1 -200 -800 -160 -760 0 FreeSans 128 0 0 0 vin2
port 4 nsew
flabel metal1 -200 -1000 -160 -960 0 FreeSans 128 0 0 0 vout
port 5 nsew
<< end >>