* NGSPICE file created from sw.ext - technology: sky130B

.subckt sky130_fd_pr__pfet_01v8_XPG7Y6 a_n50_n197# a_50_n100# w_n144_n200# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n144_n200# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_J3M27M a_50_n42# a_n108_n42# a_n50_n130# VSUBS
X0 a_50_n42# a_n50_n130# a_n108_n42# VSUBS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt sw vdd vss din vin1 vin2 vout
XXM1 din m1_942_58# w_n60_0# vdd sky130_fd_pr__pfet_01v8_XPG7Y6
XXM2 m1_942_58# m1_1356_58# w_n60_0# vdd sky130_fd_pr__pfet_01v8_XPG7Y6
XXM3 m1_942_58# vout w_n60_0# vin1 sky130_fd_pr__pfet_01v8_XPG7Y6
XXM4 m1_1356_58# vin2 w_n60_0# vout sky130_fd_pr__pfet_01v8_XPG7Y6
XXM5 m1_942_58# vss din VSUBS sky130_fd_pr__nfet_01v8_J3M27M
XXM6 m1_1356_58# vss m1_942_58# VSUBS sky130_fd_pr__nfet_01v8_J3M27M
XXM7 vout vin2 m1_942_58# VSUBS sky130_fd_pr__nfet_01v8_J3M27M
XXM8 vin1 vout m1_1356_58# VSUBS sky130_fd_pr__nfet_01v8_J3M27M
.ends

