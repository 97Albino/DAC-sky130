magic
tech sky130B
timestamp 1688376520
<< metal1 >>
rect 2187 1947 2227 1987
rect 548 1820 648 1920
rect 3275 1477 3425 1553
rect 2131 1266 2171 1306
rect 2450 1158 2490 1163
rect 2450 1128 2455 1158
rect 2485 1128 2490 1158
rect 2450 1123 2490 1128
rect 3037 951 3041 981
rect 3071 951 3077 981
rect 1350 623 1390 663
rect 3349 504 3425 1477
rect 1134 300 1156 301
rect 483 100 699 300
rect 1080 100 1156 300
rect 2450 -97 2526 403
rect 2600 150 2640 190
rect 3186 150 3226 190
rect 2450 -173 2600 -97
rect 3035 -540 3040 -510
rect 3070 -540 3075 -510
rect 2450 -778 2455 -748
rect 2485 -778 2490 -748
rect 3349 -1030 3425 -97
rect 3275 -1106 3425 -1030
rect 535 -1559 635 -1459
<< via1 >>
rect 2455 1128 2485 1158
rect 3041 951 3071 981
rect 3040 -540 3070 -510
rect 2455 -778 2485 -748
<< metal2 >>
rect 2450 1158 2490 1163
rect 2450 1128 2455 1158
rect 2485 1128 2490 1158
rect 590 623 1390 663
rect 590 -100 630 623
rect 2274 100 2350 300
rect 590 -140 1390 -100
rect 1350 -290 1390 -140
rect 2450 -748 2490 1128
rect 3035 981 3076 986
rect 3035 958 3041 981
rect 3071 958 3076 981
rect 3035 924 3039 958
rect 3073 924 3076 958
rect 3035 919 3076 924
rect 3035 835 3076 840
rect 3035 801 3039 835
rect 3073 801 3076 835
rect 3035 520 3076 801
rect 3035 -349 3075 -113
rect 3035 -383 3038 -349
rect 3072 -383 3075 -349
rect 3035 -390 3075 -383
rect 3035 -486 3075 -480
rect 3035 -520 3038 -486
rect 3072 -520 3075 -486
rect 3035 -540 3040 -520
rect 3070 -540 3075 -520
rect 3035 -545 3075 -540
rect 2450 -778 2455 -748
rect 2485 -778 2490 -748
rect 2450 -783 2490 -778
<< via2 >>
rect 3039 951 3041 958
rect 3041 951 3071 958
rect 3071 951 3073 958
rect 3039 924 3073 951
rect 3039 801 3073 835
rect 3038 -383 3072 -349
rect 3038 -510 3072 -486
rect 3038 -520 3040 -510
rect 3040 -520 3070 -510
rect 3070 -520 3072 -510
<< metal3 >>
rect 3034 958 3078 963
rect 3034 924 3039 958
rect 3073 924 3078 958
rect 3034 835 3078 924
rect 3034 801 3039 835
rect 3073 801 3078 835
rect 3034 796 3078 801
rect 3033 -349 3077 -346
rect 3033 -383 3038 -349
rect 3072 -383 3077 -349
rect 3033 -486 3077 -383
rect 3033 -520 3038 -486
rect 3072 -520 3077 -486
rect 3033 -523 3077 -520
use sw  sw_0
timestamp 1687966408
transform 1 0 2600 0 1 220
box 0 -393 860 360
use 2bit_dac  X1
timestamp 1688370130
transform 1 0 1350 0 1 1253
box -950 -953 1960 753
use 2bit_dac  X2
timestamp 1688370130
transform 1 0 1350 0 1 -653
box -950 -953 1960 753
<< labels >>
flabel metal1 548 1820 648 1920 0 FreeSans 128 0 0 0 vrefh
port 2 nsew
flabel metal1 535 -1559 635 -1459 0 FreeSans 128 0 0 0 vrefl
port 3 nsew
flabel metal1 2187 1947 2227 1987 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 1350 623 1390 663 0 FreeSans 128 0 0 0 d0
port 4 nsew
flabel metal1 2450 1123 2490 1163 0 FreeSans 128 0 0 0 d1
port 5 nsew
flabel metal1 2600 150 2640 190 0 FreeSans 128 0 0 0 d2
port 6 nsew
flabel metal1 3186 150 3226 190 0 FreeSans 128 0 0 0 vout
port 7 nsew
flabel metal1 2131 1266 2171 1306 0 FreeSans 128 0 0 0 vss
port 1 nsew
<< end >>
