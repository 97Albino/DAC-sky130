magic
tech sky130B
timestamp 1688891632
<< metal1 >>
rect 10960 17410 18020 17455
rect 10640 17320 18455 17365
rect 10825 17230 18250 17275
rect 4970 17077 8000 17153
rect 12290 17077 15320 17153
rect 19610 17077 22640 17153
rect 1801 16953 1841 16993
rect 132 16830 232 16930
rect 14041 16785 14939 17001
rect 28742 16852 28842 16952
rect 950 16571 990 16611
rect 1720 16262 1760 16302
rect 2050 16118 2090 16158
rect 2200 15145 2240 15185
rect 2200 13259 2240 13299
rect 2200 9447 2240 9487
rect 14150 1333 14830 1373
rect 12290 1230 19570 1270
rect 9830 1120 17200 1160
rect 10820 977 17009 1053
rect 2675 623 2715 663
rect 6600 658 6740 663
rect 6600 628 6605 658
rect 6635 628 6740 658
rect 6600 623 6740 628
rect 13900 623 13940 663
rect 14485 632 14525 672
rect 21240 658 21340 663
rect 21240 628 21245 658
rect 21275 628 21340 658
rect 21240 623 21340 628
rect 7285 558 7290 588
rect 7320 558 7325 588
rect 21925 558 21930 588
rect 21960 558 21965 588
rect 11126 300 17315 376
rect 6600 235 21280 240
rect 6600 205 6605 235
rect 6635 205 21245 235
rect 21275 205 21280 235
rect 6600 200 21280 205
rect 7285 135 11900 140
rect 7285 105 7290 135
rect 7320 105 11865 135
rect 11895 105 11900 135
rect 7285 100 11900 105
rect 14715 125 21965 130
rect 14715 95 14720 125
rect 14750 95 21930 125
rect 21960 95 21965 125
rect 14715 90 21965 95
<< via1 >>
rect 6605 628 6635 658
rect 21245 628 21275 658
rect 7290 558 7320 588
rect 21930 558 21960 588
rect 6605 205 6635 235
rect 21245 205 21275 235
rect 7290 105 7320 135
rect 11865 105 11895 135
rect 14720 95 14750 125
rect 21930 95 21960 125
<< metal2 >>
rect 11860 953 14335 993
rect 6600 658 6640 663
rect 6600 628 6605 658
rect 6635 628 6640 658
rect 6600 235 6640 628
rect 7285 588 7326 593
rect 7285 558 7290 588
rect 7320 558 7326 588
rect 7285 527 7326 558
rect 7285 495 7289 527
rect 7321 495 7326 527
rect 7285 488 7326 495
rect 6600 205 6605 235
rect 6635 205 6640 235
rect 6600 200 6640 205
rect 7285 296 7325 301
rect 7285 264 7289 296
rect 7321 264 7325 296
rect 7285 135 7325 264
rect 7285 105 7290 135
rect 7320 105 7325 135
rect 7285 100 7325 105
rect 11860 135 11900 953
rect 21240 658 21280 663
rect 21240 628 21245 658
rect 21275 628 21280 658
rect 11860 105 11865 135
rect 11895 105 11900 135
rect 11860 100 11900 105
rect 14715 125 14755 360
rect 21240 235 21280 628
rect 21925 588 21966 593
rect 21925 558 21930 588
rect 21960 558 21966 588
rect 21925 527 21966 558
rect 21925 495 21929 527
rect 21961 495 21966 527
rect 21925 488 21966 495
rect 21240 205 21245 235
rect 21275 205 21280 235
rect 21240 200 21280 205
rect 21925 296 21965 301
rect 21925 264 21929 296
rect 21961 264 21965 296
rect 14715 95 14720 125
rect 14750 95 14755 125
rect 14715 90 14755 95
rect 21925 125 21965 264
rect 21925 95 21930 125
rect 21960 95 21965 125
rect 21925 90 21965 95
<< via2 >>
rect 7289 495 7321 527
rect 7289 264 7321 296
rect 21929 495 21961 527
rect 21929 264 21961 296
<< metal3 >>
rect 7280 527 7330 536
rect 7280 495 7289 527
rect 7321 495 7330 527
rect 7280 296 7330 495
rect 7280 264 7289 296
rect 7321 264 7330 296
rect 7280 250 7330 264
rect 21920 527 21970 536
rect 21920 495 21929 527
rect 21961 495 21970 527
rect 21920 296 21970 495
rect 21920 264 21929 296
rect 21961 264 21970 296
rect 21920 250 21970 264
use 7bit_dac  X1
timestamp 1688567721
transform 1 0 0 0 1 0
box 0 300 14340 17455
use 7bit_dac  X2
timestamp 1688567721
transform 1 0 14640 0 1 0
box 0 300 14340 17455
use sw  X3
timestamp 1687966408
transform 1 0 13900 0 1 693
box 0 -393 860 360
<< labels >>
flabel metal1 132 16830 232 16930 0 FreeSans 128 0 0 0 vrefh
port 2 nsew
flabel metal1 28742 16852 28842 16952 0 FreeSans 128 0 0 0 vrefl
port 3 nsew
flabel metal1 1801 16953 1841 16993 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 1720 16262 1760 16302 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 950 16571 990 16611 0 FreeSans 128 0 0 0 d0
port 4 nsew
flabel metal1 2200 15145 2240 15185 0 FreeSans 128 0 0 0 d2
port 6 nsew
flabel metal1 2050 16118 2090 16158 0 FreeSans 128 0 0 0 d1
port 5 nsew
flabel metal1 14485 632 14525 672 0 FreeSans 128 0 0 0 vout
port 12 nsew
flabel metal1 13900 623 13940 663 0 FreeSans 128 0 0 0 d7
port 11 nsew
flabel metal1 2675 623 2715 663 0 FreeSans 128 0 0 0 d5
port 9 nsew
flabel metal1 6700 623 6740 663 0 FreeSans 128 0 0 0 d6
port 10 nsew
flabel metal1 2200 13259 2240 13299 0 FreeSans 128 0 0 0 d3
port 7 nsew
flabel metal1 2200 9447 2240 9487 0 FreeSans 128 0 0 0 d4
port 8 nsew
<< end >>
