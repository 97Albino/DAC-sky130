magic
tech sky130B
timestamp 1688392753
<< metal1 >>
rect 680 15424 4970 15500
rect 680 15348 756 15424
rect 4894 15348 4970 15424
rect 950 15304 990 15344
rect 1874 15335 4810 15348
rect 140 15200 240 15300
rect 1874 15285 4750 15335
rect 4800 15285 4810 15335
rect 1874 15272 4810 15285
rect 6781 15200 6881 15300
rect 950 14918 990 14958
rect 1720 14610 1760 14650
rect 2050 14465 2090 14505
rect 2200 13492 2240 13532
rect 2200 11606 2240 11646
rect 3280 11590 3855 11669
rect 3490 9642 3530 11590
rect 3320 9600 3700 9642
rect 3490 7835 3530 9600
rect 2200 7794 2240 7834
rect 2303 7799 2308 7829
rect 2338 7799 2343 7829
rect 3320 7793 3700 7835
rect 4679 7799 4684 7829
rect 4714 7799 4719 7829
rect 2786 7623 2791 7653
rect 2821 7623 2826 7653
rect 3490 5910 3530 7793
rect 4195 7623 4200 7653
rect 4230 7623 4235 7653
rect 3320 5868 3700 5910
rect 3490 4058 3530 5868
rect 3165 3979 3740 4058
rect 4005 773 4055 813
rect 2190 595 4970 600
rect 2190 565 2200 595
rect 2230 565 4935 595
rect 4965 565 4970 595
rect 2190 560 4970 565
rect 2210 363 5070 376
rect 2210 313 2220 363
rect 2270 313 5070 363
rect 2210 300 5070 313
rect 83 0 299 300
rect 680 200 756 300
rect 6264 200 6340 300
rect 680 185 6340 200
rect 680 142 3743 185
rect 3791 142 6340 185
rect 680 124 6340 142
rect 6721 0 6937 300
rect 83 -216 6937 0
rect 190 -285 6830 -280
rect 190 -315 195 -285
rect 225 -315 6795 -285
rect 6825 -315 6830 -285
rect 190 -320 6830 -315
rect 2207 -620 2676 -600
rect 2207 -660 2225 -620
rect 2265 -660 2676 -620
rect 2207 -676 2676 -660
rect 2675 -1030 2715 -990
rect 3260 -1030 3300 -990
rect 3500 -1293 3806 -1277
rect 3500 -1336 3744 -1293
rect 3792 -1336 3806 -1293
rect 3500 -1353 3806 -1336
<< via1 >>
rect 4750 15285 4800 15335
rect 2308 7799 2338 7829
rect 4684 7799 4714 7829
rect 2791 7623 2821 7653
rect 4200 7623 4230 7653
rect 2200 565 2230 595
rect 4935 565 4965 595
rect 2220 313 2270 363
rect 3743 142 3791 185
rect 195 -315 225 -285
rect 6795 -315 6825 -285
rect 2225 -660 2265 -620
rect 3744 -1336 3792 -1293
<< metal2 >>
rect 4740 15335 5070 15348
rect 4740 15285 4750 15335
rect 4800 15285 5070 15335
rect 4740 15272 5070 15285
rect 2461 7834 2493 7835
rect 2308 7830 2514 7834
rect 2308 7829 2461 7830
rect 2338 7799 2461 7829
rect 2308 7798 2461 7799
rect 2493 7798 2514 7830
rect 2308 7794 2514 7798
rect 4520 7830 4720 7835
rect 4520 7798 4527 7830
rect 4559 7829 4720 7830
rect 4559 7799 4684 7829
rect 4714 7799 4720 7829
rect 4559 7798 4720 7799
rect 2461 7793 2493 7794
rect 4520 7793 4720 7798
rect 2785 7654 2911 7659
rect 2785 7653 2874 7654
rect 2785 7623 2791 7653
rect 2821 7623 2874 7653
rect 2785 7622 2874 7623
rect 2906 7622 2911 7654
rect 2785 7617 2911 7622
rect 3425 7654 3465 7659
rect 3425 7622 3428 7654
rect 3460 7622 3465 7654
rect 190 623 990 663
rect 190 -285 230 623
rect 2050 600 2090 1123
rect 2050 595 2240 600
rect 2050 565 2200 595
rect 2230 565 2240 595
rect 2050 560 2240 565
rect 1874 363 2283 376
rect 1874 313 2220 363
rect 2270 313 2283 363
rect 1874 300 2283 313
rect 190 -315 195 -285
rect 225 -315 230 -285
rect 190 -320 230 -315
rect 2207 -620 2283 300
rect 2207 -660 2225 -620
rect 2265 -660 2283 -620
rect 2207 -676 2283 -660
rect 3425 -700 3465 7622
rect 3590 7654 3630 7660
rect 3590 7622 3595 7654
rect 3627 7622 3630 7654
rect 3590 -1253 3630 7622
rect 4136 7654 4235 7660
rect 4136 7622 4140 7654
rect 4172 7653 4235 7654
rect 4172 7623 4200 7653
rect 4230 7623 4235 7653
rect 4172 7622 4235 7623
rect 4136 7616 4235 7622
rect 4930 595 4970 1183
rect 4930 565 4935 595
rect 4965 565 4970 595
rect 4930 560 4970 565
rect 6030 540 6070 730
rect 6030 500 6830 540
rect 3530 -1293 3630 -1253
rect 3730 185 3806 200
rect 3730 142 3743 185
rect 3791 142 3806 185
rect 3730 -1293 3806 142
rect 6790 -285 6830 500
rect 6790 -315 6795 -285
rect 6825 -315 6830 -285
rect 6790 -320 6830 -315
rect 3730 -1336 3744 -1293
rect 3792 -1336 3806 -1293
rect 3730 -1353 3806 -1336
<< via2 >>
rect 2461 7798 2493 7830
rect 4527 7798 4559 7830
rect 2874 7622 2906 7654
rect 3428 7622 3460 7654
rect 3595 7622 3627 7654
rect 4140 7622 4172 7654
<< metal3 >>
rect 4770 13550 4780 13594
rect 4770 13534 4830 13550
rect 2195 13490 4830 13534
rect 2450 7830 4565 7835
rect 2450 7798 2461 7830
rect 2493 7798 4527 7830
rect 4559 7798 4565 7830
rect 2450 7793 4565 7798
rect 2867 7654 3465 7659
rect 2867 7622 2874 7654
rect 2906 7622 3428 7654
rect 3460 7622 3465 7654
rect 2867 7617 3465 7622
rect 3590 7654 4180 7660
rect 3590 7622 3595 7654
rect 3627 7622 4140 7654
rect 4172 7622 4180 7654
rect 3590 7616 4180 7622
rect 4780 2098 4830 2158
rect 2197 2054 4830 2098
use 5bit_dac  X1
timestamp 1688377021
transform 1 0 -400 0 1 7924
box 400 -7624 3720 7424
use 5bit_dac  X2
timestamp 1688377021
transform -1 0 7420 0 -1 7724
box 400 -7624 3720 7424
use sw  X3
timestamp 1687966408
transform 1 0 2675 0 1 -960
box 0 -393 860 360
<< labels >>
flabel metal1 140 15200 240 15300 0 FreeSans 128 0 0 0 vrefh
port 2 nsew
flabel metal1 6781 15200 6881 15300 0 FreeSans 128 0 0 0 vrefl
port 3 nsew
flabel metal1 950 15304 990 15344 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 1720 14610 1760 14650 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 950 14918 990 14958 0 FreeSans 128 0 0 0 d0
port 4 nsew
flabel metal1 2050 14465 2090 14505 0 FreeSans 128 0 0 0 d1
port 5 nsew
flabel metal1 2200 13492 2240 13532 0 FreeSans 128 0 0 0 d2
port 6 nsew
flabel metal1 2200 11606 2240 11646 0 FreeSans 128 0 0 0 d3
port 7 nsew
flabel metal1 2200 7794 2240 7834 0 FreeSans 128 0 0 0 d4
port 8 nsew
flabel metal1 2675 -1030 2715 -990 0 FreeSans 128 0 0 0 d5
port 9 nsew
flabel metal1 3260 -1030 3300 -990 0 FreeSans 128 0 0 0 vout
port 10 nsew
<< end >>
