* SPICE3 file created from 8bit_DAC.ext - technology: sky130A

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/corners/tt.spice
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice


X0 a_16814_1579# a_16601_1579# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1 gnd d0 a_4079_2968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_854_4021# a_1585_4331# a_1793_4331# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X3 a_11512_7066# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 a_17975_3271# a_18959_3568# a_18914_3581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X5 a_17970_4551# a_18957_4117# a_18912_4130# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X6 a_14985_138# a_16769_199# a_16989_4907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X7 a_16879_6583# a_16458_6583# a_15940_6273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_7939_5649# a_8196_5459# a_7798_6241# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X9 a_5704_753# a_5491_753# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X10 vdd d2 a_8056_3845# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X11 a_8879_2650# a_9136_2460# a_7944_2163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X12 a_14876_138# a_14663_138# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X13 a_7938_7855# a_8925_7421# a_8880_7434# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X14 a_16457_8789# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 a_1371_6537# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 a_3827_775# a_4080_762# a_2885_1196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X17 gnd a_13062_2693# a_12854_2693# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X18 a_856_3472# a_435_3472# a_119_3353# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X19 a_10148_8186# a_10148_7999# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X20 vdd d1 a_13173_1011# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X21 a_6643_1063# a_6430_1063# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X22 a_17974_4374# a_18958_4671# a_18909_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X23 a_1808_7180# a_1694_7061# a_1808_4980# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 a_433_4021# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X25 a_10678_4580# a_10465_4580# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X26 a_5911_2959# a_5490_2959# a_5175_3164# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X27 a_432_7330# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X28 a_17973_6580# a_18957_6877# a_18908_7067# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X29 a_10149_4690# a_10678_4580# a_10886_4580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X30 a_647_4575# a_434_4575# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X31 a_7803_3858# a_7988_4356# a_7943_4369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X32 gnd a_4077_7380# a_3869_7380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X33 a_6570_1574# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X34 a_3824_1506# a_4081_1316# a_2889_1019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X35 a_15205_4731# a_15205_4502# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X36 a_5174_4913# a_5174_4726# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X37 a_10465_5683# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X38 a_120_1563# a_647_1815# a_855_1815# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X39 gnd d2 a_18088_1644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X40 vdd a_3000_3804# a_2792_3804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X41 gnd d4 a_8087_4929# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X42 gnd d1 a_13172_2114# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X43 a_10149_5334# a_10677_5129# a_10885_5129# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X44 vdd a_14107_8488# a_13899_8488# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X45 a_5491_753# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X46 a_11824_5439# a_11756_5950# a_11834_7066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X47 a_6640_6578# a_6427_6578# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X48 a_13858_780# a_14111_767# a_12916_1201# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X49 a_18910_8542# a_19163_8529# a_17968_8963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X50 a_10148_6667# a_10148_6437# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X51 a_10147_8873# a_10676_8992# a_10884_8992# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X52 a_15942_2964# a_15521_2964# a_15206_2712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X53 a_6641_5475# a_6428_5475# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X54 a_6429_3269# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X55 a_13852_5369# a_14109_5179# a_12914_5613# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X56 a_10149_5564# a_10149_5334# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X57 a_16460_2171# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X58 a_119_3582# a_119_3353# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X59 a_10675_8438# a_10462_8438# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X60 a_10678_4580# a_10465_4580# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X61 a_17969_7860# a_18226_7670# a_17828_8452# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X62 a_18908_5410# a_19165_5220# a_17970_5654# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X63 a_5910_5165# a_5489_5165# a_5174_5370# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X64 a_13853_2060# a_14110_1870# a_12915_2304# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X65 a_13855_1511# a_14112_1321# a_12920_1024# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X66 a_5488_9028# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X67 a_6427_6578# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X68 a_3825_7947# a_3821_8124# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X69 a_10884_6232# a_10463_6232# a_10149_5980# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X70 a_17828_8452# a_18085_8262# a_17863_7159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X71 a_12918_5436# a_13171_5423# a_12773_6205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 a_432_8987# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X73 a_5489_7925# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X74 a_6861_2690# a_6752_2690# a_6859_4902# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X75 a_6428_5475# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X76 a_119_2020# a_647_1815# a_855_1815# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X77 gnd a_4077_9037# a_3869_9037# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X78 a_12777_6028# a_13030_6015# a_12803_7295# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X79 a_6864_7221# a_6750_7102# a_6864_5021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X80 vdd a_13032_1603# a_12824_1603# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X81 a_15940_6273# a_15519_6273# a_15205_6021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X82 a_11614_8748# a_11401_8748# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X83 a_10462_8438# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X84 gnd a_18088_1644# a_17880_1644# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X85 a_15205_4272# a_15206_3815# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X86 a_17971_3448# a_18228_3258# a_17830_4040# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X87 a_15735_3518# a_15522_3518# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X88 a_646_5124# a_433_5124# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X89 a_5704_2410# a_5491_2410# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X90 a_1725_5945# a_1512_5945# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X91 gnd a_9133_7421# a_8925_7421# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_7944_3266# a_8197_3253# a_7799_4035# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X93 a_17829_6246# a_18019_5464# a_17974_5477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X94 a_1586_2125# a_1373_2125# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X95 a_645_8987# a_432_8987# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X96 a_16670_8789# a_16457_8789# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X97 a_17969_6757# a_18956_6323# a_18911_6336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X98 vdd a_9135_1906# a_8927_1906# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X99 a_15733_6827# a_15520_6827# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X100 a_12777_6028# a_12962_6526# a_12913_6716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X101 a_13852_7026# a_14109_6836# a_12917_6539# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X102 a_16879_6583# a_16458_6583# a_15941_6827# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X103 a_5910_5165# a_5489_5165# a_5174_4913# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X104 a_8880_6331# a_9133_6318# a_7938_6752# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X105 a_15206_3815# a_15733_4067# a_15941_4067# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X106 a_6752_2690# a_6539_2690# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X107 a_1512_5945# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X108 vdd d1 a_3138_8727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X109 a_116_8638# a_644_8433# a_852_8433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X110 a_8881_5228# a_9134_5215# a_7939_5649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X111 a_5911_4616# a_5490_4616# a_5174_4497# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X112 a_10888_1271# a_10467_1271# a_10151_1381# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X113 a_14876_138# a_14663_138# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X114 a_1371_6537# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X115 a_16457_8789# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X116 a_3824_7393# a_3820_7570# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X117 a_17861_2924# a_17880_1644# a_17831_1834# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X118 a_16671_7686# a_16458_7686# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X119 a_18914_2478# a_18910_2655# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X120 a_431_8433# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X121 a_11617_2130# a_11404_2130# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X122 a_13850_8678# a_13856_7952# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X123 a_15206_3399# a_15735_3518# a_15943_3518# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X124 a_2886_7637# a_3870_7934# a_3825_7947# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X125 gnd d1 a_3139_6521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X126 a_1586_2125# a_1373_2125# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X127 a_7940_2340# a_8927_1906# a_8882_1919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X128 a_5491_2410# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X129 a_15207_963# a_15735_758# a_15943_758# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 a_3822_2055# a_3828_1329# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X131 gnd a_9133_9078# a_8925_9078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X132 a_6641_5475# a_6428_5475# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X133 a_16458_7686# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X134 a_10465_5683# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X135 a_1808_4980# a_1481_7061# a_1808_7180# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X136 a_6539_2690# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X137 a_15733_4067# a_15520_4067# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X138 a_16881_3274# a_16460_3274# a_15943_3518# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X139 vdd a_18118_2734# a_17910_2734# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X140 gnd d4 a_18118_4934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X141 a_5910_6822# a_5489_6822# a_5173_6703# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X142 a_7802_6064# a_7987_6562# a_7942_6575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X143 a_15944_1312# a_16674_1068# a_16882_1068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X144 a_12134_158# a_11713_158# a_12035_158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X145 a_10465_1820# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X146 vdd a_4080_3522# a_3872_3522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X147 a_10887_3477# a_11617_3233# a_11825_3233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X148 a_10150_3587# a_10679_3477# a_10887_3477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X149 a_5489_7925# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X150 a_6428_5475# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X151 a_2778_4901# a_3031_4888# a_2004_153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X152 vdd d2 a_18086_6056# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X153 a_8877_8165# a_8880_7434# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X154 a_11617_2130# a_11404_2130# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X155 a_1372_4331# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X156 a_8880_1547# a_8883_816# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X157 a_5172_8679# a_5700_8474# a_5908_8474# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X158 vdd d0 a_9133_6318# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X159 a_13853_2060# a_13859_1334# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X160 a_2774_5078# a_3031_4888# a_2004_153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X161 gnd d0 a_9135_3009# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X162 a_5704_2410# a_5491_2410# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X163 a_15941_5170# a_15520_5170# a_15205_5375# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X164 gnd a_3139_7624# a_2931_7624# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X165 a_10884_6232# a_10463_6232# a_10148_6437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X166 gnd a_4078_5174# a_3870_5174# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X167 gnd d1 a_8196_5459# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X168 a_18911_7439# a_19164_7426# a_17969_7860# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X169 gnd a_18229_1052# a_18021_1052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X170 gnd a_4079_4625# a_3871_4625# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X171 gnd d2 a_13030_6015# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X172 a_11544_3744# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X173 a_1792_6537# a_1725_5945# a_1803_7061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X174 vdd d1 a_18228_2155# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X175 a_3827_2432# a_4080_2419# a_2888_2122# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X176 vdd a_13029_8221# a_12821_8221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X177 a_18910_998# a_19167_808# a_17972_1242# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X178 a_17861_5124# a_17910_2734# a_17865_2747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X179 a_855_5678# a_434_5678# a_118_5788# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X180 a_7942_7678# a_8926_7975# a_8881_7988# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X181 gnd d1 a_8195_6562# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X182 a_119_3353# a_119_3123# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X183 vdd a_14111_3527# a_13903_3527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X184 a_2888_3225# a_3872_3522# a_3827_3535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X185 a_854_5124# a_1585_5434# a_1793_5434# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X186 a_16895_7226# a_16781_7107# a_16895_5026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X187 a_10467_1271# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X188 a_8883_816# a_9136_803# a_7941_1237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X189 a_10465_1820# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X190 a_10676_7335# a_10463_7335# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X191 a_11755_8156# a_11542_8156# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X192 a_6861_2690# a_6570_1574# a_6851_1063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X193 a_11933_4866# a_11512_4866# a_11834_4866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X194 a_12807_7118# a_13060_7105# a_12809_4906# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X195 a_854_4021# a_433_4021# a_118_4226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X196 a_8876_6508# a_8882_5782# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X197 a_855_2918# a_1586_3228# a_1794_3228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X198 gnd a_8196_5459# a_7988_5459# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X199 a_6864_5021# a_6537_7102# a_6864_7221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X200 a_11403_4336# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X201 gnd a_8055_6051# a_7847_6051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X202 a_117_7078# a_645_7330# a_853_7330# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X203 a_18915_1375# a_18911_1552# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X204 a_12805_5083# a_13062_4893# a_12035_158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X205 gnd a_8195_6562# a_7987_6562# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X206 a_6850_2166# a_6429_2166# a_5911_1856# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X207 a_15941_5170# a_15520_5170# a_15205_4918# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X208 a_10463_7335# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X209 gnd a_14110_4630# a_13902_4630# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X210 a_16890_7107# a_16599_5991# a_16879_6583# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X211 a_2887_4328# a_3871_4625# a_3822_4815# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X212 a_5491_2410# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X213 a_12774_3999# a_13031_3809# a_12809_2706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X214 a_13858_2437# a_14111_2424# a_12919_2127# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X215 a_7834_4942# a_8087_4929# a_7060_194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X216 a_1694_7061# a_1481_7061# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X217 a_10149_5793# a_10678_5683# a_10886_5683# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X218 vdd a_14108_9042# a_13900_9042# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X219 a_16460_3274# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X220 a_16671_7686# a_16458_7686# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X221 a_3825_6844# a_4078_6831# a_2886_6534# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X222 a_12919_3230# a_13903_3527# a_13858_3540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X223 gnd a_19164_9083# a_17972_8786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X224 a_2776_7113# a_2790_8216# a_2745_8229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X225 a_10885_6786# a_11615_6542# a_11823_6542# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X226 vout a_9566_17# a_9888_17# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X227 a_18910_2655# a_19167_2465# a_17975_2168# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X228 a_7798_6241# a_8055_6051# a_7828_7331# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X229 a_16890_4907# a_16570_2695# a_16892_2695# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X230 a_7803_3858# a_8056_3845# a_7834_2742# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X231 a_2103_153# a_1682_153# a_2004_153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X232 a_17974_4374# a_18227_4361# a_17834_3863# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X233 vdd d0 a_4079_2968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X234 gnd a_19167_3568# a_18959_3568# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X235 a_1902_4861# a_1481_4861# a_1808_4980# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X236 a_2742_6200# a_2999_6010# a_2772_7290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X237 a_10676_8992# a_10463_8992# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X238 a_6848_6578# a_6781_5986# a_6859_7102# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X239 a_117_7535# a_645_7330# a_853_7330# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X240 a_5911_5719# a_5490_5719# a_5174_5829# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X241 a_12912_8922# a_13899_8488# a_13854_8501# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X242 a_16674_1068# a_16461_1068# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X243 a_18909_5964# a_19166_5774# a_17974_5477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X244 a_16458_7686# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X245 a_17865_4947# a_17908_7146# a_17859_7336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 a_12918_4333# a_13902_4630# a_13853_4820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X247 a_16601_1579# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X248 a_11834_7066# a_11725_7066# a_11839_4985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X249 a_8881_6885# a_8877_7062# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X250 a_15941_6827# a_15520_6827# a_15204_6708# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X251 a_10886_2923# a_11617_3233# a_11825_3233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X252 a_10463_8992# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X253 a_12917_7642# a_13901_7939# a_13852_8129# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X254 a_10149_4690# a_10149_4461# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X255 gnd d4 a_3031_4888# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X256 a_18906_8719# a_18912_7993# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X257 a_647_5678# a_434_5678# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X258 gnd a_9134_7975# a_8926_7975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X259 gnd a_3000_3804# a_2792_3804# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X260 a_18907_7616# a_18912_6890# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X261 a_15522_758# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X262 a_17973_6580# a_18957_6877# a_18912_6890# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X263 a_5175_2291# a_5175_2061# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X264 a_1372_4331# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X265 gnd a_14107_8488# a_13899_8488# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X266 a_2884_3402# a_3141_3212# a_2743_3994# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X267 a_15203_8684# a_15731_8479# a_15939_8479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X268 a_10886_2923# a_10465_2923# a_10150_2671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X269 a_7834_2742# a_7848_3845# a_7803_3858# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X270 a_8881_6885# a_9134_6872# a_7942_6575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X271 a_5175_2520# a_5175_2291# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X272 a_11544_3744# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X273 a_116_9097# a_645_8987# a_853_8987# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X274 a_2881_8917# a_3138_8727# a_2745_8229# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X275 a_3820_6467# a_4077_6277# a_2882_6711# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X276 a_10675_8438# a_10462_8438# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X277 gnd d1 a_18226_6567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X278 a_433_5124# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X279 a_12916_8745# a_13169_8732# a_12776_8234# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X280 a_13855_6295# a_14108_6282# a_12913_6716# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X281 a_5173_7576# a_5701_7371# a_5909_7371# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X282 a_5176_1417# a_5705_1307# a_5913_1307# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X283 a_432_8987# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X284 gnd d1 a_8197_2150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X285 a_5172_8909# a_5172_8679# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X286 a_16878_8789# a_16811_8197# a_16895_7226# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X287 a_11403_4336# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X288 a_5173_8035# a_5173_7806# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X289 a_17972_8786# a_18225_8773# a_17832_8275# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X290 a_644_8433# a_431_8433# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X291 a_16895_5026# a_16568_7107# a_16895_7226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X292 a_12913_6716# a_13170_6526# a_12777_6028# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X293 gnd a_13032_1603# a_12824_1603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X294 a_10149_4231# a_10150_3774# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X295 gnd a_18086_6056# a_17878_6056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X296 a_10462_8438# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X297 a_12915_3407# a_13172_3217# a_12774_3999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X298 a_5911_4616# a_6641_4372# a_6849_4372# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X299 a_13855_9055# a_13851_9232# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X300 a_17975_3271# a_18228_3258# a_17830_4040# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X301 a_12914_5613# a_13171_5423# a_12773_6205# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X302 gnd a_18226_6567# a_18018_6567# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X303 vdd a_19166_1911# a_18958_1911# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X304 a_3827_2432# a_3823_2609# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X305 a_1481_7061# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X306 vdd a_9132_8524# a_8924_8524# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X307 a_12913_7819# a_13900_7385# a_13855_7398# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X308 a_10149_5564# a_10678_5683# a_10886_5683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X309 gnd d1 a_3142_1006# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X310 a_8877_5405# a_8882_4679# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X311 a_10884_6232# a_11615_6542# a_11823_6542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X312 a_3826_5741# a_3822_5918# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X313 a_5175_2061# a_5176_1604# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X314 a_11823_7645# a_11402_7645# a_10885_7889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X315 a_18913_1924# a_19166_1911# a_17971_2345# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X316 a_18915_1375# a_19168_1362# a_17976_1065# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X317 vdd d0 a_9136_3563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X318 vdd d0 a_9134_4112# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X319 vdd a_3029_7100# a_2821_7100# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X320 a_648_3472# a_435_3472# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X321 a_10150_3774# a_10677_4026# a_10885_4026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X322 a_5705_1307# a_5492_1307# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X323 a_646_4021# a_433_4021# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X324 a_117_8181# a_644_8433# a_852_8433# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X325 a_648_712# a_435_712# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X326 a_17829_6246# a_18086_6056# a_17859_7336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X327 a_8876_6508# a_9133_6318# a_7938_6752# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X328 a_7937_8958# a_8194_8768# a_7801_8270# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X329 a_16568_7107# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X330 a_7830_5119# a_8087_4929# a_7060_194# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X331 gnd d0 a_4078_7934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X332 a_15942_5724# a_15521_5724# a_15205_5834# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X333 a_8880_1547# a_9137_1357# a_7945_1060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X334 a_7943_5472# a_8196_5459# a_7798_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X335 gnd a_4079_5728# a_3871_5728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_15522_2415# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X337 a_13858_2437# a_13854_2614# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X338 a_5173_7576# a_5173_7119# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X339 a_17971_2345# a_18958_1911# a_18913_1924# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X340 a_5176_1604# a_5703_1856# a_5911_1856# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X341 vdd a_8197_3253# a_7989_3253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X342 gnd d0 a_9135_4666# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X343 a_11615_6542# a_11402_6542# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X344 a_1682_153# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X345 gnd d3 a_18118_2734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X346 a_7800_1829# a_8057_1639# a_7830_2919# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X347 a_7942_6575# a_8195_6562# a_7802_6064# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X348 a_10679_3477# a_10466_3477# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X349 a_10677_4026# a_10464_4026# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X350 a_10149_4877# a_10149_4690# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X351 a_7799_4035# a_7989_3253# a_7944_3266# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X352 a_11756_5950# a_11543_5950# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X353 a_3823_952# a_4080_762# a_2885_1196# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X354 a_10679_717# a_10466_717# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X355 a_11834_4866# a_11725_4866# a_11933_4866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X356 a_3825_5187# a_3821_5364# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X357 a_6537_7102# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X358 a_116_9097# a_116_8868# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X359 a_434_1815# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X360 a_11402_6542# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X361 a_122_818# a_648_712# a_856_712# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X362 gnd d0 a_4080_3522# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X363 a_1810_2768# a_1696_2649# a_1803_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X364 a_648_2369# a_435_2369# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X365 a_8882_5782# a_8878_5959# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X366 gnd d1 a_13173_1011# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X367 a_18911_1552# a_18914_821# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X368 gnd a_3141_3212# a_2933_3212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X369 vdd a_8085_7141# a_7877_7141# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X370 a_5703_1856# a_5490_1856# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X371 a_6568_5986# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X372 a_15520_7930# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X373 a_13857_1883# a_13853_2060# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X374 gnd a_14108_7385# a_13900_7385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X375 vdd d0 a_4079_4625# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X376 a_15204_7581# a_15732_7376# a_15940_7376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X377 vdd d4 a_3031_4888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X378 a_16879_7686# a_16811_8197# a_16895_7226# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X379 vdd d1 a_13172_2114# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X380 gnd a_9135_5769# a_8927_5769# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X381 a_5908_8474# a_5487_8474# a_5172_8679# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X382 a_6642_2166# a_6429_2166# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X383 vdd a_3140_4315# a_2932_4315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X384 a_15203_8914# a_15203_8684# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X385 a_18906_8719# a_19163_8529# a_17968_8963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X386 a_18914_821# a_19167_808# a_17972_1242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X387 a_13854_957# a_14111_767# a_12916_1201# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X388 a_11725_4866# a_11512_4866# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X389 a_15204_8040# a_15204_7811# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X390 vdd d0 a_4077_7380# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X391 a_16892_2695# a_16601_1579# a_16882_1068# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X392 a_5909_7371# a_5488_7371# a_5173_7576# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X393 a_5912_3513# a_5491_3513# a_5175_3623# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X394 a_434_1815# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X395 vdd d2 a_3000_3804# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X396 a_5910_4062# a_5489_4062# a_5174_4267# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X397 a_5490_5719# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X398 a_10679_2374# a_10466_2374# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X399 gnd d0 a_19166_3014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X400 a_5912_753# a_5491_753# a_5178_859# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 a_3823_2609# a_4080_2419# a_2888_2122# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X402 a_2743_3994# a_2933_3212# a_2884_3402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X403 a_2887_4328# a_3140_4315# a_2747_3817# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X404 a_119_2250# a_648_2369# a_856_2369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X405 a_1587_1022# a_1374_1022# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X406 a_5492_1307# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X407 a_5490_1856# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X408 a_18912_5233# a_19165_5220# a_17970_5654# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X409 a_17973_7683# a_18226_7670# a_17828_8452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X410 a_15522_2415# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X411 a_1724_8151# a_1511_8151# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X412 vdd a_9136_803# a_8928_803# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X413 a_2776_7113# a_3029_7100# a_2778_4901# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X414 a_855_2918# a_434_2918# a_119_3123# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X415 a_3827_775# a_3823_952# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X416 a_12778_3822# a_13031_3809# a_12809_2706# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 vdd a_13171_4320# a_12963_4320# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X418 a_2747_3817# a_2932_4315# a_2887_4328# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X419 a_11841_2773# a_11727_2654# a_11834_4866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X420 a_6428_4372# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X421 gnd a_14108_9042# a_13900_9042# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X422 a_18912_7993# a_18908_8170# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X423 a_17833_6069# a_18018_6567# a_17969_6757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X424 vdd d2 a_13031_3809# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X425 a_13854_2614# a_14111_2424# a_12919_2127# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X426 a_10677_5129# a_10464_5129# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X427 gnd d2 a_8055_6051# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X428 a_12774_3999# a_12964_3217# a_12915_3407# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X429 a_11756_5950# a_11543_5950# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X430 a_12918_4333# a_13171_4320# a_12778_3822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X431 gnd a_8196_4356# a_7988_4356# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X432 a_1791_8743# a_1370_8743# a_852_8433# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X433 a_15204_7581# a_15204_7124# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X434 a_10676_8992# a_10463_8992# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X435 a_11615_6542# a_11402_6542# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X436 a_6849_5475# a_6781_5986# a_6859_7102# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X437 a_5172_9138# a_5701_9028# a_5909_9028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X438 a_5910_6822# a_6640_6578# a_6848_6578# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X439 a_11618_1027# a_11405_1027# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X440 a_12912_8922# a_13899_8488# a_13850_8678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X441 a_1373_3228# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X442 a_434_5678# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X443 a_7941_1237# a_8928_803# a_8883_816# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X444 a_5489_4062# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X445 a_5911_5719# a_6641_5475# a_6849_5475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X446 a_5173_8035# a_5702_7925# a_5910_7925# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X447 a_13852_8129# a_13855_7398# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X448 a_17835_1657# a_18020_2155# a_17975_2168# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X449 a_13858_780# a_13854_957# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X450 a_10464_5129# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X451 a_12778_3822# a_12963_4320# a_12918_4333# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X452 a_11727_2654# a_11514_2654# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X453 a_15520_7930# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X454 vdd a_9136_2460# a_8928_2460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X455 a_10463_8992# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X456 a_11402_6542# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X457 a_10885_7889# a_10464_7889# a_10148_7770# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X458 a_1805_2649# a_1696_2649# a_1803_4861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X459 gnd a_4080_762# a_3872_762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X460 a_855_4575# a_434_4575# a_118_4685# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X461 a_6750_7102# a_6537_7102# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X462 a_8883_2473# a_8879_2650# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X463 a_10466_717# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X464 vdd a_9133_9078# a_8925_9078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X465 a_18911_7439# a_18907_7616# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X466 a_8883_2473# a_9136_2460# a_7944_2163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X467 a_17865_2747# a_17879_3850# a_17834_3863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X468 a_7938_7855# a_8925_7421# a_8876_7611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X469 a_16599_5991# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X470 a_116_8868# a_116_8638# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X471 vdd d0 a_14108_7385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X472 a_118_5329# a_646_5124# a_854_5124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X473 a_117_7994# a_117_7765# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X474 vdd a_4081_1316# a_3873_1316# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X475 vdd a_4079_1865# a_3871_1865# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X476 a_13851_6472# a_13857_5746# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X477 a_116_8868# a_645_8987# a_853_8987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X478 a_6537_4902# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X479 a_5175_2707# a_5175_2520# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X480 vdd d0 a_19164_7426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X481 a_6851_1063# a_6430_1063# a_5913_1307# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X482 a_15939_8479# a_15518_8479# a_15203_8684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X483 a_15205_4502# a_15734_4621# a_15942_4621# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X484 a_6847_8784# a_6426_8784# a_5908_8474# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X485 gnd a_4076_8483# a_3868_8483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X486 a_9779_17# a_9566_17# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X487 a_7944_2163# a_8928_2460# a_8883_2473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X488 a_8877_7062# a_9134_6872# a_7942_6575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X489 a_5175_3164# a_5703_2959# a_5911_2959# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X490 a_15206_2066# a_15734_1861# a_15942_1861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X491 a_15207_1422# a_15736_1312# a_15944_1312# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X492 gnd d1 a_13170_7629# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X493 a_3828_1329# a_4081_1316# a_2889_1019# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X494 a_2885_1196# a_3872_762# a_3823_952# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X495 gnd a_14111_767# a_13903_767# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X496 gnd d0 a_14109_5179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X497 a_855_4575# a_434_4575# a_118_4456# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X498 a_5176_1417# a_5176_1188# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X499 a_15734_4621# a_15521_4621# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X500 a_12809_4906# a_13062_4893# a_12035_158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X501 a_853_6227# a_432_6227# a_118_5975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X502 a_644_8433# a_431_8433# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X503 a_16880_4377# a_16459_4377# a_15942_4621# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X504 a_5173_8222# a_5173_8035# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X505 a_15734_1861# a_15521_1861# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X506 vdd a_3139_7624# a_2931_7624# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X507 vdd a_4078_5174# a_3870_5174# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X508 vdd a_19164_7426# a_18956_7426# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X509 a_10466_2374# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X510 a_8882_1919# a_8878_2096# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X511 a_10886_4580# a_11616_4336# a_11824_4336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X512 vdd a_14110_1870# a_13902_1870# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X513 a_2889_1019# a_3873_1316# a_3828_1329# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X514 a_2884_2299# a_3871_1865# a_3826_1878# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X515 gnd a_13170_7629# a_12962_7629# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X516 vdd d1 a_18229_1052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X517 gnd a_14109_5179# a_13901_5179# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X518 a_7941_8781# a_8925_9078# a_8876_9268# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X519 vdd d1 a_8195_6562# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X520 gnd a_13029_8221# a_12821_8221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X521 a_2882_6711# a_3139_6521# a_2746_6023# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X522 a_8879_2650# a_8882_1919# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X523 a_117_7535# a_117_7078# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X524 a_5703_2959# a_5490_2959# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X525 a_10147_8643# a_10148_8186# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X526 a_13859_1334# a_14112_1321# a_12920_1024# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X527 a_12916_1201# a_13903_767# a_13854_957# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X528 a_5910_5165# a_6641_5475# a_6849_5475# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X529 a_5173_7806# a_5702_7925# a_5910_7925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X530 a_13857_1883# a_14110_1870# a_12915_2304# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X531 a_15943_3518# a_15522_3518# a_15206_3399# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X532 a_15941_4067# a_15520_4067# a_15206_3815# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X533 a_1791_8743# a_1370_8743# a_853_8987# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X534 gnd a_18228_2155# a_18020_2155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X535 a_1794_2125# a_1373_2125# a_856_2369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X536 a_17861_5124# a_18118_4934# a_17091_199# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X537 a_2882_7814# a_3869_7380# a_3824_7393# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X538 a_13856_6849# a_13852_7026# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X539 a_118_4685# a_118_4456# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X540 vdd a_8195_6562# a_7987_6562# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X541 a_18911_1552# a_19168_1362# a_17976_1065# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X542 a_6642_3269# a_6429_3269# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X543 a_15203_9143# a_15732_9033# a_15940_9033# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X544 a_15941_6827# a_16671_6583# a_16879_6583# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X545 a_12915_2304# a_13902_1870# a_13857_1883# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X546 a_12920_1024# a_13904_1321# a_13859_1334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X547 a_3824_1506# a_3827_775# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X548 a_5700_8474# a_5487_8474# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X549 a_7797_8447# a_8054_8257# a_7832_7154# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X550 a_15204_8040# a_15733_7930# a_15941_7930# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X551 a_15942_5724# a_16672_5480# a_16880_5480# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X552 vdd a_4078_6831# a_3870_6831# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X553 vdd d0 a_9134_7975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X554 a_5909_9028# a_5488_9028# a_5172_9138# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X555 gnd a_8197_3253# a_7989_3253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X556 a_18907_9273# a_19164_9083# a_17972_8786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X557 a_5487_8474# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X558 a_2741_8406# a_2931_7624# a_2882_7814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X559 a_2883_5608# a_3870_5174# a_3821_5364# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X560 vdd d0 a_4078_7934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X561 a_7804_1652# a_8057_1639# a_7830_2919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X562 a_1792_7640# a_1371_7640# a_853_7330# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X563 vdd d1 a_8196_4356# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X564 a_5909_6268# a_5488_6268# a_5174_6016# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X565 a_1725_5945# a_1512_5945# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X566 a_3820_9227# a_3823_8496# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X567 a_2776_7113# a_2790_8216# a_2741_8406# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X568 a_5488_7371# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X569 a_13856_6849# a_14109_6836# a_12917_6539# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X570 a_6958_4902# a_6951_194# a_4954_133# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X571 a_12807_7118# a_12821_8221# a_12776_8234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X572 vdd a_9134_5215# a_8926_5215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X573 a_1808_7180# a_1511_8151# a_1792_7640# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X574 a_16882_1068# a_16814_1579# a_16892_2695# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X575 a_15942_1861# a_16673_2171# a_16881_2171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X576 vdd a_19167_3568# a_18959_3568# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X577 a_5490_2959# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X578 a_7799_4035# a_7989_3253# a_7940_3443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X579 a_16781_7107# a_16568_7107# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X580 a_7943_4369# a_8196_4356# a_7803_3858# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X581 a_2746_6023# a_2999_6010# a_2772_7290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X582 a_18912_6890# a_19165_6877# a_17973_6580# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X583 a_1584_6537# a_1371_6537# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X584 a_1805_2649# a_1514_1533# a_1795_1022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X585 a_5178_859# a_5704_753# a_5912_753# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X586 a_1794_2125# a_1373_2125# a_855_1815# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X587 a_1512_5945# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X588 a_13855_1511# a_13858_780# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X589 a_5911_2959# a_6642_3269# a_6850_3269# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X590 a_16881_3274# a_16813_3785# a_16897_2814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X591 a_13855_6295# a_13851_6472# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X592 a_8880_9091# a_10147_9102# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X593 a_118_4226# a_119_3769# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X594 a_6568_5986# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X595 a_6847_8784# a_6426_8784# a_5909_9028# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X596 a_854_5124# a_433_5124# a_118_5329# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X597 a_16673_2171# a_16460_2171# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X598 a_10678_5683# a_10465_5683# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X599 a_12916_8745# a_13900_9042# a_13855_9055# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X600 vdd d0 a_14107_8488# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X601 a_11836_2654# a_11545_1538# a_11826_1027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X602 a_6569_3780# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X603 vdd a_2998_8216# a_2790_8216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X604 a_15204_8227# a_15204_8040# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X605 gnd d2 a_3000_3804# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X606 vdd a_3031_4888# a_2823_4888# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X607 gnd d0 a_14110_2973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X608 a_10148_6437# a_10676_6232# a_10884_6232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X609 a_10885_4026# a_11616_4336# a_11824_4336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X610 a_6848_7681# a_6427_7681# a_5909_7371# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X611 a_6781_5986# a_6568_5986# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X612 a_10150_3128# a_10150_2671# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X613 a_16813_3785# a_16600_3785# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X614 a_10148_6896# a_10148_6667# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X615 vdd d1 a_18226_6567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X616 a_15521_1861# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X617 a_15523_1312# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X618 a_12912_8922# a_13169_8732# a_12776_8234# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X619 gnd a_4080_2419# a_3872_2419# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X620 a_13851_6472# a_14108_6282# a_12913_6716# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X621 a_435_3472# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X622 a_16882_1068# a_16461_1068# a_15943_758# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X623 gnd a_9136_803# a_8928_803# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X624 a_435_712# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X625 a_10887_3477# a_10466_3477# a_10150_3358# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X626 a_15521_5724# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X627 a_15204_7811# a_15733_7930# a_15941_7930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X628 a_15941_5170# a_16672_5480# a_16880_5480# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X629 a_11725_7066# a_11512_7066# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X630 vdd d0 a_14109_4076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X631 a_16459_4377# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X632 a_17968_8963# a_18225_8773# a_17832_8275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X633 a_12917_6539# a_13170_6526# a_12777_6028# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X634 a_7942_7678# a_8926_7975# a_8877_8165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X635 a_15203_8914# a_15732_9033# a_15940_9033# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X636 a_15940_6273# a_16671_6583# a_16879_6583# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X637 vdd a_18226_6567# a_18018_6567# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X638 a_6569_3780# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X639 gnd d2 a_13031_3809# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X640 a_118_4872# a_118_4685# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X641 a_2004_153# a_2823_4888# a_2778_4901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X642 a_118_5788# a_647_5678# a_855_5678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X643 a_854_6781# a_1584_6537# a_1792_6537# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X644 a_645_6227# a_432_6227# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X645 a_15731_8479# a_15518_8479# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X646 vdd d0 a_9135_1906# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X647 a_5175_2520# a_5704_2410# a_5912_2410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X648 a_11512_7066# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X649 a_10151_1568# a_10678_1820# a_10886_1820# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X650 a_647_1815# a_434_1815# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X651 vdd a_13031_3809# a_12823_3809# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X652 a_2778_2701# a_2792_3804# a_2747_3817# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X653 vdd d0 a_19165_7980# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X654 gnd a_14111_2424# a_13903_2424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X655 a_2888_2122# a_3872_2419# a_3823_2609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X656 a_17972_1242# a_18959_808# a_18914_821# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X657 a_7060_194# a_6951_194# a_4954_133# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X658 a_13857_5746# a_13853_5923# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X659 a_8884_1370# a_9137_1357# a_7945_1060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X660 a_7941_1237# a_8928_803# a_8879_993# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X661 a_8878_3199# a_8883_2473# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X662 gnd d0 a_14110_5733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X663 a_8882_1919# a_9135_1906# a_7940_2340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_17974_5477# a_18227_5464# a_17829_6246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X665 a_10148_6437# a_10149_5980# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X666 a_6866_2809# a_6752_2690# a_6859_4902# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X667 a_1793_4331# a_1726_3739# a_1810_2768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X668 vdd a_13060_7105# a_12852_7105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X669 a_12134_158# a_14876_138# a_9888_17# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X670 a_854_6781# a_433_6781# a_117_6662# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X671 gnd a_8056_3845# a_7848_3845# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X672 a_1584_6537# a_1371_6537# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X673 a_1805_2649# a_1514_1533# a_1794_2125# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X674 a_15518_8479# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X675 a_5701_7371# a_5488_7371# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X676 a_435_2369# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X677 a_10150_3774# a_10150_3587# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X678 a_120_1376# a_649_1266# a_857_1266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X679 a_857_1266# a_1587_1022# a_1795_1022# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X680 vdd a_4079_5728# a_3871_5728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X681 a_10885_7889# a_10464_7889# a_10148_7999# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X682 vdd a_19165_7980# a_18957_7980# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X683 a_16811_8197# a_16598_8197# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X684 a_12035_158# a_12854_4893# a_12809_4906# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X685 a_1803_7061# a_1694_7061# a_1808_4980# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X686 a_3823_8496# a_3819_8673# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X687 a_8881_4125# a_9134_4112# a_7939_4546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X688 a_18914_2478# a_19167_2465# a_17975_2168# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X689 gnd a_14110_5733# a_13902_5733# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X690 a_17859_7336# a_17878_6056# a_17829_6246# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X691 vdd d0 a_4077_9037# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X692 a_3821_8124# a_3824_7393# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X693 vdd d3 a_18118_2734# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X694 a_7938_6752# a_8195_6562# a_7802_6064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X695 a_10678_1820# a_10465_1820# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X696 a_12809_2706# a_12823_3809# a_12778_3822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X697 a_12919_2127# a_13903_2424# a_13854_2614# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X698 a_647_1815# a_434_1815# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X699 a_10150_2025# a_10678_1820# a_10886_1820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X700 a_649_1266# a_436_1266# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X701 a_16599_5991# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X702 a_8880_9091# a_8876_9268# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X703 a_6951_194# a_6738_194# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X704 a_7940_2340# a_8197_2150# a_7804_1652# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X705 a_1793_5434# a_1372_5434# a_854_5124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X706 a_10678_5683# a_10465_5683# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X707 a_6752_2690# a_6539_2690# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X708 a_1514_1533# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X709 a_10149_4877# a_10677_5129# a_10885_5129# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X710 a_117_8181# a_117_7994# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X711 a_11824_4336# a_11757_3744# a_11841_2773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X712 a_1726_3739# a_1513_3739# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X713 a_5174_5829# a_5703_5719# a_5911_5719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X714 a_6640_6578# a_6427_6578# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X715 a_17975_2168# a_18959_2465# a_18914_2478# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X716 a_11836_2654# a_11545_1538# a_11825_2130# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X717 a_10150_2255# a_10150_2025# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X718 a_3826_2981# a_4079_2968# a_2884_3402# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X719 a_2778_4901# a_2821_7100# a_2776_7113# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X720 vdd d0 a_4080_3522# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X721 a_13856_5192# a_13852_5369# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X722 a_10149_5980# a_10676_6232# a_10884_6232# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X723 a_6848_7681# a_6427_7681# a_5910_7925# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X724 vdd a_3141_3212# a_2933_3212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X725 a_3820_6467# a_3826_5741# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X726 a_2885_1196# a_3142_1006# a_2744_1788# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X727 a_16769_199# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X728 vdd a_4076_8483# a_3868_8483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X729 a_15943_3518# a_16673_3274# a_16881_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X730 a_8883_816# a_8879_993# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X731 a_5488_9028# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X732 a_6427_6578# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X733 a_2887_5431# a_3871_5728# a_3822_5918# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X734 a_18913_1924# a_18909_2101# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X735 a_10678_1820# a_10465_1820# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X736 a_3821_4261# a_4078_4071# a_2883_4505# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X737 a_5488_6268# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 vdd a_9135_5769# a_8927_5769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X739 a_117_6662# a_117_6432# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X740 gnd d1 a_18229_1052# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X741 gnd d0 a_4079_4625# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X742 gnd d0 a_4076_8483# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X743 a_2744_1788# a_3001_1598# a_2774_2878# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X744 a_5175_2291# a_5704_2410# a_5912_2410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X745 a_11757_3744# a_11544_3744# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X746 a_6859_7102# a_6750_7102# a_6864_5021# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X747 a_15940_6273# a_15519_6273# a_15204_6478# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X748 gnd a_3138_8727# a_2930_8727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X749 gnd a_4077_6277# a_3869_6277# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X750 a_18910_2655# a_18913_1924# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X751 a_8879_8537# a_8875_8714# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X752 a_118_5559# a_118_5329# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X753 a_15735_3518# a_15522_3518# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X754 a_646_5124# a_433_5124# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X755 vdd d0 a_19166_3014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X756 a_10149_5793# a_10149_5564# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X757 a_15735_758# a_15522_758# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X758 a_2743_3994# a_2933_3212# a_2888_3225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X759 a_10885_4026# a_10464_4026# a_10150_3774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X760 a_853_6227# a_1584_6537# a_1792_6537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X761 a_12916_1201# a_13173_1011# a_12775_1793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X762 a_16673_3274# a_16460_3274# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X763 a_13852_4266# a_14109_4076# a_12914_4510# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X764 a_7834_4942# a_7877_7141# a_7832_7154# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X765 a_5911_4616# a_5490_4616# a_5174_4726# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X766 a_15205_5605# a_15205_5375# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X767 a_7801_8270# a_8054_8257# a_7832_7154# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X768 a_1794_3228# a_1726_3739# a_1810_2768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X769 gnd a_19166_1911# a_18958_1911# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X770 gnd d0 a_19167_3568# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X771 gnd d0 a_19165_4117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X772 a_14985_138# a_14876_138# a_9888_17# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X773 a_5911_1856# a_5490_1856# a_5176_1604# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X774 a_5913_1307# a_5492_1307# a_5176_1188# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X775 a_854_6781# a_433_6781# a_117_6891# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X776 a_17833_6069# a_18018_6567# a_17973_6580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X777 a_12913_7819# a_13900_7385# a_13851_7575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X778 a_3825_6844# a_3821_7021# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X779 a_12919_2127# a_13172_2114# a_12779_1616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X780 vdd d0 a_14108_9042# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X781 a_15732_7376# a_15519_7376# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 a_17831_1834# a_18021_1052# a_17976_1065# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X783 a_16811_8197# a_16598_8197# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X784 a_17863_7159# a_18116_7146# a_17865_4947# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X785 a_15521_2964# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X786 a_12774_3999# a_12964_3217# a_12919_3230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X787 a_7943_5472# a_8927_5769# a_8878_5959# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X788 a_10148_6896# a_10677_6786# a_10885_6786# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X789 a_15209_864# a_15735_758# a_15943_758# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X790 vdd d0 a_19166_4671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X791 a_856_3472# a_435_3472# a_119_3582# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X792 a_10149_5334# a_10149_4877# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X793 a_11822_8748# a_11401_8748# a_10883_8438# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X794 a_6951_194# a_6738_194# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X795 a_856_712# a_435_712# a_122_818# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X796 a_15519_7376# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X797 a_1514_1533# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X798 a_11825_3233# a_11757_3744# a_11841_2773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X799 a_1726_3739# a_1513_3739# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X800 a_5910_6822# a_5489_6822# a_5173_6932# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X801 a_17971_2345# a_18958_1911# a_18909_2101# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X802 a_18908_7067# a_19165_6877# a_17973_6580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X803 a_15943_758# a_16674_1068# a_16882_1068# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X804 a_12134_158# a_11713_158# a_11933_4866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X805 vdd a_4080_762# a_3872_762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X806 a_1795_1022# a_1374_1022# a_856_712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X807 vdd a_18227_4361# a_18019_4361# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X808 a_7060_194# a_7879_4929# a_7834_4942# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X809 a_5489_5165# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X810 a_12916_8745# a_13900_9042# a_13851_9232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X811 a_16769_199# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X812 a_7945_1060# a_8929_1357# a_8884_1370# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X813 a_646_6781# a_433_6781# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X814 a_3824_6290# a_3820_6467# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X815 a_15942_2964# a_15521_2964# a_15206_3169# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X816 gnd d0 a_14107_8488# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X817 a_15205_4918# a_15205_4731# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X818 a_6781_5986# a_6568_5986# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X819 a_15206_3399# a_15206_3169# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X820 a_11757_3744# a_11544_3744# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X821 a_2885_8740# a_3869_9037# a_3824_9050# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X822 a_5701_9028# a_5488_9028# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X823 a_856_2369# a_435_2369# a_119_2250# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X824 a_16890_7107# a_16781_7107# a_16895_5026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X825 a_10467_1271# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X826 a_5702_7925# a_5489_7925# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X827 a_6861_2690# a_6570_1574# a_6850_2166# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X828 a_2885_1196# a_3872_762# a_3827_775# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X829 vdd a_14111_767# a_13903_767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X830 vdd d1 a_13170_7629# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X831 vdd d0 a_14110_2973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X832 a_11933_4866# a_11512_4866# a_11839_4985# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X833 vdd d0 a_14109_5179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X834 a_11826_1027# a_11405_1027# a_10887_717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X835 a_10149_5980# a_10149_5793# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X836 a_1803_4861# a_1483_2649# a_1805_2649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X837 a_5489_5165# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X838 a_432_6227# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X839 vdd a_4080_2419# a_3872_2419# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X840 gnd a_19163_8529# a_18955_8529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X841 gnd a_3140_4315# a_2932_4315# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X842 gnd d0 a_4077_7380# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X843 a_6850_2166# a_6429_2166# a_5912_2410# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X844 a_7834_2742# a_8087_2729# a_7830_5119# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X845 vdd a_13170_7629# a_12962_7629# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X846 vdd a_14109_5179# a_13901_5179# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X847 a_7941_8781# a_8925_9078# a_8880_9091# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X848 a_15206_2525# a_15735_2415# a_15943_2415# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X849 a_16600_3785# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X850 a_1694_7061# a_1481_7061# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X851 a_16892_2695# a_16783_2695# a_16890_4907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X852 a_11713_158# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X853 a_16460_3274# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X854 gnd a_13031_3809# a_12823_3809# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X855 a_2778_2701# a_2792_3804# a_2743_3994# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X856 a_2886_6534# a_3139_6521# a_2746_6023# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 a_17972_1242# a_18959_808# a_18910_998# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 a_12916_1201# a_13903_767# a_13858_780# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X859 a_18909_3204# a_18914_2478# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X860 a_10464_4026# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X861 a_10148_6667# a_10677_6786# a_10885_6786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X862 a_5053_133# a_4632_133# a_4954_133# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X863 a_2103_153# a_1682_153# a_1902_4861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X864 a_1481_4861# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X865 a_2881_8917# a_3868_8483# a_3819_8673# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X866 vdd a_14111_2424# a_13903_2424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X867 a_2888_2122# a_3872_2419# a_3827_2432# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X868 vdd d1 a_8197_3253# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X869 vdd d0 a_14109_6836# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X870 a_119_3123# a_647_2918# a_855_2918# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X871 a_11822_8748# a_11401_8748# a_10884_8992# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X872 gnd a_13171_4320# a_12963_4320# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X873 a_2747_3817# a_2932_4315# a_2883_4505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X874 a_17970_5654# a_18227_5464# a_17829_6246# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X875 a_5489_6822# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X876 a_16783_2695# a_16570_2695# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X877 gnd d0 a_4077_9037# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X878 a_2741_8406# a_2931_7624# a_2886_7637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X879 a_17969_7860# a_18956_7426# a_18911_7439# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X880 a_2883_5608# a_3870_5174# a_3825_5187# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X881 a_15941_6827# a_15520_6827# a_15204_6937# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X882 a_17971_2345# a_18228_2155# a_17835_1657# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X883 a_15942_4621# a_15521_4621# a_15205_4502# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X884 a_12809_2706# a_12823_3809# a_12774_3999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X885 vdd a_14109_6836# a_13901_6836# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X886 a_3826_1878# a_3822_2055# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X887 a_647_5678# a_434_5678# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X888 a_12772_8411# a_12962_7629# a_12913_7819# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X889 gnd a_9133_6318# a_8925_6318# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X890 a_12914_5613# a_13901_5179# a_13852_5369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X891 vdd d3 a_13060_7105# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X892 a_1793_5434# a_1372_5434# a_855_5678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X893 a_11823_7645# a_11402_7645# a_10884_7335# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X894 a_6429_2166# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X895 a_119_3123# a_119_2666# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X896 a_6641_4372# a_6428_4372# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X897 a_11512_4866# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X898 a_13851_9232# a_13854_8501# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X899 a_12807_7118# a_12821_8221# a_12772_8411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X900 gnd a_9134_5215# a_8926_5215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X901 a_11839_7185# a_11542_8156# a_11823_7645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X902 a_646_6781# a_433_6781# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X903 a_12919_2127# a_13903_2424# a_13858_2437# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X904 a_3823_2609# a_3826_1878# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X905 a_5702_7925# a_5489_7925# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X906 a_10150_3358# a_10679_3477# a_10887_3477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X907 a_12778_3822# a_12963_4320# a_12914_4510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X908 a_1371_7640# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X909 a_10151_922# a_10679_717# a_10887_717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X910 gnd a_9136_2460# a_8928_2460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X911 a_18914_821# a_18910_998# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X912 gnd d1 a_3141_3212# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X913 a_3822_3158# a_4079_2968# a_2884_3402# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X914 a_6850_3269# a_6782_3780# a_6866_2809# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X915 a_5173_8222# a_5700_8474# a_5908_8474# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X916 gnd d1 a_3139_7624# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X917 a_1374_1022# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X918 a_1586_3228# a_1373_3228# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X919 a_15732_9033# a_15519_9033# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X920 a_16671_6583# a_16458_6583# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X921 a_7937_8958# a_8924_8524# a_8875_8714# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X922 a_433_5124# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X923 a_3822_3158# a_3827_2432# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X924 a_5173_7119# a_5701_7371# a_5909_7371# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X925 a_15733_7930# a_15520_7930# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X926 a_5176_1188# a_5705_1307# a_5913_1307# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X927 a_16672_5480# a_16459_5480# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X928 a_2886_6534# a_3870_6831# a_3825_6844# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X929 a_15206_2296# a_15735_2415# a_15943_2415# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X930 gnd d0 a_14108_7385# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X931 a_1803_4861# a_1483_2649# a_1810_2768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X932 gnd a_4081_1316# a_3873_1316# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X933 gnd a_4079_1865# a_3871_1865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X934 a_2748_1611# a_3001_1598# a_2774_2878# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X935 a_13854_2614# a_13857_1883# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X936 vdd d1 a_3140_4315# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X937 a_5910_4062# a_6641_4372# a_6849_4372# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X938 a_7797_8447# a_7987_7665# a_7942_7678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X939 gnd d0 a_19164_7426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X940 a_7939_5649# a_8926_5215# a_8881_5228# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X941 a_15519_9033# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X942 a_16458_6583# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X943 a_7944_2163# a_8928_2460# a_8879_2650# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X944 gnd a_2998_8216# a_2790_8216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X945 a_7832_7154# a_7846_8257# a_7801_8270# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X946 a_15206_3628# a_15206_3399# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X947 vdd d0 a_4076_8483# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X948 a_16459_5480# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X949 a_6782_3780# a_6569_3780# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X950 a_11617_3233# a_11404_3233# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X951 a_6849_4372# a_6782_3780# a_6866_2809# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_10150_2484# a_10679_2374# a_10887_2374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X953 a_119_3769# a_119_3582# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X954 a_8881_5228# a_8877_5405# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X955 a_13853_3163# a_13858_2437# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X956 vdd d0 a_9133_7421# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X957 a_5705_1307# a_5492_1307# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X958 a_5053_133# a_4632_133# a_2103_153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X959 a_5172_9138# a_5172_8909# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X960 gnd a_19164_7426# a_18956_7426# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X961 a_8877_7062# a_8880_6331# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X962 a_10884_7335# a_10463_7335# a_10148_7540# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X963 vdd d0 a_9136_803# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X964 a_5174_4267# a_5702_4062# a_5910_4062# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X965 a_648_712# a_435_712# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X966 gnd a_14110_1870# a_13902_1870# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X967 a_2889_1019# a_3873_1316# a_3824_1506# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X968 a_2884_2299# a_3871_1865# a_3822_2055# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X969 gnd d0 a_14111_3527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X970 a_1696_2649# a_1483_2649# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X971 gnd d0 a_14109_4076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X972 a_16568_7107# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X973 gnd d0 a_14108_9042# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X974 a_17831_1834# a_18021_1052# a_17972_1242# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X975 a_18911_6336# a_19164_6323# a_17969_6757# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X976 a_10465_2923# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X977 gnd d0 a_4078_5174# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X978 a_16881_2171# a_16460_2171# a_15942_1861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X979 gnd a_18907_9273# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X980 a_436_1266# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X981 gnd d0 a_19164_9083# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X982 a_1682_153# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X983 vdd d0 a_14110_4630# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X984 a_6782_3780# a_6569_3780# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X985 vdd d4 a_13062_4893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X986 a_10676_6232# a_10463_6232# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X987 vdd d2 a_18087_3850# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X988 a_2882_7814# a_3869_7380# a_3820_7570# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X989 gnd a_13172_3217# a_12964_3217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X990 a_15206_3169# a_15206_2712# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X991 vdd d0 a_14110_5733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X992 a_855_1815# a_1586_2125# a_1794_2125# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X993 a_15205_5834# a_15734_5724# a_15942_5724# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X994 a_5704_3513# a_5491_3513# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X995 a_5702_4062# a_5489_4062# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X996 a_10679_717# a_10466_717# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X997 a_12920_1024# a_13904_1321# a_13855_1511# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X998 a_6850_3269# a_6429_3269# a_5911_2959# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X999 a_12915_2304# a_13902_1870# a_13853_2060# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1000 a_17834_3863# a_18087_3850# a_17865_2747# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1001 gnd a_8087_4929# a_7879_4929# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1002 a_433_6781# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1003 a_7941_1237# a_8198_1047# a_7800_1829# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1004 a_6864_5021# a_6750_4902# a_6958_4902# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1005 gnd a_4078_6831# a_3870_6831# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1006 gnd a_19164_9083# a_18956_9083# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1007 gnd d0 a_9134_7975# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1008 vdd d0 a_9136_2460# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1009 a_5172_8679# a_5173_8222# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1010 a_15733_7930# a_15520_7930# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1011 a_648_2369# a_435_2369# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1012 a_16672_5480# a_16459_5480# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1013 a_3825_7947# a_4078_7934# a_2886_7637# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1014 a_10463_6232# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1015 gnd d0 a_4080_762# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1016 a_8877_4302# a_9134_4112# a_7939_4546# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1017 vdd a_14110_5733# a_13902_5733# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1018 gnd d2 a_8056_3845# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1019 a_17834_3863# a_18019_4361# a_17974_4374# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1020 a_8877_4302# a_8883_3576# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1021 a_15732_9033# a_15519_9033# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1022 a_13854_8501# a_13850_8678# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1023 a_16671_6583# a_16458_6583# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1024 a_15204_8227# a_15731_8479# a_15939_8479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1025 a_10886_2923# a_10465_2923# a_10150_3128# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1026 a_2774_2878# a_3031_2688# a_2774_5078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1027 a_15204_7124# a_15732_7376# a_15940_7376# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1028 a_16459_5480# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1029 a_18910_8542# a_18906_8719# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1030 a_13852_8129# a_14109_7939# a_12917_7642# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1031 a_856_2369# a_1586_2125# a_1794_2125# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1032 vdd d0 a_4081_1316# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1033 vdd d0 a_4079_1865# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1034 vdd a_18087_3850# a_17879_3850# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1035 a_3822_5918# a_3825_5187# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1036 a_18908_8170# a_18911_7439# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1037 a_11824_5439# a_11403_5439# a_10885_5129# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1038 a_2885_8740# a_3869_9037# a_3820_9227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1039 a_16892_2695# a_16601_1579# a_16881_2171# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1040 a_6750_4902# a_6537_4902# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1041 a_117_6432# a_645_6227# a_853_6227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1042 a_5491_3513# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1043 a_15519_9033# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1044 a_16458_6583# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1045 a_7803_3858# a_7988_4356# a_7939_4546# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1046 a_10679_2374# a_10466_2374# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1047 a_5912_753# a_5491_753# a_5176_958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1048 a_12809_4906# a_12852_7105# a_12807_7118# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1049 a_9888_17# a_9779_17# vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1050 a_4632_133# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1051 gnd d2 a_18086_6056# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1052 a_15206_3815# a_15206_3628# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1053 gnd d1 a_13169_8732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1054 a_11617_3233# a_11404_3233# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1055 a_6958_4902# a_6537_4902# a_6864_5021# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1056 a_2887_5431# a_3871_5728# a_3826_5741# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1057 a_17973_7683# a_18957_7980# a_18912_7993# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1058 a_12805_2883# a_13062_2693# a_12805_5083# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1059 a_17865_2747# a_18118_2734# a_17861_5124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1060 a_5913_1307# a_6643_1063# a_6851_1063# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1061 gnd a_9134_6872# a_8926_6872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1062 a_3825_4084# a_4078_4071# a_2883_4505# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1063 a_12918_5436# a_13902_5733# a_13853_5923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1064 a_18907_6513# a_18913_5787# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1065 a_15203_9143# a_15203_8914# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1066 a_3824_9050# a_5172_9138# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1067 a_11836_2654# a_11727_2654# a_11834_4866# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1068 vdd a_3138_8727# a_2930_8727# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1069 vdd a_4077_6277# a_3869_6277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1070 gnd d1 a_18228_2155# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1071 a_1696_2649# a_1483_2649# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1072 a_10886_4580# a_10465_4580# a_10149_4690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1073 a_11542_8156# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1074 a_2884_2299# a_3141_2109# a_2748_1611# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1075 a_3820_7570# a_4077_7380# a_2882_7814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1076 gnd a_13169_8732# a_12961_8732# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1077 gnd a_14108_6282# a_13900_6282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1078 a_15942_4621# a_16672_4377# a_16880_4377# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1079 a_8882_4679# a_8878_4856# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1080 a_10677_5129# a_10464_5129# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1081 a_1895_153# a_1682_153# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1082 a_5703_5719# a_5490_5719# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1083 a_3822_4815# a_4079_4625# a_2887_4328# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1084 a_12920_1024# a_13173_1011# a_12775_1793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1085 a_8880_6331# a_8876_6508# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1086 gnd d1 a_8197_3253# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1087 a_17865_4947# a_18118_4934# a_17091_199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1088 a_5909_6268# a_6640_6578# a_6848_6578# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1089 a_8878_5959# a_8881_5228# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1090 a_5172_8909# a_5701_9028# a_5909_9028# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1091 gnd d0 a_4079_5728# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1092 a_10676_6232# a_10463_6232# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1093 a_434_5678# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1094 a_5174_5600# a_5174_5370# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1095 a_5173_6473# a_5701_6268# a_5909_6268# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1096 a_5489_4062# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1097 a_13856_4089# a_14109_4076# a_12914_4510# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1098 a_2881_8917# a_3868_8483# a_3823_8496# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1099 vdd d0 a_19167_3568# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1100 a_1791_8743# a_1724_8151# a_1808_7180# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1101 a_5173_6932# a_5173_6703# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1102 vdd d0 a_19165_4117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1103 a_10464_5129# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1104 gnd a_3140_5418# a_2932_5418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1105 a_15736_1312# a_15523_1312# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1106 a_3827_3535# a_3823_3712# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1107 a_11727_2654# a_11514_2654# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1108 a_433_6781# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1109 gnd a_9135_1906# a_8927_1906# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1110 a_10886_4580# a_10465_4580# a_10149_4461# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1111 gnd a_18085_8262# a_17877_8262# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1112 a_12915_2304# a_13172_2114# a_12779_1616# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1113 a_16879_6583# a_16812_5991# a_16890_7107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1114 vdd a_13030_6015# a_12822_6015# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1115 vdd a_14112_1321# a_13904_1321# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1116 gnd d0 a_19165_7980# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1117 a_15520_5170# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1118 a_7943_5472# a_8927_5769# a_8882_5782# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1119 a_10463_6232# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1120 a_16672_4377# a_16459_4377# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1121 a_15203_8684# a_15204_8227# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1122 a_10884_7335# a_11615_7645# a_11823_7645# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1123 a_855_1815# a_434_1815# a_119_2020# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1124 a_6750_7102# a_6537_7102# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1125 a_2745_8229# a_2930_8727# a_2881_8917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1126 a_7802_6064# a_8055_6051# a_7828_7331# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1127 a_18913_3027# a_19166_3014# a_17971_3448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1128 a_18912_6890# a_18908_7067# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1129 vdd a_9133_6318# a_8925_6318# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1130 vdd a_18228_3258# a_18020_3258# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1131 gnd d0 a_19166_4671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1132 a_17831_1834# a_18088_1644# a_17861_2924# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1133 a_5912_2410# a_5491_2410# a_5175_2291# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1134 a_118_4872# a_646_5124# a_854_5124# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1135 a_8876_7611# a_9133_7421# a_7938_7855# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1136 vdd d3 a_8085_7141# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1137 gnd a_19165_7980# a_18957_7980# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1138 a_16570_2695# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1139 a_13858_3540# a_13854_3717# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1140 a_6430_1063# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1141 a_7945_1060# a_8929_1357# a_8880_1547# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1142 a_7940_2340# a_8927_1906# a_8878_2096# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1143 vdd d2 a_8057_1639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1144 a_1810_2768# a_1513_3739# a_1794_3228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1145 a_15207_1609# a_15734_1861# a_15942_1861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1146 a_15207_1193# a_15736_1312# a_15944_1312# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1147 gnd d0 a_9135_5769# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1148 a_9566_17# d7 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1149 a_15520_5170# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1150 a_2772_7290# a_2791_6010# a_2746_6023# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1151 a_4632_133# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1152 a_6859_4902# a_6539_2690# a_6866_2809# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1153 a_857_1266# a_436_1266# a_120_1147# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1154 a_855_1815# a_434_1815# a_120_1563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1155 a_853_6227# a_432_6227# a_117_6432# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1156 vdd a_8197_2150# a_7989_2150# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1157 a_15734_1861# a_15521_1861# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1158 a_17975_2168# a_18959_2465# a_18910_2655# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1159 a_16989_4907# a_16568_4907# a_16895_5026# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1160 a_10677_6786# a_10464_6786# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1161 a_11825_2130# a_11404_2130# a_10887_2374# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1162 a_7832_7154# a_7846_8257# a_7797_8447# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1163 a_7804_1652# a_7989_2150# a_7944_2163# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1164 a_6864_7221# a_6567_8192# a_6848_7681# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1165 a_16880_4377# a_16813_3785# a_16897_2814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1166 a_13855_9055# a_15203_9143# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1167 a_7801_8270# a_7986_8768# a_7937_8958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1168 a_5176_1188# a_5176_958# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1169 vdd a_3001_1598# a_2793_1598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1170 vdd a_3142_1006# a_2934_1006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1171 gnd d0 a_4080_2419# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1172 a_120_1147# a_120_917# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1173 a_15943_3518# a_15522_3518# a_15206_3628# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1174 a_10464_6786# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1175 a_15941_4067# a_15520_4067# a_15205_4272# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1176 a_5174_4913# a_5702_5165# a_5910_5165# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1177 gnd d0 a_9136_803# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1178 a_15734_5724# a_15521_5724# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1179 a_15943_758# a_15522_758# a_15209_864# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1180 vdd a_19163_8529# a_18955_8529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1181 a_18908_5410# a_18913_4684# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1182 a_2744_1788# a_2934_1006# a_2889_1019# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1183 a_15520_6827# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1184 a_6642_3269# a_6429_3269# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1185 a_120_1376# a_120_1147# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1186 vdd d2 a_13029_8221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1187 a_7830_2919# a_8087_2729# a_7830_5119# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1188 a_15204_6478# a_15732_6273# a_15940_6273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1189 a_434_2918# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1190 a_11825_2130# a_11404_2130# a_10886_1820# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1191 a_16813_3785# a_16600_3785# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1192 a_7828_7331# a_7847_6051# a_7802_6064# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1193 a_15204_6937# a_15204_6708# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1194 a_116_8638# a_117_8181# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1195 a_117_6891# a_646_6781# a_854_6781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1196 a_5909_6268# a_5488_6268# a_5173_6473# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1197 a_5912_2410# a_5491_2410# a_5175_2520# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1198 a_18907_6513# a_19164_6323# a_17969_6757# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1199 a_1808_7180# a_1511_8151# a_1791_8743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1200 gnd a_3029_7100# a_2821_7100# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1201 a_16781_7107# a_16568_7107# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1202 a_17972_1242# a_18229_1052# a_17831_1834# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1203 a_5174_5370# a_5702_5165# a_5910_5165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1204 vdd a_19167_808# a_18959_808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1205 a_17833_6069# a_18086_6056# a_17859_7336# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1206 a_7945_1060# a_8198_1047# a_7800_1829# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1207 a_5173_6703# a_5173_6473# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1208 a_6537_4902# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1209 a_5174_5829# a_5174_5600# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1210 a_17973_6580# a_18226_6567# a_17833_6069# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1211 a_10885_5129# a_10464_5129# a_10149_4877# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1212 vdd d3 a_18116_7146# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1213 a_5176_958# a_5178_859# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1214 a_18908_4307# a_18914_3581# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1215 a_17968_8963# a_18955_8529# a_18906_8719# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1216 vdd a_13062_4893# a_12854_4893# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1217 a_120_917# a_122_818# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1218 a_1810_2768# a_1513_3739# a_1793_4331# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1219 a_3821_8124# a_4078_7934# a_2886_7637# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1220 a_11615_7645# a_11402_7645# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1221 a_12772_8411# a_12962_7629# a_12917_7642# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1222 a_2778_2701# a_3031_2688# a_2774_5078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1223 a_12914_5613# a_13901_5179# a_13856_5192# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1224 a_119_3582# a_648_3472# a_856_3472# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1225 a_12779_1616# a_12964_2114# a_12915_2304# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1226 a_18913_5787# a_18909_5964# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1227 gnd d0 a_19166_5774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1228 a_8878_3199# a_9135_3009# a_7940_3443# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1229 a_11824_5439# a_11403_5439# a_10886_5683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1230 vdd a_18116_7146# a_17908_7146# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1231 vdd d3 a_3031_2688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1232 a_15522_3518# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1233 a_15520_4067# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1234 a_5175_2707# a_5703_2959# a_5911_2959# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1235 a_10677_6786# a_10464_6786# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1236 a_1373_2125# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1237 vref a_116_9097# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1238 a_5173_6932# a_5702_6822# a_5910_6822# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1239 a_11402_7645# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1240 vdd a_19167_2465# a_18959_2465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1241 a_13852_7026# a_13855_6295# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1242 vdd d1 a_3141_3212# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1243 gnd a_18227_4361# a_18019_4361# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1244 a_10150_2484# a_10150_2255# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1245 a_6864_7221# a_6567_8192# a_6847_8784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1246 vdd d1 a_3139_7624# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1247 gnd a_19166_5774# a_18958_5774# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 gnd a_8085_7141# a_7877_7141# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1249 a_5174_5370# a_5174_4913# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1250 a_7937_8958# a_8924_8524# a_8879_8537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1251 a_16882_1068# a_16461_1068# a_15944_1312# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1252 a_12809_2706# a_13062_2693# a_12805_5083# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1253 a_8883_3576# a_9136_3563# a_7944_3266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1254 a_435_712# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1255 a_15521_5724# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1256 a_10464_6786# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1257 a_7834_2742# a_7848_3845# a_7799_4035# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1258 a_10151_1381# a_10680_1271# a_10888_1271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1259 a_10888_1271# a_11618_1027# a_11826_1027# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1260 a_15205_4918# a_15733_5170# a_15941_5170# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1261 a_12917_6539# a_13901_6836# a_13856_6849# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1262 a_7938_6752# a_8925_6318# a_8876_6508# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1263 a_15207_1422# a_15207_1193# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1264 a_2888_2122# a_3141_2109# a_2748_1611# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1265 a_5703_2959# a_5490_2959# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1266 a_18913_4684# a_18909_4861# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1267 vdd a_9134_6872# a_8926_6872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1268 a_11404_2130# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1269 a_117_6891# a_117_6662# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1270 a_1373_2125# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1271 a_1585_4331# a_1372_4331# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1272 a_18912_5233# a_18908_5410# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1273 a_118_5559# a_647_5678# a_855_5678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1274 a_7797_8447# a_7987_7665# a_7938_7855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1275 a_7939_5649# a_8926_5215# a_8877_5405# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1276 a_8878_4856# a_9135_4666# a_7943_4369# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1277 a_8877_8165# a_9134_7975# a_7942_7678# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1278 a_7828_7331# a_8085_7141# a_7834_4942# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1279 a_15206_3169# a_15734_2964# a_15942_2964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1280 a_645_6227# a_432_6227# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1281 a_8876_9268# a_8879_8537# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1282 gnd a_13062_4893# a_12854_4893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1283 gnd d0 a_9132_8524# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1284 a_117_6662# a_646_6781# a_854_6781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1285 a_15734_2964# a_15521_2964# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1286 a_8882_5782# a_9135_5769# a_7943_5472# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1287 a_10150_2025# a_10151_1568# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1288 a_5700_8474# a_5487_8474# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1289 vdd d0 a_14111_3527# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1290 a_10680_1271# a_10467_1271# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1291 a_15205_5375# a_15733_5170# a_15941_5170# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1292 a_5701_7371# a_5488_7371# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1293 a_16880_5480# a_16812_5991# a_16890_7107# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1294 a_435_2369# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1295 vdd d1 a_8195_7665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1296 vdd a_3139_6521# a_2931_6521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1297 a_856_712# a_1587_1022# a_1795_1022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1298 vdd d0 a_9134_5215# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1299 a_120_1147# a_649_1266# a_857_1266# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1300 a_15204_6708# a_15204_6478# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1301 a_11404_2130# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1302 vdd d0 a_4078_5174# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1303 a_15205_5834# a_15205_5605# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1304 a_11616_4336# a_11403_4336# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1305 a_5174_6016# a_5174_5829# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1306 a_16989_4907# a_16982_199# a_14985_138# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1307 vdd a_3140_5418# a_2932_5418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1308 a_5490_2959# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1309 a_5053_133# a_9779_17# vout gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1310 a_13857_2986# a_14110_2973# a_12915_3407# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1311 vdd d4 a_8087_4929# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1312 vdd d0 a_19164_9083# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1313 a_7830_5119# a_7879_2729# a_7830_2919# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1314 vdd d0 a_9137_1357# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1315 a_5174_4726# a_5703_4616# a_5911_4616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1316 vdd d3 a_3029_7100# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1317 a_649_1266# a_436_1266# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1318 vdd a_13172_3217# a_12964_3217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1319 gnd d0 a_14109_6836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1320 a_117_6432# a_118_5975# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1321 gnd a_18228_3258# a_18020_3258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1322 gnd d0 a_14110_4630# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1323 a_12775_1793# a_13032_1603# a_12805_2883# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1324 a_17835_1657# a_18088_1644# a_17861_2924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1325 vdd a_8195_7665# a_7987_7665# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1326 vdd d1 a_18227_4361# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1327 a_16461_1068# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1328 vdd a_8054_8257# a_7846_8257# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1329 a_5174_5600# a_5703_5719# a_5911_5719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1330 a_17835_1657# a_18020_2155# a_17971_2345# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1331 a_10466_3477# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1332 a_6849_4372# a_6428_4372# a_5910_4062# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1333 vdd a_19164_9083# a_18956_9083# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1334 a_17969_7860# a_18956_7426# a_18907_7616# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1335 gnd d2 a_8057_1639# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1336 a_11839_4985# a_11512_7066# a_11834_7066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1337 gnd a_19168_1362# a_18960_1362# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1338 vdd d0 a_4080_762# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1339 gnd a_14109_6836# a_13901_6836# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1340 a_118_4226# a_646_4021# a_854_4021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1341 a_15204_6937# a_15733_6827# a_15941_6827# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1342 a_13856_7952# a_14109_7939# a_12917_7642# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1343 a_15942_2964# a_16673_3274# a_16881_3274# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1344 a_3820_9227# a_4077_9037# a_2885_8740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1345 vdd d0 a_4078_6831# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1346 a_5703_4616# a_5490_4616# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1347 a_1792_6537# a_1371_6537# a_853_6227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1348 a_15205_5375# a_15205_4918# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1349 a_16878_8789# a_16457_8789# a_15939_8479# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1350 vdd a_8087_4929# a_7879_4929# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1351 a_5488_6268# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1352 a_1794_3228# a_1373_3228# a_855_2918# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1353 vdd a_9137_1357# a_8929_1357# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1354 a_1370_8743# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1355 vdd a_8057_1639# a_7849_1639# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1356 a_13853_5923# a_13856_5192# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1357 gnd a_3001_1598# a_2793_1598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1358 a_15735_758# a_15522_758# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1359 a_1585_4331# a_1372_4331# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1360 a_17976_1065# a_18960_1362# a_18911_1552# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1361 a_10887_3477# a_10466_3477# a_10150_3587# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1362 a_10885_4026# a_10464_4026# a_10149_4231# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1363 a_10886_5683# a_10465_5683# a_10149_5564# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1364 a_10887_717# a_10466_717# a_10153_823# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1365 a_1808_4980# a_1694_4861# a_1902_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1366 a_17972_8786# a_18956_9083# a_18907_9273# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1367 a_2886_6534# a_3870_6831# a_3821_7021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1368 vdd d1 a_13169_8732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1369 a_7830_2919# a_7849_1639# a_7804_1652# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1370 a_16673_3274# a_16460_3274# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1371 vdd d0 a_4080_2419# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1372 a_8883_3576# a_8879_3753# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1373 a_17861_2924# a_18118_2734# a_17861_5124# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1374 a_10148_7083# a_10148_6896# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1375 a_5176_1604# a_5176_1417# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1376 gnd d1 a_3140_4315# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1377 gnd d0 a_19163_8529# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1378 a_12918_5436# a_13902_5733# a_13857_5746# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1379 a_5490_4616# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1380 a_6850_2166# a_6783_1574# a_6861_2690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1381 a_1694_4861# a_1481_4861# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1382 a_3821_4261# a_3827_3535# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1383 a_5913_1307# a_5492_1307# a_5176_1417# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1384 a_5911_1856# a_5490_1856# a_5175_2061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1385 a_118_5788# a_118_5559# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1386 a_3823_8496# a_4076_8483# a_2881_8917# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1387 a_15731_8479# a_15518_8479# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1388 vdd a_13169_8732# a_12961_8732# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1389 vdd a_14108_6282# a_13900_6282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1390 a_15732_7376# a_15519_7376# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1391 vdd d1 a_18226_7670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1392 a_9779_17# a_9566_17# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1393 a_11616_4336# a_11403_4336# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1394 vdd d0 a_19165_5220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1395 a_13851_7575# a_14108_7385# a_12913_7819# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1396 a_6848_6578# a_6427_6578# a_5909_6268# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1397 a_17091_199# a_16982_199# a_14985_138# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1398 a_5174_4497# a_5174_4267# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1399 vdd d2 a_2998_8216# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1400 gnd d0 a_9133_7421# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1401 a_15205_6021# a_15205_5834# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1402 a_5912_2410# a_6642_2166# a_6850_2166# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1403 a_17976_1065# a_18229_1052# a_17831_1834# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1404 gnd d1 a_13171_5423# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1405 a_3826_4638# a_4079_4625# a_2887_4328# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1406 a_6849_5475# a_6428_5475# a_5910_5165# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1407 gnd a_19167_808# a_18959_808# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1408 vdd d0 a_4079_5728# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1409 a_6426_8784# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1410 a_15518_8479# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1411 vdd d0 a_19166_1911# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1412 a_856_712# a_435_712# a_120_917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1413 a_10883_8438# a_10462_8438# a_10148_8186# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1414 a_12917_7642# a_13170_7629# a_12772_8411# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1415 a_15519_7376# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1416 a_10887_2374# a_10466_2374# a_10150_2255# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1417 vdd a_18226_7670# a_18018_7670# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1418 a_6783_1574# a_6570_1574# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1419 vdd a_19165_5220# a_18957_5220# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1420 a_13852_4266# a_13858_3540# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1421 a_16600_3785# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1422 a_16897_2814# a_16783_2695# a_16890_4907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1423 vdd a_18085_8262# a_17877_8262# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1424 a_11822_8748# a_11755_8156# a_11839_7185# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1425 gnd a_13171_5423# a_12963_5423# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1426 a_7942_6575# a_8926_6872# a_8877_7062# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1427 a_1795_1022# a_1374_1022# a_857_1266# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1428 a_16982_199# a_16769_199# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1429 gnd a_13030_6015# a_12822_6015# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1430 a_2745_8229# a_2930_8727# a_2885_8740# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1431 a_18909_3204# a_19166_3014# a_17971_3448# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1432 gnd a_18227_5464# a_18019_5464# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1433 a_118_5329# a_118_4872# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1434 a_1803_7061# a_1512_5945# a_1792_6537# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1435 a_8882_3022# a_9135_3009# a_7940_3443# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1436 gnd d3 a_3031_2688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1437 a_12776_8234# a_12961_8732# a_12912_8922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1438 a_12913_6716# a_13900_6282# a_13851_6472# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1439 a_16878_8789# a_16457_8789# a_15940_9033# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1440 a_1792_6537# a_1371_6537# a_854_6781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1441 a_15735_2415# a_15522_2415# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1442 gnd d0 a_9133_9078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1443 a_3826_4638# a_3822_4815# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1444 a_8879_8537# a_9132_8524# a_7937_8958# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1445 a_854_7884# a_433_7884# a_117_7765# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1446 a_1584_7640# a_1371_7640# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1447 vdd a_8198_1047# a_7990_1047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1448 gnd d0 a_9136_2460# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1449 a_16568_4907# d4 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1450 vdd a_3031_2688# a_2823_2688# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1451 a_11933_4866# a_11926_158# a_12134_158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1452 a_5701_9028# a_5488_9028# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1453 a_1370_8743# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1454 a_16783_2695# a_16570_2695# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1455 a_856_2369# a_435_2369# a_119_2479# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1456 a_17834_3863# a_18019_4361# a_17970_4551# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1457 a_18914_3581# a_19167_3568# a_17975_3271# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1458 a_18912_4130# a_19165_4117# a_17970_4551# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1459 a_5701_6268# a_5488_6268# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1460 a_10150_2671# a_10150_2484# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1461 a_11826_1027# a_11405_1027# a_10888_1271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1462 a_17865_2747# a_17879_3850# a_17830_4040# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1463 a_10151_1152# a_10151_922# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1464 vdd d0 a_9135_5769# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1465 a_7938_7855# a_8195_7665# a_7797_8447# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1466 a_6958_4902# a_6537_4902# a_6859_4902# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1467 a_2742_6200# a_2932_5418# a_2883_5608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1468 a_10150_3128# a_10678_2923# a_10886_2923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1469 a_647_2918# a_434_2918# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1470 a_16879_7686# a_16458_7686# a_15940_7376# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1471 a_10886_5683# a_10465_5683# a_10149_5793# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1472 a_3821_7021# a_3824_6290# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1473 a_16812_5991# a_16599_5991# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1474 a_2772_7290# a_2791_6010# a_2742_6200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1475 a_17863_7159# a_17877_8262# a_17828_8452# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1476 a_432_6227# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1477 a_12803_7295# a_12822_6015# a_12777_6028# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1478 gnd d0 a_4081_1316# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1479 gnd d0 a_4079_1865# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1480 a_11834_4866# a_11514_2654# a_11836_2654# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1481 a_10151_1381# a_10151_1152# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1482 a_13857_4643# a_13853_4820# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1483 a_1371_7640# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1484 a_18909_4861# a_19166_4671# a_17974_4374# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1485 a_2774_5078# a_2823_2688# a_2778_2701# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1486 a_1511_8151# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1487 a_10148_7083# a_10676_7335# a_10884_7335# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1488 a_7799_4035# a_8056_3845# a_7834_2742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1489 a_6849_5475# a_6428_5475# a_5911_5719# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1490 a_7801_8270# a_7986_8768# a_7941_8781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1491 a_7938_6752# a_8925_6318# a_8880_6331# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1492 a_11713_158# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1493 a_3825_4084# a_3821_4261# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1494 a_118_5975# a_118_5788# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1495 a_10464_4026# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1496 a_17973_7683# a_18957_7980# a_18908_8170# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1497 vdd d0 a_4078_4071# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1498 vdd a_3141_2109# a_2933_2109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1499 a_10678_2923# a_10465_2923# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1500 a_1481_4861# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1501 vdd d2 a_3001_1598# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1502 gnd a_3031_4888# a_2823_4888# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1503 a_4954_133# a_6738_194# a_7060_194# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1504 a_6426_8784# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1505 gnd d1 a_13172_3217# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1506 a_6640_7681# a_6427_7681# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1507 a_3824_7393# a_4077_7380# a_2882_7814# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1508 a_5489_6822# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1509 a_15521_2964# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1510 a_10148_7770# a_10148_7540# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1511 gnd d2 a_13029_8221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1512 a_12805_5083# a_12854_2693# a_12809_2706# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1513 vdd a_2999_6010# a_2791_6010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1514 a_10151_922# a_10153_823# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1515 a_119_2250# a_119_2020# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1516 a_15942_4621# a_15521_4621# a_15205_4731# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1517 gnd d1 a_8194_8768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1518 a_13856_4089# a_13852_4266# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1519 a_853_7330# a_1584_7640# a_1792_7640# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1520 a_15735_2415# a_15522_2415# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1521 gnd d0 a_4077_6277# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1522 a_13850_8678# a_14107_8488# a_12912_8922# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1523 a_15942_1861# a_15521_1861# a_15207_1609# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1524 a_15944_1312# a_15523_1312# a_15207_1193# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1525 a_16982_199# a_16769_199# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1526 a_5174_4726# a_5174_4497# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1527 a_12779_1616# a_13032_1603# a_12805_2883# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1528 a_1902_4861# a_1895_153# a_2103_153# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1529 a_2748_1611# a_2933_2109# a_2888_2122# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1530 vdd d1 a_13171_4320# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1531 a_6429_2166# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1532 a_6641_4372# a_6428_4372# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1533 a_6427_7681# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1534 a_13853_3163# a_14110_2973# a_12915_3407# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1535 a_11512_4866# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1536 a_11405_1027# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1537 a_119_2479# a_119_2250# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1538 a_10884_7335# a_10463_7335# a_10148_7083# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1539 gnd a_8054_8257# a_7846_8257# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1540 a_11839_7185# a_11542_8156# a_11822_8748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1541 gnd a_13060_7105# a_12852_7105# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1542 vdd d2 a_13032_1603# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1543 gnd a_19166_3014# a_18958_3014# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1544 a_17969_6757# a_18226_6567# a_17833_6069# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1545 gnd a_8194_8768# a_7986_8768# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1546 a_5911_2959# a_5490_2959# a_5175_2707# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1547 a_5175_3623# a_5704_3513# a_5912_3513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1548 a_15940_7376# a_15519_7376# a_15204_7124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1549 a_10153_823# a_10679_717# a_10887_717# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1550 a_5702_5165# a_5489_5165# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1551 a_17828_8452# a_18018_7670# a_17973_7683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1552 gnd a_14112_1321# a_13904_1321# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1553 gnd d1 a_8196_4356# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1554 a_14663_138# d6 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1555 a_17968_8963# a_18955_8529# a_18910_8542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1556 a_10148_7999# a_10677_7889# a_10885_7889# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1557 a_1374_1022# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1558 a_1586_3228# a_1373_3228# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1559 vdd a_18118_4934# a_17910_4934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1560 a_3824_9050# a_4077_9037# a_2885_8740# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1561 a_10884_8992# a_11614_8748# a_11822_8748# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1562 vdd a_19168_1362# a_18960_1362# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1563 a_15732_6273# a_15519_6273# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1564 a_7944_2163# a_8197_2150# a_7804_1652# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1565 vdd d2 a_8054_8257# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1566 a_12779_1616# a_12964_2114# a_12919_2127# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1567 vdd d0 a_19166_5774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1568 a_16879_7686# a_16458_7686# a_15941_7930# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1569 a_12803_7295# a_13060_7105# a_12809_4906# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1570 a_2741_8406# a_2998_8216# a_2776_7113# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1571 a_8880_7434# a_9133_7421# a_7938_7855# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1572 vdd a_8055_6051# a_7847_6051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1573 a_5174_4267# a_5175_3810# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1574 a_6859_4902# a_6750_4902# a_6958_4902# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1575 a_18908_8170# a_19165_7980# a_17973_7683# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1576 gnd a_8057_1639# a_7849_1639# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1577 a_17971_3448# a_18958_3014# a_18909_3204# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1578 a_2778_4901# a_2821_7100# a_2772_7290# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1579 a_10884_8992# a_10463_8992# a_10147_8873# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1580 a_18907_9273# a_18910_8542# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1581 a_119_2020# a_120_1563# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1582 a_11926_158# a_11713_158# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1583 a_5702_5165# a_5489_5165# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1584 a_15519_6273# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1585 a_13857_5746# a_14110_5733# a_12918_5436# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1586 vdd a_19166_5774# a_18958_5774# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1587 a_2889_1019# a_3142_1006# a_2744_1788# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1588 a_18914_3581# a_18910_3758# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1589 a_7830_2919# a_7849_1639# a_7800_1829# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1590 a_10886_1820# a_11617_2130# a_11825_2130# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1591 a_10150_2255# a_10679_2374# a_10887_2374# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1592 a_17091_199# a_17910_4934# a_17865_4947# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1593 a_8879_3753# a_9136_3563# a_7944_3266# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1594 a_646_7884# a_433_7884# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1595 a_17976_1065# a_18960_1362# a_18915_1375# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1596 a_1585_5434# a_1372_5434# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1597 a_15521_4621# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1598 a_11514_2654# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1599 a_5175_3810# a_5702_4062# a_5910_4062# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1600 gnd d0 a_14111_767# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1601 a_4954_133# a_6738_194# a_6958_4902# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1602 a_5910_7925# a_5489_7925# a_5173_7806# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1603 a_6640_7681# a_6427_7681# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1604 a_8880_9091# a_9133_9078# a_7941_8781# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1605 a_1372_5434# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 gnd d0 a_14108_6282# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1607 a_17865_4947# a_17908_7146# a_17863_7159# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1608 a_9888_17# a_14663_138# a_14985_138# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1609 a_16881_2171# a_16460_2171# a_15943_2415# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1610 a_15206_2296# a_15206_2066# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1611 a_8882_4679# a_9135_4666# a_7943_4369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1612 a_3819_8673# a_4076_8483# a_2881_8917# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1613 a_436_1266# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1614 vdd d0 a_9132_8524# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1615 a_119_2666# a_647_2918# a_855_2918# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1616 gnd d1 a_18225_8773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1617 a_10887_2374# a_11617_2130# a_11825_2130# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1618 a_5702_6822# a_5489_6822# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1619 vdd d0 a_14110_1870# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1620 vdd d0 a_14112_1321# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1621 vdd d1 a_13170_6526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1622 a_10883_8438# a_10462_8438# a_10147_8643# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1623 a_15205_5605# a_15734_5724# a_15942_5724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1624 a_16814_1579# a_16601_1579# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1625 a_6738_194# d5 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1626 a_15206_2525# a_15206_2296# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1627 a_8878_5959# a_9135_5769# a_7943_5472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1628 a_5704_3513# a_5491_3513# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1629 a_6427_7681# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1630 a_7834_4942# a_7877_7141# a_7828_7331# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1631 a_5702_4062# a_5489_4062# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1632 vdd d1 a_13171_5423# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1633 a_17974_5477# a_18958_5774# a_18909_5964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1634 a_6850_3269# a_6429_3269# a_5912_3513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1635 a_16897_2814# a_16600_3785# a_16880_4377# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1636 a_5704_753# a_5491_753# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1637 gnd d0 a_9137_1357# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1638 a_3827_3535# a_4080_3522# a_2888_3225# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1639 gnd d0 a_9135_1906# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1640 vdd d1 a_18228_3258# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1641 gnd a_18225_8773# a_18017_8773# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1642 gnd d1 a_8195_7665# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1643 gnd a_3139_6521# a_2931_6521# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1644 gnd d0 a_9134_5215# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1645 vdd a_13170_6526# a_12962_6526# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1646 a_14663_138# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1647 a_15733_5170# a_15520_5170# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1648 a_2886_7637# a_3139_7624# a_2741_8406# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1649 a_3825_5187# a_4078_5174# a_2883_5608# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1650 a_7830_5119# a_7879_2729# a_7834_2742# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1651 a_6643_1063# a_6430_1063# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1652 vdd a_13171_5423# a_12963_5423# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1653 a_8876_7611# a_8881_6885# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1654 a_7942_6575# a_8926_6872# a_8881_6885# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1655 a_12772_8411# a_13029_8221# a_12807_7118# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1656 a_433_4021# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1657 a_10883_8438# a_11614_8748# a_11822_8748# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1658 a_8881_4125# a_8877_4302# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1659 a_854_7884# a_433_7884# a_117_7994# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1660 vdd a_18227_5464# a_18019_5464# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1661 a_6570_1574# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1662 gnd a_8195_7665# a_7987_7665# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1663 gnd a_8198_1047# a_7990_1047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1664 gnd a_3031_2688# a_2823_2688# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1665 a_118_4456# a_647_4575# a_855_4575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1666 vdd d1 a_8197_2150# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1667 a_118_5975# a_645_6227# a_853_6227# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1668 a_5491_3513# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1669 a_13858_3540# a_14111_3527# a_12919_3230# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1670 a_2882_6711# a_3869_6277# a_3820_6467# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1671 a_15206_2066# a_15207_1609# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1672 vdd a_9135_3009# a_8927_3009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1673 vdd a_18086_6056# a_17878_6056# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1674 a_16890_4907# a_16781_4907# a_16989_4907# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1675 a_5491_753# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1676 a_10885_7889# a_11615_7645# a_11823_7645# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1677 gnd a_9137_1357# a_8929_1357# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1678 a_15733_5170# a_15520_5170# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1679 a_16812_5991# a_16599_5991# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1680 a_2746_6023# a_2931_6521# a_2886_6534# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1681 a_6429_3269# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1682 a_6847_8784# a_6780_8192# a_6864_7221# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1683 a_16460_2171# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1684 a_5910_7925# a_5489_7925# a_5173_8035# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1685 vdd d1 a_3142_1006# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1686 a_5912_753# a_6643_1063# a_6851_1063# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1687 a_2742_6200# a_2932_5418# a_2887_5431# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1688 a_13851_9232# a_14108_9042# a_12916_8745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1689 a_3823_3712# a_3826_2981# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1690 a_13853_4820# a_14110_4630# a_12918_4333# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1691 a_11823_6542# a_11402_6542# a_10884_6232# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1692 a_2774_5078# a_2823_2688# a_2774_2878# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1693 gnd a_9136_3563# a_8928_3563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1694 gnd a_9134_4112# a_8926_4112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1695 gnd a_19167_2465# a_18959_2465# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1696 a_16570_2695# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1697 a_118_4685# a_647_4575# a_855_4575# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1698 vdd a_8196_4356# a_7988_4356# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1699 a_11542_8156# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1700 a_10886_1820# a_10465_1820# a_10150_2025# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1701 a_15940_9033# a_15519_9033# a_15203_8914# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1702 a_11401_8748# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1703 a_7940_3443# a_8927_3009# a_8882_3022# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1704 a_11834_7066# a_11543_5950# a_11824_5439# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1705 a_15941_4067# a_16672_4377# a_16880_4377# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1706 a_1895_153# a_1682_153# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1707 a_5703_5719# a_5490_5719# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1708 a_15941_7930# a_15520_7930# a_15204_7811# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1709 a_9888_17# a_14663_138# a_12134_158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1710 gnd a_3141_2109# a_2933_2109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1711 a_16880_5480# a_16459_5480# a_15941_5170# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1712 a_6859_4902# a_6539_2690# a_6861_2690# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1713 a_17972_8786# a_18956_9083# gnd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1714 a_1793_4331# a_1372_4331# a_854_4021# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1715 a_3822_2055# a_4079_1865# a_2884_2299# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1716 vdd a_9135_4666# a_8927_4666# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1717 gnd d2 a_3001_1598# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1718 gnd a_4079_2968# a_3871_2968# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1719 vdd d0 a_19163_8529# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1720 a_12917_6539# a_13901_6836# a_13852_7026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1721 a_5175_3394# a_5175_3164# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1722 a_5174_6016# a_5701_6268# a_5909_6268# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1723 a_13854_3717# a_13857_2986# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1724 a_15733_6827# a_15520_6827# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1725 a_6738_194# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1726 a_10465_2923# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1727 a_1792_7640# a_1724_8151# a_1808_7180# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1728 a_15736_1312# a_15523_1312# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1729 a_12805_5083# a_12854_2693# a_12805_2883# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1730 a_7944_3266# a_8928_3563# a_8879_3753# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1731 a_7939_4546# a_8926_4112# a_8877_4302# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1732 a_8881_7988# a_9134_7975# a_7942_7678# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1733 vdd d0 a_19167_808# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1734 a_15205_4272# a_15733_4067# a_15941_4067# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1735 a_10888_1271# a_10467_1271# a_10151_1152# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1736 gnd d0 a_19164_6323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1737 a_10886_1820# a_10465_1820# a_10151_1568# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1738 a_13854_8501# a_14107_8488# a_12912_8922# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1739 a_16672_4377# a_16459_4377# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1740 vdd a_4078_4071# a_3870_4071# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1741 a_2748_1611# a_2933_2109# a_2884_2299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1742 gnd d1 a_18226_7670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1743 gnd d0 a_19165_5220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1744 a_7798_6241# a_7988_5459# a_7943_5472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1745 gnd d2 a_2998_8216# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1746 a_11824_4336# a_11403_4336# a_10885_4026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1747 a_11841_2773# a_11544_3744# a_11825_3233# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1748 a_7943_4369# a_8927_4666# a_8882_4679# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1749 gnd d2 a_13032_1603# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1750 a_119_2666# a_119_2479# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1751 a_15206_3628# a_15735_3518# a_15943_3518# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1752 gnd a_14110_2973# a_13902_2973# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1753 a_2884_3402# a_3871_2968# a_3822_3158# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1754 a_12913_7819# a_13170_7629# a_12772_8411# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1755 vdd d2 a_2999_6010# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1756 gnd a_19164_6323# a_18956_6323# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1757 a_2774_2878# a_2793_1598# a_2748_1611# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1758 vdd a_13173_1011# a_12965_1011# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1759 a_6430_1063# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1760 gnd d0 a_14111_2424# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1761 gnd a_18226_7670# a_18018_7670# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1762 gnd a_19165_5220# a_18957_5220# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1763 a_10148_7770# a_10677_7889# a_10885_7889# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1764 a_1808_4980# a_1481_7061# a_1803_7061# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1765 a_15733_4067# a_15520_4067# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1766 a_16881_3274# a_16460_3274# a_15942_2964# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1767 a_17832_8275# a_18017_8773# a_17968_8963# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1768 a_4845_133# a_4632_133# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1769 a_17975_2168# a_18228_2155# a_17835_1657# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1770 a_10465_4580# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1771 vdd a_14109_4076# a_13901_4076# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1772 a_2883_4505# a_3870_4071# a_3825_4084# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1773 a_16895_5026# a_16781_4907# a_16989_4907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1774 a_1794_2125# a_1727_1533# a_1805_2649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1775 gnd d2 a_8054_8257# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1776 vdd d0 a_19167_2465# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1777 gnd d3 a_13060_7105# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1778 a_857_1266# a_436_1266# a_120_1376# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1779 gnd d1 a_18227_4361# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1780 a_12776_8234# a_12961_8732# a_12916_8745# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1781 a_6848_7681# a_6780_8192# a_6864_7221# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1782 a_12913_6716# a_13900_6282# a_13855_6295# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1783 a_8878_4856# a_8881_4125# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1784 vdd d0 a_9133_9078# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1785 a_5909_9028# a_6639_8784# a_6847_8784# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1786 a_8875_8714# a_9132_8524# a_7937_8958# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1787 a_12915_3407# a_13902_2973# a_13853_3163# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1788 a_11834_7066# a_11543_5950# a_11823_6542# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1789 gnd a_13172_2114# a_12964_2114# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1790 a_853_8987# a_1583_8743# a_1791_8743# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1791 a_433_7884# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1792 vdd d0 a_14109_7939# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1793 a_15941_7930# a_15520_7930# a_15204_8040# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1794 a_16880_5480# a_16459_5480# a_15942_5724# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1795 a_10884_8992# a_10463_8992# a_10147_9102# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1796 gnd a_4078_7934# a_3870_7934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1797 a_11823_6542# a_11402_6542# a_10885_6786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1798 a_12805_2883# a_12824_1603# a_12779_1616# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1799 a_2772_7290# a_3029_7100# a_2778_4901# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1800 a_12775_1793# a_12965_1011# a_12920_1024# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1801 vout a_9566_17# a_5053_133# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1802 a_18910_3758# a_19167_3568# a_17975_3271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1803 a_18908_4307# a_19165_4117# a_17970_4551# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1804 a_15940_9033# a_15519_9033# a_15203_9143# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1805 gnd d0 a_9134_6872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1806 a_11401_8748# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1807 a_855_5678# a_434_5678# a_118_5559# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1808 a_646_7884# a_433_7884# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1809 gnd d0 a_4078_6831# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1810 a_10465_4580# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1811 a_16781_4907# a_16568_4907# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1812 a_1585_5434# a_1372_5434# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1813 a_11615_7645# a_11402_7645# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1814 a_12914_4510# a_13901_4076# a_13856_4089# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1815 a_17970_5654# a_18957_5220# a_18912_5233# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1816 a_1727_1533# a_1514_1533# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1817 a_11825_2130# a_11758_1538# a_11836_2654# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1818 a_7942_7678# a_8195_7665# a_7797_8447# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1819 a_17863_7159# a_17877_8262# a_17832_8275# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1820 vdd a_14109_7939# a_13901_7939# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1821 a_5173_6473# a_5174_6016# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1822 a_3826_2981# a_3822_3158# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1823 a_15734_5724# a_15521_5724# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1824 a_15943_758# a_15522_758# a_15207_963# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1825 a_3826_5741# a_4079_5728# a_2887_5431# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1826 vdd d2 a_8055_6051# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1827 a_11755_8156# a_11542_8156# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1828 a_1793_4331# a_1372_4331# a_855_4575# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1829 a_10886_5683# a_11616_5439# a_11824_5439# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1830 a_12773_6205# a_12963_5423# a_12914_5613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1831 a_854_4021# a_433_4021# a_119_3769# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1832 a_856_3472# a_1586_3228# a_1794_3228# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1833 a_15520_6827# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1834 a_12803_7295# a_12822_6015# a_12773_6205# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1835 a_6864_5021# a_6537_7102# a_6859_7102# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1836 a_16568_4907# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1837 a_8881_7988# a_8877_8165# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1838 a_18913_4684# a_19166_4671# a_17974_4374# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1839 a_15205_6021# a_15732_6273# a_15940_6273# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1840 a_1372_5434# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1841 a_11402_7645# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1842 a_18908_7067# a_18911_6336# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1843 a_6539_2690# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1844 a_648_3472# a_435_3472# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1845 a_7939_4546# a_8196_4356# a_7803_3858# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1846 a_6567_8192# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1847 gnd d3 a_8087_2729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1848 vdd d3 a_13062_2693# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1849 gnd d1 a_3140_5418# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1850 a_11758_1538# a_11545_1538# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1851 a_1513_3739# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1852 gnd d0 a_4078_4071# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1853 gnd d2 a_18085_8262# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1854 a_13857_2986# a_13853_3163# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1855 a_15206_2712# a_15206_2525# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1856 a_11841_2773# a_11544_3744# a_11824_4336# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1857 a_11824_4336# a_11403_4336# a_10886_4580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1858 a_10149_4461# a_10149_4231# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1859 a_852_8433# a_431_8433# a_117_8181# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1860 a_3821_5364# a_3826_4638# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1861 a_5175_3623# a_5175_3394# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1862 vdd a_4077_7380# a_3869_7380# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1863 vdd d1 a_13172_3217# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1864 gnd d1 a_18228_3258# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1865 a_1902_4861# a_1481_4861# a_1803_4861# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1866 a_10885_5129# a_10464_5129# a_10149_5334# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1867 a_16674_1068# a_16461_1068# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1868 a_5911_5719# a_5490_5719# a_5174_5600# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1869 a_13855_7398# a_14108_7385# a_12913_7819# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1870 vdd d1 a_8194_8768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1871 a_18910_998# a_15209_864# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1872 a_10679_3477# a_10466_3477# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1873 a_18912_4130# a_18908_4307# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1874 gnd a_2999_6010# a_2791_6010# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1875 gnd a_18118_4934# a_17910_4934# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1876 vdd d0 a_4077_6277# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1877 a_4845_133# a_4632_133# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1878 a_8880_7434# a_8876_7611# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1879 a_16601_1579# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1880 a_11839_7185# a_11725_7066# a_11839_4985# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1881 a_1795_1022# a_1727_1533# a_1805_2649# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1882 a_10676_7335# a_10463_7335# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1883 gnd d0 a_19166_1911# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1884 gnd d0 a_19168_1362# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1885 a_11543_5950# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1886 gnd a_8087_2729# a_7879_2729# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1887 a_2743_3994# a_3000_3804# a_2778_2701# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1888 a_15522_3518# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1889 a_15520_4067# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1890 a_11545_1538# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1891 vdd a_19166_3014# a_18958_3014# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1892 a_5908_8474# a_6639_8784# a_6847_8784# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1893 vdd a_8194_8768# a_7986_8768# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1894 a_15522_758# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1895 a_852_8433# a_1583_8743# a_1791_8743# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1896 a_15940_9033# a_16670_8789# a_16878_8789# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1897 gnd a_9135_3009# a_8927_3009# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1898 a_5173_6703# a_5702_6822# a_5910_6822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1899 a_15943_2415# a_15522_2415# a_15206_2296# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1900 a_17828_8452# a_18018_7670# a_17969_7860# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1901 a_10463_7335# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1902 a_2004_153# a_2823_4888# a_2774_5078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1903 a_5175_3164# a_5175_2707# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1904 a_5908_8474# a_5487_8474# a_5173_8222# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1905 gnd d0 a_19165_6877# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1906 a_13855_9055# a_14108_9042# a_12916_8745# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1907 a_1727_1533# a_1514_1533# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1908 a_11826_1027# a_11758_1538# a_11836_2654# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1909 a_5910_7925# a_6640_7681# a_6848_7681# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1910 vdd a_9133_7421# a_8925_7421# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1911 gnd a_19165_4117# a_18957_4117# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1912 a_10887_717# a_11618_1027# a_11826_1027# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1913 a_10151_1152# a_10680_1271# a_10888_1271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1914 a_15204_6478# a_15205_6021# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1915 a_2745_8229# a_2998_8216# a_2776_7113# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1916 a_16890_4907# a_16570_2695# a_16897_2814# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1917 a_1803_7061# a_1512_5945# a_1793_5434# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1918 a_17971_3448# a_18958_3014# a_18913_3027# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1919 a_1583_8743# a_1370_8743# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1920 vdd a_18228_2155# a_18020_2155# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1921 a_17830_4040# a_18020_3258# a_17975_3271# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1922 a_7940_3443# a_8927_3009# a_8878_3199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1923 a_16895_5026# a_16568_7107# a_16890_7107# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1924 a_13853_5923# a_14110_5733# a_12918_5436# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1925 gnd a_19165_6877# a_18957_6877# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1926 a_12809_4906# a_12852_7105# a_12803_7295# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1927 a_8878_2096# a_9135_1906# a_7940_2340# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1928 vdd a_19166_4671# a_18958_4671# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1929 a_6567_8192# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1930 a_1481_7061# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1931 a_855_2918# a_434_2918# a_119_2666# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1932 vdd a_8056_3845# a_7848_3845# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1933 a_16598_8197# d2 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1934 a_853_7330# a_432_7330# a_117_7535# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1935 a_10885_6786# a_10464_6786# a_10148_6667# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1936 a_9566_17# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1937 a_11758_1538# a_11545_1538# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1938 a_15207_1193# a_15207_963# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1939 a_1513_3739# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1940 a_17975_3271# a_18959_3568# a_18910_3758# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1941 a_17970_4551# a_18957_4117# a_18908_4307# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1942 a_10677_7889# a_10464_7889# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1943 a_434_2918# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1944 a_11616_5439# a_11403_5439# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1945 a_10680_1271# a_10467_1271# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1946 a_13851_7575# a_13856_6849# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1947 gnd d0 a_19167_808# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1948 vdd d0 a_14111_767# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1949 vdd a_4079_2968# a_3871_2968# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1950 a_10149_4231# a_10677_4026# a_10885_4026# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1951 a_646_4021# a_433_4021# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1952 a_7060_194# a_7879_4929# a_7830_5119# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1953 a_18911_6336# a_18907_6513# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1954 a_18909_5964# a_18912_5233# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1955 a_8876_9268# a_9133_9078# a_7941_8781# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1956 a_5175_3810# a_5175_3623# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1957 a_11543_5950# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1958 a_10147_8643# a_10675_8438# a_10883_8438# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1959 vdd d0 a_14108_6282# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1960 a_120_1563# a_120_1376# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1961 a_17974_4374# a_18958_4671# a_18913_4684# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1962 a_15942_5724# a_15521_5724# a_15205_5605# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1963 a_10147_9102# a_10147_8873# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1964 a_6750_4902# a_6537_4902# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1965 a_11403_5439# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1966 a_10464_7889# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1967 a_5174_4497# a_5703_4616# a_5911_4616# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1968 vdd d1 a_18225_8773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1969 vdd d0 a_19164_6323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1970 a_6859_7102# a_6568_5986# a_6849_5475# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1971 a_5175_2061# a_5703_1856# a_5911_1856# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1972 a_853_7330# a_432_7330# a_117_7078# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1973 a_6639_8784# a_6426_8784# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1974 gnd d1 a_13170_6526# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1975 a_15943_2415# a_15522_2415# a_15206_2525# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1976 a_17974_5477# a_18958_5774# a_18913_5787# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1977 a_16461_1068# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1978 a_2774_2878# a_2793_1598# a_2744_1788# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1979 a_11545_1538# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1980 a_8882_3022# a_8878_3199# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1981 vdd a_14110_2973# a_13902_2973# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1982 a_2884_3402# a_3871_2968# a_3826_2981# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1983 a_10677_4026# a_10464_4026# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1984 a_6866_2809# a_6569_3780# a_6849_4372# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1985 a_6849_4372# a_6428_4372# a_5911_4616# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1986 a_1793_5434# a_1725_5945# a_1803_7061# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1987 a_3823_3712# a_4080_3522# a_2888_3225# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1988 a_11825_3233# a_11404_3233# a_10886_2923# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1989 a_5173_7119# a_5173_6932# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1990 a_11839_4985# a_11512_7066# a_11839_7185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1991 a_15939_8479# a_16670_8789# a_16878_8789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1992 vdd a_18225_8773# a_18017_8773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1993 a_11839_4985# a_11725_4866# a_11933_4866# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1994 a_434_4575# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1995 vdd a_19164_6323# a_18956_6323# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1996 a_6537_7102# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1997 a_119_3353# a_648_3472# a_856_3472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1998 a_119_3769# a_646_4021# a_854_4021# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X1999 gnd d2 a_18087_3850# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2000 a_117_7994# a_646_7884# a_854_7884# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2001 a_2882_7814# a_3139_7624# a_2741_8406# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2002 a_3821_5364# a_4078_5174# a_2883_5608# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2003 a_18907_7616# a_19164_7426# a_17969_7860# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2004 a_15204_6708# a_15733_6827# a_15941_6827# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2005 vdd d1 a_8198_1047# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2006 vdd d0 a_14111_2424# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2007 a_120_917# a_648_712# a_856_712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2008 a_8879_3753# a_8882_3022# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2009 gnd a_13170_6526# a_12962_6526# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2010 a_18909_4861# a_18912_4130# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2011 gnd d1 a_13171_4320# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2012 gnd d1 a_18227_5464# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2013 a_15207_963# a_15209_864# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2014 a_5703_4616# a_5490_4616# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2015 a_13856_5192# a_14109_5179# a_12914_5613# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2016 a_12776_8234# a_13029_8221# a_12807_7118# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2017 a_5703_1856# a_5490_1856# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2018 a_433_7884# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2019 a_1794_3228# a_1373_3228# a_856_3472# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2020 a_15939_8479# a_15518_8479# a_15204_8227# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2021 a_5173_7806# a_5173_7576# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2022 a_5909_7371# a_6640_7681# a_6848_7681# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2023 a_2887_5431# a_3140_5418# a_2742_6200# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2024 gnd d3 a_8085_7141# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2025 a_15941_7930# a_16671_7686# a_16879_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2026 a_12805_2883# a_12824_1603# a_12775_1793# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2027 a_17832_8275# a_18085_8262# a_17863_7159# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2028 a_853_8987# a_432_8987# a_116_8868# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2029 a_12915_3407# a_13902_2973# a_13857_2986# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2030 a_13854_3717# a_14111_3527# a_12919_3230# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2031 a_12773_6205# a_13030_6015# a_12803_7295# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2032 a_1583_8743# a_1370_8743# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2033 a_2882_6711# a_3869_6277# a_3824_6290# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2034 a_6866_2809# a_6569_3780# a_6850_3269# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2035 vdd a_4078_7934# a_3870_7934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2036 a_6642_2166# a_6429_2166# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2037 a_11725_4866# a_11512_4866# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2038 a_434_4575# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2039 a_8878_2096# a_8884_1370# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2040 a_5909_7371# a_5488_7371# a_5173_7119# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2041 a_5912_3513# a_5491_3513# a_5175_3394# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2042 a_5910_4062# a_5489_4062# a_5175_3810# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2043 a_1803_4861# a_1694_4861# a_1902_4861# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2044 a_10887_717# a_10466_717# a_10151_922# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2045 a_5490_5719# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2046 a_10885_5129# a_11616_5439# a_11824_5439# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2047 gnd a_18087_3850# a_17879_3850# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2048 a_16895_7226# a_16598_8197# a_16879_7686# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2049 vdd d0 a_9134_6872# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2050 gnd a_8197_2150# a_7989_2150# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2051 a_2746_6023# a_2931_6521# a_2882_6711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2052 a_16598_8197# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2053 a_3821_7021# a_4078_6831# a_2886_6534# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2054 a_12777_6028# a_12962_6526# a_12917_6539# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2055 a_10885_6786# a_10464_6786# a_10148_6896# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2056 a_119_2479# a_648_2369# a_856_2369# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2057 a_18912_7993# a_19165_7980# a_17973_7683# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2058 a_5490_4616# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2059 a_1584_7640# a_1371_7640# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2060 a_6851_1063# a_6783_1574# a_6861_2690# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2061 a_13857_4643# a_14110_4630# a_12918_4333# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2062 a_15206_2712# a_15734_2964# a_15942_2964# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2063 vdd a_9136_3563# a_8928_3563# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2064 vdd a_9134_4112# a_8926_4112# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2065 a_1694_4861# a_1481_4861# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2066 a_12773_6205# a_12963_5423# a_12918_5436# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2067 a_1587_1022# a_1374_1022# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2068 a_5490_1856# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2069 a_5492_1307# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2070 a_17970_4551# a_18227_4361# a_17834_3863# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2071 a_7804_1652# a_7989_2150# a_7940_2340# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2072 a_8877_5405# a_9134_5215# a_7939_5649# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2073 a_3823_952# a_122_818# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2074 a_1724_8151# a_1511_8151# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2075 gnd d1 a_3138_8727# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2076 a_10150_3587# a_10150_3358# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2077 a_6428_4372# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2078 gnd a_3142_1006# a_2934_1006# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2079 a_6848_6578# a_6427_6578# a_5910_6822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2080 gnd d3 a_13062_2693# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2081 a_15734_2964# a_15521_2964# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2082 a_3819_8673# a_3825_7947# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2083 vdd d1 a_3141_2109# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2084 a_5911_1856# a_6642_2166# a_6850_2166# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2085 a_3822_4815# a_3825_4084# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2086 a_117_7078# a_117_6891# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2087 vdd d1 a_3139_6521# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2088 a_852_8433# a_431_8433# a_116_8638# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2089 a_17859_7336# a_17878_6056# a_17833_6069# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2090 a_7800_1829# a_7990_1047# a_7945_1060# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2091 a_16781_4907# a_16568_4907# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2092 gnd a_9135_4666# a_8927_4666# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2093 a_2744_1788# a_2934_1006# a_2885_1196# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2094 vdd d1 a_3140_5418# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2095 a_6639_8784# a_6426_8784# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2096 a_5487_8474# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2097 a_10887_2374# a_10466_2374# a_10150_2484# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2098 a_6783_1574# a_6570_1574# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2099 vdd a_9134_7975# a_8926_7975# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2100 a_7944_3266# a_8928_3563# a_8883_3576# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2101 a_11618_1027# a_11405_1027# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2102 a_7939_4546# a_8926_4112# a_8881_4125# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2103 a_6780_8192# a_6567_8192# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2104 a_1373_3228# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2105 a_7798_6241# a_7988_5459# a_7939_5649# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2106 a_10148_7540# a_10676_7335# a_10884_7335# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2107 a_13854_957# a_10153_823# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2108 a_11823_7645# a_11755_8156# a_11839_7185# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2109 a_11825_3233# a_11404_3233# a_10887_3477# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2110 a_7828_7331# a_7847_6051# a_7798_6241# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2111 a_645_7330# a_432_7330# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2112 a_10147_8873# a_10147_8643# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2113 a_10148_7999# a_10148_7770# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2114 vdd a_13062_2693# a_12854_2693# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2115 gnd a_18118_2734# a_17910_2734# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2116 a_15204_7124# a_15204_6937# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2117 a_7802_6064# a_7987_6562# a_7938_6752# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2118 gnd d0 a_14112_1321# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2119 gnd d0 a_14110_1870# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2120 gnd a_4080_3522# a_3872_3522# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2121 gnd a_4078_4071# a_3870_4071# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2122 a_2747_3817# a_3000_3804# a_2778_2701# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2123 a_13853_4820# a_13856_4089# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2124 a_10466_3477# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2125 vdd d4 a_18118_4934# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2126 gnd d4 a_13062_4893# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2127 a_10466_717# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2128 a_7943_4369# a_8927_4666# a_8878_4856# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2129 vdd d0 a_19168_1362# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2130 a_3828_1329# a_3824_1506# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2131 a_15204_7811# a_15204_7581# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2132 a_12035_158# a_11926_158# a_12134_158# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2133 gnd d2 a_2999_6010# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2134 vdd a_4079_4625# a_3871_4625# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2135 a_15940_7376# a_16671_7686# a_16879_7686# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2136 a_11404_3233# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2137 vdd d2 a_13030_6015# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2138 gnd d3 a_18116_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2139 vdd d2 a_18088_1644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2140 gnd a_13173_1011# a_12965_1011# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2141 a_5701_6268# a_5488_6268# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2142 a_17832_8275# a_18017_8773# a_17972_8786# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2143 a_854_7884# a_1584_7640# a_1792_7640# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2144 a_645_7330# a_432_7330# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2145 a_17861_5124# a_17910_2734# a_17861_2924# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2146 a_6851_1063# a_6430_1063# a_5912_753# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2147 a_13856_7952# a_13852_8129# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2148 gnd a_14111_3527# a_13903_3527# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2149 a_2888_3225# a_3872_3522# a_3823_3712# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2150 gnd a_14109_4076# a_13901_4076# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2151 a_15205_4731# a_15734_4621# a_15942_4621# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2152 vdd d1 a_8196_5459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2153 a_10147_9102# a_10676_8992# a_10884_8992# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2154 gnd d0 a_14109_7939# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2155 a_1483_2649# d3 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2156 a_2883_4505# a_3870_4071# a_3821_4261# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2157 a_11834_4866# a_11514_2654# a_11841_2773# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2158 a_16895_7226# a_16598_8197# a_16878_8789# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2159 a_10148_7540# a_10148_7083# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2160 gnd a_18116_7146# a_17908_7146# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2161 vdd d0 a_19165_6877# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2162 vdd a_13172_2114# a_12964_2114# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2163 a_17830_4040# a_18020_3258# a_17971_3448# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2164 a_15734_4621# a_15521_4621# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2165 a_13859_1334# a_13855_1511# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2166 a_16880_4377# a_16459_4377# a_15941_4067# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2167 a_18909_2101# a_19166_1911# a_17971_2345# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2168 a_1511_8151# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2169 a_435_3472# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2170 vdd a_14110_4630# a_13902_4630# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2171 a_118_4456# a_118_4226# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2172 a_2887_4328# a_3871_4625# a_3826_4638# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2173 vdd a_8196_5459# a_7988_5459# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2174 gnd a_14109_7939# a_13901_7939# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2175 a_10466_2374# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2176 a_12775_1793# a_12965_1011# a_12916_1201# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2177 a_17829_6246# a_18019_5464# a_17970_5654# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2178 vdd a_4077_9037# a_3869_9037# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2179 a_17969_6757# a_18956_6323# a_18907_6513# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2180 vdd a_19165_6877# a_18957_6877# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2181 vdd a_18088_1644# a_17880_1644# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2182 a_12919_3230# a_13903_3527# a_13854_3717# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2183 a_12914_4510# a_13901_4076# a_13852_4266# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2184 a_17970_5654# a_18957_5220# a_18908_5410# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2185 a_10677_7889# a_10464_7889# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2186 a_11616_5439# a_11403_5439# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2187 a_3822_5918# a_4079_5728# a_2887_5431# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2188 a_17859_7336# a_18116_7146# a_17865_4947# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2189 a_7940_3443# a_8197_3253# a_7799_4035# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2190 a_645_8987# a_432_8987# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2191 a_13855_7398# a_13851_7575# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2192 a_10148_8186# a_10675_8438# a_10883_8438# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2193 a_15207_1609# a_15207_1422# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2194 a_10150_3358# a_10150_3128# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2195 a_6780_8192# a_6567_8192# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2196 a_18913_5787# a_19166_5774# a_17974_5477# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2197 a_7832_7154# a_8085_7141# a_7834_4942# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2198 a_12918_4333# a_13902_4630# a_13857_4643# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2199 a_10464_7889# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2200 a_11403_5439# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2201 vdd d3 a_8087_2729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2202 a_3820_7570# a_3825_6844# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2203 a_15942_1861# a_15521_1861# a_15206_2066# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2204 a_15944_1312# a_15523_1312# a_15207_1422# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2205 a_3826_1878# a_4079_1865# a_2884_2299# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2206 a_2886_7637# a_3870_7934# a_3821_8124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2207 a_2103_153# a_4845_133# a_5053_133# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2208 a_6859_7102# a_6568_5986# a_6848_6578# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2209 a_2004_153# a_1895_153# a_2103_153# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2210 a_17861_2924# a_17880_1644# a_17835_1657# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2211 a_855_4575# a_1585_4331# a_1793_4331# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2212 a_5909_9028# a_5488_9028# a_5172_8909# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2213 a_11405_1027# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2214 a_14985_138# a_16769_199# a_17091_199# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2215 vdd d2 a_18085_8262# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2216 a_18913_3027# a_18909_3204# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2217 a_15205_4502# a_15205_4272# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2218 a_431_8433# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2219 a_5488_7371# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2220 a_16881_2171# a_16814_1579# a_16892_2695# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2221 a_15943_2415# a_16673_2171# a_16881_2171# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2222 a_117_7765# a_117_7535# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2223 a_5175_3394# a_5704_3513# a_5912_3513# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2224 a_13852_5369# a_13857_4643# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2225 a_15940_7376# a_15519_7376# a_15204_7581# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2226 a_12917_7642# a_13901_7939# a_13856_7952# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2227 a_18910_3758# a_18913_3027# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2228 a_5176_958# a_5704_753# a_5912_753# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2229 a_117_7765# a_646_7884# a_854_7884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2230 vdd a_14108_7385# a_13900_7385# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2231 gnd d1 a_8198_1047# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2232 a_2888_3225# a_3141_3212# a_2743_3994# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2233 a_11404_3233# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2234 a_8879_993# a_5178_859# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2235 a_5912_3513# a_6642_3269# a_6850_3269# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2236 gnd d3 a_3029_7100# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2237 a_3824_6290# a_4077_6277# a_2882_6711# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2238 a_15732_6273# a_15519_6273# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2239 a_2885_8740# a_3138_8727# a_2745_8229# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2240 vdd a_8087_2729# a_7879_2729# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2241 gnd d0 a_9133_6318# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2242 a_1483_2649# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2243 a_854_5124# a_433_5124# a_118_4872# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2244 vdd d1 a_18227_5464# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2245 a_2883_4505# a_3140_4315# a_2747_3817# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2246 a_16897_2814# a_16600_3785# a_16881_3274# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2247 a_853_8987# a_432_8987# a_116_9097# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2248 a_8875_8714# a_8881_7988# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2249 a_16673_2171# a_16460_2171# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2250 a_3824_9050# a_3820_9227# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2251 a_18909_2101# a_18915_1375# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2252 a_2883_5608# a_3140_5418# a_2742_6200# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2253 a_11926_158# a_11713_158# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2254 vdd d0 a_9135_3009# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2255 a_10150_2671# a_10678_2923# a_10886_2923# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2256 a_647_2918# a_434_2918# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2257 a_15519_6273# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2258 a_12919_3230# a_13172_3217# a_12774_3999# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2259 vdd a_18229_1052# a_18021_1052# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2260 gnd d0 a_19167_2465# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2261 a_12035_158# a_12854_4893# a_12805_5083# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2262 a_15521_4621# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2263 gnd a_9132_8524# a_8924_8524# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2264 vdd a_19165_4117# a_18957_4117# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2265 a_11823_6542# a_11756_5950# a_11834_7066# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2266 a_1792_7640# a_1371_7640# a_854_7884# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2267 a_8879_993# a_9136_803# a_7941_1237# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2268 a_855_5678# a_1585_5434# a_1793_5434# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2269 a_15521_1861# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2270 a_15523_1312# d0 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2271 a_11514_2654# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2272 a_16989_4907# a_16568_4907# a_16890_4907# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2273 a_17091_199# a_17910_4934# a_17861_5124# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2274 a_12914_4510# a_13171_4320# a_12778_3822# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2275 gnd d0 a_9136_3563# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2276 gnd d0 a_9134_4112# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2277 a_11725_7066# a_11512_7066# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2278 a_16459_4377# d1 gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2279 a_11614_8748# a_11401_8748# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2280 a_10151_1568# a_10151_1381# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2281 a_10678_2923# a_10465_2923# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2282 a_8884_1370# a_8880_1547# gnd sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2283 a_7941_8781# a_8194_8768# a_7801_8270# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2284 gnd d1 a_3141_2109# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2285 a_16890_7107# a_16599_5991# a_16880_5480# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2286 gnd a_19166_4671# a_18958_4671# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2287 a_16670_8789# a_16457_8789# gnd gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2288 a_17830_4040# a_18087_3850# a_17865_2747# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2289 a_432_7330# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2290 a_5702_6822# a_5489_6822# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2291 a_7800_1829# a_7990_1047# a_7941_1237# gnd sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2292 vdd d0 a_9135_4666# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2293 a_4954_133# a_4845_133# a_5053_133# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2294 a_10149_4461# a_10678_4580# a_10886_4580# vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
X2295 a_647_4575# a_434_4575# vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
C0 a_12777_6028# vdd 0.0273f
C1 a_15206_2525# a_15206_2296# 0.539f
C2 a_3823_2609# vdd 0.311f
C3 a_5172_8679# a_5700_8474# 0.194f
C4 a_1895_153# a_2004_153# 0.117f
C5 a_4080_762# a_3827_775# 0.125f
C6 a_15204_8227# a_15204_8040# 0.0622f
C7 a_6850_2166# vdd 0.0373f
C8 a_1795_1022# a_1374_1022# 0.0104f
C9 a_15732_9033# a_15203_9143# 0.194f
C10 a_1726_3739# a_1513_3739# 0.448f
C11 a_7801_8270# a_7986_8768# 0.231f
C12 a_13852_5369# a_13901_5179# 0.218f
C13 a_6429_2166# d1 0.0235f
C14 a_8883_2473# a_7944_2163# 0.278f
C15 a_2823_4888# a_2774_5078# 0.203f
C16 a_10678_2923# a_10886_2923# 0.3f
C17 a_6864_5021# a_6750_4902# 0.178f
C18 a_2886_6534# vdd 0.0951f
C19 a_12774_3999# vdd 0.0316f
C20 a_8882_1919# a_8879_2650# 0.0292f
C21 a_1481_7061# d3 0.0235f
C22 a_13855_9055# d0 0.00533f
C23 a_18229_1052# a_17976_1065# 0.11f
C24 a_3824_1506# a_2889_1019# 0.254f
C25 a_2793_1598# a_2744_1788# 0.22f
C26 a_6864_7221# a_6537_7102# 0.0467f
C27 a_13853_2060# a_13902_1870# 0.218f
C28 a_432_8987# a_116_9097# 0.0467f
C29 a_2884_3402# a_3141_3212# 0.0467f
C30 a_10148_7999# a_10148_7770# 0.539f
C31 a_645_7330# a_432_7330# 0.448f
C32 a_12778_3822# a_12918_4333# 0.206f
C33 a_2774_5078# vdd 0.0323f
C34 a_3869_7380# a_2882_7814# 0.283f
C35 a_17865_4947# a_17908_7146# 0.208f
C36 a_7834_4942# vdd 0.0264f
C37 a_2103_153# a_2004_153# 0.527f
C38 a_12803_7295# a_13030_6015# 0.0192f
C39 a_5173_6703# a_5910_6822# 0.426f
C40 a_117_7078# a_646_6781# 0.0185f
C41 a_856_2369# a_648_2369# 0.291f
C42 a_8878_5959# a_7939_5649# 0.112f
C43 a_645_7330# a_853_7330# 0.3f
C44 a_15941_6827# vdd 0.454f
C45 a_14108_6282# a_12913_6716# 0.0192f
C46 a_10885_4026# a_11403_4336# 0.11f
C47 a_11824_4336# a_11616_4336# 0.26f
C48 a_16890_7107# a_16781_7107# 0.117f
C49 a_16890_4907# a_16568_4907# 0.11f
C50 a_1803_4861# a_1483_2649# 0.0104f
C51 a_3822_3158# a_3872_2419# 0.011f
C52 a_5174_4726# a_5911_4616# 0.277f
C53 a_11822_8748# a_10884_8992# 0.133f
C54 a_9132_8524# vdd 0.183f
C55 a_10148_7083# vdd 0.143f
C56 a_117_7535# a_645_7330# 0.194f
C57 a_119_2020# vdd 0.312f
C58 a_16672_4377# a_16880_4377# 0.26f
C59 a_15940_6273# a_16458_6583# 0.11f
C60 a_10679_2374# a_10150_2484# 0.194f
C61 a_18957_5220# vdd 0.0325f
C62 a_10150_3128# a_10150_2671# 0.519f
C63 a_5705_1307# a_5913_1307# 0.291f
C64 a_3870_5174# a_3821_5364# 0.218f
C65 a_2823_4888# a_2883_5608# 0.0121f
C66 a_16892_2695# vdd 0.0269f
C67 a_5175_2520# a_5491_2410# 0.0467f
C68 a_10466_2374# vdd 0.178f
C69 a_11404_3233# d1 0.0235f
C70 a_3870_5174# a_4078_5174# 0.448f
C71 a_15521_4621# a_15734_4621# 0.448f
C72 a_3824_1506# vdd 0.311f
C73 a_19166_4671# a_18909_4861# 0.0467f
C74 a_5703_5719# a_5174_5829# 0.194f
C75 a_18957_5220# a_18912_5233# 0.154f
C76 a_7798_6241# vdd 0.0316f
C77 a_10151_1381# a_10678_1820# 0.011f
C78 a_15205_5834# a_15942_5724# 0.277f
C79 a_9779_17# vdd 0.0342f
C80 a_9888_17# vout 0.348f
C81 a_647_5678# a_118_5788# 0.194f
C82 a_2887_5431# a_3822_5918# 0.254f
C83 a_8926_4112# vdd 0.0325f
C84 d0 a_118_5559# 0.0138f
C85 a_8925_6318# a_8876_6508# 0.218f
C86 a_3872_2419# a_3827_2432# 0.151f
C87 a_1584_6537# vdd 0.0342f
C88 a_17835_1657# a_18020_2155# 0.231f
C89 a_120_1376# a_649_1266# 0.194f
C90 a_2883_5608# vdd 0.439f
C91 a_19167_3568# a_17975_3271# 0.0192f
C92 a_16989_4907# a_16568_4907# 0.0104f
C93 a_5704_3513# vdd 0.0342f
C94 a_6430_1063# a_5913_1307# 0.0467f
C95 a_15204_6708# a_15941_6827# 0.426f
C96 a_18909_3204# a_18914_2478# 0.0625f
C97 a_8926_7975# a_7942_7678# 0.292f
C98 a_15733_5170# a_15205_4918# 0.14f
C99 a_11618_1027# a_10888_1271# 0.219f
C100 a_10149_4690# vdd 0.323f
C101 a_13852_5369# vdd 0.314f
C102 vdd a_18908_5410# 0.314f
C103 a_19165_4117# d0 0.0233f
C104 a_16881_2171# a_15942_1861# 0.302f
C105 a_16461_1068# d1 0.0235f
C106 a_15206_3169# a_15943_3518# 0.112f
C107 a_18227_5464# vdd 0.183f
C108 a_18912_5233# a_18908_5410# 0.559f
C109 a_10679_717# a_10887_717# 0.3f
C110 a_5489_7925# a_5173_8035# 0.0467f
C111 a_3826_4638# a_4079_4625# 0.11f
C112 a_18021_1052# vdd 0.0325f
C113 a_8197_2150# a_7944_2163# 0.11f
C114 a_431_8433# d0 0.0235f
C115 a_10153_823# a_13854_957# 0.884f
C116 a_1795_1022# a_1805_2649# 0.206f
C117 a_2792_3804# a_2747_3817# 0.157f
C118 a_434_4575# a_118_4685# 0.0467f
C119 a_11544_3744# a_11825_3233# 0.11f
C120 a_853_7330# a_432_7330# 0.0104f
C121 a_15523_1312# a_15207_1193# 0.125f
C122 a_15204_7124# a_15733_6827# 0.0185f
C123 a_4080_762# vdd 0.183f
C124 a_8928_3563# a_8877_4302# 0.011f
C125 d0 a_18911_7439# 0.0138f
C126 a_856_3472# a_855_2918# 0.498f
C127 d0 a_120_1147# 0.0138f
C128 a_117_7535# a_432_7330# 0.0467f
C129 a_118_5975# a_647_5678# 0.0185f
C130 a_10886_1820# a_11825_2130# 0.302f
C131 a_16783_2695# a_16897_2814# 0.193f
C132 a_2882_6711# vdd 0.439f
C133 a_8928_2460# a_8879_2650# 0.218f
C134 a_15205_4272# a_15733_4067# 0.194f
C135 a_5702_7925# a_5489_7925# 0.448f
C136 a_854_4021# a_433_4021# 0.0104f
C137 a_8878_4856# a_9135_4666# 0.0467f
C138 a_11834_4866# a_11839_4985# 0.498f
C139 a_117_7535# a_853_7330# 0.255f
C140 a_12918_4333# a_14110_4630# 0.0192f
C141 d4 a_13062_4893# 0.0233f
C142 a_10678_4580# a_10465_4580# 0.448f
C143 a_16459_4377# a_15942_4621# 0.0467f
C144 a_13901_6836# a_13856_6849# 0.151f
C145 a_10153_823# a_10679_717# 0.187f
C146 vdd a_13854_3717# 0.311f
C147 a_8884_1370# vdd 0.135f
C148 a_14111_767# vdd 0.183f
C149 a_18912_4130# d0 0.0138f
C150 a_18956_9083# a_19164_9083# 0.448f
C151 a_4079_1865# a_3822_2055# 0.0467f
C152 a_118_5975# a_432_6227# 0.11f
C153 a_435_712# d0 0.0235f
C154 a_16897_2814# a_16673_3274# 0.0774f
C155 a_6537_4902# vdd 0.178f
C156 a_6639_8784# a_6847_8784# 0.26f
C157 a_7834_2742# a_7879_2729# 0.128f
C158 a_10150_2484# a_10886_2923# 0.155f
C159 a_17973_7683# a_17828_8452# 0.326f
C160 a_18226_6567# d1 0.0233f
C161 a_118_4685# a_855_4575# 0.277f
C162 a_7804_1652# a_7944_2163# 0.206f
C163 a_4079_1865# vdd 0.183f
C164 a_8878_2096# vdd 0.314f
C165 a_8087_4929# a_7830_5119# 0.0467f
C166 a_13857_1883# vdd 0.133f
C167 a_6859_7102# vdd 0.0269f
C168 a_10677_4026# a_10150_3774# 0.14f
C169 d0 a_3824_7393# 0.0138f
C170 a_644_8433# a_852_8433# 0.3f
C171 a_2790_8216# a_2745_8229# 0.157f
C172 a_18907_7616# vdd 0.314f
C173 a_7879_4929# a_7834_4942# 0.128f
C174 a_2745_8229# a_2930_8727# 0.231f
C175 a_18913_1924# a_18910_2655# 0.0292f
C176 a_5173_8222# vdd 0.135f
C177 a_15207_1193# a_15207_1422# 0.539f
C178 a_118_4872# d0 0.00888f
C179 a_19166_1911# a_18913_1924# 0.125f
C180 a_122_818# vdd 0.0985f
C181 a_1585_5434# a_1793_5434# 0.241f
C182 a_10677_6786# vdd 0.0342f
C183 a_5172_9138# a_5909_9028# 0.277f
C184 a_3820_7570# a_3824_7393# 0.559f
C185 a_10883_8438# a_10147_8643# 0.255f
C186 a_118_4685# vdd 0.323f
C187 d0 a_433_5124# 0.0235f
C188 a_5912_2410# a_5704_2410# 0.291f
C189 a_7988_5459# a_7943_5472# 0.181f
C190 a_10151_1568# vdd 0.135f
C191 a_15204_7811# a_15520_7930# 0.125f
C192 a_8927_1906# a_8884_1370# 0.0185f
C193 a_17908_7146# a_17863_7159# 0.128f
C194 a_18913_3027# a_19166_3014# 0.125f
C195 a_2741_8406# a_2776_7113# 0.298f
C196 a_18907_6513# a_18956_6323# 0.218f
C197 a_2931_7624# a_2741_8406# 0.251f
C198 a_2887_4328# a_2883_4505# 0.518f
C199 a_6643_1063# a_5913_1307# 0.219f
C200 a_16458_6583# a_15941_6827# 0.0467f
C201 a_15733_7930# a_15204_7811# 0.143f
C202 a_119_3123# vdd 0.312f
C203 a_11727_2654# a_11836_2654# 0.117f
C204 a_5909_7371# vdd 0.1f
C205 a_13858_3540# a_14111_3527# 0.11f
C206 a_18913_1924# d0 0.0138f
C207 a_2934_1006# a_2744_1788# 0.251f
C208 a_10151_1381# a_10151_1152# 0.539f
C209 a_8927_1906# a_8878_2096# 0.218f
C210 a_12779_1616# vdd 0.0273f
C211 a_15735_758# vdd 0.0342f
C212 a_3826_5741# a_3820_6467# 0.0622f
C213 a_5490_5719# a_5703_5719# 0.448f
C214 a_6848_6578# a_5910_6822# 0.133f
C215 a_8196_4356# a_7943_4369# 0.11f
C216 a_5172_8909# vdd 0.128f
C217 a_854_6781# vdd 0.454f
C218 a_5174_4726# a_5910_5165# 0.155f
C219 a_13171_4320# vdd 0.183f
C220 a_17865_2747# a_17910_2734# 0.128f
C221 a_19166_5774# vdd 0.183f
C222 a_7942_7678# vdd 0.0799f
C223 a_11725_4866# a_10886_4580# 0.0121f
C224 a_12917_7642# a_13856_7952# 0.278f
C225 a_10150_2484# a_10466_2374# 0.0467f
C226 a_12807_7118# vdd 0.0269f
C227 a_11826_1027# a_11758_1538# 0.146f
C228 a_1810_2768# a_1483_2649# 0.0467f
C229 a_1805_2649# a_1483_2649# 0.11f
C230 a_19164_6323# a_17969_6757# 0.0192f
C231 a_12809_4906# a_12805_5083# 0.518f
C232 a_2887_4328# a_2932_4315# 0.181f
C233 a_16895_7226# a_16890_7107# 0.464f
C234 a_17877_8262# a_17863_7159# 0.19f
C235 a_6866_2809# a_5911_2959# 0.0355f
C236 a_6568_5986# vdd 0.178f
C237 a_11542_8156# a_11823_7645# 0.11f
C238 a_17969_7860# a_19164_7426# 0.0192f
C239 a_15733_6827# vdd 0.0342f
C240 a_433_7884# d0 0.0235f
C241 a_15205_5375# a_15205_5605# 0.0292f
C242 a_5176_958# a_5913_1307# 0.112f
C243 a_15735_758# a_15943_758# 0.3f
C244 a_10150_2025# a_10678_1820# 0.194f
C245 d0 a_10466_3477# 0.0235f
C246 a_15521_5724# a_15205_5605# 0.125f
C247 a_8195_7665# a_7942_7678# 0.11f
C248 a_5909_6268# a_5910_6822# 0.498f
C249 a_120_1563# d0 0.00888f
C250 a_4080_2419# a_3872_2419# 0.448f
C251 a_3826_4638# vdd 0.146f
C252 a_15732_6273# a_15205_6021# 0.14f
C253 a_13853_3163# a_12915_3407# 0.316f
C254 a_18226_7670# a_17969_7860# 0.0467f
C255 a_16897_2814# a_16600_3785# 0.0104f
C256 a_10677_5129# vdd 0.0342f
C257 a_855_1815# vdd 0.0799f
C258 a_9134_4112# vdd 0.183f
C259 a_16895_7226# a_16878_8789# 0.14f
C260 a_6849_4372# vdd 0.0373f
C261 a_16783_2695# a_16892_2695# 0.117f
C262 a_18227_4361# a_17974_4374# 0.11f
C263 a_1793_5434# a_855_5678# 0.322f
C264 a_18909_5964# vdd 0.311f
C265 a_3138_8727# vdd 0.183f
C266 a_17877_8262# a_17828_8452# 0.22f
C267 a_16814_1579# a_16892_2695# 0.198f
C268 a_646_6781# vdd 0.0342f
C269 a_8056_3845# d2 0.0233f
C270 a_6750_4902# a_5911_4616# 0.0121f
C271 a_853_6227# a_118_5788# 0.155f
C272 a_1794_2125# vdd 0.0373f
C273 a_7877_7141# a_8085_7141# 0.448f
C274 a_18909_5964# a_18912_5233# 0.0292f
C275 a_8883_816# a_9136_803# 0.125f
C276 a_18118_2734# d3 0.0233f
C277 a_15204_6708# a_15733_6827# 0.143f
C278 a_3824_1506# a_3873_1316# 0.218f
C279 a_119_2666# vdd 0.143f
C280 a_8883_816# a_8879_993# 0.559f
C281 a_10147_8873# a_10147_9102# 0.539f
C282 a_11933_4866# a_12134_158# 0.174f
C283 a_855_4575# a_1793_4331# 0.133f
C284 a_14876_138# vdd 0.0342f
C285 a_8926_6872# a_9134_6872# 0.448f
C286 a_2823_4888# a_2004_153# 0.282f
C287 a_7834_2742# a_7803_3858# 0.206f
C288 a_18907_6513# a_18911_6336# 0.559f
C289 a_17974_5477# a_18958_5774# 0.292f
C290 a_12920_1024# a_13855_1511# 0.254f
C291 a_2886_6534# a_2931_6521# 0.181f
C292 a_7942_6575# a_8877_7062# 0.254f
C293 a_6847_8784# a_5908_8474# 0.302f
C294 d0 a_18913_3027# 0.0138f
C295 a_13857_2986# a_12915_3407# 0.426f
C296 a_3826_1878# a_2884_2299# 0.426f
C297 a_122_818# a_856_712# 1.07f
C298 a_17973_7683# a_18957_7980# 0.292f
C299 a_16461_1068# a_16882_1068# 0.0104f
C300 a_12914_4510# a_12963_4320# 0.243f
C301 a_11725_7066# a_11839_7185# 0.178f
C302 a_2884_3402# a_2933_3212# 0.219f
C303 a_12920_1024# a_13173_1011# 0.11f
C304 a_13032_1603# d2 0.0233f
C305 a_6866_2809# vdd 0.038f
C306 a_16458_7686# vdd 0.178f
C307 a_647_2918# vdd 0.0342f
C308 a_2004_153# vdd 0.0211f
C309 a_1793_4331# vdd 0.0373f
C310 a_12821_8221# a_12772_8411# 0.22f
C311 a_854_7884# vdd 0.455f
C312 a_11404_2130# d1 0.0235f
C313 a_18913_3027# a_18910_3758# 0.0292f
C314 a_13851_6472# a_13857_5746# 0.0622f
C315 a_15205_5834# a_15205_5605# 0.539f
C316 a_118_5975# a_117_6432# 0.519f
C317 a_2882_7814# vdd 0.439f
C318 a_7830_5119# a_6958_4902# 0.0189f
C319 a_10148_7540# vdd 0.312f
C320 a_1371_7640# a_1792_7640# 0.0104f
C321 a_17833_6069# a_17878_6056# 0.157f
C322 a_6570_1574# a_6850_2166# 0.0467f
C323 a_6738_194# a_6958_4902# 0.0467f
C324 a_14985_138# a_14876_138# 0.117f
C325 a_10150_3587# a_10885_4026# 0.155f
C326 a_6569_3780# a_6849_4372# 0.0467f
C327 a_16989_4907# a_16982_199# 0.178f
C328 a_8054_8257# vdd 0.183f
C329 a_11823_7645# vdd 0.0273f
C330 a_12779_1616# a_12964_2114# 0.231f
C331 a_10153_823# a_11933_4866# 0.247f
C332 a_853_6227# a_118_5975# 0.279f
C333 a_18913_5787# a_19166_5774# 0.11f
C334 a_5702_4062# a_5175_3810# 0.14f
C335 a_2103_153# a_4845_133# 0.194f
C336 a_17865_2747# a_17830_4040# 0.298f
C337 a_8880_1547# vdd 0.311f
C338 a_12776_8234# vdd 0.0273f
C339 a_17861_2924# a_18088_1644# 0.0192f
C340 a_5911_5719# a_5174_5370# 0.112f
C341 a_4078_7934# vdd 0.183f
C342 a_1794_3228# a_855_2918# 0.206f
C343 a_18960_1362# a_18909_2101# 0.011f
C344 a_15204_6478# a_15205_6021# 0.519f
C345 a_19165_7980# vdd 0.183f
C346 a_15207_963# a_15209_864# 0.519f
C347 a_15206_3399# a_15735_3518# 0.143f
C348 a_6426_8784# d1 0.0235f
C349 a_16811_8197# a_16878_8789# 0.195f
C350 a_8880_7434# a_8876_7611# 0.559f
C351 a_434_4575# a_647_4575# 0.448f
C352 a_5910_6822# a_6750_7102# 0.0126f
C353 a_10884_6232# a_10463_6232# 0.0104f
C354 a_5490_5719# d0 0.0235f
C355 a_9136_3563# d0 0.0233f
C356 a_13903_767# a_13854_957# 0.218f
C357 a_1586_3228# a_1810_2768# 0.0774f
C358 a_5175_2061# vdd 0.312f
C359 a_13854_957# a_13858_780# 0.559f
C360 a_6866_2809# a_6569_3780# 0.0104f
C361 a_10676_6232# a_10149_5980# 0.14f
C362 a_6851_1063# a_5913_1307# 0.322f
C363 a_435_2369# a_648_2369# 0.448f
C364 a_16674_1068# a_16882_1068# 0.241f
C365 a_8882_1919# d0 0.0138f
C366 a_7940_3443# a_8879_3753# 0.112f
C367 a_116_8868# a_853_8987# 0.426f
C368 a_18957_6877# a_18908_7067# 0.218f
C369 d4 a_6537_4902# 0.0235f
C370 a_8879_993# a_5178_859# 0.884f
C371 a_18909_5964# a_18913_5787# 0.539f
C372 a_1895_153# a_1902_4861# 0.178f
C373 a_3819_8673# a_3823_8496# 0.559f
C374 a_9136_2460# a_7944_2163# 0.0192f
C375 a_16568_7107# a_16890_7107# 0.11f
C376 a_5173_7806# a_5173_7576# 0.0292f
C377 a_6642_2166# a_6429_2166# 0.448f
C378 vdd a_15206_2066# 0.312f
C379 a_434_5678# a_118_5788# 0.0467f
C380 a_3139_6521# d1 0.0233f
C381 a_5488_9028# vdd 0.178f
C382 a_435_2369# d0 0.0235f
C383 a_646_4021# vdd 0.0342f
C384 a_15206_3628# a_15733_4067# 0.011f
C385 a_855_4575# a_647_4575# 0.291f
C386 a_10677_4026# vdd 0.0342f
C387 a_3870_6831# a_3820_7570# 0.011f
C388 a_8879_8537# a_9132_8524# 0.125f
C389 a_15205_5375# vdd 0.312f
C390 a_10677_7889# vdd 0.0342f
C391 a_1793_4331# a_1513_3739# 0.0467f
C392 a_12805_2883# a_12809_2706# 0.484f
C393 a_10463_8992# vdd 0.178f
C394 a_15209_864# d0 0.00888f
C395 a_6859_7102# a_6537_7102# 0.11f
C396 a_3823_2609# a_3827_2432# 0.539f
C397 a_3825_5187# vdd 0.133f
C398 a_15521_5724# vdd 0.178f
C399 a_2931_6521# a_2882_6711# 0.243f
C400 a_18228_3258# a_17971_3448# 0.0467f
C401 a_17971_3448# a_18020_3258# 0.219f
C402 a_16459_5480# a_15941_5170# 0.11f
C403 a_12035_158# a_11933_4866# 7.78f
C404 a_2103_153# a_1902_4861# 0.174f
C405 a_2774_2878# a_2744_1788# 0.14f
C406 a_647_4575# vdd 0.0342f
C407 a_7938_7855# a_8876_7611# 0.316f
C408 a_431_8433# a_852_8433# 0.0104f
C409 a_15206_2296# a_15943_2415# 0.426f
C410 a_6864_5021# a_5910_6822# 0.132f
C411 a_2998_8216# d2 0.0233f
C412 a_12962_6526# vdd 0.0325f
C413 a_15940_7376# a_16671_7686# 0.169f
C414 a_16890_4907# vdd 0.0264f
C415 a_17833_6069# a_18086_6056# 0.11f
C416 a_12914_5613# a_12809_4906# 0.0518f
C417 a_3825_6844# a_3869_7380# 0.0185f
C418 a_11544_3744# d2 0.0235f
C419 a_10885_6786# a_11839_4985# 0.132f
C420 a_12824_1603# a_12775_1793# 0.22f
C421 a_11725_7066# a_11839_4985# 0.342f
C422 a_856_3472# vdd 0.455f
C423 a_11403_5439# vdd 0.178f
C424 d2 a_18085_8262# 0.0233f
C425 a_12773_6205# a_13171_5423# 0.0192f
C426 a_17832_8275# a_18017_8773# 0.231f
C427 a_13852_4266# a_13901_4076# 0.218f
C428 a_15203_8914# a_15203_9143# 0.539f
C429 a_9133_6318# d0 0.0233f
C430 a_15206_3815# a_15735_3518# 0.0185f
C431 a_3821_4261# vdd 0.314f
C432 a_16897_2814# a_16570_2695# 0.0467f
C433 a_3869_6277# a_3820_6467# 0.218f
C434 a_6428_4372# a_6849_4372# 0.0104f
C435 a_5173_7806# d0 0.0138f
C436 a_5173_8035# vdd 0.323f
C437 a_10466_717# d0 0.0235f
C438 a_6951_194# a_7060_194# 0.117f
C439 a_11545_1538# vdd 0.178f
C440 a_10885_4026# a_10149_4231# 0.255f
C441 a_16989_4907# vdd 0.0369f
C442 a_7942_6575# vdd 0.0951f
C443 a_1511_8151# a_1791_8743# 0.0467f
C444 a_2774_5078# a_2774_2878# 0.176f
C445 a_12134_158# vdd 0.39f
C446 a_1794_2125# a_1514_1533# 0.0467f
C447 a_18229_1052# vdd 0.183f
C448 a_13852_4266# vdd 0.314f
C449 a_17865_2747# a_17861_2924# 0.484f
C450 a_10887_717# vdd 0.021f
C451 a_10149_4690# a_10886_4580# 0.277f
C452 a_10148_7999# a_10677_7889# 0.194f
C453 a_11405_1027# a_11826_1027# 0.0104f
C454 a_13855_9055# a_15203_9143# 0.036f
C455 a_11834_4866# a_11824_4336# 0.0928f
C456 a_2823_2688# a_2774_5078# 0.333f
C457 a_15205_5834# vdd 0.323f
C458 a_17834_3863# a_18227_4361# 0.0192f
C459 a_5702_7925# vdd 0.0342f
C460 a_5175_3810# d0 0.00888f
C461 a_5176_1604# a_5176_1417# 0.0622f
C462 a_2886_7637# vdd 0.0799f
C463 a_8882_5782# vdd 0.135f
C464 a_10464_5129# a_10885_5129# 0.0104f
C465 a_14111_2424# a_13858_2437# 0.11f
C466 a_17971_2345# vdd 0.439f
C467 a_14112_1321# vdd 0.183f
C468 a_3141_2109# a_2888_2122# 0.11f
C469 a_18227_4361# vdd 0.183f
C470 a_5173_6703# a_5489_6822# 0.125f
C471 vdd a_11615_7645# 0.0342f
C472 a_11542_8156# a_11839_7185# 0.0104f
C473 a_3141_2109# a_2884_2299# 0.0467f
C474 a_9133_9078# a_7941_8781# 0.0192f
C475 a_16989_4907# a_14985_138# 0.133f
C476 a_6567_8192# d2 0.0235f
C477 a_12919_2127# a_13858_2437# 0.278f
C478 a_15734_1861# a_15207_1422# 0.011f
C479 a_13060_7105# a_12809_4906# 0.0192f
C480 a_5912_2410# a_6429_2166# 0.0467f
C481 a_8926_5215# vdd 0.0325f
C482 a_19163_8529# d0 0.0233f
C483 a_5489_4062# vdd 0.178f
C484 a_7830_2919# vdd 0.0323f
C485 a_14985_138# a_12134_158# 0.498f
C486 a_16769_199# a_16982_199# 0.448f
C487 a_854_5124# a_118_5329# 0.255f
C488 a_16881_2171# vdd 0.0373f
C489 a_8056_3845# a_7848_3845# 0.448f
C490 d0 a_19166_3014# 0.0233f
C491 a_117_7994# a_646_7884# 0.194f
C492 a_117_8181# vdd 0.135f
C493 a_6641_4372# vdd 0.0342f
C494 a_7846_8257# a_7832_7154# 0.19f
C495 a_10153_823# vdd 0.0985f
C496 a_10150_3774# a_10464_4026# 0.11f
C497 a_15734_2964# a_15521_2964# 0.448f
C498 a_3140_5418# a_2883_5608# 0.0467f
C499 a_7830_5119# a_8087_2729# 0.0192f
C500 a_10149_4461# a_10149_4231# 0.0292f
C501 a_11824_5439# a_11834_7066# 0.206f
C502 a_18958_4671# a_17974_4374# 0.292f
C503 a_13172_3217# a_12919_3230# 0.11f
C504 a_5488_7371# a_5173_7119# 0.11f
C505 a_12777_6028# a_12917_6539# 0.206f
C506 a_10887_3477# a_11841_2773# 0.205f
C507 a_5173_6932# a_5910_6822# 0.277f
C508 a_6641_5475# a_5910_5165# 0.169f
C509 a_10883_8438# a_11614_8748# 0.169f
C510 a_13852_5369# a_12918_4333# 0.155f
C511 a_6958_4902# a_5178_859# 0.247f
C512 a_14111_3527# a_12919_3230# 0.0192f
C513 a_11617_2130# a_11825_2130# 0.26f
C514 a_15520_6827# vdd 0.178f
C515 a_10150_3128# a_10886_2923# 0.255f
C516 a_10884_6232# a_10148_6437# 0.255f
C517 d3 a_8087_2729# 0.0233f
C518 a_6780_8192# a_6848_7681# 0.146f
C519 a_5490_4616# a_5174_4497# 0.125f
C520 a_11841_2773# a_11825_3233# 0.348f
C521 a_11933_4866# a_11839_4985# 0.214f
C522 a_3870_7934# vdd 0.0325f
C523 a_17861_5124# vdd 0.0323f
C524 a_13856_6849# vdd 0.145f
C525 a_5489_4062# a_5174_4267# 0.0467f
C526 a_6427_6578# a_5910_6822# 0.0467f
C527 a_11615_6542# a_10885_6786# 0.195f
C528 a_17975_2168# vdd 0.0951f
C529 a_7846_8257# a_7797_8447# 0.22f
C530 a_18019_4361# a_17974_4374# 0.181f
C531 a_11617_2130# a_10886_1820# 0.169f
C532 a_19167_3568# a_18959_3568# 0.448f
C533 a_1372_5434# vdd 0.178f
C534 a_3001_1598# vdd 0.183f
C535 a_11836_2654# a_11826_1027# 0.206f
C536 a_6849_5475# a_5911_5719# 0.322f
C537 a_3823_3712# a_3826_2981# 0.0292f
C538 a_3819_8673# a_3825_7947# 0.0622f
C539 a_9133_6318# a_8880_6331# 0.125f
C540 a_13901_7939# a_13856_7952# 0.151f
C541 a_12913_6716# vdd 0.439f
C542 a_6427_7681# d1 0.0235f
C543 a_15520_6827# a_15204_6708# 0.125f
C544 a_14111_767# a_12916_1201# 0.0192f
C545 a_3823_8496# d0 0.0138f
C546 a_434_1815# a_647_1815# 0.448f
C547 a_10464_6786# a_10677_6786# 0.448f
C548 a_16570_2695# a_16892_2695# 0.11f
C549 a_4080_2419# a_3823_2609# 0.0467f
C550 a_10887_2374# vdd 0.454f
C551 a_3138_8727# a_2930_8727# 0.448f
C552 a_15205_4918# vdd 0.144f
C553 a_17972_8786# a_19164_9083# 0.0192f
C554 a_117_7994# a_117_7765# 0.539f
C555 a_18225_8773# a_17832_8275# 0.0192f
C556 a_19166_1911# d0 0.0233f
C557 a_11839_7185# vdd 0.0369f
C558 a_6851_1063# a_6850_2166# 0.504f
C559 a_15518_8479# a_15203_8684# 0.0467f
C560 a_5175_2291# vdd 0.128f
C561 a_9133_9078# vdd 0.183f
C562 a_12035_158# vdd 0.0211f
C563 a_4845_133# vdd 0.0342f
C564 a_6539_2690# a_6861_2690# 0.11f
C565 a_3031_2688# vdd 0.183f
C566 a_7834_4942# a_7060_194# 0.448f
C567 a_5704_753# a_5178_859# 0.187f
C568 a_15734_1861# a_15521_1861# 0.448f
C569 a_3001_1598# a_2793_1598# 0.448f
C570 a_18228_2155# vdd 0.183f
C571 a_5174_5600# a_5911_5719# 0.426f
C572 a_3823_3712# vdd 0.311f
C573 a_10883_8438# vdd 0.0799f
C574 a_1373_2125# vdd 0.178f
C575 a_8925_6318# a_8882_5782# 0.0185f
C576 a_18907_9273# vdd 0.311f
C577 a_13903_2424# a_13858_2437# 0.151f
C578 a_16890_4907# a_16783_2695# 0.218f
C579 a_11824_5439# a_10885_5129# 0.206f
C580 a_8878_4856# a_7939_4546# 0.112f
C581 a_7939_5649# a_7988_5459# 0.219f
C582 a_12915_2304# a_13902_1870# 0.283f
C583 a_11616_5439# vdd 0.0342f
C584 a_120_917# vdd 0.312f
C585 a_436_1266# a_649_1266# 0.448f
C586 a_4079_2968# a_2884_3402# 0.0192f
C587 a_11542_8156# a_11755_8156# 0.448f
C588 a_15941_7930# a_16879_7686# 0.322f
C589 a_16769_199# vdd 0.178f
C590 a_8883_2473# vdd 0.145f
C591 a_10149_5793# vdd 0.323f
C592 a_1682_153# d5 0.0235f
C593 a_9136_803# a_7941_1237# 0.0192f
C594 a_13171_4320# a_12918_4333# 0.11f
C595 a_12916_8745# a_13169_8732# 0.11f
C596 a_9133_9078# a_8925_9078# 0.448f
C597 a_433_4021# d0 0.0235f
C598 a_10887_3477# a_11404_3233# 0.0467f
C599 a_8879_993# a_7941_1237# 0.316f
C600 a_15205_4272# a_15205_4502# 0.0292f
C601 a_1794_3228# vdd 0.0273f
C602 a_15942_4621# a_15734_4621# 0.291f
C603 a_15518_8479# d0 0.0235f
C604 a_6850_3269# a_5911_2959# 0.206f
C605 a_18959_2465# a_18910_2655# 0.218f
C606 a_5703_1856# a_5490_1856# 0.448f
C607 a_855_4575# a_1902_4861# 0.0863f
C608 vdd a_18017_8773# 0.0325f
C609 a_3029_7100# vdd 0.183f
C610 a_5910_5165# a_5702_5165# 0.3f
C611 a_17973_7683# a_19165_7980# 0.0192f
C612 a_10147_8643# a_10148_8186# 0.519f
C613 a_8057_1639# vdd 0.183f
C614 a_2885_8740# a_3820_9227# 0.254f
C615 a_8878_5959# a_9135_5769# 0.0467f
C616 a_11404_3233# a_11825_3233# 0.0104f
C617 a_856_3472# a_1373_3228# 0.0467f
C618 a_12775_1793# vdd 0.0316f
C619 a_17971_3448# vdd 0.439f
C620 a_8876_7611# vdd 0.314f
C621 a_15736_1312# a_15523_1312# 0.448f
C622 a_2743_3994# a_2884_3402# 0.133f
C623 a_6539_2690# a_6752_2690# 0.448f
C624 a_16769_199# a_14985_138# 0.0104f
C625 a_7943_4369# a_8877_5405# 0.155f
C626 a_15205_4731# a_15205_4918# 0.0625f
C627 a_3869_6277# a_2882_6711# 0.283f
C628 a_17973_6580# a_18912_6890# 0.278f
C629 a_4079_2968# a_3871_2968# 0.448f
C630 a_4080_3522# vdd 0.183f
C631 a_8876_9268# a_7941_8781# 0.254f
C632 a_3139_7624# d1 0.0233f
C633 a_1902_4861# vdd 0.0369f
C634 a_4077_7380# a_3869_7380# 0.448f
C635 a_10883_8438# a_10148_7999# 0.155f
C636 a_2742_6200# a_2883_5608# 0.133f
C637 a_5702_6822# vdd 0.0342f
C638 a_5700_8474# a_5173_8222# 0.14f
C639 a_12805_5083# a_13062_4893# 0.0467f
C640 a_1511_8151# vdd 0.178f
C641 a_13030_6015# vdd 0.183f
C642 a_6780_8192# a_6847_8784# 0.195f
C643 a_13853_2060# a_13857_1883# 0.559f
C644 a_17831_1834# a_17976_1065# 0.326f
C645 a_16881_3274# a_15942_2964# 0.206f
C646 a_12773_6205# a_12822_6015# 0.22f
C647 a_5487_8474# vdd 0.178f
C648 a_15940_9033# vdd 0.454f
C649 a_17910_4934# a_17970_5654# 0.0121f
C650 a_19167_808# a_18914_821# 0.125f
C651 a_8194_8768# d1 0.0233f
C652 a_6641_4372# a_6428_4372# 0.448f
C653 a_8884_1370# a_7945_1060# 0.278f
C654 a_12809_4906# a_12852_7105# 0.208f
C655 a_9135_3009# vdd 0.183f
C656 a_6864_7221# a_6750_7102# 0.178f
C657 a_10884_7335# a_10885_7889# 0.498f
C658 a_648_712# vdd 0.0342f
C659 a_3871_1865# a_3826_1878# 0.154f
C660 a_3825_6844# vdd 0.145f
C661 a_16881_2171# a_16814_1579# 0.195f
C662 a_8878_2096# a_7945_1060# 0.155f
C663 a_3828_1329# a_2889_1019# 0.278f
C664 a_645_6227# a_432_6227# 0.448f
C665 a_15521_4621# vdd 0.178f
C666 a_857_1266# vdd 0.455f
C667 a_2999_6010# vdd 0.183f
C668 a_11839_4985# vdd 0.0369f
C669 a_5175_2520# a_5912_2410# 0.277f
C670 a_9888_17# a_9779_17# 0.117f
C671 d2 a_18087_3850# 0.0233f
C672 a_10149_5793# a_10465_5683# 0.0467f
C673 a_2745_8229# a_2776_7113# 0.206f
C674 a_15736_1312# a_15207_1422# 0.194f
C675 a_8880_6331# d0 0.0138f
C676 a_6850_3269# vdd 0.0273f
C677 a_11755_8156# vdd 0.0342f
C678 a_14109_5179# a_13852_5369# 0.0467f
C679 a_8198_1047# a_7941_1237# 0.0467f
C680 a_7800_1829# a_7830_2919# 0.14f
C681 a_6951_194# a_4954_133# 0.299f
C682 a_8197_2150# vdd 0.183f
C683 a_17835_1657# vdd 0.0273f
C684 a_119_2020# a_119_2250# 0.0292f
C685 a_8877_4302# a_8881_4125# 0.559f
C686 a_6848_7681# a_6847_8784# 0.498f
C687 a_10150_2484# a_10887_2374# 0.277f
C688 a_10149_5334# vdd 0.312f
C689 a_13858_2437# vdd 0.145f
C690 a_13031_3809# vdd 0.183f
C691 a_10464_4026# vdd 0.178f
C692 a_5173_7119# a_5701_7371# 0.14f
C693 a_3828_1329# a_3822_2055# 0.0622f
C694 a_116_8638# a_852_8433# 0.255f
C695 a_118_5788# vdd 0.323f
C696 a_18958_4671# vdd 0.0325f
C697 a_1584_7640# vdd 0.0342f
C698 a_120_917# a_856_712# 0.255f
C699 a_1794_3228# a_1513_3739# 0.11f
C700 d0 a_3825_7947# 0.00533f
C701 a_3828_1329# vdd 0.135f
C702 a_6850_3269# a_6429_3269# 0.0104f
C703 a_3822_2055# a_2884_2299# 0.316f
C704 a_10467_1271# a_10151_1152# 0.125f
C705 a_18907_6513# a_17969_6757# 0.316f
C706 a_13903_767# vdd 0.0325f
C707 d0 a_13855_7398# 0.0138f
C708 a_11841_2773# a_11514_2654# 0.0467f
C709 a_9137_1357# vdd 0.183f
C710 a_13901_4076# a_13858_3540# 0.0185f
C711 a_15731_8479# vdd 0.0342f
C712 a_17969_7860# vdd 0.439f
C713 a_2888_2122# vdd 0.0951f
C714 a_5176_1604# a_5703_1856# 0.14f
C715 a_11545_1538# a_11758_1538# 0.448f
C716 a_18116_7146# a_17859_7336# 0.0467f
C717 a_16890_7107# a_15941_6827# 0.28f
C718 a_2884_2299# vdd 0.439f
C719 a_13900_7385# a_13856_6849# 0.0185f
C720 a_7801_8270# a_7832_7154# 0.206f
C721 a_10462_8438# a_10675_8438# 0.448f
C722 a_13858_780# vdd 0.133f
C723 a_18019_4361# a_17834_3863# 0.231f
C724 a_3000_3804# a_2792_3804# 0.448f
C725 a_17861_5124# a_17910_2734# 0.333f
C726 a_6864_5021# a_6864_7221# 0.176f
C727 a_853_8987# a_432_8987# 0.0104f
C728 a_18019_4361# vdd 0.0325f
C729 a_7847_6051# a_7798_6241# 0.22f
C730 a_8876_9268# vdd 0.311f
C731 a_118_4456# a_118_4685# 0.539f
C732 a_15733_5170# a_15941_5170# 0.3f
C733 a_3872_3522# vdd 0.0325f
C734 a_12805_5083# a_12774_3999# 0.198f
C735 a_13858_3540# vdd 0.135f
C736 a_2883_4505# a_2932_4315# 0.243f
C737 a_18908_8170# vdd 0.311f
C738 a_7804_1652# vdd 0.0273f
C739 a_6850_3269# a_6569_3780# 0.11f
C740 a_1808_4980# vdd 0.0369f
C741 a_18116_7146# d3 0.0233f
C742 a_10149_5980# d0 0.00888f
C743 a_3824_6290# a_3820_6467# 0.559f
C744 d6 vdd 0.089f
C745 a_7938_6752# a_8877_7062# 0.112f
C746 a_7801_8270# a_7797_8447# 0.524f
C747 a_118_5975# vdd 0.135f
C748 a_2887_4328# a_4079_4625# 0.0192f
C749 a_15732_6273# a_15519_6273# 0.448f
C750 a_18907_9273# a_18910_8542# 0.0292f
C751 a_1585_5434# a_1372_5434# 0.448f
C752 a_15521_4621# a_15205_4731# 0.0467f
C753 a_18225_8773# vdd 0.183f
C754 a_18911_6336# d0 0.0138f
C755 a_15939_8479# vdd 0.0799f
C756 a_8927_3009# a_8883_2473# 0.0185f
C757 a_18958_5774# vdd 0.0325f
C758 a_2931_7624# a_3139_7624# 0.448f
C759 a_648_712# a_856_712# 0.3f
C760 a_1724_8151# a_1791_8743# 0.195f
C761 a_12807_7118# a_13029_8221# 0.0192f
C762 a_13170_6526# vdd 0.183f
C763 a_18914_821# a_18911_1552# 0.0292f
C764 a_15522_758# a_15209_864# 0.113f
C765 a_18227_5464# d1 0.0233f
C766 a_15734_2964# a_15942_2964# 0.3f
C767 a_3826_2981# a_2884_3402# 0.426f
C768 a_434_1815# a_119_2020# 0.0467f
C769 a_8925_9078# a_8876_9268# 0.218f
C770 a_16897_2814# a_16880_4377# 0.14f
C771 a_11615_6542# vdd 0.0342f
C772 a_857_1266# a_856_712# 0.498f
C773 a_10676_8992# vdd 0.0342f
C774 a_3871_4625# a_4079_4625# 0.448f
C775 a_10883_8438# a_11401_8748# 0.11f
C776 a_17971_3448# a_17975_3271# 0.518f
C777 a_3141_3212# a_2933_3212# 0.448f
C778 a_6639_8784# vdd 0.0342f
C779 a_120_1376# vdd 0.323f
C780 a_17879_3850# a_17834_3863# 0.157f
C781 a_7803_3858# a_7939_4546# 0.345f
C782 a_11841_2773# a_11544_3744# 0.0104f
C783 a_2774_5078# a_1803_4861# 0.409f
C784 a_10151_1381# a_10467_1271# 0.0467f
C785 a_12805_2883# a_12854_2693# 0.203f
C786 a_3870_4071# a_2883_4505# 0.283f
C787 a_13854_8501# d0 0.0138f
C788 a_10680_1271# a_10151_1152# 0.143f
C789 a_3825_4084# d0 0.0138f
C790 a_17879_3850# vdd 0.0325f
C791 a_18914_821# vdd 0.133f
C792 a_2821_7100# vdd 0.0325f
C793 a_15941_5170# a_15942_5724# 0.498f
C794 a_1481_7061# vdd 0.178f
C795 a_3871_2968# a_3826_2981# 0.154f
C796 a_645_6227# a_117_6432# 0.194f
C797 a_18019_5464# a_17974_5477# 0.181f
C798 a_10885_6786# a_11834_7066# 0.28f
C799 a_7944_3266# a_7799_4035# 0.326f
C800 a_2884_3402# vdd 0.439f
C801 a_11725_7066# a_11834_7066# 0.117f
C802 a_15733_7930# a_15520_7930# 0.448f
C803 a_13852_7026# a_14109_6836# 0.0467f
C804 a_117_7078# a_645_7330# 0.14f
C805 a_8927_3009# a_9135_3009# 0.448f
C806 a_15520_5170# d0 0.0235f
C807 a_11512_4866# a_11834_4866# 0.11f
C808 a_7945_1060# a_8880_1547# 0.254f
C809 a_18957_4117# a_18908_4307# 0.218f
C810 a_1794_3228# a_1373_3228# 0.0104f
C811 a_7801_8270# a_8194_8768# 0.0192f
C812 a_15204_7811# vdd 0.128f
C813 a_11542_8156# a_11822_8748# 0.0467f
C814 a_853_6227# a_645_6227# 0.3f
C815 a_1372_5434# a_855_5678# 0.0467f
C816 a_19165_5220# d0 0.0233f
C817 a_8057_1639# a_7800_1829# 0.0467f
C818 a_17861_5124# a_17830_4040# 0.198f
C819 a_8876_6508# a_8927_5769# 0.011f
C820 a_11614_8748# a_11822_8748# 0.26f
C821 a_8882_3022# a_8879_3753# 0.0292f
C822 a_15943_3518# a_15735_3518# 0.291f
C823 a_8926_5215# a_8881_5228# 0.154f
C824 a_15204_6478# a_15519_6273# 0.0467f
C825 a_17971_3448# a_17910_2734# 0.0126f
C826 a_18911_6336# a_18908_7067# 0.0292f
C827 a_5488_7371# a_5701_7371# 0.448f
C828 a_7834_2742# a_8056_3845# 0.0192f
C829 a_8197_3253# a_7799_4035# 0.0192f
C830 a_1902_4861# a_1694_4861# 0.337f
C831 d0 a_10149_5564# 0.0138f
C832 a_10147_8643# a_10884_8992# 0.112f
C833 a_8085_7141# a_7832_7154# 0.11f
C834 a_10149_4461# d0 0.0138f
C835 a_12915_2304# a_13854_2614# 0.112f
C836 a_1726_3739# a_1810_2768# 0.263f
C837 a_7828_7331# a_8055_6051# 0.0192f
C838 a_1795_1022# a_1587_1022# 0.241f
C839 a_15940_7376# a_16458_7686# 0.11f
C840 a_8882_4679# a_8926_5215# 0.0185f
C841 a_18911_6336# a_18956_6323# 0.154f
C842 a_12809_2706# a_12854_2693# 0.128f
C843 a_3821_4261# a_4078_4071# 0.0467f
C844 a_3871_2968# vdd 0.0325f
C845 a_13855_1511# a_13859_1334# 0.539f
C846 a_11933_4866# a_11713_158# 0.0467f
C847 a_10148_6667# a_10148_6896# 0.539f
C848 d0 a_5490_1856# 0.0235f
C849 a_6864_5021# a_6859_4902# 0.498f
C850 a_1694_7061# a_854_6781# 0.0126f
C851 a_4078_5174# d0 0.0233f
C852 a_8881_6885# d0 0.00533f
C853 a_10676_6232# a_10463_6232# 0.448f
C854 a_7944_3266# vdd 0.0799f
C855 a_7943_4369# a_9135_4666# 0.0192f
C856 a_5174_4726# a_5702_5165# 0.011f
C857 a_19164_9083# d0 0.0233f
C858 a_18913_5787# a_18958_5774# 0.151f
C859 a_15940_6273# a_15732_6273# 0.3f
C860 a_1793_5434# a_1512_5945# 0.11f
C861 a_2746_6023# vdd 0.0273f
C862 a_16890_4907# a_16570_2695# 0.0104f
C863 a_9888_17# a_14876_138# 0.335f
C864 a_1370_8743# a_852_8433# 0.11f
C865 a_3823_8496# a_3820_9227# 0.0292f
C866 a_12917_6539# a_12962_6526# 0.181f
C867 a_6848_6578# a_6859_7102# 0.328f
C868 a_12807_7118# a_12962_7629# 0.0267f
C869 a_12913_7819# a_13852_8129# 0.112f
C870 a_13029_8221# a_12776_8234# 0.11f
C871 a_9135_5769# a_8927_5769# 0.448f
C872 a_18118_4934# a_17091_199# 0.0192f
C873 a_12914_4510# a_13901_4076# 0.283f
C874 a_13171_4320# d1 0.0233f
C875 a_13902_2973# a_13858_2437# 0.0185f
C876 a_2887_4328# vdd 0.0988f
C877 a_10465_4580# vdd 0.178f
C878 a_3870_5174# a_2883_5608# 0.283f
C879 a_13851_7575# a_13855_7398# 0.559f
C880 a_18912_4130# a_18909_4861# 0.0292f
C881 a_117_7078# a_432_7330# 0.11f
C882 a_17970_4551# a_19165_4117# 0.0192f
C883 a_17972_1242# a_18959_808# 0.283f
C884 d0 a_15205_6021# 0.00888f
C885 a_12916_8745# a_12961_8732# 0.181f
C886 a_8197_3253# vdd 0.183f
C887 a_18910_998# a_18914_821# 0.559f
C888 a_646_4021# a_118_4226# 0.194f
C889 a_18914_3581# a_19167_3568# 0.11f
C890 a_4077_7380# vdd 0.183f
C891 a_5700_8474# a_5173_8035# 0.011f
C892 a_10151_1381# a_10680_1271# 0.194f
C893 a_6640_6578# vdd 0.0342f
C894 a_5491_753# a_5704_753# 0.448f
C895 a_7938_6752# vdd 0.439f
C896 a_13855_9055# a_14108_9042# 0.11f
C897 a_8878_3199# a_8928_2460# 0.011f
C898 a_3828_1329# a_3873_1316# 0.151f
C899 a_8880_7434# a_8925_7421# 0.154f
C900 a_13857_2986# d0 0.0138f
C901 a_117_7078# a_853_7330# 0.279f
C902 a_2998_8216# a_2741_8406# 0.0467f
C903 a_12918_5436# a_13851_6472# 0.155f
C904 a_5173_6932# a_5489_6822# 0.0467f
C905 a_17861_2924# a_17971_2345# 0.249f
C906 a_117_7078# a_117_7535# 0.519f
C907 a_15207_963# a_15522_758# 0.0467f
C908 a_12914_4510# vdd 0.439f
C909 a_15520_4067# vdd 0.178f
C910 a_5175_3394# a_5175_3164# 0.0292f
C911 a_6849_5475# a_6781_5986# 0.146f
C912 a_2823_4888# a_2778_4901# 0.128f
C913 a_10464_7889# vdd 0.178f
C914 a_5908_8474# vdd 0.0799f
C915 a_13904_1321# a_13855_1511# 0.218f
C916 a_11822_8748# vdd 0.0373f
C917 a_3871_4625# vdd 0.0325f
C918 a_2791_6010# a_2772_7290# 0.255f
C919 a_3001_1598# a_2774_2878# 0.0192f
C920 a_5913_1307# a_5176_1417# 0.277f
C921 a_16459_5480# a_15942_5724# 0.0467f
C922 a_7846_8257# a_8054_8257# 0.448f
C923 a_2887_5431# vdd 0.0799f
C924 a_16882_1068# a_16892_2695# 0.206f
C925 a_3820_6467# a_3871_5728# 0.011f
C926 a_10151_922# a_10887_717# 0.255f
C927 a_7828_7331# vdd 0.0321f
C928 a_2778_4901# vdd 0.0264f
C929 a_3138_8727# d1 0.0233f
C930 a_8926_7975# a_9134_7975# 0.448f
C931 a_6848_6578# a_6568_5986# 0.0467f
C932 a_13856_4089# a_13901_4076# 0.154f
C933 a_433_6781# a_854_6781# 0.0104f
C934 a_12916_8745# a_13855_9055# 0.278f
C935 a_9136_2460# vdd 0.183f
C936 a_119_3582# a_854_4021# 0.155f
C937 a_18118_4934# a_17865_4947# 0.11f
C938 a_10462_8438# d0 0.0235f
C939 a_14108_6282# a_13855_6295# 0.125f
C940 a_1808_4980# a_1694_4861# 0.178f
C941 a_7804_1652# a_7800_1829# 0.518f
C942 a_5174_5600# a_5174_5370# 0.0292f
C943 a_17970_4551# a_18912_4130# 0.426f
C944 a_17971_3448# a_17830_4040# 0.133f
C945 a_16598_8197# vdd 0.178f
C946 a_118_4456# a_647_4575# 0.143f
C947 a_6864_5021# a_7834_4942# 0.233f
C948 a_8877_7062# a_9134_6872# 0.0467f
C949 a_5176_1604# d0 0.00888f
C950 a_3824_6290# a_2882_6711# 0.426f
C951 a_18913_1924# a_18909_2101# 0.559f
C952 a_13850_8678# a_12912_8922# 0.316f
C953 a_18908_4307# vdd 0.314f
C954 a_8087_4929# vdd 0.183f
C955 a_17861_5124# a_17861_2924# 0.176f
C956 a_3827_3535# d0 0.00533f
C957 a_15204_6478# a_15940_6273# 0.255f
C958 a_17910_4934# a_17091_199# 0.282f
C959 a_10148_6667# a_10885_6786# 0.426f
C960 a_11405_1027# a_10887_717# 0.11f
C961 a_9136_803# vdd 0.183f
C962 a_15522_758# d0 0.0235f
C963 a_16458_7686# d1 0.0235f
C964 a_2774_2878# a_3031_2688# 0.0467f
C965 a_10153_823# a_10151_922# 0.519f
C966 a_7938_7855# a_8925_7421# 0.283f
C967 a_14663_138# vdd 0.178f
C968 a_17972_8786# a_17968_8963# 0.518f
C969 a_13856_4089# vdd 0.133f
C970 a_434_1815# a_855_1815# 0.0104f
C971 a_8879_993# vdd 0.314f
C972 a_18913_1924# a_18958_1911# 0.154f
C973 a_15521_2964# a_15942_2964# 0.0104f
C974 a_2823_2688# a_3031_2688# 0.448f
C975 a_13851_9232# a_12912_8922# 0.112f
C976 a_10678_1820# vdd 0.0342f
C977 a_1724_8151# vdd 0.0342f
C978 a_434_2918# a_119_3123# 0.0467f
C979 a_13856_7952# d0 0.00533f
C980 a_12773_6205# a_12809_4906# 0.181f
C981 a_15944_1312# vdd 0.455f
C982 a_10148_7999# a_10464_7889# 0.0467f
C983 a_12917_6539# a_13856_6849# 0.278f
C984 a_10884_7335# a_10676_7335# 0.3f
C985 a_11824_4336# vdd 0.0373f
C986 a_16670_8789# vdd 0.0342f
C987 a_433_6781# a_646_6781# 0.448f
C988 a_16881_2171# a_16460_2171# 0.0104f
C989 a_13903_3527# a_13854_3717# 0.218f
C990 a_11404_2130# a_11825_2130# 0.0104f
C991 a_12920_1024# a_13859_1334# 0.278f
C992 a_13852_5369# a_12914_5613# 0.316f
C993 a_5175_3394# a_5175_3623# 0.539f
C994 a_12824_1603# a_12805_2883# 0.255f
C995 a_17973_7683# a_17969_7860# 0.518f
C996 a_8928_3563# vdd 0.0325f
C997 a_14985_138# a_14663_138# 0.11f
C998 a_9566_17# d7 0.0235f
C999 a_18910_2655# a_18914_2478# 0.539f
C1000 a_11756_5950# a_11823_6542# 0.195f
C1001 a_12913_6716# a_12917_6539# 0.518f
C1002 a_15207_1609# a_15942_1861# 0.279f
C1003 a_855_5678# a_118_5788# 0.277f
C1004 a_6859_7102# a_6750_7102# 0.117f
C1005 a_9566_17# vdd 0.178f
C1006 a_12775_1793# a_12916_1201# 0.133f
C1007 a_5172_8679# a_5909_9028# 0.112f
C1008 a_12774_3999# a_12915_3407# 0.133f
C1009 a_11404_2130# a_10886_1820# 0.11f
C1010 a_15204_8040# a_15731_8479# 0.011f
C1011 a_18957_6877# a_17973_6580# 0.292f
C1012 a_646_7884# a_433_7884# 0.448f
C1013 a_15944_1312# a_15943_758# 0.498f
C1014 a_17910_4934# a_17865_4947# 0.128f
C1015 a_117_7994# a_854_7884# 0.277f
C1016 a_8881_7988# a_7942_7678# 0.278f
C1017 a_10148_8186# vdd 0.135f
C1018 a_11836_2654# a_11545_1538# 0.0104f
C1019 a_8925_6318# a_7938_6752# 0.283f
C1020 a_15205_4502# d0 0.0138f
C1021 a_118_5329# vdd 0.312f
C1022 a_2887_4328# a_2747_3817# 0.206f
C1023 a_4081_1316# a_2889_1019# 0.0192f
C1024 a_17973_7683# a_18908_8170# 0.254f
C1025 a_5911_5719# vdd 0.455f
C1026 a_7834_4942# a_8085_7141# 0.0192f
C1027 a_16459_4377# vdd 0.178f
C1028 a_11402_6542# a_10885_6786# 0.0467f
C1029 d0 a_18914_2478# 0.00533f
C1030 a_11713_158# vdd 0.178f
C1031 a_16813_3785# vdd 0.0342f
C1032 a_7940_2340# a_8879_2650# 0.112f
C1033 a_11727_2654# a_11514_2654# 0.448f
C1034 a_13857_4643# d0 0.00533f
C1035 a_10676_6232# a_10148_6437# 0.194f
C1036 a_645_7330# vdd 0.0342f
C1037 a_12919_3230# vdd 0.0799f
C1038 a_6642_2166# a_6850_2166# 0.26f
C1039 a_8198_1047# vdd 0.183f
C1040 a_15523_1312# d0 0.0235f
C1041 a_5489_5165# a_5174_5370# 0.0467f
C1042 a_9888_17# a_12134_158# 0.714f
C1043 d0 a_14109_6836# 0.0233f
C1044 a_3826_4638# a_3870_5174# 0.0185f
C1045 a_13904_1321# a_12920_1024# 0.292f
C1046 a_12821_8221# vdd 0.0325f
C1047 a_18118_2734# vdd 0.183f
C1048 a_17091_199# a_15209_864# 0.252f
C1049 a_8883_816# a_7941_1237# 0.426f
C1050 a_7937_8958# a_8924_8524# 0.283f
C1051 a_3821_8124# a_3824_7393# 0.0292f
C1052 a_9134_7975# vdd 0.183f
C1053 a_1793_4331# a_1803_4861# 0.0928f
C1054 a_8876_9268# a_8879_8537# 0.0292f
C1055 a_13169_8732# a_12776_8234# 0.0192f
C1056 a_3822_3158# a_2888_2122# 0.155f
C1057 a_3031_4888# a_2823_4888# 0.448f
C1058 a_17831_1834# vdd 0.0316f
C1059 a_14109_7939# a_13852_8129# 0.0467f
C1060 a_4081_1316# vdd 0.183f
C1061 a_119_2666# a_434_2918# 0.11f
C1062 a_10886_5683# a_10149_5564# 0.426f
C1063 a_17908_7146# a_17969_7860# 0.0126f
C1064 a_7802_6064# a_7798_6241# 0.518f
C1065 a_15939_8479# a_15204_8040# 0.155f
C1066 a_117_6432# a_432_6227# 0.0467f
C1067 a_6864_5021# a_6537_4902# 0.0467f
C1068 a_7944_3266# a_7989_3253# 0.181f
C1069 a_19166_4671# a_18958_4671# 0.448f
C1070 a_15206_3628# a_15735_3518# 0.194f
C1071 a_15941_7930# a_16895_7226# 0.168f
C1072 a_855_2918# a_119_2479# 0.155f
C1073 a_15734_5724# a_15205_6021# 0.0185f
C1074 a_6850_2166# a_6783_1574# 0.195f
C1075 a_1793_5434# a_1725_5945# 0.146f
C1076 a_6859_7102# a_6864_5021# 0.594f
C1077 a_16881_3274# vdd 0.0273f
C1078 a_5175_2291# a_5491_2410# 0.125f
C1079 a_15940_9033# a_16457_8789# 0.0467f
C1080 a_8878_5959# a_8882_5782# 0.539f
C1081 d0 a_13859_1334# 0.00533f
C1082 a_853_6227# a_432_6227# 0.0104f
C1083 a_3031_4888# vdd 0.183f
C1084 a_3827_2432# a_2888_2122# 0.278f
C1085 a_5912_753# a_5913_1307# 0.498f
C1086 a_434_2918# a_647_2918# 0.448f
C1087 a_12772_8411# a_12913_7819# 0.133f
C1088 a_8087_4929# a_7879_4929# 0.448f
C1089 a_6861_2690# a_6859_4902# 0.206f
C1090 a_11403_5439# d1 0.0235f
C1091 a_10148_7999# a_10148_8186# 0.0622f
C1092 a_9135_1906# vdd 0.183f
C1093 a_433_7884# a_117_7765# 0.125f
C1094 a_3871_1865# a_3822_2055# 0.218f
C1095 a_11834_7066# vdd 0.0269f
C1096 a_17829_6246# a_17859_7336# 0.14f
C1097 a_1371_7640# a_854_7884# 0.0467f
C1098 a_11617_3233# vdd 0.0342f
C1099 a_7989_3253# a_8197_3253# 0.448f
C1100 a_18907_7616# a_18912_6890# 0.0625f
C1101 a_120_1563# a_647_1815# 0.14f
C1102 a_15204_6478# a_15941_6827# 0.112f
C1103 a_13903_767# a_12916_1201# 0.283f
C1104 a_3141_2109# a_2748_1611# 0.0192f
C1105 a_3871_1865# vdd 0.0325f
C1106 a_10463_8992# a_10147_9102# 0.0467f
C1107 a_13858_780# a_12916_1201# 0.426f
C1108 a_6958_4902# vdd 0.0369f
C1109 a_2776_7113# a_2882_7814# 0.423f
C1110 a_14110_1870# vdd 0.183f
C1111 a_10151_1152# vdd 0.128f
C1112 a_12912_8922# vdd 0.439f
C1113 a_7939_5649# a_7943_5472# 0.518f
C1114 a_5911_4616# a_6859_4902# 0.0518f
C1115 a_9134_6872# vdd 0.183f
C1116 a_2931_7624# a_2882_7814# 0.219f
C1117 a_18959_2465# a_18914_2478# 0.151f
C1118 a_18019_5464# a_17829_6246# 0.251f
C1119 a_2881_8917# vdd 0.439f
C1120 vdd a_432_7330# 0.178f
C1121 a_117_6662# a_854_6781# 0.426f
C1122 a_17974_4374# a_18913_4684# 0.278f
C1123 a_10149_4877# d0 0.00888f
C1124 a_11757_3744# a_11824_4336# 0.195f
C1125 a_16601_1579# vdd 0.178f
C1126 a_2774_2878# a_2884_2299# 0.249f
C1127 a_15519_7376# a_15204_7124# 0.11f
C1128 a_8883_3576# a_8926_4112# 0.0185f
C1129 a_18908_4307# a_17975_3271# 0.155f
C1130 a_853_7330# vdd 0.1f
C1131 a_18229_1052# d1 0.0233f
C1132 a_8198_1047# a_7990_1047# 0.448f
C1133 a_8927_1906# a_9135_1906# 0.448f
C1134 a_8926_6872# a_8877_7062# 0.218f
C1135 a_6426_8784# a_5909_9028# 0.0467f
C1136 a_117_7535# vdd 0.312f
C1137 a_11401_8748# a_11822_8748# 0.0104f
C1138 a_3821_7021# a_2886_6534# 0.254f
C1139 a_5700_8474# a_5487_8474# 0.448f
C1140 a_2746_6023# a_2931_6521# 0.231f
C1141 a_12919_2127# a_13172_2114# 0.11f
C1142 a_2743_3994# a_3141_3212# 0.0192f
C1143 a_17879_3850# a_17830_4040# 0.22f
C1144 a_9135_4666# d0 0.0233f
C1145 a_12915_3407# a_13854_3717# 0.112f
C1146 a_15204_8040# a_15204_7811# 0.539f
C1147 a_17861_2924# a_17835_1657# 0.347f
C1148 a_11836_2654# a_10887_2374# 0.276f
C1149 a_5175_2707# a_5175_3164# 0.519f
C1150 a_18227_4361# d1 0.0233f
C1151 a_7940_2340# a_8882_1919# 0.426f
C1152 a_15732_7376# a_15519_7376# 0.448f
C1153 a_5912_2410# a_6850_2166# 0.133f
C1154 a_6850_2166# a_6861_2690# 0.328f
C1155 a_16890_4907# a_16781_4907# 0.117f
C1156 a_7937_8958# a_7941_8781# 0.518f
C1157 a_2881_8917# a_4076_8483# 0.0192f
C1158 a_13852_8129# vdd 0.311f
C1159 a_6752_2690# a_6859_4902# 0.218f
C1160 a_10884_7335# a_10148_7083# 0.279f
C1161 a_434_5678# a_647_5678# 0.448f
C1162 a_16897_2814# a_15943_3518# 0.205f
C1163 a_5490_4616# vdd 0.178f
C1164 a_11826_1027# a_10888_1271# 0.322f
C1165 a_15206_2525# a_15943_2415# 0.277f
C1166 a_117_6662# a_646_6781# 0.143f
C1167 a_7801_8270# a_8054_8257# 0.11f
C1168 a_856_2369# a_119_2020# 0.112f
C1169 a_8087_4929# d4 0.0233f
C1170 a_10147_8873# d0 0.0138f
C1171 a_11614_8748# a_10884_8992# 0.195f
C1172 a_3822_3158# a_2884_3402# 0.316f
C1173 a_4078_5174# a_3821_5364# 0.0467f
C1174 a_7830_2919# a_7879_2729# 0.203f
C1175 a_12807_7118# a_13060_7105# 0.11f
C1176 a_16880_5480# a_15941_5170# 0.206f
C1177 a_11616_4336# vdd 0.0342f
C1178 a_16989_4907# a_16781_4907# 0.337f
C1179 a_5704_753# vdd 0.0342f
C1180 a_17975_2168# a_18909_3204# 0.155f
C1181 a_15939_8479# a_16457_8789# 0.11f
C1182 a_7942_6575# a_8195_6562# 0.11f
C1183 d0 a_10150_2671# 0.00888f
C1184 a_13852_4266# a_14109_4076# 0.0467f
C1185 a_1794_2125# a_1805_2649# 0.328f
C1186 a_10885_5129# vdd 0.104f
C1187 a_2932_5418# vdd 0.0325f
C1188 a_853_8987# a_116_8638# 0.112f
C1189 a_119_3582# a_648_3472# 0.194f
C1190 a_19165_5220# a_17970_5654# 0.0192f
C1191 a_3870_5174# a_3825_5187# 0.154f
C1192 a_15941_5170# vdd 0.104f
C1193 a_7834_2742# a_7848_3845# 0.19f
C1194 a_19163_8529# a_17968_8963# 0.0192f
C1195 a_5173_6932# a_5909_7371# 0.155f
C1196 a_11512_4866# a_11933_4866# 0.0104f
C1197 a_15521_1861# d0 0.0235f
C1198 a_2885_8740# a_2745_8229# 0.206f
C1199 a_8925_7421# vdd 0.0325f
C1200 a_1372_5434# d1 0.0235f
C1201 a_5173_6703# a_5702_6822# 0.143f
C1202 a_15734_2964# vdd 0.0342f
C1203 a_10151_1381# vdd 0.323f
C1204 a_13857_2986# a_13853_3163# 0.559f
C1205 a_15520_4067# a_15941_4067# 0.0104f
C1206 a_13857_1883# a_12915_2304# 0.426f
C1207 a_2887_5431# a_3826_5741# 0.278f
C1208 a_117_7994# a_117_8181# 0.0622f
C1209 a_853_6227# a_1371_6537# 0.11f
C1210 a_3871_2968# a_3822_3158# 0.218f
C1211 a_7987_7665# a_7938_7855# 0.219f
C1212 a_5175_3394# vdd 0.128f
C1213 a_9137_1357# a_7945_1060# 0.0192f
C1214 a_1793_4331# a_1810_2768# 0.14f
C1215 a_15942_4621# vdd 0.454f
C1216 a_12805_2883# vdd 0.0323f
C1217 a_10150_2255# d0 0.0138f
C1218 a_15519_7376# vdd 0.178f
C1219 a_5491_753# a_5178_859# 0.113f
C1220 a_853_6227# a_117_6432# 0.255f
C1221 a_10465_1820# a_10886_1820# 0.0104f
C1222 a_5175_2707# a_5703_2959# 0.14f
C1223 a_5175_2707# a_5490_2959# 0.11f
C1224 a_7988_5459# a_7798_6241# 0.251f
C1225 a_5173_7119# vdd 0.143f
C1226 a_118_4685# a_646_5124# 0.011f
C1227 a_10887_3477# a_10886_2923# 0.498f
C1228 a_11402_7645# vdd 0.178f
C1229 a_2742_6200# a_2999_6010# 0.0467f
C1230 a_8877_4302# vdd 0.314f
C1231 a_10148_6667# vdd 0.128f
C1232 a_3871_2968# a_3827_2432# 0.0185f
C1233 a_2823_2688# a_2884_3402# 0.0126f
C1234 a_435_3472# a_119_3353# 0.125f
C1235 a_3821_7021# a_2882_6711# 0.112f
C1236 a_16890_4907# a_16880_4377# 0.0928f
C1237 a_16568_4907# a_16895_5026# 0.0467f
C1238 a_12915_2304# a_12779_1616# 0.345f
C1239 a_5174_6016# a_5173_6473# 0.519f
C1240 a_9134_5215# vdd 0.183f
C1241 a_1696_2649# vdd 0.0342f
C1242 a_4080_2419# a_2888_2122# 0.0192f
C1243 a_7937_8958# vdd 0.439f
C1244 a_10465_4580# a_10886_4580# 0.0104f
C1245 a_11825_3233# a_10886_2923# 0.206f
C1246 a_4632_133# a_4845_133# 0.448f
C1247 a_10884_8992# vdd 0.454f
C1248 a_18228_2155# d1 0.0233f
C1249 a_5173_7806# a_5910_7925# 0.426f
C1250 a_5176_1604# a_5490_1856# 0.11f
C1251 a_9136_803# a_8928_803# 0.448f
C1252 a_18018_7670# a_17863_7159# 0.0267f
C1253 a_2103_153# a_5178_859# 0.0416f
C1254 a_5175_2520# a_5704_2410# 0.194f
C1255 a_8879_993# a_8928_803# 0.218f
C1256 a_12917_6539# a_13170_6526# 0.11f
C1257 a_8198_1047# a_7800_1829# 0.0192f
C1258 a_1373_2125# d1 0.0235f
C1259 a_3822_5918# vdd 0.311f
C1260 a_7830_5119# a_7799_4035# 0.198f
C1261 a_4077_6277# vdd 0.183f
C1262 a_4081_1316# a_3873_1316# 0.448f
C1263 a_8880_9091# a_7941_8781# 0.278f
C1264 a_2931_7624# a_2886_7637# 0.181f
C1265 a_15203_8684# a_15204_8227# 0.519f
C1266 a_18118_2734# a_17910_2734# 0.448f
C1267 a_10463_6232# d0 0.0235f
C1268 a_645_6227# vdd 0.0342f
C1269 a_12035_158# a_12805_5083# 0.177f
C1270 a_17969_6757# a_18908_7067# 0.112f
C1271 a_12809_2706# vdd 0.0269f
C1272 a_8878_3199# a_7940_3443# 0.316f
C1273 a_15205_4731# a_15941_5170# 0.155f
C1274 a_10884_6232# a_10149_5793# 0.155f
C1275 a_8926_6872# vdd 0.0325f
C1276 a_16881_3274# a_16673_3274# 0.241f
C1277 d4 a_3031_4888# 0.0233f
C1278 a_1808_7180# a_1792_7640# 0.348f
C1279 vout a_5053_133# 0.134f
C1280 a_18018_7670# a_17828_8452# 0.251f
C1281 a_6780_8192# vdd 0.0342f
C1282 a_16895_7226# a_16879_7686# 0.348f
C1283 a_8087_2729# vdd 0.183f
C1284 a_16880_5480# a_16459_5480# 0.0104f
C1285 a_17969_6757# a_18956_6323# 0.283f
C1286 a_13852_4266# a_13903_3527# 0.011f
C1287 a_13851_9232# a_13900_9042# 0.218f
C1288 a_5911_1856# vdd 0.0799f
C1289 a_15940_9033# a_15732_9033# 0.291f
C1290 a_1481_4861# vdd 0.178f
C1291 a_17859_7336# vdd 0.0321f
C1292 a_18909_3204# a_17971_3448# 0.316f
C1293 d0 a_18912_7993# 0.00533f
C1294 a_11402_6542# vdd 0.178f
C1295 a_15205_4731# a_15942_4621# 0.277f
C1296 a_1682_153# a_2004_153# 0.11f
C1297 a_436_1266# vdd 0.178f
C1298 a_16601_1579# a_16814_1579# 0.448f
C1299 a_1803_7061# vdd 0.0269f
C1300 a_16459_5480# vdd 0.178f
C1301 a_11826_1027# a_11825_2130# 0.504f
C1302 a_8882_3022# d0 0.0138f
C1303 a_7830_5119# vdd 0.0323f
C1304 a_12914_4510# a_12918_4333# 0.518f
C1305 a_645_8987# vdd 0.0342f
C1306 a_18019_5464# vdd 0.0325f
C1307 a_6738_194# vdd 0.178f
C1308 a_1791_8743# a_1583_8743# 0.26f
C1309 a_19166_1911# a_18909_2101# 0.0467f
C1310 a_15941_4067# a_16459_4377# 0.11f
C1311 a_15206_2296# a_15206_2066# 0.0292f
C1312 a_3868_8483# a_3819_8673# 0.218f
C1313 a_8929_1357# vdd 0.0325f
C1314 a_7834_2742# a_7940_3443# 0.392f
C1315 a_7830_2919# a_7849_1639# 0.255f
C1316 a_18913_4684# vdd 0.146f
C1317 a_15204_8227# d0 0.00888f
C1318 a_3141_3212# vdd 0.183f
C1319 d3 vdd 0.712f
C1320 a_18911_7439# a_18907_7616# 0.559f
C1321 a_7943_4369# a_7939_4546# 0.518f
C1322 a_2887_5431# a_3140_5418# 0.11f
C1323 a_19166_1911# a_18958_1911# 0.448f
C1324 a_6848_7681# vdd 0.0273f
C1325 a_855_5678# a_118_5329# 0.112f
C1326 a_16813_3785# a_16600_3785# 0.448f
C1327 a_856_3472# a_1810_2768# 0.205f
C1328 a_120_1563# a_119_2020# 0.519f
C1329 a_8927_5769# a_8882_5782# 0.151f
C1330 a_6866_2809# a_6642_3269# 0.0774f
C1331 a_5910_7925# a_5173_7576# 0.112f
C1332 a_16881_2171# a_16882_1068# 0.504f
C1333 a_2748_1611# vdd 0.0273f
C1334 a_5910_4062# a_6849_4372# 0.302f
C1335 a_10886_4580# a_11824_4336# 0.133f
C1336 a_4954_133# a_4845_133# 0.117f
C1337 a_12961_8732# a_12776_8234# 0.231f
C1338 a_15940_9033# a_16878_8789# 0.133f
C1339 a_15941_7930# a_16671_7686# 0.219f
C1340 a_15734_1861# a_15206_2066# 0.194f
C1341 a_14110_4630# d0 0.0233f
C1342 a_856_2369# a_855_1815# 0.498f
C1343 a_15519_9033# vdd 0.178f
C1344 a_12772_8411# vdd 0.0316f
C1345 a_1793_5434# a_1792_6537# 0.504f
C1346 a_119_2479# vdd 0.323f
C1347 a_1727_1533# vdd 0.0342f
C1348 a_13172_2114# vdd 0.183f
C1349 a_8880_9091# vdd 0.00337f
C1350 a_10678_4580# vdd 0.0342f
C1351 a_12775_1793# a_12965_1011# 0.251f
C1352 a_7939_5649# a_8877_5405# 0.316f
C1353 a_12807_7118# a_12852_7105# 0.128f
C1354 a_10150_2025# vdd 0.312f
C1355 a_15518_8479# a_15204_8227# 0.11f
C1356 a_8197_2150# d1 0.0233f
C1357 a_11512_4866# vdd 0.178f
C1358 a_122_818# a_435_712# 0.113f
C1359 a_856_2369# a_1794_2125# 0.133f
C1360 a_18085_8262# a_17863_7159# 0.0192f
C1361 a_16811_8197# a_16879_7686# 0.146f
C1362 a_5175_2707# a_5911_2959# 0.279f
C1363 a_853_8987# a_1370_8743# 0.0467f
C1364 a_5176_1188# vdd 0.128f
C1365 a_5488_7371# vdd 0.178f
C1366 a_16881_3274# a_16600_3785# 0.11f
C1367 a_18911_6336# a_17969_6757# 0.426f
C1368 a_2743_3994# a_2933_3212# 0.251f
C1369 a_10464_5129# vdd 0.178f
C1370 a_5701_9028# vdd 0.0342f
C1371 a_11617_2130# a_11404_2130# 0.448f
C1372 a_2793_1598# a_2748_1611# 0.157f
C1373 a_15207_1609# vdd 0.135f
C1374 a_118_4685# a_118_4872# 0.0625f
C1375 a_5700_8474# a_5908_8474# 0.3f
C1376 a_117_8181# a_644_8433# 0.14f
C1377 a_18088_1644# d2 0.0233f
C1378 a_15521_2964# vdd 0.178f
C1379 a_17973_6580# a_18908_7067# 0.254f
C1380 a_2881_8917# a_2930_8727# 0.243f
C1381 a_10884_7335# a_10148_7540# 0.255f
C1382 a_5911_4616# a_6849_4372# 0.133f
C1383 a_1902_4861# a_1803_4861# 0.814f
C1384 a_649_1266# vdd 0.0342f
C1385 a_17828_8452# a_18085_8262# 0.0467f
C1386 a_11933_4866# a_11834_4866# 0.814f
C1387 a_1808_4980# a_1694_7061# 0.342f
C1388 a_2998_8216# a_2745_8229# 0.11f
C1389 a_6567_8192# a_6864_7221# 0.0104f
C1390 a_15519_6273# d0 0.0235f
C1391 a_10678_5683# vdd 0.0342f
C1392 a_8925_9078# a_8880_9091# 0.151f
C1393 a_5174_5370# vdd 0.312f
C1394 a_10884_7335# a_11823_7645# 0.206f
C1395 a_15205_5834# a_15732_6273# 0.011f
C1396 a_10467_1271# a_10680_1271# 0.448f
C1397 a_16457_8789# a_16670_8789# 0.448f
C1398 a_8883_816# vdd 0.133f
C1399 a_8876_7611# a_9133_7421# 0.0467f
C1400 a_2883_4505# vdd 0.439f
C1401 a_17974_5477# a_17829_6246# 0.326f
C1402 a_13900_9042# vdd 0.0325f
C1403 a_9133_6318# a_8876_6508# 0.0467f
C1404 a_6781_5986# vdd 0.0342f
C1405 a_6866_2809# a_6861_2690# 0.586f
C1406 a_18958_3014# vdd 0.0325f
C1407 a_16673_2171# a_15943_2415# 0.195f
C1408 a_13855_6295# vdd 0.133f
C1409 a_7942_6575# a_7802_6064# 0.206f
C1410 a_3029_7100# a_2776_7113# 0.11f
C1411 a_854_4021# a_1793_4331# 0.302f
C1412 a_117_7765# d0 0.0138f
C1413 a_4632_133# d6 0.0235f
C1414 a_18225_8773# d1 0.0233f
C1415 a_7879_4929# a_7830_5119# 0.203f
C1416 a_2886_6534# a_3870_6831# 0.292f
C1417 a_2746_6023# a_2742_6200# 0.518f
C1418 a_5175_2707# vdd 0.143f
C1419 a_10465_1820# d0 0.0235f
C1420 a_2932_4315# vdd 0.0325f
C1421 a_10463_6232# a_10149_5980# 0.11f
C1422 a_853_8987# a_116_9097# 0.277f
C1423 a_7987_7665# vdd 0.0325f
C1424 d0 a_14108_9042# 0.0233f
C1425 a_11618_1027# a_11826_1027# 0.241f
C1426 a_4078_6831# vdd 0.183f
C1427 a_3824_9050# vdd 0.00337f
C1428 a_10463_7335# vdd 0.178f
C1429 a_19167_2465# a_18910_2655# 0.0467f
C1430 a_15939_8479# a_16878_8789# 0.302f
C1431 d1 a_13170_6526# 0.0233f
C1432 a_5174_4497# vdd 0.128f
C1433 a_11401_8748# a_10884_8992# 0.0467f
C1434 a_10884_6232# a_11615_6542# 0.169f
C1435 a_12854_4893# vdd 0.0325f
C1436 a_12914_5613# a_12035_158# 0.137f
C1437 a_3868_8483# a_3823_8496# 0.154f
C1438 a_15520_7930# vdd 0.178f
C1439 a_12774_3999# a_12964_3217# 0.251f
C1440 a_17833_6069# a_18226_6567# 0.0192f
C1441 a_7987_7665# a_8195_7665# 0.448f
C1442 a_12964_2114# a_13172_2114# 0.448f
C1443 a_8057_1639# a_7849_1639# 0.448f
C1444 a_18956_9083# a_18907_9273# 0.218f
C1445 a_5175_2061# a_5912_2410# 0.112f
C1446 a_15733_7930# vdd 0.0342f
C1447 a_6847_8784# vdd 0.0373f
C1448 a_10148_6896# a_10885_6786# 0.277f
C1449 a_1481_7061# a_1694_7061# 0.448f
C1450 a_18957_6877# a_18907_7616# 0.011f
C1451 a_12963_4320# vdd 0.0325f
C1452 a_19167_2465# d0 0.0233f
C1453 a_8196_4356# a_7939_4546# 0.0467f
C1454 a_8087_4929# a_7060_194# 0.0192f
C1455 a_6866_2809# a_6752_2690# 0.193f
C1456 a_647_5678# vdd 0.0342f
C1457 a_2887_5431# a_2742_6200# 0.326f
C1458 a_10465_5683# a_10678_5683# 0.448f
C1459 a_12773_6205# a_12777_6028# 0.518f
C1460 a_1792_6537# a_1584_6537# 0.26f
C1461 a_2742_6200# a_2778_4901# 0.181f
C1462 a_5174_4267# a_5174_4497# 0.0292f
C1463 d4 a_1481_4861# 0.0235f
C1464 a_1584_7640# a_1371_7640# 0.448f
C1465 a_5178_859# vdd 0.0974f
C1466 a_10677_4026# a_10150_3587# 0.011f
C1467 a_1481_4861# a_1694_4861# 0.448f
C1468 a_10676_8992# a_10147_9102# 0.194f
C1469 a_17861_2924# a_18118_2734# 0.0467f
C1470 a_1808_4980# a_1803_4861# 0.498f
C1471 a_857_1266# a_1374_1022# 0.0467f
C1472 a_2882_7814# a_3824_7393# 0.426f
C1473 a_3870_4071# vdd 0.0325f
C1474 a_18020_2155# vdd 0.0325f
C1475 a_15734_4621# vdd 0.0342f
C1476 a_15941_4067# a_15942_4621# 0.498f
C1477 a_12803_7295# vdd 0.0321f
C1478 a_646_4021# a_854_4021# 0.3f
C1479 a_11824_5439# vdd 0.0273f
C1480 a_17861_2924# a_17831_1834# 0.14f
C1481 a_8927_4666# vdd 0.0325f
C1482 a_432_6227# vdd 0.178f
C1483 d2 a_11543_5950# 0.0235f
C1484 a_5489_6822# d0 0.0235f
C1485 a_11727_2654# a_11841_2773# 0.193f
C1486 a_855_1815# a_120_1563# 0.279f
C1487 a_5174_5370# a_5174_4913# 0.519f
C1488 a_1583_8743# vdd 0.0342f
C1489 a_18116_7146# vdd 0.183f
C1490 a_7942_6575# a_7987_6562# 0.181f
C1491 a_10886_4580# a_11616_4336# 0.195f
C1492 a_16881_3274# a_16460_3274# 0.0104f
C1493 a_7944_2163# vdd 0.0951f
C1494 a_117_6891# a_854_6781# 0.277f
C1495 a_3822_5918# a_3826_5741# 0.539f
C1496 a_1514_1533# a_1727_1533# 0.448f
C1497 a_1794_3228# a_1810_2768# 0.348f
C1498 a_19167_3568# d0 0.0233f
C1499 a_5491_3513# a_5912_3513# 0.0104f
C1500 a_5492_1307# a_5176_1188# 0.125f
C1501 a_2883_4505# a_2747_3817# 0.345f
C1502 a_5173_6473# vdd 0.312f
C1503 d3 a_6537_7102# 0.0235f
C1504 a_13902_4630# vdd 0.0325f
C1505 a_8878_2096# a_8882_1919# 0.559f
C1506 a_8198_1047# a_7945_1060# 0.11f
C1507 a_19167_3568# a_18910_3758# 0.0467f
C1508 a_18908_4307# a_18959_3568# 0.011f
C1509 a_18959_2465# a_19167_2465# 0.448f
C1510 a_16674_1068# a_16461_1068# 0.448f
C1511 a_5172_9138# a_5172_8909# 0.539f
C1512 a_10884_7335# a_11615_7645# 0.169f
C1513 a_433_7884# a_854_7884# 0.0104f
C1514 a_13172_3217# vdd 0.183f
C1515 a_8882_3022# a_7940_3443# 0.426f
C1516 a_5489_4062# a_5910_4062# 0.0104f
C1517 a_854_5124# vdd 0.104f
C1518 a_14111_3527# vdd 0.183f
C1519 a_17833_6069# a_17969_6757# 0.345f
C1520 a_17976_1065# a_19168_1362# 0.0192f
C1521 a_7937_8958# a_8879_8537# 0.426f
C1522 a_16671_7686# a_16879_7686# 0.241f
C1523 d4 a_11512_4866# 0.0235f
C1524 a_8881_4125# vdd 0.133f
C1525 a_3142_1006# a_2885_1196# 0.0467f
C1526 a_15523_1312# a_15207_1422# 0.0467f
C1527 a_9888_17# a_14663_138# 0.0104f
C1528 a_11834_4866# vdd 0.0264f
C1529 a_6641_4372# a_5910_4062# 0.169f
C1530 a_2932_4315# a_2747_3817# 0.231f
C1531 a_8197_3253# d1 0.0233f
C1532 a_2933_3212# vdd 0.0325f
C1533 a_11725_7066# a_10885_6786# 0.0126f
C1534 a_15942_5724# a_15205_5605# 0.426f
C1535 a_2885_8740# a_3138_8727# 0.11f
C1536 vdd a_5701_7371# 0.0342f
C1537 d0 a_10148_7770# 0.0138f
C1538 a_10151_1568# a_10886_1820# 0.279f
C1539 a_5491_3513# d0 0.0235f
C1540 a_117_6891# a_646_6781# 0.194f
C1541 a_5704_3513# a_5175_3810# 0.0185f
C1542 a_13858_3540# a_13903_3527# 0.151f
C1543 a_1895_153# a_2103_153# 0.335f
C1544 a_16895_5026# vdd 0.0369f
C1545 a_7938_7855# a_8880_7434# 0.426f
C1546 a_7804_1652# a_7849_1639# 0.157f
C1547 a_15205_4731# a_15734_4621# 0.194f
C1548 a_18956_7426# a_18907_7616# 0.218f
C1549 a_7828_7331# a_7847_6051# 0.255f
C1550 a_13853_2060# a_14110_1870# 0.0467f
C1551 a_10151_922# a_10151_1152# 0.0292f
C1552 a_2932_5418# a_3140_5418# 0.448f
C1553 a_3821_8124# a_3825_7947# 0.539f
C1554 a_5704_753# a_5176_958# 0.194f
C1555 a_16895_7226# a_16781_7107# 0.178f
C1556 a_17091_199# a_17970_5654# 0.137f
C1557 a_10148_6667# a_10464_6786# 0.125f
C1558 a_119_3769# vdd 0.135f
C1559 a_118_4872# a_647_4575# 0.0185f
C1560 a_10149_5980# a_10148_6437# 0.519f
C1561 a_5703_2959# a_5175_3164# 0.194f
C1562 a_5490_2959# a_5175_3164# 0.0467f
C1563 a_13032_1603# a_12779_1616# 0.11f
C1564 a_855_4575# a_1585_4331# 0.195f
C1565 a_8881_5228# a_9134_5215# 0.125f
C1566 a_6849_5475# vdd 0.0273f
C1567 a_12821_8221# a_13029_8221# 0.448f
C1568 a_2821_7100# a_2776_7113# 0.128f
C1569 a_9888_17# a_9566_17# 0.11f
C1570 a_1793_4331# a_1372_4331# 0.0104f
C1571 a_1792_6537# a_854_6781# 0.133f
C1572 a_17974_5477# vdd 0.0799f
C1573 a_6848_6578# a_6640_6578# 0.26f
C1574 a_13899_8488# a_12912_8922# 0.283f
C1575 a_9135_5769# d0 0.0233f
C1576 a_15735_758# a_15209_864# 0.187f
C1577 a_5705_1307# a_5176_1188# 0.143f
C1578 a_6958_4902# a_7060_194# 7.78f
C1579 a_19164_7426# vdd 0.183f
C1580 a_10677_4026# a_10149_4231# 0.194f
C1581 a_3868_8483# a_3825_7947# 0.0185f
C1582 a_1585_4331# vdd 0.0342f
C1583 a_117_8181# a_431_8433# 0.11f
C1584 a_18228_3258# a_18020_3258# 0.448f
C1585 a_5911_4616# a_6641_4372# 0.195f
C1586 a_13857_4643# a_13853_4820# 0.539f
C1587 a_14108_6282# vdd 0.183f
C1588 a_8876_6508# a_7943_5472# 0.155f
C1589 a_13904_1321# a_13859_1334# 0.151f
C1590 a_13902_5733# vdd 0.0325f
C1591 a_853_8987# a_852_8433# 0.498f
C1592 a_16671_6583# vdd 0.0342f
C1593 a_2886_6534# a_2772_7290# 0.0437f
C1594 a_1371_6537# vdd 0.178f
C1595 a_18226_7670# vdd 0.183f
C1596 a_16598_8197# a_16878_8789# 0.0467f
C1597 a_2886_6534# a_3820_7570# 0.155f
C1598 a_5173_6932# a_5702_6822# 0.194f
C1599 a_17908_7146# a_17859_7336# 0.218f
C1600 a_1682_153# a_1902_4861# 0.0467f
C1601 a_5909_6268# a_6640_6578# 0.169f
C1602 a_5174_5600# vdd 0.128f
C1603 a_12919_2127# a_14111_2424# 0.0192f
C1604 a_15733_5170# vdd 0.0342f
C1605 a_12778_3822# a_12823_3809# 0.157f
C1606 a_7938_6752# a_8195_6562# 0.0467f
C1607 a_12914_4510# a_14109_4076# 0.0192f
C1608 a_5704_3513# a_5912_3513# 0.291f
C1609 a_119_3353# vdd 0.128f
C1610 a_17865_4947# a_17970_5654# 0.0518f
C1611 a_855_1815# a_1586_2125# 0.169f
C1612 a_117_6432# vdd 0.312f
C1613 a_13902_1870# a_13859_1334# 0.0185f
C1614 a_10148_7083# d0 0.00888f
C1615 a_17976_1065# a_18911_1552# 0.254f
C1616 a_9132_8524# d0 0.0233f
C1617 a_15944_1312# a_15207_1193# 0.426f
C1618 a_3826_1878# a_3822_2055# 0.559f
C1619 a_853_6227# vdd 0.0799f
C1620 a_10888_1271# a_10887_717# 0.498f
C1621 a_1794_2125# a_1586_2125# 0.26f
C1622 d0 a_10466_2374# 0.0235f
C1623 a_2778_2701# a_2792_3804# 0.19f
C1624 a_3826_1878# vdd 0.133f
C1625 a_5909_9028# a_5172_8909# 0.426f
C1626 a_8880_6331# a_8876_6508# 0.559f
C1627 a_2887_5431# a_4079_5728# 0.0192f
C1628 a_16878_8789# a_16670_8789# 0.26f
C1629 a_9135_5769# a_7943_5472# 0.0192f
C1630 a_5912_2410# a_5175_2291# 0.426f
C1631 a_1373_2125# a_856_2369# 0.0467f
C1632 a_12772_8411# a_13170_7629# 0.0192f
C1633 a_17833_6069# a_17973_6580# 0.206f
C1634 a_15942_2964# vdd 0.1f
C1635 a_435_3472# vdd 0.178f
C1636 a_19166_4671# a_18913_4684# 0.11f
C1637 a_15203_8914# a_15940_9033# 0.426f
C1638 a_5703_2959# a_5490_2959# 0.448f
C1639 a_18913_1924# a_17971_2345# 0.426f
C1640 a_12854_2693# vdd 0.0325f
C1641 a_13901_5179# a_13856_5192# 0.154f
C1642 a_8883_816# a_8928_803# 0.154f
C1643 a_17976_1065# vdd 0.0799f
C1644 a_15206_3815# a_15520_4067# 0.11f
C1645 a_16459_4377# d1 0.0235f
C1646 a_8877_8165# a_7942_7678# 0.254f
C1647 a_13856_4089# a_14109_4076# 0.125f
C1648 a_18226_6567# a_17969_6757# 0.0467f
C1649 a_10467_1271# vdd 0.178f
C1650 a_5703_1856# a_5175_2061# 0.194f
C1651 a_15522_2415# vdd 0.178f
C1652 a_10147_8643# vdd 0.312f
C1653 a_16880_5480# a_15942_5724# 0.322f
C1654 a_10678_4580# a_10886_4580# 0.291f
C1655 a_6750_4902# a_6859_4902# 0.117f
C1656 a_8198_1047# d1 0.0233f
C1657 a_17974_5477# a_18913_5787# 0.278f
C1658 a_5172_9138# a_5488_9028# 0.0467f
C1659 a_6850_3269# a_6642_3269# 0.241f
C1660 a_15519_6273# a_15205_6021# 0.11f
C1661 a_15942_5724# vdd 0.455f
C1662 a_5911_5719# a_6428_5475# 0.0467f
C1663 a_16879_6583# a_15940_6273# 0.302f
C1664 a_4080_762# d0 0.0233f
C1665 a_13851_6472# a_13900_6282# 0.218f
C1666 a_15942_1861# vdd 0.0799f
C1667 a_5490_4616# a_5703_4616# 0.448f
C1668 a_15733_5170# a_15205_4731# 0.011f
C1669 a_2776_7113# a_2778_4901# 0.206f
C1670 a_2778_2701# a_2774_5078# 0.685f
C1671 a_13901_6836# vdd 0.0325f
C1672 a_17976_1065# a_18915_1375# 0.278f
C1673 a_13854_957# vdd 0.314f
C1674 a_10148_6896# vdd 0.323f
C1675 a_5909_7371# a_5173_7576# 0.255f
C1676 a_2774_2878# a_2748_1611# 0.347f
C1677 a_16568_7107# a_16781_7107# 0.448f
C1678 a_6568_5986# d2 0.0235f
C1679 a_7943_5472# a_7798_6241# 0.326f
C1680 a_2932_5418# a_2742_6200# 0.251f
C1681 a_3825_4084# a_3822_4815# 0.0292f
C1682 a_5489_5165# vdd 0.178f
C1683 a_2882_6711# a_2772_7290# 0.285f
C1684 a_5911_2959# a_5175_3164# 0.255f
C1685 a_7941_1237# vdd 0.439f
C1686 a_3142_1006# a_2744_1788# 0.0192f
C1687 a_120_917# a_120_1147# 0.0292f
C1688 a_8882_3022# a_8878_3199# 0.559f
C1689 a_8884_1370# d0 0.00533f
C1690 a_6640_7681# a_5910_7925# 0.219f
C1691 a_4077_6277# a_3869_6277# 0.448f
C1692 a_15735_758# a_15207_963# 0.194f
C1693 a_14111_767# d0 0.0233f
C1694 a_16568_4907# vdd 0.178f
C1695 a_18118_4934# a_17861_5124# 0.0467f
C1696 a_14111_2424# a_13903_2424# 0.448f
C1697 a_15204_7581# a_15204_7811# 0.0292f
C1698 a_10679_717# vdd 0.0342f
C1699 a_14107_8488# a_12912_8922# 0.0192f
C1700 a_15204_8040# a_15520_7930# 0.0467f
C1701 a_3821_7021# a_3825_6844# 0.539f
C1702 a_4079_1865# d0 0.0233f
C1703 a_13856_5192# vdd 0.133f
C1704 a_13857_1883# d0 0.0138f
C1705 a_12919_2127# a_13903_2424# 0.292f
C1706 a_15733_7930# a_15204_8040# 0.194f
C1707 a_5173_8222# d0 0.00888f
C1708 a_434_5678# vdd 0.178f
C1709 a_16671_6583# a_16458_6583# 0.448f
C1710 a_122_818# d0 0.00888f
C1711 a_15519_7376# a_15940_7376# 0.0104f
C1712 a_3827_3535# a_2888_3225# 0.278f
C1713 a_120_917# a_435_712# 0.0467f
C1714 a_7877_7141# a_7832_7154# 0.128f
C1715 a_5176_958# a_5176_1188# 0.0292f
C1716 a_5489_7925# vdd 0.178f
C1717 a_856_3472# a_648_3472# 0.291f
C1718 a_8196_5459# vdd 0.183f
C1719 a_10151_1568# d0 0.00888f
C1720 a_855_5678# a_647_5678# 0.291f
C1721 a_8194_8768# a_7986_8768# 0.448f
C1722 a_854_5124# a_1585_5434# 0.169f
C1723 a_17865_2747# a_18087_3850# 0.0192f
C1724 a_16570_2695# d3 0.0235f
C1725 a_16458_7686# a_15941_7930# 0.0467f
C1726 a_5174_6016# vdd 0.135f
C1727 a_11825_2130# a_11545_1538# 0.0467f
C1728 a_3824_9050# a_4077_9037# 0.11f
C1729 a_10680_1271# vdd 0.0342f
C1730 a_10676_6232# a_10149_5793# 0.011f
C1731 a_11823_6542# a_11543_5950# 0.0467f
C1732 a_17833_6069# a_18018_6567# 0.231f
C1733 a_5175_3164# vdd 0.312f
C1734 a_8880_7434# vdd 0.133f
C1735 d0 a_5172_8909# 0.0138f
C1736 a_118_5559# a_118_5788# 0.539f
C1737 d0 a_19166_5774# 0.0233f
C1738 a_13857_4643# a_14110_4630# 0.11f
C1739 a_3872_762# a_2885_1196# 0.283f
C1740 a_855_2918# vdd 0.1f
C1741 a_8929_1357# a_7945_1060# 0.292f
C1742 a_7990_1047# a_7941_1237# 0.219f
C1743 a_11756_5950# a_11543_5950# 0.448f
C1744 a_7830_5119# a_7060_194# 0.177f
C1745 a_6427_7681# a_6640_7681# 0.448f
C1746 a_12822_6015# a_12777_6028# 0.157f
C1747 a_8054_8257# d2 0.0233f
C1748 a_1895_153# vdd 0.0342f
C1749 a_17973_6580# a_18226_6567# 0.11f
C1750 a_5491_753# vdd 0.178f
C1751 a_6738_194# a_7060_194# 0.11f
C1752 a_857_1266# a_120_1147# 0.426f
C1753 a_5703_2959# a_5911_2959# 0.3f
C1754 a_5490_2959# a_5911_2959# 0.0104f
C1755 a_4079_2968# a_3826_2981# 0.125f
C1756 a_13169_8732# a_12912_8922# 0.0467f
C1757 a_16811_8197# a_16895_7226# 0.263f
C1758 a_12913_7819# vdd 0.439f
C1759 a_10885_6786# vdd 0.454f
C1760 a_17861_5124# a_17910_4934# 0.203f
C1761 a_5488_9028# a_5909_9028# 0.0104f
C1762 a_11725_7066# vdd 0.0342f
C1763 a_15944_1312# a_16882_1068# 0.322f
C1764 a_3869_7380# vdd 0.0325f
C1765 a_4078_4071# a_2883_4505# 0.0192f
C1766 a_15940_6273# a_15205_6021# 0.279f
C1767 a_3826_4638# d0 0.00533f
C1768 a_16989_4907# a_15209_864# 0.247f
C1769 a_648_712# a_435_712# 0.448f
C1770 a_11512_7066# a_11839_7185# 0.0467f
C1771 a_6866_2809# a_5912_3513# 0.205f
C1772 a_119_2666# a_648_2369# 0.0185f
C1773 a_9134_4112# d0 0.0233f
C1774 a_7988_4356# vdd 0.0325f
C1775 a_13855_1511# a_14112_1321# 0.0467f
C1776 a_11824_4336# a_11403_4336# 0.0104f
C1777 a_16879_6583# a_15941_6827# 0.133f
C1778 a_2103_153# vdd 0.39f
C1779 a_12134_158# a_15209_864# 0.0416f
C1780 a_3141_2109# vdd 0.183f
C1781 a_8881_7988# a_9134_7975# 0.11f
C1782 a_16459_4377# a_16880_4377# 0.0104f
C1783 a_17972_8786# a_18907_9273# 0.254f
C1784 a_5489_5165# a_5174_4913# 0.11f
C1785 a_16813_3785# a_16880_4377# 0.195f
C1786 a_18228_3258# vdd 0.183f
C1787 a_18020_3258# vdd 0.0325f
C1788 a_17969_7860# a_18911_7439# 0.426f
C1789 a_854_5124# a_855_5678# 0.498f
C1790 a_12963_4320# a_12918_4333# 0.181f
C1791 a_14111_2424# vdd 0.183f
C1792 a_119_2666# d0 0.00888f
C1793 a_17908_7146# a_18116_7146# 0.448f
C1794 a_7938_7855# vdd 0.439f
C1795 a_4079_2968# vdd 0.183f
C1796 a_6958_4902# a_4954_133# 0.133f
C1797 a_13903_3527# a_12919_3230# 0.292f
C1798 a_9779_17# a_5053_133# 0.178f
C1799 a_8883_2473# a_8879_2650# 0.539f
C1800 a_12919_2127# vdd 0.0951f
C1801 a_17834_3863# a_17974_4374# 0.206f
C1802 a_10465_2923# vdd 0.178f
C1803 a_12824_1603# vdd 0.0325f
C1804 a_5173_7806# a_5173_8035# 0.539f
C1805 a_3819_8673# a_2886_7637# 0.155f
C1806 a_16673_3274# a_15942_2964# 0.169f
C1807 a_18907_6513# a_18958_5774# 0.011f
C1808 a_8875_8714# a_9132_8524# 0.0467f
C1809 a_7938_6752# a_7802_6064# 0.345f
C1810 a_5175_3623# vdd 0.323f
C1811 a_117_7078# vdd 0.143f
C1812 a_10150_3774# vdd 0.135f
C1813 a_1791_8743# vdd 0.0373f
C1814 a_13852_7026# a_13856_6849# 0.539f
C1815 a_18911_7439# a_18908_8170# 0.0292f
C1816 a_17974_4374# vdd 0.0988f
C1817 a_8927_4666# a_8882_4679# 0.151f
C1818 a_10678_2923# a_10465_2923# 0.448f
C1819 a_5703_2959# vdd 0.0342f
C1820 a_17832_8275# vdd 0.0273f
C1821 a_5490_2959# vdd 0.178f
C1822 a_17972_8786# a_18017_8773# 0.181f
C1823 a_17829_6246# vdd 0.0316f
C1824 a_8195_7665# a_7938_7855# 0.0467f
C1825 a_11402_7645# d1 0.0235f
C1826 a_16568_7107# a_16895_7226# 0.0467f
C1827 a_16881_3274# a_16880_4377# 0.498f
C1828 a_2741_8406# a_2745_8229# 0.524f
C1829 a_8883_3576# a_7944_3266# 0.278f
C1830 a_10466_717# a_10887_717# 0.0104f
C1831 a_13902_5733# a_14110_5733# 0.448f
C1832 a_12772_8411# a_13029_8221# 0.0467f
C1833 a_6750_4902# a_6537_4902# 0.448f
C1834 a_5176_958# a_5178_859# 0.519f
C1835 a_1371_7640# a_853_7330# 0.11f
C1836 a_12913_6716# a_13852_7026# 0.112f
C1837 a_2743_3994# vdd 0.0316f
C1838 a_5702_7925# a_5173_7806# 0.143f
C1839 a_7828_7331# a_8085_7141# 0.0467f
C1840 a_8924_8524# vdd 0.0325f
C1841 a_10887_2374# a_11825_2130# 0.133f
C1842 a_3820_7570# a_2882_7814# 0.316f
C1843 a_116_8868# a_645_8987# 0.143f
C1844 a_7828_7331# a_7802_6064# 0.347f
C1845 a_11834_4866# a_10886_4580# 0.0518f
C1846 a_6427_6578# a_6640_6578# 0.448f
C1847 a_11841_2773# a_10886_2923# 0.0355f
C1848 a_117_8181# a_116_8638# 0.519f
C1849 a_12805_5083# a_12805_2883# 0.176f
C1850 a_15732_7376# a_15204_7124# 0.14f
C1851 a_18914_3581# a_18908_4307# 0.0622f
C1852 a_17973_6580# a_17969_6757# 0.518f
C1853 a_2887_5431# a_3871_5728# 0.292f
C1854 a_7989_2150# a_7940_2340# 0.243f
C1855 a_4078_7934# d0 0.0233f
C1856 a_19165_5220# a_18957_5220# 0.448f
C1857 a_18226_7670# a_17973_7683# 0.11f
C1858 a_19167_2465# a_18914_2478# 0.11f
C1859 a_11933_4866# vdd 0.0369f
C1860 a_3819_8673# a_3870_7934# 0.011f
C1861 d0 a_19165_7980# 0.0233f
C1862 a_5702_4062# a_5489_4062# 0.448f
C1863 a_13853_4820# a_14110_4630# 0.0467f
C1864 a_12918_4333# a_13902_4630# 0.292f
C1865 a_3870_4071# a_4078_4071# 0.448f
C1866 a_10464_4026# a_10149_4231# 0.0467f
C1867 a_17971_3448# a_18913_3027# 0.426f
C1868 a_10886_1820# a_10887_2374# 0.498f
C1869 a_19168_1362# a_18911_1552# 0.0467f
C1870 a_10153_823# a_10466_717# 0.113f
C1871 d2 a_11545_1538# 0.0235f
C1872 a_120_1376# a_120_1147# 0.539f
C1873 a_10883_8438# a_10675_8438# 0.3f
C1874 a_19167_808# vdd 0.183f
C1875 a_8877_7062# vdd 0.311f
C1876 a_15205_5605# vdd 0.128f
C1877 a_3824_9050# a_3869_9037# 0.151f
C1878 a_11618_1027# a_10887_717# 0.169f
C1879 a_18226_6567# a_18018_6567# 0.448f
C1880 a_7800_1829# a_7941_1237# 0.133f
C1881 a_13850_8678# vdd 0.314f
C1882 a_16781_4907# a_15942_4621# 0.0121f
C1883 a_17091_199# a_17865_4947# 0.448f
C1884 a_5489_4062# a_5175_3810# 0.11f
C1885 a_16568_4907# d4 0.0235f
C1886 a_10147_9102# a_10884_8992# 0.277f
C1887 a_19165_5220# a_18908_5410# 0.0467f
C1888 a_7834_4942# a_7877_7141# 0.208f
C1889 a_11926_158# a_12134_158# 0.335f
C1890 a_1803_7061# a_1694_7061# 0.117f
C1891 a_4079_4625# vdd 0.183f
C1892 a_3823_952# a_3872_762# 0.218f
C1893 a_16601_1579# a_16882_1068# 0.11f
C1894 a_19168_1362# vdd 0.183f
C1895 a_11402_6542# d1 0.0235f
C1896 a_10884_6232# a_11402_6542# 0.11f
C1897 a_18957_4117# vdd 0.0325f
C1898 a_11512_7066# a_11839_4985# 0.0104f
C1899 a_5488_9028# d0 0.0235f
C1900 a_10149_4461# a_10149_4690# 0.539f
C1901 a_9133_7421# a_8925_7421# 0.448f
C1902 a_16459_5480# d1 0.0235f
C1903 a_12805_5083# a_12809_2706# 0.685f
C1904 a_13851_9232# vdd 0.311f
C1905 a_119_2250# a_119_2479# 0.539f
C1906 a_12803_7295# a_12917_6539# 0.0437f
C1907 a_7879_2729# a_8087_2729# 0.448f
C1908 a_16982_199# vdd 0.0342f
C1909 a_12963_5423# vdd 0.0325f
C1910 a_12917_7642# a_13852_8129# 0.254f
C1911 a_8926_7975# vdd 0.0325f
C1912 a_12920_1024# a_14112_1321# 0.0192f
C1913 a_1373_2125# a_1586_2125# 0.448f
C1914 a_15732_9033# a_15519_9033# 0.448f
C1915 a_2741_8406# a_3139_7624# 0.0192f
C1916 a_3821_5364# a_2883_5608# 0.316f
C1917 a_10463_8992# d0 0.0235f
C1918 a_4078_5174# a_2883_5608# 0.0192f
C1919 a_15521_5724# d0 0.0235f
C1920 a_3825_5187# d0 0.0138f
C1921 a_2887_4328# a_3140_4315# 0.11f
C1922 a_12919_2127# a_12964_2114# 0.181f
C1923 a_17972_1242# a_18021_1052# 0.219f
C1924 a_7938_6752# a_7987_6562# 0.243f
C1925 a_13903_2424# vdd 0.0325f
C1926 a_3141_3212# d1 0.0233f
C1927 a_3827_775# vdd 0.133f
C1928 a_1803_4861# a_1696_2649# 0.218f
C1929 a_15204_6937# a_15941_6827# 0.277f
C1930 a_15204_7124# vdd 0.143f
C1931 a_10153_823# a_11926_158# 0.0111f
C1932 a_6850_2166# a_6429_2166# 0.0104f
C1933 a_7944_3266# a_8879_3753# 0.254f
C1934 a_4079_5728# a_3822_5918# 0.0467f
C1935 a_7830_5119# a_7879_2729# 0.333f
C1936 a_6864_5021# a_6958_4902# 0.214f
C1937 a_7941_8781# vdd 0.021f
C1938 a_19168_1362# a_18915_1375# 0.11f
C1939 a_14109_7939# vdd 0.183f
C1940 a_12772_8411# a_12962_7629# 0.251f
C1941 a_16458_7686# a_16879_7686# 0.0104f
C1942 a_14985_138# a_16982_199# 0.299f
C1943 a_646_4021# a_433_4021# 0.448f
C1944 a_7060_194# a_5178_859# 0.252f
C1945 a_11542_8156# vdd 0.178f
C1946 a_12915_3407# a_12919_3230# 0.518f
C1947 a_11614_8748# vdd 0.0342f
C1948 a_18228_3258# a_17975_3271# 0.11f
C1949 a_7828_7331# a_7987_6562# 0.0774f
C1950 a_18020_3258# a_17975_3271# 0.181f
C1951 a_434_4575# a_855_4575# 0.0104f
C1952 a_5174_4497# a_5703_4616# 0.143f
C1953 a_8055_6051# vdd 0.183f
C1954 a_12775_1793# a_13173_1011# 0.0192f
C1955 d1 a_13172_2114# 0.0233f
C1956 a_18957_5220# a_17970_5654# 0.283f
C1957 a_8928_803# a_7941_1237# 0.283f
C1958 a_15732_7376# vdd 0.0342f
C1959 a_13901_5179# vdd 0.0325f
C1960 a_17880_1644# a_18088_1644# 0.448f
C1961 a_12775_1793# a_13032_1603# 0.0467f
C1962 a_12774_3999# a_12823_3809# 0.22f
C1963 a_16673_2171# a_16892_2695# 0.0267f
C1964 a_8928_3563# a_8883_3576# 0.151f
C1965 a_855_2918# a_1373_3228# 0.11f
C1966 a_6539_2690# a_6859_4902# 0.0104f
C1967 a_18225_8773# a_17972_8786# 0.11f
C1968 a_18910_2655# a_17971_2345# 0.112f
C1969 a_5489_6822# a_5910_6822# 0.0104f
C1970 a_12913_7819# a_13900_7385# 0.283f
C1971 a_5911_2959# vdd 0.1f
C1972 a_13902_5733# a_13857_5746# 0.151f
C1973 a_18910_998# a_19167_808# 0.0467f
C1974 a_11404_3233# a_10886_2923# 0.11f
C1975 a_3001_1598# d2 0.0233f
C1976 a_11616_4336# a_11403_4336# 0.448f
C1977 a_434_4575# vdd 0.178f
C1978 a_19166_1911# a_17971_2345# 0.0192f
C1979 a_2743_3994# a_2747_3817# 0.524f
C1980 a_8875_8714# a_7942_7678# 0.155f
C1981 a_15942_4621# a_16880_4377# 0.133f
C1982 a_18906_8719# vdd 0.314f
C1983 a_1481_4861# a_1803_4861# 0.11f
C1984 a_17969_6757# a_18018_6567# 0.243f
C1985 a_7799_4035# vdd 0.0316f
C1986 a_8925_9078# a_7941_8781# 0.292f
C1987 a_17970_5654# a_18908_5410# 0.316f
C1988 a_2889_1019# a_3822_2055# 0.155f
C1989 a_4078_7934# a_3825_7947# 0.11f
C1990 a_3826_2981# vdd 0.133f
C1991 a_6429_3269# a_5911_2959# 0.11f
C1992 a_18227_5464# a_17970_5654# 0.0467f
C1993 a_120_1376# a_120_1563# 0.0622f
C1994 d0 a_8882_5782# 0.00533f
C1995 a_854_7884# a_1808_7180# 0.168f
C1996 d0 a_14112_1321# 0.0233f
C1997 a_646_5124# a_118_5329# 0.194f
C1998 a_2889_1019# vdd 0.0799f
C1999 a_3825_6844# a_3870_6831# 0.151f
C2000 a_8880_9091# a_10147_9102# 0.034f
C2001 a_18911_1552# vdd 0.311f
C2002 a_13901_4076# vdd 0.0325f
C2003 a_5489_4062# d0 0.0235f
C2004 a_4077_6277# a_3824_6290# 0.125f
C2005 a_18909_3204# a_18958_3014# 0.218f
C2006 a_12035_158# a_11926_158# 0.117f
C2007 a_117_8181# d0 0.00888f
C2008 a_13857_2986# a_13854_3717# 0.0292f
C2009 a_855_5678# a_434_5678# 0.0104f
C2010 a_10153_823# d0 0.00888f
C2011 a_12809_4906# a_13062_4893# 0.11f
C2012 a_16781_7107# a_15941_6827# 0.0126f
C2013 a_855_4575# vdd 0.454f
C2014 a_2823_4888# vdd 0.0325f
C2015 a_8883_2473# a_8928_2460# 0.151f
C2016 a_7937_8958# a_7801_8270# 0.345f
C2017 a_16880_5480# vdd 0.0273f
C2018 a_5488_6268# a_5173_6473# 0.0467f
C2019 a_6738_194# a_4954_133# 0.0104f
C2020 a_17975_2168# a_18910_2655# 0.254f
C2021 a_19165_4117# a_18908_4307# 0.0467f
C2022 a_1795_1022# a_1794_2125# 0.504f
C2023 a_17834_3863# vdd 0.0273f
C2024 d7 vdd 0.0445f
C2025 a_5173_6703# a_5173_6473# 0.0292f
C2026 a_15520_6827# d0 0.0235f
C2027 a_4077_7380# a_3824_7393# 0.125f
C2028 a_3822_2055# vdd 0.314f
C2029 a_17970_4551# a_18909_4861# 0.112f
C2030 a_10464_6786# a_10148_6896# 0.0467f
C2031 a_18958_1911# a_18909_2101# 0.218f
C2032 a_13858_780# a_13855_1511# 0.0292f
C2033 a_15520_4067# a_15205_4272# 0.0467f
C2034 a_18912_5233# vdd 0.133f
C2035 a_18911_1552# a_18915_1375# 0.539f
C2036 d0 a_13856_6849# 0.00533f
C2037 a_10678_2923# vdd 0.0342f
C2038 a_7834_4942# a_7939_5649# 0.0518f
C2039 a_13854_957# a_12916_1201# 0.316f
C2040 a_8878_4856# a_8927_4666# 0.218f
C2041 a_12773_6205# a_13030_6015# 0.0467f
C2042 a_18018_7670# a_17969_7860# 0.219f
C2043 a_119_3769# a_118_4226# 0.519f
C2044 a_10463_6232# a_10148_6437# 0.0467f
C2045 a_12961_8732# a_12912_8922# 0.243f
C2046 a_6848_6578# a_6781_5986# 0.195f
C2047 a_18956_7426# a_17969_7860# 0.283f
C2048 a_7943_5472# a_8882_5782# 0.278f
C2049 a_6429_3269# vdd 0.178f
C2050 a_8195_7665# vdd 0.183f
C2051 a_3872_762# a_4080_762# 0.448f
C2052 a_118_5329# a_118_5559# 0.0292f
C2053 a_8928_3563# a_8879_3753# 0.218f
C2054 a_10679_2374# a_10150_2671# 0.0185f
C2055 a_14985_138# vdd 0.0212f
C2056 a_17971_3448# a_19166_3014# 0.0192f
C2057 a_15943_758# vdd 0.021f
C2058 a_16460_3274# a_15942_2964# 0.11f
C2059 a_8057_1639# d2 0.0233f
C2060 a_12915_2304# a_14110_1870# 0.0192f
C2061 a_15734_2964# a_15206_2712# 0.14f
C2062 a_8927_1906# vdd 0.0325f
C2063 a_5174_4267# vdd 0.312f
C2064 a_15204_6708# vdd 0.128f
C2065 a_3826_4638# a_3821_5364# 0.0625f
C2066 a_4076_8483# vdd 0.183f
C2067 a_1808_4980# a_1792_6537# 0.122f
C2068 a_18908_4307# a_18912_4130# 0.559f
C2069 a_18915_1375# vdd 0.135f
C2070 a_7939_5649# a_7798_6241# 0.133f
C2071 a_19165_6877# vdd 0.183f
C2072 a_12920_1024# a_12775_1793# 0.326f
C2073 a_2793_1598# vdd 0.0325f
C2074 a_15519_7376# a_15204_7581# 0.0467f
C2075 d0 a_15205_4918# 0.00888f
C2076 a_8925_9078# vdd 0.0325f
C2077 a_15943_2415# a_16892_2695# 0.276f
C2078 a_1696_2649# a_1810_2768# 0.193f
C2079 a_16880_5480# a_16812_5991# 0.146f
C2080 a_11836_2654# a_11834_4866# 0.206f
C2081 a_1805_2649# a_1696_2649# 0.117f
C2082 a_6640_7681# a_5909_7371# 0.169f
C2083 a_17865_4947# a_17863_7159# 0.206f
C2084 a_9133_9078# d0 0.0233f
C2085 a_5175_2291# d0 0.0138f
C2086 a_6569_3780# vdd 0.178f
C2087 a_12854_4893# a_12805_5083# 0.203f
C2088 a_15521_5724# a_15734_5724# 0.448f
C2089 a_1511_8151# d2 0.0235f
C2090 a_13030_6015# d2 0.0233f
C2091 a_12913_7819# a_13170_7629# 0.0467f
C2092 a_13852_5369# a_13857_4643# 0.0625f
C2093 a_10679_2374# a_10150_2255# 0.143f
C2094 a_10148_7999# vdd 0.323f
C2095 a_15736_1312# a_15944_1312# 0.291f
C2096 a_10148_7770# a_10885_7889# 0.426f
C2097 a_16812_5991# vdd 0.0342f
C2098 a_15204_6937# a_15733_6827# 0.194f
C2099 a_8878_4856# a_8881_4125# 0.0292f
C2100 a_17973_6580# a_18018_6567# 0.181f
C2101 a_7990_1047# vdd 0.0325f
C2102 a_12772_8411# a_12917_7642# 0.326f
C2103 a_10465_5683# vdd 0.178f
C2104 a_5701_6268# a_5173_6473# 0.194f
C2105 a_9779_17# vout 0.305f
C2106 a_18228_3258# a_17830_4040# 0.0192f
C2107 a_15205_4731# vdd 0.323f
C2108 a_17830_4040# a_18020_3258# 0.251f
C2109 d2 a_2999_6010# 0.0233f
C2110 a_17975_2168# a_18959_2465# 0.292f
C2111 a_18910_998# vdd 0.314f
C2112 a_2886_7637# a_3825_7947# 0.278f
C2113 a_1513_3739# vdd 0.178f
C2114 a_15735_758# a_15522_758# 0.448f
C2115 a_15940_9033# a_15203_8684# 0.112f
C2116 a_10677_4026# a_10885_4026# 0.3f
C2117 a_8883_2473# d0 0.00533f
C2118 a_10464_6786# a_10885_6786# 0.0104f
C2119 a_18913_5787# vdd 0.135f
C2120 a_13901_6836# a_12917_6539# 0.292f
C2121 d2 a_13031_3809# 0.0233f
C2122 a_856_712# vdd 0.021f
C2123 a_646_7884# a_117_7765# 0.143f
C2124 a_11825_3233# a_11824_4336# 0.498f
C2125 a_12964_2114# vdd 0.0325f
C2126 a_18906_8719# a_18910_8542# 0.559f
C2127 a_18909_5964# a_17970_5654# 0.112f
C2128 a_9136_2460# a_8879_2650# 0.0467f
C2129 a_5174_4913# vdd 0.144f
C2130 a_4079_2968# a_3822_3158# 0.0467f
C2131 a_8925_6318# vdd 0.0325f
C2132 a_5173_7119# a_5173_6932# 0.0625f
C2133 a_10886_2923# a_10150_2671# 0.279f
C2134 a_118_4872# a_118_5329# 0.519f
C2135 a_7879_4929# vdd 0.0325f
C2136 a_11403_5439# a_10886_5683# 0.0467f
C2137 a_6782_3780# a_6849_4372# 0.195f
C2138 a_11614_8748# a_11401_8748# 0.448f
C2139 a_15205_5834# a_15734_5724# 0.194f
C2140 a_11757_3744# vdd 0.0342f
C2141 a_3029_7100# a_2772_7290# 0.0467f
C2142 a_13172_3217# d1 0.0233f
C2143 a_118_5329# a_433_5124# 0.0467f
C2144 a_1803_7061# a_1512_5945# 0.0104f
C2145 a_5910_7925# a_6864_7221# 0.168f
C2146 a_2747_3817# vdd 0.0273f
C2147 a_4080_3522# d0 0.0233f
C2148 a_10149_4877# a_10149_4690# 0.0625f
C2149 a_18906_8719# a_18955_8529# 0.218f
C2150 a_8879_8537# a_8924_8524# 0.154f
C2151 a_15520_5170# a_15205_5375# 0.0467f
C2152 a_5175_2061# a_5490_1856# 0.0467f
C2153 a_16895_5026# a_16890_7107# 0.594f
C2154 a_6850_3269# a_5912_3513# 0.322f
C2155 a_3870_7934# a_3825_7947# 0.151f
C2156 a_16460_2171# a_15942_1861# 0.11f
C2157 a_9136_3563# a_7944_3266# 0.0192f
C2158 a_16458_6583# vdd 0.178f
C2159 a_5491_753# a_5176_958# 0.0467f
C2160 a_6958_4902# a_5911_4616# 0.0863f
C2161 a_17971_3448# a_18910_3758# 0.112f
C2162 a_10679_717# a_10151_922# 0.194f
C2163 a_7989_3253# a_7799_4035# 0.251f
C2164 a_10150_2484# vdd 0.323f
C2165 a_7945_1060# a_7941_1237# 0.518f
C2166 a_12915_2304# a_12805_2883# 0.249f
C2167 a_5704_2410# a_5175_2291# 0.143f
C2168 a_12809_2706# a_12915_3407# 0.392f
C2169 a_2778_2701# a_3031_2688# 0.11f
C2170 a_17878_6056# a_17859_7336# 0.255f
C2171 a_15203_8684# a_15731_8479# 0.194f
C2172 a_3822_5918# a_3871_5728# 0.218f
C2173 a_5487_8474# d0 0.0235f
C2174 a_6639_8784# a_5909_9028# 0.195f
C2175 vdd a_17975_3271# 0.0799f
C2176 a_19166_4671# a_17974_4374# 0.0192f
C2177 a_3821_4261# a_3825_4084# 0.559f
C2178 d0 a_9135_3009# 0.0233f
C2179 a_15522_2415# a_15735_2415# 0.448f
C2180 a_5911_5719# a_5174_5829# 0.277f
C2181 a_10150_2484# a_10678_2923# 0.011f
C2182 a_8883_3576# a_8877_4302# 0.0622f
C2183 a_2889_1019# a_3873_1316# 0.292f
C2184 a_6866_2809# a_6782_3780# 0.263f
C2185 a_3825_6844# d0 0.00533f
C2186 a_8927_3009# vdd 0.0325f
C2187 a_1805_2649# a_1727_1533# 0.198f
C2188 a_2934_1006# a_2889_1019# 0.181f
C2189 a_5492_1307# vdd 0.178f
C2190 a_12805_5083# a_11834_4866# 0.409f
C2191 a_18910_8542# vdd 0.133f
C2192 a_15521_4621# d0 0.0235f
C2193 a_16881_3274# a_15943_3518# 0.322f
C2194 a_6428_4372# vdd 0.178f
C2195 a_3825_6844# a_3820_7570# 0.0625f
C2196 a_13060_7105# d3 0.0233f
C2197 a_6427_7681# a_5910_7925# 0.0467f
C2198 a_1514_1533# vdd 0.178f
C2199 a_2999_6010# a_2772_7290# 0.0192f
C2200 a_17877_8262# a_17832_8275# 0.157f
C2201 a_16783_2695# vdd 0.0342f
C2202 a_3825_5187# a_3821_5364# 0.559f
C2203 a_645_8987# a_432_8987# 0.448f
C2204 a_11933_4866# a_10886_4580# 0.0863f
C2205 a_3825_5187# a_4078_5174# 0.125f
C2206 a_5909_6268# a_5173_6473# 0.255f
C2207 a_6859_7102# a_5910_6822# 0.28f
C2208 a_855_4575# a_1694_4861# 0.0121f
C2209 a_18955_8529# vdd 0.0325f
C2210 a_16814_1579# vdd 0.0342f
C2211 a_18960_1362# a_17976_1065# 0.292f
C2212 a_3873_1316# a_3822_2055# 0.011f
C2213 a_16671_6583# a_16890_7107# 0.0267f
C2214 d0 a_13858_2437# 0.00533f
C2215 a_13851_7575# a_13856_6849# 0.0625f
C2216 a_13902_2973# vdd 0.0325f
C2217 a_10464_4026# d0 0.0235f
C2218 a_7989_3253# vdd 0.0325f
C2219 a_13901_7939# a_13852_8129# 0.218f
C2220 a_5490_4616# a_5911_4616# 0.0104f
C2221 a_3873_1316# vdd 0.0325f
C2222 a_10887_3477# a_11617_3233# 0.219f
C2223 a_15939_8479# a_15203_8684# 0.255f
C2224 d4 vdd 0.356f
C2225 a_8085_7141# d3 0.0233f
C2226 a_6849_5475# a_6428_5475# 0.0104f
C2227 a_13900_7385# vdd 0.0325f
C2228 a_11617_2130# a_10887_2374# 0.195f
C2229 a_3828_1329# d0 0.00533f
C2230 a_16673_3274# vdd 0.0342f
C2231 a_2934_1006# vdd 0.0325f
C2232 a_6642_2166# a_5911_1856# 0.169f
C2233 a_1694_4861# vdd 0.0342f
C2234 a_12778_3822# a_12774_3999# 0.524f
C2235 a_9137_1357# d0 0.0233f
C2236 a_11401_8748# vdd 0.178f
C2237 a_1371_6537# d1 0.0235f
C2238 a_7800_1829# vdd 0.0316f
C2239 a_18226_7670# d1 0.0233f
C2240 a_17910_2734# vdd 0.0325f
C2241 a_11617_3233# a_11825_3233# 0.241f
C2242 a_10150_2255# a_10466_2374# 0.125f
C2243 a_13858_780# d0 0.0138f
C2244 a_6848_6578# a_6849_5475# 0.504f
C2245 a_1373_3228# vdd 0.178f
C2246 a_5911_5719# a_5910_5165# 0.498f
C2247 a_10884_7335# a_11402_7645# 0.11f
C2248 a_18957_7980# a_18912_7993# 0.151f
C2249 a_16781_4907# a_16895_5026# 0.178f
C2250 a_2741_8406# a_2882_7814# 0.133f
C2251 a_6537_7102# vdd 0.178f
C2252 a_18229_1052# a_17972_1242# 0.0467f
C2253 a_10888_1271# a_10151_1152# 0.426f
C2254 a_5176_1604# a_5175_2061# 0.519f
C2255 a_1587_1022# a_857_1266# 0.219f
C2256 a_15521_2964# a_15206_2712# 0.11f
C2257 a_8881_6885# a_7942_6575# 0.278f
C2258 a_1585_5434# vdd 0.0342f
C2259 a_18906_8719# a_17973_7683# 0.155f
C2260 a_15941_7930# a_15204_7811# 0.426f
C2261 a_856_2369# a_1696_2649# 0.0126f
C2262 a_17828_8452# a_17863_7159# 0.298f
C2263 d0 a_13858_3540# 0.00533f
C2264 a_12916_8745# a_14108_9042# 0.0192f
C2265 a_5488_6268# a_5174_6016# 0.11f
C2266 a_5172_8679# a_5173_8222# 0.519f
C2267 a_12914_5613# a_12854_4893# 0.0121f
C2268 a_7938_6752# a_9133_6318# 0.0192f
C2269 a_118_5975# d0 0.00888f
C2270 a_14109_5179# a_13856_5192# 0.125f
C2271 a_13857_1883# a_13902_1870# 0.154f
C2272 a_15940_6273# a_15519_6273# 0.0104f
C2273 a_5705_1307# vdd 0.0342f
C2274 a_18086_6056# a_17859_7336# 0.0192f
C2275 a_15518_8479# a_15731_8479# 0.448f
C2276 a_2931_6521# vdd 0.0325f
C2277 a_117_6891# a_645_7330# 0.011f
C2278 a_15734_1861# a_15207_1609# 0.14f
C2279 a_2886_6534# a_3139_6521# 0.11f
C2280 a_12807_7118# a_12809_4906# 0.206f
C2281 a_6866_2809# a_6539_2690# 0.0467f
C2282 a_3823_2609# a_3872_2419# 0.218f
C2283 a_5053_133# a_4845_133# 0.33f
C2284 a_12913_6716# a_13900_6282# 0.283f
C2285 a_117_8181# a_852_8433# 0.279f
C2286 a_8928_3563# a_9136_3563# 0.448f
C2287 a_10886_1820# a_10678_1820# 0.3f
C2288 a_10150_3128# a_10465_2923# 0.0467f
C2289 a_10149_5793# a_10149_5980# 0.0622f
C2290 a_6430_1063# vdd 0.178f
C2291 a_14110_5733# vdd 0.183f
C2292 a_15205_5834# a_15205_6021# 0.0622f
C2293 a_3826_5741# vdd 0.135f
C2294 a_5909_9028# a_5908_8474# 0.498f
C2295 a_15203_8914# a_15519_9033# 0.125f
C2296 a_11758_1538# vdd 0.0342f
C2297 a_11512_7066# a_11834_7066# 0.11f
C2298 a_8928_803# vdd 0.0325f
C2299 a_5172_8679# a_5172_8909# 0.0292f
C2300 a_6570_1574# vdd 0.178f
C2301 a_10677_5129# a_10149_4877# 0.14f
C2302 a_12915_2304# a_13172_2114# 0.0467f
C2303 a_2790_8216# vdd 0.0325f
C2304 a_7800_1829# a_7990_1047# 0.251f
C2305 a_15941_4067# vdd 0.0799f
C2306 a_17973_7683# vdd 0.0799f
C2307 a_2930_8727# vdd 0.0325f
C2308 a_8877_5405# a_8926_5215# 0.218f
C2309 a_10148_8186# a_10675_8438# 0.14f
C2310 a_5911_1856# a_5176_1417# 0.155f
C2311 a_5911_5719# a_5490_5719# 0.0104f
C2312 a_12805_5083# a_12854_2693# 0.333f
C2313 a_13903_3527# a_14111_3527# 0.448f
C2314 a_16600_3785# vdd 0.178f
C2315 a_3823_952# a_2885_1196# 0.316f
C2316 a_7797_8447# a_7832_7154# 0.298f
C2317 a_3822_3158# a_3826_2981# 0.559f
C2318 a_15939_8479# a_15518_8479# 0.0104f
C2319 a_15204_8040# vdd 0.323f
C2320 a_15520_5170# a_15205_4918# 0.11f
C2321 a_11616_5439# a_10886_5683# 0.219f
C2322 a_15205_4272# a_15942_4621# 0.112f
C2323 a_5912_2410# a_5911_1856# 0.498f
C2324 a_18914_821# d0 0.0138f
C2325 a_855_5678# vdd 0.455f
C2326 a_3821_4261# a_3827_3535# 0.0622f
C2327 a_10149_5793# a_10886_5683# 0.277f
C2328 a_17834_3863# a_17830_4040# 0.524f
C2329 a_1511_8151# a_1808_7180# 0.0104f
C2330 a_2821_7100# a_2772_7290# 0.218f
C2331 a_10151_1381# a_10888_1271# 0.277f
C2332 a_2881_8917# a_2885_8740# 0.518f
C2333 a_17830_4040# vdd 0.0316f
C2334 a_9136_2460# a_8928_2460# 0.448f
C2335 a_8879_8537# vdd 0.133f
C2336 a_1803_7061# a_1725_5945# 0.198f
C2337 a_15204_7811# d0 0.0138f
C2338 a_2744_1788# a_2885_1196# 0.133f
C2339 vdd a_13170_7629# 0.183f
C2340 a_117_6891# a_853_7330# 0.155f
C2341 a_854_7884# a_1792_7640# 0.322f
C2342 a_5704_753# a_5912_753# 0.3f
C2343 a_16881_2171# a_16673_2171# 0.26f
C2344 a_15520_6827# a_15204_6937# 0.0467f
C2345 a_5701_6268# a_5174_6016# 0.14f
C2346 a_15522_3518# vdd 0.178f
C2347 a_3822_3158# vdd 0.314f
C2348 a_856_2369# a_119_2479# 0.277f
C2349 a_18959_808# a_18914_821# 0.154f
C2350 a_10886_4580# vdd 0.454f
C2351 a_436_1266# a_120_1147# 0.125f
C2352 a_17908_7146# vdd 0.0325f
C2353 a_4077_9037# vdd 0.183f
C2354 a_15943_2415# a_15206_2066# 0.112f
C2355 a_8196_5459# d1 0.0233f
C2356 a_12822_6015# a_13030_6015# 0.448f
C2357 a_13060_7105# a_12803_7295# 0.0467f
C2358 a_18955_8529# a_18910_8542# 0.154f
C2359 a_3139_6521# a_2882_6711# 0.0467f
C2360 a_1586_3228# a_856_3472# 0.219f
C2361 a_16598_8197# d2 0.0235f
C2362 a_13850_8678# a_13899_8488# 0.218f
C2363 a_10464_6786# vdd 0.178f
C2364 a_8881_5228# vdd 0.133f
C2365 a_12964_3217# a_12919_3230# 0.181f
C2366 a_8882_1919# a_9135_1906# 0.125f
C2367 a_19166_4671# vdd 0.183f
C2368 a_3827_2432# vdd 0.145f
C2369 a_5176_1188# a_5176_1417# 0.539f
C2370 a_10149_5793# a_10149_5564# 0.539f
C2371 a_6643_1063# vdd 0.0342f
C2372 a_13855_9055# a_13900_9042# 0.151f
C2373 a_2741_8406# a_2886_7637# 0.326f
C2374 a_2746_6023# a_2772_7290# 0.347f
C2375 a_18907_9273# a_19164_9083# 0.0467f
C2376 a_11823_6542# a_11839_4985# 0.122f
C2377 a_8882_4679# vdd 0.146f
C2378 a_12916_1201# vdd 0.439f
C2379 a_10465_4580# d0 0.0235f
C2380 a_15520_4067# a_15733_4067# 0.448f
C2381 a_12778_3822# a_13171_4320# 0.0192f
C2382 a_17877_8262# vdd 0.0325f
C2383 a_5911_5719# a_5703_5719# 0.291f
C2384 a_12962_7629# a_12913_7819# 0.219f
C2385 a_12918_4333# vdd 0.0988f
C2386 a_1795_1022# a_857_1266# 0.322f
C2387 a_4077_7380# d0 0.0233f
C2388 a_16568_4907# a_16781_4907# 0.448f
C2389 a_3140_5418# vdd 0.183f
C2390 a_2774_2878# vdd 0.0323f
C2391 a_10148_7540# a_10885_7889# 0.112f
C2392 a_2883_4505# a_3140_4315# 0.0467f
C2393 a_17973_6580# a_18907_7616# 0.155f
C2394 a_1808_4980# a_1808_7180# 0.176f
C2395 a_10149_5334# a_10886_5683# 0.112f
C2396 a_10884_6232# a_10885_6786# 0.498f
C2397 a_11544_3744# a_11824_4336# 0.0467f
C2398 a_2778_2701# a_2884_3402# 0.392f
C2399 a_3824_1506# a_2885_1196# 0.112f
C2400 a_119_2020# a_647_1815# 0.194f
C2401 a_11823_7645# a_10885_7889# 0.322f
C2402 a_13857_5746# vdd 0.135f
C2403 a_2823_2688# vdd 0.0325f
C2404 a_4077_7380# a_3820_7570# 0.0467f
C2405 a_7940_3443# a_9135_3009# 0.0192f
C2406 a_15520_4067# d0 0.0235f
C2407 a_10464_4026# a_10885_4026# 0.0104f
C2408 a_5176_958# vdd 0.312f
C2409 d0 a_10464_7889# 0.0235f
C2410 a_5705_1307# a_5492_1307# 0.448f
C2411 a_16457_8789# vdd 0.178f
C2412 a_8881_6885# a_8876_7611# 0.0625f
C2413 a_3141_2109# d1 0.0233f
C2414 a_2881_8917# a_3819_8673# 0.316f
C2415 a_15944_1312# a_15207_963# 0.112f
C2416 a_2103_153# a_4632_133# 0.0467f
C2417 a_3140_4315# a_2932_4315# 0.448f
C2418 a_14110_2973# vdd 0.183f
C2419 a_18228_3258# d1 0.0233f
C2420 a_13172_3217# a_12915_3407# 0.0467f
C2421 a_3821_7021# a_4078_6831# 0.0467f
C2422 a_10884_7335# a_10463_7335# 0.0104f
C2423 a_4078_4071# vdd 0.183f
C2424 a_9136_2460# d0 0.0233f
C2425 a_8877_8165# a_9134_7975# 0.0467f
C2426 a_2778_4901# a_2772_7290# 0.681f
C2427 a_7939_5649# a_8926_5215# 0.283f
C2428 a_5909_6268# a_5174_6016# 0.279f
C2429 a_7834_4942# a_7832_7154# 0.206f
C2430 a_10883_8438# a_10462_8438# 0.0104f
C2431 a_2793_1598# a_2774_2878# 0.255f
C2432 a_11713_158# a_11926_158# 0.448f
C2433 a_8878_2096# a_7940_2340# 0.316f
C2434 a_17861_2924# vdd 0.0323f
C2435 a_649_1266# a_120_1147# 0.143f
C2436 a_117_6432# a_117_6662# 0.0292f
C2437 a_16460_3274# vdd 0.178f
C2438 a_15940_7376# a_15204_7124# 0.279f
C2439 a_3827_3535# a_3823_3712# 0.539f
C2440 a_4080_762# a_2885_1196# 0.0192f
C2441 a_16881_2171# a_15943_2415# 0.133f
C2442 a_9136_803# d0 0.0233f
C2443 a_13859_1334# a_14112_1321# 0.11f
C2444 a_7834_2742# a_7830_2919# 0.484f
C2445 a_13856_4089# d0 0.0138f
C2446 a_15736_1312# a_15207_1609# 0.0185f
C2447 a_18960_1362# a_19168_1362# 0.448f
C2448 a_10149_5334# a_10149_5564# 0.0292f
C2449 a_5173_6932# a_5701_7371# 0.011f
C2450 a_17975_2168# a_18914_2478# 0.278f
C2451 a_10463_8992# a_10147_8873# 0.125f
C2452 a_5700_8474# vdd 0.0342f
C2453 a_16570_2695# vdd 0.178f
C2454 a_12917_6539# vdd 0.0951f
C2455 a_1481_7061# a_1808_7180# 0.0467f
C2456 a_17830_4040# a_17975_3271# 0.326f
C2457 a_10885_7889# a_10677_7889# 0.291f
C2458 a_10148_7083# a_10676_7335# 0.14f
C2459 a_14109_6836# a_13856_6849# 0.11f
C2460 a_10151_922# vdd 0.312f
C2461 a_13853_2060# vdd 0.314f
C2462 a_12913_7819# a_14108_7385# 0.0192f
C2463 a_8880_7434# a_9133_7421# 0.125f
C2464 a_10151_1381# a_10886_1820# 0.155f
C2465 a_15732_7376# a_15940_7376# 0.3f
C2466 a_10150_3128# vdd 0.312f
C2467 a_118_5559# a_647_5678# 0.143f
C2468 a_13853_3163# a_13858_2437# 0.0625f
C2469 a_11615_6542# a_11823_6542# 0.26f
C2470 a_5174_4497# a_5911_4616# 0.426f
C2471 a_15521_1861# a_15206_2066# 0.0467f
C2472 a_434_4575# a_118_4456# 0.125f
C2473 a_3869_6277# vdd 0.0325f
C2474 a_10150_3128# a_10678_2923# 0.194f
C2475 a_17879_3850# a_18087_3850# 0.448f
C2476 a_15940_6273# a_15941_6827# 0.498f
C2477 a_854_5124# a_646_5124# 0.3f
C2478 a_7945_1060# vdd 0.0799f
C2479 a_3869_9037# vdd 0.0325f
C2480 a_855_4575# a_118_4226# 0.112f
C2481 a_434_2918# a_855_2918# 0.0104f
C2482 a_13857_1883# a_13854_2614# 0.0292f
C2483 a_5909_7371# a_5910_7925# 0.498f
C2484 a_14109_5179# a_13901_5179# 0.448f
C2485 a_7938_6752# a_8880_6331# 0.426f
C2486 a_13899_8488# vdd 0.0325f
C2487 a_6859_7102# a_6864_7221# 0.464f
C2488 a_2791_6010# a_2999_6010# 0.448f
C2489 a_5491_2410# vdd 0.178f
C2490 a_13850_8678# a_14107_8488# 0.0467f
C2491 a_16460_2171# vdd 0.178f
C2492 a_11405_1027# vdd 0.178f
C2493 a_12805_2883# a_13032_1603# 0.0192f
C2494 a_11512_7066# d3 0.0235f
C2495 a_10148_8186# d0 0.00888f
C2496 a_13904_1321# a_14112_1321# 0.448f
C2497 a_10679_2374# a_10466_2374# 0.448f
C2498 a_7060_194# vdd 0.0211f
C2499 a_15206_2712# a_15942_2964# 0.279f
C2500 a_4080_3522# a_3827_3535# 0.11f
C2501 a_118_4226# vdd 0.312f
C2502 a_16601_1579# d2 0.0235f
C2503 a_4080_2419# vdd 0.183f
C2504 a_2103_153# a_4954_133# 0.498f
C2505 a_6851_1063# vdd 0.0273f
C2506 a_118_4456# a_855_4575# 0.426f
C2507 a_12805_5083# a_11933_4866# 0.0189f
C2508 a_1585_5434# a_855_5678# 0.219f
C2509 a_10151_1568# a_10465_1820# 0.11f
C2510 a_8878_3199# a_8883_2473# 0.0625f
C2511 a_5703_1856# a_5911_1856# 0.3f
C2512 a_12852_7105# a_12803_7295# 0.218f
C2513 a_12918_5436# a_13902_5733# 0.292f
C2514 a_5488_6268# vdd 0.178f
C2515 a_15206_2296# a_15522_2415# 0.125f
C2516 a_3000_3804# a_2743_3994# 0.0467f
C2517 a_16897_2814# a_16892_2695# 0.586f
C2518 a_7938_7855# a_9133_7421# 0.0192f
C2519 a_9134_7975# d0 0.0233f
C2520 a_5173_6703# vdd 0.128f
C2521 a_6850_3269# a_6782_3780# 0.146f
C2522 a_19165_7980# a_18912_7993# 0.11f
C2523 a_118_4456# vdd 0.128f
C2524 a_2742_6200# vdd 0.0316f
C2525 a_15735_2415# vdd 0.0342f
C2526 a_2933_2109# a_2888_2122# 0.181f
C2527 a_12914_5613# a_13856_5192# 0.426f
C2528 a_13029_8221# vdd 0.183f
C2529 a_2933_2109# a_2884_2299# 0.243f
C2530 a_4081_1316# d0 0.0233f
C2531 a_10885_7889# a_11615_7645# 0.219f
C2532 a_15940_7376# vdd 0.1f
C2533 a_1586_3228# a_1794_3228# 0.241f
C2534 a_12917_7642# a_12913_7819# 0.518f
C2535 a_649_1266# a_120_1563# 0.0185f
C2536 a_7988_4356# a_7803_3858# 0.231f
C2537 a_18960_1362# a_18911_1552# 0.218f
C2538 a_15940_9033# a_15203_9143# 0.277f
C2539 a_12915_3407# a_12854_2693# 0.0126f
C2540 a_16598_8197# a_16879_7686# 0.11f
C2541 a_2881_8917# a_3823_8496# 0.426f
C2542 vdd a_5703_4616# 0.0342f
C2543 a_7847_6051# a_8055_6051# 0.448f
C2544 a_13853_5923# a_13902_5733# 0.218f
C2545 a_16880_5480# a_16599_5991# 0.11f
C2546 a_646_7884# a_854_7884# 0.291f
C2547 a_7990_1047# a_7945_1060# 0.181f
C2548 a_6427_7681# a_5909_7371# 0.11f
C2549 d0 a_9135_1906# 0.0233f
C2550 a_14109_5179# vdd 0.183f
C2551 a_17972_1242# a_18914_821# 0.426f
C2552 a_7939_4546# a_8926_4112# 0.283f
C2553 a_11836_2654# vdd 0.0269f
C2554 a_3820_6467# a_2882_6711# 0.316f
C2555 a_18959_3568# vdd 0.0325f
C2556 a_13031_3809# a_12823_3809# 0.448f
C2557 a_5704_3513# a_5491_3513# 0.448f
C2558 a_16599_5991# vdd 0.178f
C2559 a_5910_5165# a_5174_5370# 0.255f
C2560 a_16989_4907# a_17091_199# 7.78f
C2561 a_18960_1362# vdd 0.0325f
C2562 a_12809_2706# a_12964_3217# 0.0267f
C2563 a_855_1815# a_647_1815# 0.3f
C2564 a_5174_4726# a_5490_4616# 0.0467f
C2565 a_9888_17# vdd 0.022f
C2566 a_12809_4906# a_12035_158# 0.448f
C2567 a_15734_1861# a_15942_1861# 0.3f
C2568 d0 a_14110_1870# 0.0233f
C2569 d0 a_10151_1152# 0.0138f
C2570 a_9134_6872# d0 0.0233f
C2571 d0 a_432_7330# 0.0235f
C2572 a_8878_3199# a_9135_3009# 0.0467f
C2573 a_1803_7061# a_1792_6537# 0.328f
C2574 a_8878_4856# vdd 0.311f
C2575 a_116_8868# vdd 0.128f
C2576 a_8878_5959# vdd 0.311f
C2577 a_7846_8257# vdd 0.0325f
C2578 a_3823_952# a_4080_762# 0.0467f
C2579 a_8881_7988# a_8924_8524# 0.0185f
C2580 a_15521_4621# a_15205_4502# 0.125f
C2581 a_5172_9138# a_5701_9028# 0.194f
C2582 a_18913_3027# a_18958_3014# 0.154f
C2583 a_3827_3535# a_3872_3522# 0.151f
C2584 a_7944_3266# a_7940_3443# 0.518f
C2585 a_119_3769# a_854_4021# 0.279f
C2586 a_15734_2964# a_15206_3169# 0.194f
C2587 a_13902_2973# a_14110_2973# 0.448f
C2588 a_119_2250# vdd 0.128f
C2589 a_18907_6513# a_17974_5477# 0.155f
C2590 a_19164_6323# vdd 0.183f
C2591 a_9888_17# a_14985_138# 0.307f
C2592 a_1810_2768# a_855_2918# 0.0355f
C2593 a_15732_9033# vdd 0.0342f
C2594 a_18960_1362# a_18915_1375# 0.151f
C2595 a_7879_4929# a_7060_194# 0.282f
C2596 a_5175_2520# a_5175_2291# 0.539f
C2597 a_16880_5480# a_16890_7107# 0.206f
C2598 a_5701_6268# vdd 0.0342f
C2599 a_7797_8447# a_7942_7678# 0.326f
C2600 a_6537_4902# a_6859_4902# 0.11f
C2601 a_854_4021# a_1585_4331# 0.169f
C2602 a_6430_1063# a_6643_1063# 0.448f
C2603 a_1724_8151# a_1808_7180# 0.263f
C2604 a_10886_1820# a_10150_2025# 0.255f
C2605 a_7834_4942# a_7798_6241# 0.181f
C2606 a_7940_3443# a_8197_3253# 0.0467f
C2607 a_854_7884# a_117_7765# 0.426f
C2608 a_10885_7889# a_11839_7185# 0.168f
C2609 a_11514_2654# d3 0.0235f
C2610 a_435_2369# a_119_2479# 0.0467f
C2611 a_5912_753# a_5178_859# 1.07f
C2612 a_12805_2883# a_13062_2693# 0.0467f
C2613 a_5490_4616# d0 0.0235f
C2614 a_7847_6051# vdd 0.0325f
C2615 a_16783_2695# a_16570_2695# 0.448f
C2616 a_14107_8488# vdd 0.183f
C2617 a_16890_7107# vdd 0.0269f
C2618 a_2885_8740# a_3824_9050# 0.278f
C2619 a_16673_3274# a_16460_3274# 0.448f
C2620 a_17861_2924# a_17910_2734# 0.203f
C2621 a_1694_7061# vdd 0.0342f
C2622 a_16458_7686# a_16671_7686# 0.448f
C2623 a_854_5124# a_118_4872# 0.279f
C2624 a_12962_7629# vdd 0.0325f
C2625 a_10149_4461# a_10465_4580# 0.125f
C2626 a_5175_3394# a_5912_3513# 0.426f
C2627 a_18909_3204# vdd 0.314f
C2628 a_16812_5991# a_16599_5991# 0.448f
C2629 a_5173_7119# a_5173_7576# 0.519f
C2630 a_5702_6822# a_5910_6822# 0.291f
C2631 a_3823_952# a_122_818# 0.884f
C2632 a_854_5124# a_433_5124# 0.0104f
C2633 a_3138_8727# a_2745_8229# 0.0192f
C2634 a_18911_7439# a_19164_7426# 0.125f
C2635 a_17861_5124# a_17091_199# 0.177f
C2636 d1 vdd 2.85f
C2637 a_10884_6232# vdd 0.0799f
C2638 a_4632_133# vdd 0.178f
C2639 a_15207_1193# vdd 0.128f
C2640 a_11727_2654# a_10887_2374# 0.0126f
C2641 a_3826_4638# a_3822_4815# 0.539f
C2642 a_14110_5733# a_13857_5746# 0.11f
C2643 a_2887_4328# a_3821_5364# 0.155f
C2644 a_1511_8151# a_1792_7640# 0.11f
C2645 a_3821_8124# a_2882_7814# 0.112f
C2646 a_8881_7988# a_8926_7975# 0.151f
C2647 a_13850_8678# a_12917_7642# 0.155f
C2648 a_5172_9138# a_3824_9050# 0.036f
C2649 a_10887_2374# a_10150_2255# 0.426f
C2650 a_5174_4913# a_5703_4616# 0.0185f
C2651 a_16878_8789# vdd 0.0373f
C2652 a_2886_6534# a_2882_6711# 0.518f
C2653 a_13852_7026# a_13855_6295# 0.0292f
C2654 a_18957_5220# a_18908_5410# 0.218f
C2655 a_6429_3269# d1 0.0235f
C2656 a_11404_2130# a_10887_2374# 0.0467f
C2657 a_7879_2729# vdd 0.0325f
C2658 a_8195_7665# d1 0.0233f
C2659 a_15206_3399# vdd 0.128f
C2660 a_6428_5475# vdd 0.178f
C2661 a_7944_2163# a_8879_2650# 0.254f
C2662 a_10885_4026# a_11824_4336# 0.302f
C2663 a_12805_5083# vdd 0.0323f
C2664 a_5175_3394# d0 0.0138f
C2665 a_14109_4076# a_13901_4076# 0.448f
C2666 a_8054_8257# a_7832_7154# 0.0192f
C2667 a_9566_17# a_5053_133# 0.0467f
C2668 a_12809_2706# a_13062_2693# 0.11f
C2669 a_4078_7934# a_3821_8124# 0.0467f
C2670 a_6848_6578# vdd 0.0373f
C2671 a_13853_5923# a_13856_5192# 0.0292f
C2672 a_2791_6010# a_2746_6023# 0.157f
C2673 a_3871_4625# a_3821_5364# 0.011f
C2674 a_10150_3358# vdd 0.128f
C2675 a_15519_7376# d0 0.0235f
C2676 a_3822_3158# a_3827_2432# 0.0625f
C2677 a_7800_1829# a_7945_1060# 0.326f
C2678 a_119_3582# a_646_4021# 0.011f
C2679 a_12809_4906# a_11839_4985# 0.233f
C2680 a_10147_9102# vdd 0.323f
C2681 a_18909_2101# a_17971_2345# 0.316f
C2682 a_434_1815# vdd 0.178f
C2683 a_5173_7119# d0 0.00888f
C2684 a_117_7994# vdd 0.323f
C2685 a_5172_8679# a_5487_8474# 0.0467f
C2686 a_16769_199# d5 0.0235f
C2687 a_10884_7335# a_10148_6896# 0.155f
C2688 a_10676_7335# a_10148_7540# 0.194f
C2689 a_433_6781# vdd 0.178f
C2690 a_12916_8745# a_12776_8234# 0.206f
C2691 a_1682_153# a_1895_153# 0.448f
C2692 a_10148_6667# d0 0.0138f
C2693 a_16812_5991# a_16890_7107# 0.198f
C2694 a_13169_8732# vdd 0.183f
C2695 a_17861_5124# a_17865_4947# 0.518f
C2696 a_10149_4877# a_10149_5334# 0.519f
C2697 a_12965_1011# vdd 0.0325f
C2698 d0 a_9134_5215# 0.0233f
C2699 a_18958_1911# a_17971_2345# 0.283f
C2700 a_14109_4076# vdd 0.183f
C2701 a_17880_1644# a_17835_1657# 0.157f
C2702 a_3000_3804# vdd 0.183f
C2703 a_855_4575# a_1803_4861# 0.0518f
C2704 a_6849_4372# a_6859_4902# 0.0928f
C2705 a_4078_6831# a_3870_6831# 0.448f
C2706 a_1584_7640# a_1792_7640# 0.241f
C2707 a_7828_7331# a_7877_7141# 0.218f
C2708 a_5701_9028# a_5909_9028# 0.291f
C2709 a_5910_7925# a_5173_8035# 0.277f
C2710 a_3821_4261# a_2888_3225# 0.155f
C2711 a_12917_7642# a_14109_7939# 0.0192f
C2712 a_8054_8257# a_7797_8447# 0.0467f
C2713 a_16781_4907# vdd 0.0342f
C2714 a_5909_6268# vdd 0.0799f
C2715 a_18959_3568# a_17975_3271# 0.292f
C2716 a_8195_6562# vdd 0.183f
C2717 a_6750_4902# a_6958_4902# 0.337f
C2718 a_4079_5728# vdd 0.183f
C2719 a_6641_5475# a_5911_5719# 0.219f
C2720 a_7943_4369# a_8927_4666# 0.292f
C2721 a_119_3582# a_856_3472# 0.277f
C2722 a_7801_8270# a_7941_8781# 0.206f
C2723 a_14108_7385# vdd 0.183f
C2724 a_7989_2150# a_8197_2150# 0.448f
C2725 a_1726_3739# a_1793_4331# 0.195f
C2726 a_4077_6277# d0 0.0233f
C2727 a_17970_4551# a_18227_4361# 0.0467f
C2728 a_1682_153# a_2103_153# 0.0104f
C2729 a_7940_2340# a_7830_2919# 0.249f
C2730 a_17878_6056# a_17829_6246# 0.22f
C2731 a_9134_4112# a_7939_4546# 0.0192f
C2732 a_1803_4861# vdd 0.0264f
C2733 a_17091_199# a_16769_199# 0.11f
C2734 a_6567_8192# a_6780_8192# 0.448f
C2735 d3 a_13062_2693# 0.0233f
C2736 a_10148_7083# a_10677_6786# 0.0185f
C2737 a_117_8181# a_646_7884# 0.0185f
C2738 a_7803_3858# a_7799_4035# 0.524f
C2739 a_5702_7925# a_5910_7925# 0.291f
C2740 a_3826_5741# a_3869_6277# 0.0185f
C2741 a_12914_5613# a_12963_5423# 0.219f
C2742 a_4954_133# vdd 0.021f
C2743 a_9133_7421# vdd 0.183f
C2744 a_6866_2809# a_6859_4902# 0.583f
C2745 a_5174_5600# a_5174_5829# 0.539f
C2746 a_434_5678# a_118_5559# 0.125f
C2747 a_13852_8129# a_13855_7398# 0.0292f
C2748 a_15943_3518# a_15942_2964# 0.498f
C2749 a_15206_3815# vdd 0.135f
C2750 a_16672_4377# a_16459_4377# 0.448f
C2751 a_434_2918# vdd 0.178f
C2752 a_11841_2773# a_11824_4336# 0.14f
C2753 a_1371_7640# vdd 0.178f
C2754 a_11823_6542# a_11834_7066# 0.328f
C2755 a_6849_5475# a_5910_5165# 0.206f
C2756 a_3139_7624# a_2882_7814# 0.0467f
C2757 a_436_1266# d0 0.0235f
C2758 a_15206_2525# a_15734_2964# 0.011f
C2759 a_18907_9273# a_17968_8963# 0.112f
C2760 a_2776_7113# vdd 0.0269f
C2761 a_3870_5174# vdd 0.0325f
C2762 a_2931_7624# vdd 0.0325f
C2763 a_10148_7540# a_10148_7770# 0.0292f
C2764 a_8881_7988# vdd 0.135f
C2765 a_6851_1063# a_6430_1063# 0.0104f
C2766 a_6567_8192# a_6848_7681# 0.11f
C2767 a_7989_2150# a_7804_1652# 0.231f
C2768 a_11756_5950# a_11834_7066# 0.198f
C2769 a_5488_7371# a_5173_7576# 0.0467f
C2770 a_15941_6827# a_15733_6827# 0.291f
C2771 a_2823_2688# a_2774_2878# 0.203f
C2772 a_16458_6583# d1 0.0235f
C2773 a_12915_2304# a_12919_2127# 0.518f
C2774 d0 a_18913_4684# 0.00533f
C2775 a_6851_1063# a_6570_1574# 0.11f
C2776 a_7803_3858# vdd 0.0273f
C2777 a_18958_3014# a_19166_3014# 0.448f
C2778 a_12914_5613# a_13901_5179# 0.283f
C2779 a_3824_6290# vdd 0.133f
C2780 a_15206_3169# a_15521_2964# 0.0467f
C2781 a_1584_6537# a_854_6781# 0.195f
C2782 a_10467_1271# a_10888_1271# 0.0104f
C2783 a_1374_1022# vdd 0.178f
C2784 a_648_2369# a_119_2479# 0.194f
C2785 a_15204_7581# a_15204_7124# 0.519f
C2786 a_16880_4377# vdd 0.0373f
C2787 a_5909_9028# a_6847_8784# 0.133f
C2788 a_7988_5459# a_8196_5459# 0.448f
C2789 a_1585_4331# a_1372_4331# 0.448f
C2790 a_12917_7642# vdd 0.0799f
C2791 a_13854_8501# a_12912_8922# 0.426f
C2792 a_18957_4117# a_18914_3581# 0.0185f
C2793 a_17972_1242# a_17831_1834# 0.133f
C2794 a_855_1815# a_119_2020# 0.255f
C2795 a_17968_8963# a_18017_8773# 0.243f
C2796 a_13903_3527# vdd 0.0325f
C2797 a_8884_1370# a_8878_2096# 0.0622f
C2798 a_3821_8124# a_2886_7637# 0.254f
C2799 a_6750_7102# vdd 0.0342f
C2800 a_7849_1639# vdd 0.0325f
C2801 a_7801_8270# vdd 0.0273f
C2802 d0 a_15519_9033# 0.0235f
C2803 a_6428_4372# d1 0.0235f
C2804 a_8880_9091# d0 0.00533f
C2805 a_15732_7376# a_15204_7581# 0.194f
C2806 a_9134_4112# a_8926_4112# 0.448f
C2807 a_16672_5480# a_15941_5170# 0.169f
C2808 a_18086_6056# a_17829_6246# 0.0467f
C2809 a_16882_1068# vdd 0.0273f
C2810 a_4077_9037# a_3869_9037# 0.448f
C2811 a_18957_7980# a_19165_7980# 0.448f
C2812 a_15941_7930# a_15520_7930# 0.0104f
C2813 a_2004_153# a_2774_5078# 0.177f
C2814 a_5176_1188# d0 0.0138f
C2815 a_11403_4336# vdd 0.178f
C2816 a_5488_7371# d0 0.0235f
C2817 a_10147_8873# a_10676_8992# 0.143f
C2818 a_12778_3822# a_13031_3809# 0.11f
C2819 a_8927_5769# vdd 0.0325f
C2820 a_15733_7930# a_15941_7930# 0.291f
C2821 a_119_3769# a_648_3472# 0.0185f
C2822 a_11836_2654# a_11758_1538# 0.198f
C2823 a_3000_3804# a_2747_3817# 0.11f
C2824 a_12773_6205# a_12803_7295# 0.14f
C2825 a_10677_5129# a_10149_4690# 0.011f
C2826 a_5175_3623# a_5910_4062# 0.155f
C2827 a_12852_7105# a_12913_7819# 0.0126f
C2828 a_10464_5129# d0 0.0235f
C2829 a_15207_1609# d0 0.00888f
C2830 a_11401_8748# d1 0.0235f
C2831 a_16890_4907# a_16897_2814# 0.583f
C2832 a_10148_7770# a_10677_7889# 0.143f
C2833 a_13172_3217# a_12964_3217# 0.448f
C2834 a_18956_9083# vdd 0.0325f
C2835 a_10148_8186# a_10462_8438# 0.11f
C2836 a_1373_3228# d1 0.0235f
C2837 a_15521_2964# d0 0.0235f
C2838 a_16882_1068# a_15943_758# 0.206f
C2839 a_10148_7083# a_10148_7540# 0.519f
C2840 a_3823_3712# a_2888_3225# 0.254f
C2841 a_10885_4026# a_11616_4336# 0.169f
C2842 a_8882_3022# a_9135_3009# 0.125f
C2843 a_5174_4726# a_5174_4497# 0.539f
C2844 a_3821_8124# a_3870_7934# 0.218f
C2845 a_11514_2654# a_11834_4866# 0.0104f
C2846 a_11841_2773# a_11617_3233# 0.0774f
C2847 a_12914_5613# vdd 0.439f
C2848 a_11826_1027# a_11545_1538# 0.11f
C2849 a_645_8987# a_116_9097# 0.194f
C2850 a_10885_5129# a_10886_5683# 0.498f
C2851 a_12918_5436# a_12963_5423# 0.181f
C2852 a_4080_2419# a_3827_2432# 0.11f
C2853 a_117_6662# vdd 0.128f
C2854 a_8881_6885# a_9134_6872# 0.11f
C2855 a_15205_5834# a_15940_6273# 0.155f
C2856 a_6851_1063# a_6643_1063# 0.241f
C2857 a_8883_816# d0 0.0138f
C2858 a_10150_3774# a_10150_3587# 0.0622f
C2859 a_6864_5021# vdd 0.0369f
C2860 a_2004_153# a_2883_5608# 0.137f
C2861 a_7802_6064# a_8055_6051# 0.11f
C2862 a_644_8433# vdd 0.0342f
C2863 a_7944_2163# a_8928_2460# 0.292f
C2864 a_11826_1027# a_10887_717# 0.206f
C2865 a_5174_5600# a_5490_5719# 0.125f
C2866 d0 a_13855_6295# 0.0138f
C2867 a_17975_2168# a_19167_2465# 0.0192f
C2868 a_6859_7102# a_6568_5986# 0.0104f
C2869 a_1805_2649# vdd 0.0269f
C2870 a_1810_2768# vdd 0.038f
C2871 a_6640_6578# a_5910_6822# 0.195f
C2872 a_119_3353# a_648_3472# 0.143f
C2873 a_18912_6890# vdd 0.145f
C2874 a_10680_1271# a_10888_1271# 0.291f
C2875 a_1512_5945# vdd 0.178f
C2876 a_5175_2707# d0 0.00888f
C2877 a_5174_6016# a_5174_5829# 0.0622f
C2878 a_1374_1022# a_856_712# 0.11f
C2879 a_15204_7581# vdd 0.312f
C2880 a_18958_4671# a_18909_4861# 0.218f
C2881 a_5910_5165# a_5489_5165# 0.0104f
C2882 a_18956_7426# a_19164_7426# 0.448f
C2883 a_3869_7380# a_3824_7393# 0.154f
C2884 a_15206_2712# vdd 0.143f
C2885 a_15944_1312# a_16461_1068# 0.0467f
C2886 a_13855_9055# a_13851_9232# 0.539f
C2887 a_1371_6537# a_1792_6537# 0.0104f
C2888 a_4078_6831# d0 0.0233f
C2889 a_2881_8917# a_3820_9227# 0.112f
C2890 a_15520_5170# a_15941_5170# 0.0104f
C2891 a_7937_8958# a_7986_8768# 0.243f
C2892 a_15206_2296# vdd 0.128f
C2893 a_12777_6028# a_12962_6526# 0.231f
C2894 a_3824_9050# d0 0.00533f
C2895 a_10463_7335# d0 0.0235f
C2896 a_18018_7670# a_18226_7670# 0.448f
C2897 a_6430_1063# d1 0.0235f
C2898 a_5174_4497# d0 0.0138f
C2899 a_12913_6716# a_13851_6472# 0.316f
C2900 a_6567_8192# a_6847_8784# 0.0467f
C2901 a_15732_6273# vdd 0.0342f
C2902 a_3872_2419# a_2888_2122# 0.292f
C2903 a_3139_7624# a_2886_7637# 0.11f
C2904 a_4080_3522# a_2888_3225# 0.0192f
C2905 a_8876_6508# a_8882_5782# 0.0622f
C2906 a_2742_6200# a_3140_5418# 0.0192f
C2907 a_15523_1312# a_15944_1312# 0.0104f
C2908 a_435_3472# a_648_3472# 0.448f
C2909 a_15204_8227# a_15731_8479# 0.14f
C2910 a_13060_7105# vdd 0.183f
C2911 a_14108_7385# a_13900_7385# 0.448f
C2912 a_15520_7930# d0 0.0235f
C2913 a_18908_8170# a_18912_7993# 0.539f
C2914 a_17878_6056# vdd 0.0325f
C2915 a_1803_4861# a_1694_4861# 0.117f
C2916 a_19165_6877# a_18912_6890# 0.11f
C2917 a_7937_8958# a_8875_8714# 0.316f
C2918 a_18914_3581# vdd 0.135f
C2919 a_853_6227# a_1792_6537# 0.302f
C2920 a_1803_7061# a_1808_7180# 0.464f
C2921 a_16672_5480# a_16459_5480# 0.448f
C2922 a_8197_2150# a_7940_2340# 0.0467f
C2923 a_6642_3269# a_5911_2959# 0.169f
C2924 a_16672_4377# a_15942_4621# 0.195f
C2925 a_18225_8773# a_17968_8963# 0.0467f
C2926 a_15734_1861# vdd 0.0342f
C2927 a_10147_8643# a_10675_8438# 0.194f
C2928 a_8878_5959# a_8881_5228# 0.0292f
C2929 a_6426_8784# a_6639_8784# 0.448f
C2930 a_432_8987# vdd 0.178f
C2931 a_12915_3407# vdd 0.439f
C2932 a_8085_7141# vdd 0.183f
C2933 a_5491_753# a_5912_753# 0.0104f
C2934 a_5172_8679# a_5908_8474# 0.255f
C2935 a_7802_6064# vdd 0.0273f
C2936 a_119_2666# a_119_3123# 0.519f
C2937 a_8878_4856# a_8882_4679# 0.539f
C2938 a_8881_6885# a_8925_7421# 0.0185f
C2939 a_12962_7629# a_13170_7629# 0.448f
C2940 d0 a_5178_859# 0.00888f
C2941 a_10679_2374# a_10887_2374# 0.291f
C2942 a_854_6781# a_646_6781# 0.291f
C2943 a_1372_5434# a_1793_5434# 0.0104f
C2944 a_5173_6932# vdd 0.323f
C2945 a_18909_5964# a_19166_5774# 0.0467f
C2946 a_18957_4117# a_19165_4117# 0.448f
C2947 a_122_818# a_2004_153# 0.252f
C2948 a_3871_5728# vdd 0.0325f
C2949 a_8884_1370# a_8880_1547# 0.539f
C2950 a_16890_4907# a_16892_2695# 0.206f
C2951 a_12914_4510# a_13853_4820# 0.112f
C2952 a_3825_5187# a_2883_5608# 0.426f
C2953 a_9135_5769# a_8882_5782# 0.11f
C2954 a_1682_153# vdd 0.178f
C2955 d1 a_13170_7629# 0.0233f
C2956 a_13850_8678# a_13901_7939# 0.011f
C2957 a_15939_8479# a_15204_8227# 0.279f
C2958 a_11402_6542# a_11823_6542# 0.0104f
C2959 a_16674_1068# a_15944_1312# 0.219f
C2960 a_15944_1312# a_15207_1422# 0.277f
C2961 d0 a_432_6227# 0.0235f
C2962 a_1513_3739# a_1810_2768# 0.0104f
C2963 a_119_3123# a_647_2918# 0.194f
C2964 a_13901_6836# a_13852_7026# 0.218f
C2965 a_11617_3233# a_11404_3233# 0.448f
C2966 a_5174_5600# a_5703_5719# 0.143f
C2967 a_10885_7889# a_10464_7889# 0.0104f
C2968 a_5173_7576# a_5701_7371# 0.194f
C2969 a_9566_17# vout 0.0104f
C2970 a_12918_5436# vdd 0.0799f
C2971 a_18019_4361# a_17970_4551# 0.243f
C2972 a_6427_6578# vdd 0.178f
C2973 a_6642_2166# vdd 0.0342f
C2974 a_12961_8732# vdd 0.0325f
C2975 a_5175_2707# a_5704_2410# 0.0185f
C2976 a_1724_8151# a_1792_7640# 0.146f
C2977 a_7804_1652# a_7940_2340# 0.345f
C2978 a_4079_5728# a_3826_5741# 0.11f
C2979 a_12035_158# a_13062_4893# 0.0192f
C2980 a_10150_3774# a_10149_4231# 0.519f
C2981 a_11725_7066# a_11512_7066# 0.448f
C2982 a_15203_8914# vdd 0.128f
C2983 a_8883_3576# vdd 0.135f
C2984 a_17861_5124# a_17865_2747# 0.685f
C2985 a_12915_2304# vdd 0.439f
C2986 a_13854_2614# a_13858_2437# 0.539f
C2987 a_1370_8743# a_1583_8743# 0.448f
C2988 a_15204_6478# vdd 0.312f
C2989 a_6642_3269# vdd 0.0342f
C2990 a_16598_8197# a_16895_7226# 0.0104f
C2991 a_15206_3399# a_15522_3518# 0.125f
C2992 a_1794_2125# a_855_1815# 0.302f
C2993 a_3001_1598# a_2744_1788# 0.0467f
C2994 a_6783_1574# vdd 0.0342f
C2995 a_646_5124# vdd 0.0342f
C2996 a_16814_1579# a_16882_1068# 0.146f
C2997 a_13853_5923# vdd 0.311f
C2998 a_7800_1829# a_7849_1639# 0.22f
C2999 a_8877_5405# a_9134_5215# 0.0467f
C3000 a_18957_4117# a_18912_4130# 0.154f
C3001 a_3872_3522# a_2888_3225# 0.292f
C3002 a_13856_4089# a_13853_4820# 0.0292f
C3003 a_13856_7952# a_13852_8129# 0.539f
C3004 d0 a_14111_3527# 0.0233f
C3005 a_13901_7939# a_14109_7939# 0.448f
C3006 a_10150_3774# a_10679_3477# 0.0185f
C3007 a_7830_5119# a_7940_3443# 0.132f
C3008 a_18086_6056# vdd 0.183f
C3009 a_6642_3269# a_6429_3269# 0.448f
C3010 a_8881_4125# d0 0.0138f
C3011 a_11725_4866# a_11839_4985# 0.178f
C3012 a_6537_7102# a_6750_7102# 0.448f
C3013 a_1696_2649# a_1483_2649# 0.448f
C3014 a_13855_9055# vdd 0.00337f
C3015 a_12807_7118# a_12776_8234# 0.206f
C3016 a_6866_2809# a_6849_4372# 0.14f
C3017 a_17972_8786# a_17832_8275# 0.206f
C3018 a_8881_6885# a_8926_6872# 0.151f
C3019 a_10149_5980# a_10678_5683# 0.0185f
C3020 a_1726_3739# a_1794_3228# 0.146f
C3021 a_15206_3815# a_15941_4067# 0.279f
C3022 a_3140_5418# d1 0.0233f
C3023 a_17969_7860# a_17863_7159# 0.423f
C3024 a_12913_6716# a_12777_6028# 0.345f
C3025 a_16881_2171# a_16892_2695# 0.328f
C3026 a_1795_1022# a_1727_1533# 0.146f
C3027 a_15520_6827# a_15941_6827# 0.0104f
C3028 a_5911_1856# a_5490_1856# 0.0104f
C3029 a_15204_6478# a_15204_6708# 0.0292f
C3030 a_118_4456# a_118_4226# 0.0292f
C3031 a_18229_1052# a_18021_1052# 0.448f
C3032 a_5489_6822# a_5702_6822# 0.448f
C3033 a_2790_8216# a_2776_7113# 0.19f
C3034 a_5910_4062# vdd 0.0799f
C3035 a_119_2666# a_647_2918# 0.14f
C3036 a_12778_3822# a_12914_4510# 0.345f
C3037 a_7987_6562# vdd 0.0325f
C3038 a_7988_4356# a_7943_4369# 0.181f
C3039 a_18088_1644# a_17835_1657# 0.11f
C3040 a_10884_7335# vdd 0.1f
C3041 a_16457_8789# d1 0.0235f
C3042 a_119_3769# d0 0.00888f
C3043 a_3821_7021# vdd 0.311f
C3044 a_1805_2649# a_1514_1533# 0.0104f
C3045 a_856_2369# vdd 0.454f
C3046 a_3140_4315# vdd 0.183f
C3047 a_2746_6023# a_3139_6521# 0.0192f
C3048 a_118_4685# a_647_4575# 0.194f
C3049 a_6426_8784# a_5908_8474# 0.11f
C3050 a_117_6891# a_117_7078# 0.0625f
C3051 a_5176_1417# vdd 0.323f
C3052 a_17880_1644# a_17831_1834# 0.22f
C3053 a_855_4575# a_854_4021# 0.498f
C3054 a_5488_9028# a_5172_8909# 0.125f
C3055 a_15206_3169# a_15942_2964# 0.255f
C3056 a_16878_8789# a_16457_8789# 0.0104f
C3057 a_17969_7860# a_17828_8452# 0.133f
C3058 a_118_5559# vdd 0.128f
C3059 a_10886_5683# a_10678_5683# 0.291f
C3060 a_12916_1201# a_12965_1011# 0.219f
C3061 a_15941_4067# a_16880_4377# 0.302f
C3062 a_10679_717# a_10466_717# 0.448f
C3063 a_10150_3587# vdd 0.323f
C3064 d0 a_19164_7426# 0.0233f
C3065 a_5912_2410# vdd 0.454f
C3066 a_16598_8197# a_16811_8197# 0.448f
C3067 a_18907_6513# vdd 0.314f
C3068 a_6861_2690# vdd 0.0269f
C3069 a_1725_5945# vdd 0.0342f
C3070 a_18914_3581# a_17975_3271# 0.278f
C3071 a_5174_4267# a_5910_4062# 0.255f
C3072 a_5173_8222# a_5173_8035# 0.0622f
C3073 a_6864_5021# a_6537_7102# 0.0104f
C3074 a_14108_6282# d0 0.0233f
C3075 a_16600_3785# a_16880_4377# 0.0467f
C3076 a_13062_2693# a_12854_2693# 0.448f
C3077 a_16460_3274# d1 0.0235f
C3078 a_854_4021# vdd 0.0799f
C3079 a_856_3472# a_119_3123# 0.112f
C3080 a_19165_4117# vdd 0.183f
C3081 a_8879_3753# vdd 0.311f
C3082 a_10678_4580# a_10149_4461# 0.143f
C3083 a_119_3769# a_433_4021# 0.11f
C3084 a_2774_5078# a_3031_2688# 0.0192f
C3085 a_5173_7806# a_5489_7925# 0.125f
C3086 a_2883_4505# a_3825_4084# 0.426f
C3087 a_2888_3225# a_2884_3402# 0.518f
C3088 a_120_1376# a_647_1815# 0.011f
C3089 a_431_8433# vdd 0.178f
C3090 a_12852_7105# vdd 0.0325f
C3091 a_5911_4616# vdd 0.454f
C3092 a_10887_2374# a_10466_2374# 0.0104f
C3093 a_5174_5600# d0 0.0138f
C3094 a_13901_7939# vdd 0.0325f
C3095 d3 a_1483_2649# 0.0235f
C3096 a_119_3353# d0 0.0138f
C3097 a_13900_6282# a_13855_6295# 0.154f
C3098 a_12915_2304# a_12964_2114# 0.243f
C3099 a_7988_5459# vdd 0.0325f
C3100 a_17865_2747# a_17971_3448# 0.392f
C3101 a_5702_7925# a_5173_8222# 0.0185f
C3102 a_18911_7439# vdd 0.133f
C3103 a_1792_7640# a_853_7330# 0.206f
C3104 a_120_1147# vdd 0.128f
C3105 a_2778_2701# a_2933_3212# 0.0267f
C3106 a_11713_158# d5 0.0235f
C3107 a_15205_4502# a_15942_4621# 0.426f
C3108 a_12917_7642# a_13170_7629# 0.11f
C3109 a_5703_5719# a_5174_6016# 0.0185f
C3110 a_17833_6069# a_17859_7336# 0.347f
C3111 a_5911_1856# a_6429_2166# 0.11f
C3112 a_18019_5464# a_17970_5654# 0.219f
C3113 a_5176_1604# a_5911_1856# 0.279f
C3114 a_12809_2706# a_12823_3809# 0.19f
C3115 a_13899_8488# a_14107_8488# 0.448f
C3116 d0 a_3826_1878# 0.0138f
C3117 a_13902_2973# a_12915_3407# 0.283f
C3118 a_10149_5564# a_10678_5683# 0.143f
C3119 a_435_3472# d0 0.0235f
C3120 a_5174_4267# a_5911_4616# 0.112f
C3121 a_12824_1603# a_13032_1603# 0.448f
C3122 a_2933_2109# a_2748_1611# 0.231f
C3123 a_435_712# vdd 0.178f
C3124 a_18912_4130# vdd 0.133f
C3125 a_13902_1870# a_14110_1870# 0.448f
C3126 a_6640_7681# a_6848_7681# 0.241f
C3127 a_15736_1312# vdd 0.0342f
C3128 a_16460_2171# d1 0.0235f
C3129 a_11405_1027# d1 0.0235f
C3130 a_6752_2690# vdd 0.0342f
C3131 a_5701_6268# a_5488_6268# 0.448f
C3132 a_12777_6028# a_13030_6015# 0.11f
C3133 a_15205_4272# vdd 0.312f
C3134 a_5053_133# a_5178_859# 1.05f
C3135 a_8877_8165# a_8880_7434# 0.0292f
C3136 a_3824_7393# vdd 0.133f
C3137 a_10150_3128# a_10150_3358# 0.0292f
C3138 a_15943_3518# vdd 0.455f
C3139 a_15522_2415# d0 0.0235f
C3140 a_10467_1271# d0 0.0235f
C3141 a_7939_5649# a_9134_5215# 0.0192f
C3142 a_118_4872# vdd 0.144f
C3143 a_10676_6232# vdd 0.0342f
C3144 a_1902_4861# a_2774_5078# 0.0189f
C3145 a_433_5124# vdd 0.178f
C3146 a_12822_6015# a_12803_7295# 0.255f
C3147 a_11824_5439# a_11823_6542# 0.504f
C3148 a_10887_3477# vdd 0.455f
C3149 a_11824_5439# a_10886_5683# 0.322f
C3150 a_10886_4580# a_11403_4336# 0.0467f
C3151 a_10888_1271# vdd 0.455f
C3152 a_10149_4877# a_10885_5129# 0.279f
C3153 a_2886_6534# a_3825_6844# 0.278f
C3154 a_18907_6513# a_18913_5787# 0.0622f
C3155 a_11756_5950# a_11824_5439# 0.146f
C3156 a_18913_1924# vdd 0.133f
C3157 a_11825_3233# vdd 0.0273f
C3158 a_3870_4071# a_3825_4084# 0.154f
C3159 a_3140_4315# a_2747_3817# 0.0192f
C3160 a_5174_5829# vdd 0.323f
C3161 a_5489_5165# d0 0.0235f
C3162 a_10149_4231# vdd 0.312f
C3163 a_8196_4356# a_7988_4356# 0.448f
C3164 a_12134_158# a_14876_138# 0.194f
C3165 a_18118_4934# vdd 0.183f
C3166 a_5702_4062# a_5175_3623# 0.011f
C3167 a_17970_4551# a_18908_4307# 0.316f
C3168 a_12774_3999# a_13031_3809# 0.0467f
C3169 a_15520_6827# a_15733_6827# 0.448f
C3170 a_16890_7107# a_16599_5991# 0.0104f
C3171 a_3823_2609# a_2888_2122# 0.254f
C3172 a_3823_2609# a_2884_2299# 0.112f
C3173 a_5702_5165# a_5174_5370# 0.194f
C3174 a_433_7884# vdd 0.178f
C3175 a_8877_8165# a_7938_7855# 0.112f
C3176 a_6641_4372# a_6849_4372# 0.26f
C3177 a_6428_4372# a_5910_4062# 0.11f
C3178 a_15203_9143# a_15519_9033# 0.0467f
C3179 a_5912_753# vdd 0.021f
C3180 a_18957_7980# a_18908_8170# 0.218f
C3181 a_5175_3164# a_5912_3513# 0.112f
C3182 a_13856_5192# d0 0.0138f
C3183 a_10466_3477# vdd 0.178f
C3184 a_120_1563# vdd 0.135f
C3185 a_10679_3477# vdd 0.0342f
C3186 a_5175_3623# a_5175_3810# 0.0622f
C3187 d0 a_434_5678# 0.0235f
C3188 a_7834_2742# a_8087_2729# 0.11f
C3189 a_5492_1307# a_5176_1417# 0.0467f
C3190 a_3826_5741# a_3871_5728# 0.151f
C3191 a_17972_8786# vdd 0.021f
C3192 a_8879_2650# vdd 0.311f
C3193 a_16895_5026# a_16879_6583# 0.122f
C3194 a_15206_2525# a_15942_2964# 0.155f
C3195 a_5489_7925# d0 0.0235f
C3196 a_3824_9050# a_3820_9227# 0.539f
C3197 a_2882_7814# a_2886_7637# 0.518f
C3198 a_5909_6268# a_5488_6268# 0.0104f
C3199 d3 a_6539_2690# 0.0235f
C3200 a_16982_199# a_15209_864# 0.0111f
C3201 a_12918_5436# a_14110_5733# 0.0192f
C3202 a_5910_5165# vdd 0.104f
C3203 a_435_712# a_856_712# 0.0104f
C3204 d0 a_5174_6016# 0.00888f
C3205 a_4954_133# a_7060_194# 0.294f
C3206 a_855_4575# a_1372_4331# 0.0467f
C3207 a_11512_7066# vdd 0.178f
C3208 a_7834_2742# a_7830_5119# 0.685f
C3209 a_122_818# a_120_917# 0.519f
C3210 a_15206_2525# a_15522_2415# 0.0467f
C3211 a_3824_1506# a_3828_1329# 0.539f
C3212 a_11823_7645# a_11615_7645# 0.241f
C3213 a_852_8433# a_1583_8743# 0.169f
C3214 a_18957_6877# vdd 0.0325f
C3215 a_8880_7434# d0 0.0138f
C3216 a_18913_3027# vdd 0.133f
C3217 a_4078_7934# a_2886_7637# 0.0192f
C3218 a_2885_8740# vdd 0.021f
C3219 a_1372_4331# vdd 0.178f
C3220 a_3869_6277# a_3824_6290# 0.154f
C3221 a_117_6891# vdd 0.323f
C3222 a_5911_4616# a_6428_4372# 0.0467f
C3223 a_12777_6028# a_13170_6526# 0.0192f
C3224 a_18085_8262# a_17832_8275# 0.11f
C3225 a_11402_7645# a_10885_7889# 0.0467f
C3226 a_2887_4328# a_3822_4815# 0.254f
C3227 a_7828_7331# a_7832_7154# 0.606f
C3228 a_13853_5923# a_14110_5733# 0.0467f
C3229 a_17910_4934# vdd 0.0325f
C3230 a_5491_753# d0 0.0235f
C3231 a_8927_4666# a_8877_5405# 0.011f
C3232 a_18958_4671# a_18908_5410# 0.011f
C3233 a_8056_3845# a_7799_4035# 0.0467f
C3234 a_6849_5475# a_6641_5475# 0.241f
C3235 a_10147_8873# a_10884_8992# 0.426f
C3236 a_6570_1574# a_6783_1574# 0.448f
C3237 a_17879_3850# a_17865_2747# 0.19f
C3238 a_16671_6583# a_16879_6583# 0.26f
C3239 a_10465_1820# a_10678_1820# 0.448f
C3240 a_7943_4369# vdd 0.0988f
C3241 a_122_818# a_1902_4861# 0.247f
C3242 a_5172_9138# vdd 0.323f
C3243 a_5175_3623# a_5912_3513# 0.277f
C3244 a_8196_5459# a_7943_5472# 0.11f
C3245 a_18957_6877# a_19165_6877# 0.448f
C3246 a_12773_6205# a_12963_5423# 0.251f
C3247 a_11933_4866# a_11926_158# 0.178f
C3248 a_5173_8222# a_5487_8474# 0.11f
C3249 a_3869_7380# a_3820_7570# 0.218f
C3250 a_11757_3744# a_11825_3233# 0.146f
C3251 a_3871_4625# a_3822_4815# 0.218f
C3252 a_12775_1793# a_12779_1616# 0.518f
C3253 a_5705_1307# a_5176_1417# 0.194f
C3254 a_5703_1856# vdd 0.0342f
C3255 a_1373_2125# a_855_1815# 0.11f
C3256 a_14108_6282# a_13900_6282# 0.448f
C3257 a_4078_7934# a_3870_7934# 0.448f
C3258 a_16890_4907# a_16989_4907# 0.814f
C3259 a_122_818# a_648_712# 0.187f
C3260 a_11825_2130# vdd 0.0373f
C3261 a_5490_5719# vdd 0.178f
C3262 a_14111_2424# d0 0.0233f
C3263 a_9136_3563# vdd 0.183f
C3264 a_8877_8165# a_8926_7975# 0.218f
C3265 a_18958_3014# a_18914_2478# 0.0185f
C3266 a_15521_5724# a_15205_5834# 0.0467f
C3267 a_7940_2340# a_9135_1906# 0.0192f
C3268 a_11841_2773# a_11834_4866# 0.583f
C3269 a_10675_8438# vdd 0.0342f
C3270 a_1373_2125# a_1794_2125# 0.0104f
C3271 a_6428_5475# d1 0.0235f
C3272 a_648_3472# vdd 0.0342f
C3273 a_4079_2968# d0 0.0233f
C3274 a_8056_3845# vdd 0.183f
C3275 d0 a_10465_2923# 0.0235f
C3276 a_13852_7026# vdd 0.311f
C3277 a_2887_5431# a_3820_6467# 0.155f
C3278 a_8882_1919# vdd 0.133f
C3279 a_8884_1370# a_9137_1357# 0.11f
C3280 a_3870_4071# a_3827_3535# 0.0185f
C3281 a_13903_767# a_14111_767# 0.448f
C3282 a_5701_6268# a_5909_6268# 0.3f
C3283 a_117_7078# d0 0.00888f
C3284 a_10150_3774# d0 0.00888f
C3285 a_10886_1820# vdd 0.0799f
C3286 a_13855_1511# vdd 0.311f
C3287 a_11823_7645# a_11839_7185# 0.348f
C3288 a_16672_5480# a_15942_5724# 0.219f
C3289 a_2774_5078# a_2884_3402# 0.132f
C3290 a_10149_4877# a_10678_4580# 0.0185f
C3291 a_7938_6752# a_8876_6508# 0.316f
C3292 a_5490_2959# d0 0.0235f
C3293 a_15734_5724# a_15942_5724# 0.291f
C3294 a_13173_1011# vdd 0.183f
C3295 a_13858_780# a_14111_767# 0.125f
C3296 a_15520_5170# a_15733_5170# 0.448f
C3297 a_3870_6831# vdd 0.0325f
C3298 a_13032_1603# vdd 0.183f
C3299 a_435_2369# vdd 0.178f
C3300 a_4079_1865# a_2884_2299# 0.0192f
C3301 a_13169_8732# d1 0.0233f
C3302 a_15207_1609# a_15207_1422# 0.0622f
C3303 a_1792_6537# vdd 0.0373f
C3304 a_1586_2125# vdd 0.0342f
C3305 a_17969_7860# a_18907_7616# 0.316f
C3306 a_6570_1574# a_6861_2690# 0.0104f
C3307 a_17969_6757# a_17859_7336# 0.285f
C3308 a_16673_3274# a_15943_3518# 0.219f
C3309 a_1370_8743# a_1791_8743# 0.0104f
C3310 a_18018_7670# vdd 0.0325f
C3311 a_5702_7925# a_5173_8035# 0.194f
C3312 a_5910_5165# a_5174_4913# 0.279f
C3313 a_15209_864# vdd 0.0974f
C3314 a_13858_3540# a_13854_3717# 0.539f
C3315 a_13851_7575# a_13901_6836# 0.011f
C3316 a_14110_2973# a_12915_3407# 0.0192f
C3317 a_10149_4877# a_10464_5129# 0.11f
C3318 a_10148_7770# a_10464_7889# 0.125f
C3319 a_18956_7426# vdd 0.0325f
C3320 a_116_9097# vref 0.034f
C3321 a_8927_1906# a_8882_1919# 0.154f
C3322 a_855_5678# a_118_5559# 0.426f
C3323 a_8195_6562# d1 0.0233f
C3324 a_6864_5021# a_7060_194# 0.0424f
C3325 a_12918_5436# a_13857_5746# 0.278f
C3326 a_11542_8156# d2 0.0235f
C3327 a_3819_8673# vdd 0.314f
C3328 a_11514_2654# vdd 0.178f
C3329 a_12964_3217# vdd 0.0325f
C3330 a_2886_6534# a_2746_6023# 0.206f
C3331 a_5175_2061# a_5175_2291# 0.0292f
C3332 a_15206_3628# vdd 0.323f
C3333 a_1794_3228# a_1793_4331# 0.498f
C3334 d2 a_8055_6051# 0.0233f
C3335 a_6738_194# d5 0.0235f
C3336 a_10148_7999# a_10675_8438# 0.011f
C3337 a_116_8638# vdd 0.312f
C3338 a_16890_4907# a_17861_5124# 0.409f
C3339 a_18906_8719# a_19163_8529# 0.0467f
C3340 a_15209_864# a_15943_758# 1.07f
C3341 a_12778_3822# a_12809_2706# 0.206f
C3342 a_19167_808# d0 0.0233f
C3343 a_15205_4502# a_15734_4621# 0.143f
C3344 a_9133_6318# vdd 0.183f
C3345 a_12963_5423# a_13171_5423# 0.448f
C3346 a_18118_4934# d4 0.0233f
C3347 d0 a_15205_5605# 0.0138f
C3348 a_10153_823# a_12134_158# 0.53f
C3349 a_4632_133# a_4954_133# 0.11f
C3350 a_10466_717# vdd 0.178f
C3351 a_6848_6578# a_5909_6268# 0.302f
C3352 a_5173_7806# vdd 0.128f
C3353 a_10153_823# a_10887_717# 1.07f
C3354 a_13853_5923# a_13857_5746# 0.539f
C3355 a_7801_8270# a_7846_8257# 0.157f
C3356 a_15205_5375# a_15205_4918# 0.519f
C3357 a_12913_6716# a_12962_6526# 0.243f
C3358 a_2004_153# a_1902_4861# 7.78f
C3359 a_6850_3269# a_6849_4372# 0.498f
C3360 a_5702_4062# vdd 0.0342f
C3361 a_18088_1644# a_17831_1834# 0.0467f
C3362 a_4079_4625# d0 0.0233f
C3363 a_5909_9028# vdd 0.454f
C3364 a_1371_7640# d1 0.0235f
C3365 a_12913_7819# a_13855_7398# 0.426f
C3366 a_4076_8483# a_3819_8673# 0.0467f
C3367 a_5703_5719# vdd 0.0342f
C3368 a_19168_1362# d0 0.0233f
C3369 a_17970_5654# a_17974_5477# 0.518f
C3370 a_8878_3199# a_7944_2163# 0.155f
C3371 a_12773_6205# vdd 0.0316f
C3372 a_10677_5129# a_10149_5334# 0.194f
C3373 a_16989_4907# a_17861_5124# 0.0189f
C3374 a_17972_1242# a_17976_1065# 0.518f
C3375 a_1808_4980# a_854_6781# 0.132f
C3376 a_117_7535# a_117_7765# 0.0292f
C3377 a_15941_4067# a_15205_4272# 0.255f
C3378 a_14109_5179# a_12914_5613# 0.0192f
C3379 a_8878_5959# a_8927_5769# 0.218f
C3380 a_5175_3810# vdd 0.135f
C3381 a_8928_2460# vdd 0.0325f
C3382 a_8877_8165# vdd 0.311f
C3383 a_19167_808# a_18959_808# 0.448f
C3384 a_5911_2959# a_5912_3513# 0.498f
C3385 a_2886_7637# a_3870_7934# 0.292f
C3386 a_3827_775# d0 0.0138f
C3387 a_12854_4893# a_12809_4906# 0.128f
C3388 a_15940_7376# a_15204_7581# 0.255f
C3389 a_15206_2712# a_15735_2415# 0.0185f
C3390 a_12917_7642# a_12962_7629# 0.181f
C3391 a_8196_4356# vdd 0.183f
C3392 a_2778_2701# a_2743_3994# 0.298f
C3393 a_15204_7124# d0 0.00888f
C3394 a_1374_1022# d1 0.0235f
C3395 a_6850_3269# a_6866_2809# 0.348f
C3396 a_15206_2296# a_15735_2415# 0.143f
C3397 a_5702_4062# a_5174_4267# 0.194f
C3398 a_15207_1609# a_15521_1861# 0.11f
C3399 a_18910_998# a_15209_864# 0.884f
C3400 a_19163_8529# vdd 0.183f
C3401 a_10150_2025# a_10150_2255# 0.0292f
C3402 a_17975_2168# a_17971_2345# 0.518f
C3403 a_2774_5078# a_2778_4901# 0.518f
C3404 a_15941_7930# vdd 0.455f
C3405 a_11618_1027# vdd 0.0342f
C3406 a_7828_7331# a_7834_4942# 0.681f
C3407 a_13857_4643# a_13902_4630# 0.151f
C3408 a_16895_5026# a_16781_7107# 0.342f
C3409 a_12916_8745# a_12912_8922# 0.518f
C3410 a_18958_5774# a_19166_5774# 0.448f
C3411 a_19166_3014# vdd 0.183f
C3412 a_16813_3785# a_16897_2814# 0.263f
C3413 a_14109_7939# d0 0.0233f
C3414 a_10465_4580# a_10149_4690# 0.0467f
C3415 a_17865_4947# a_17859_7336# 0.681f
C3416 a_5175_2520# a_5175_2707# 0.0625f
C3417 d2 vdd 1.42f
C3418 a_2881_8917# a_2745_8229# 0.345f
C3419 a_13851_7575# a_12913_7819# 0.316f
C3420 a_2998_8216# vdd 0.183f
C3421 a_13853_2060# a_12915_2304# 0.316f
C3422 a_11926_158# vdd 0.0342f
C3423 a_2881_8917# a_3868_8483# 0.283f
C3424 a_12920_1024# vdd 0.0799f
C3425 a_11544_3744# vdd 0.178f
C3426 a_5174_4267# a_5175_3810# 0.519f
C3427 a_1584_7640# a_854_7884# 0.219f
C3428 a_11823_7645# a_11755_8156# 0.146f
C3429 a_18085_8262# vdd 0.183f
C3430 a_17973_6580# a_17859_7336# 0.0437f
C3431 a_15206_3169# vdd 0.312f
C3432 a_12035_158# a_12134_158# 0.527f
C3433 a_7828_7331# a_7798_6241# 0.14f
C3434 a_11616_5439# a_11403_5439# 0.448f
C3435 a_8087_4929# a_7834_4942# 0.11f
C3436 a_6430_1063# a_5912_753# 0.11f
C3437 a_6951_194# a_6958_4902# 0.178f
C3438 a_2746_6023# a_2882_6711# 0.345f
C3439 a_434_4575# d0 0.0235f
C3440 a_11403_4336# d1 0.0235f
C3441 a_13062_2693# vdd 0.183f
C3442 a_2887_5431# a_2883_5608# 0.518f
C3443 a_5173_7576# vdd 0.312f
C3444 a_12809_4906# a_12803_7295# 0.681f
C3445 a_15203_8684# vdd 0.312f
C3446 a_11823_6542# a_10885_6786# 0.133f
C3447 a_15943_3518# a_15522_3518# 0.0104f
C3448 a_5174_4726# vdd 0.323f
C3449 a_2883_5608# a_2778_4901# 0.0518f
C3450 a_15207_963# vdd 0.312f
C3451 a_856_3472# a_1794_3228# 0.322f
C3452 a_5173_6703# a_5173_6932# 0.539f
C3453 a_16881_3274# a_16897_2814# 0.348f
C3454 a_18909_4861# a_18913_4684# 0.539f
C3455 a_2103_153# a_5053_133# 0.152f
C3456 a_18909_5964# a_18958_5774# 0.218f
C3457 a_1791_8743# a_1808_7180# 0.14f
C3458 a_9137_1357# a_8880_1547# 0.0467f
C3459 d0 a_3826_2981# 0.0138f
C3460 a_16568_7107# d3 0.0235f
C3461 a_5912_3513# vdd 0.455f
C3462 a_18914_3581# a_18959_3568# 0.151f
C3463 a_8877_7062# a_8880_6331# 0.0292f
C3464 a_18228_2155# a_17971_2345# 0.0467f
C3465 a_16989_4907# a_16769_199# 0.0467f
C3466 a_1808_4980# a_2004_153# 0.0424f
C3467 a_5173_6473# a_5910_6822# 0.112f
C3468 a_8925_6318# a_9133_6318# 0.448f
C3469 a_9135_4666# a_8927_4666# 0.448f
C3470 a_3823_8496# vdd 0.133f
C3471 a_120_1376# a_855_1815# 0.155f
C3472 a_10153_823# a_12035_158# 0.252f
C3473 a_13171_5423# vdd 0.183f
C3474 a_18910_2655# vdd 0.311f
C3475 a_15733_4067# vdd 0.0342f
C3476 a_6569_3780# d2 0.0235f
C3477 a_17865_2747# a_18118_2734# 0.11f
C3478 a_10147_8643# a_10462_8438# 0.0467f
C3479 a_6851_1063# a_6783_1574# 0.146f
C3480 a_853_8987# a_645_8987# 0.291f
C3481 a_648_2369# vdd 0.0342f
C3482 a_19166_1911# vdd 0.183f
C3483 a_6429_3269# a_5912_3513# 0.0467f
C3484 a_6567_8192# vdd 0.178f
C3485 a_15207_963# a_15943_758# 0.255f
C3486 a_16673_2171# a_15942_1861# 0.169f
C3487 a_10148_6667# a_10148_6437# 0.0292f
C3488 a_6958_4902# a_6859_4902# 0.814f
C3489 a_7942_6575# a_8876_7611# 0.155f
C3490 a_116_8868# a_432_8987# 0.125f
C3491 a_6859_7102# a_6640_6578# 0.0267f
C3492 a_10886_4580# a_10149_4231# 0.112f
C3493 a_7989_2150# a_7944_2163# 0.181f
C3494 a_12774_3999# a_12919_3230# 0.326f
C3495 a_5702_5165# a_5489_5165# 0.448f
C3496 a_18908_8170# a_19165_7980# 0.0467f
C3497 d0 vdd 5.7f
C3498 a_10677_4026# a_10464_4026# 0.448f
C3499 a_2931_7624# a_2776_7113# 0.0267f
C3500 a_2885_8740# a_2930_8727# 0.181f
C3501 a_1513_3739# d2 0.0235f
C3502 d0 a_18912_5233# 0.0138f
C3503 a_2772_7290# vdd 0.0321f
C3504 a_10150_3774# a_10885_4026# 0.279f
C3505 a_4076_8483# a_3823_8496# 0.125f
C3506 a_17975_2168# a_18228_2155# 0.11f
C3507 a_11834_7066# a_11543_5950# 0.0104f
C3508 a_3820_7570# vdd 0.314f
C3509 a_9566_17# a_9779_17# 0.448f
C3510 a_5173_8222# a_5908_8474# 0.279f
C3511 a_18910_3758# vdd 0.311f
C3512 a_6848_6578# a_6864_5021# 0.122f
C3513 a_1370_8743# vdd 0.178f
C3514 a_15734_5724# a_15205_5605# 0.143f
C3515 a_8057_1639# a_7830_2919# 0.0192f
C3516 a_117_6662# a_433_6781# 0.125f
C3517 a_6780_8192# a_6864_7221# 0.263f
C3518 a_11617_3233# a_10886_2923# 0.169f
C3519 a_13853_4820# a_13902_4630# 0.218f
C3520 a_117_7994# a_644_8433# 0.011f
C3521 a_5912_2410# a_5491_2410# 0.0104f
C3522 a_6643_1063# a_5912_753# 0.169f
C3523 a_2888_3225# a_3141_3212# 0.11f
C3524 a_433_4021# vdd 0.178f
C3525 a_2821_7100# a_2882_7814# 0.0126f
C3526 a_4076_8483# d0 0.0233f
C3527 d0 a_18915_1375# 0.00533f
C3528 a_8875_8714# a_8924_8524# 0.218f
C3529 a_15204_6708# d0 0.0138f
C3530 a_7847_6051# a_7802_6064# 0.157f
C3531 a_6848_7681# a_5910_7925# 0.322f
C3532 a_19165_6877# d0 0.0233f
C3533 a_18959_808# vdd 0.0325f
C3534 a_15518_8479# vdd 0.178f
C3535 a_11757_3744# a_11544_3744# 0.448f
C3536 a_3031_4888# a_2774_5078# 0.0467f
C3537 a_11825_2130# a_11758_1538# 0.195f
C3538 a_12914_4510# a_13171_4320# 0.0467f
C3539 a_12778_3822# a_12963_4320# 0.231f
C3540 a_854_4021# a_118_4226# 0.255f
C3541 a_18018_6567# a_17859_7336# 0.0774f
C3542 a_6851_1063# a_6861_2690# 0.206f
C3543 a_1587_1022# vdd 0.0342f
C3544 a_17859_7336# a_17863_7159# 0.606f
C3545 a_6426_8784# a_6847_8784# 0.0104f
C3546 a_16460_3274# a_15943_3518# 0.0467f
C3547 a_3824_1506# a_4081_1316# 0.0467f
C3548 a_3826_4638# a_2887_4328# 0.278f
C3549 a_5174_4726# a_5174_4913# 0.0625f
C3550 a_17861_5124# a_17971_3448# 0.132f
C3551 a_7943_5472# vdd 0.0799f
C3552 a_2885_8740# a_4077_9037# 0.0192f
C3553 a_16895_5026# a_16895_7226# 0.176f
C3554 a_15203_8914# a_15732_9033# 0.143f
C3555 a_12919_2127# a_13853_3163# 0.155f
C3556 a_19163_8529# a_18910_8542# 0.125f
C3557 a_6848_7681# a_6864_7221# 0.348f
C3558 a_18959_2465# vdd 0.0325f
C3559 a_1791_8743# a_852_8433# 0.302f
C3560 a_17835_1657# a_17971_2345# 0.345f
C3561 a_1805_2649# a_1803_4861# 0.206f
C3562 a_5176_958# a_5912_753# 0.255f
C3563 a_1803_4861# a_1810_2768# 0.583f
C3564 a_7799_4035# a_7848_3845# 0.22f
C3565 d0 a_10465_5683# 0.0235f
C3566 a_18908_7067# vdd 0.311f
C3567 a_7938_7855# a_7877_7141# 0.0126f
C3568 a_12805_5083# a_12915_3407# 0.132f
C3569 a_13850_8678# a_13854_8501# 0.559f
C3570 a_2778_2701# vdd 0.0269f
C3571 a_15943_2415# a_15522_2415# 0.0104f
C3572 a_3821_4261# a_3872_3522# 0.011f
C3573 a_116_9097# vdd 0.323f
C3574 a_19163_8529# a_18955_8529# 0.448f
C3575 a_10151_1568# a_10678_1820# 0.14f
C3576 a_3826_4638# a_3871_4625# 0.151f
C3577 a_6427_6578# d1 0.0235f
C3578 a_10463_8992# a_10676_8992# 0.448f
C3579 a_5704_2410# vdd 0.0342f
C3580 a_1514_1533# d2 0.0235f
C3581 a_18021_1052# a_17831_1834# 0.251f
C3582 a_18018_7670# a_17973_7683# 0.181f
C3583 a_18956_6323# vdd 0.0325f
C3584 a_11727_2654# a_11834_4866# 0.218f
C3585 a_10150_3128# a_10887_3477# 0.112f
C3586 a_15206_2525# vdd 0.323f
C3587 a_3141_2109# a_2933_2109# 0.448f
C3588 a_18913_5787# d0 0.00533f
C3589 a_12962_6526# a_13170_6526# 0.448f
C3590 a_10151_922# a_10888_1271# 0.112f
C3591 a_13901_6836# a_14109_6836# 0.448f
C3592 a_13854_8501# a_13851_9232# 0.0292f
C3593 a_5175_3394# a_5491_3513# 0.125f
C3594 a_16601_1579# a_16892_2695# 0.0104f
C3595 a_15943_2415# a_15942_1861# 0.498f
C3596 a_13852_4266# a_13858_3540# 0.0622f
C3597 a_8926_7975# a_8875_8714# 0.011f
C3598 a_8880_6331# vdd 0.133f
C3599 a_15733_7930# a_15204_8227# 0.0185f
C3600 a_5176_1188# a_5913_1307# 0.426f
C3601 a_4077_6277# a_3820_6467# 0.0467f
C3602 a_7941_8781# a_7986_8768# 0.181f
C3603 a_12919_3230# a_13854_3717# 0.254f
C3604 a_5911_4616# a_5703_4616# 0.291f
C3605 a_6427_7681# a_6848_7681# 0.0104f
C3606 a_10465_1820# a_10150_2025# 0.0467f
C3607 a_15941_4067# a_15206_3628# 0.155f
C3608 d0 a_5174_4913# 0.00888f
C3609 a_18019_4361# a_18227_4361# 0.448f
C3610 a_2889_1019# a_3142_1006# 0.11f
C3611 a_16879_7686# vdd 0.0273f
C3612 a_19165_6877# a_18908_7067# 0.0467f
C3613 a_7943_4369# a_8882_4679# 0.278f
C3614 a_856_2369# a_119_2250# 0.426f
C3615 a_17975_2168# a_17835_1657# 0.206f
C3616 a_17972_1242# a_19167_808# 0.0192f
C3617 a_7848_3845# vdd 0.0325f
C3618 a_4077_7380# a_2882_7814# 0.0192f
C3619 a_18910_998# a_18959_808# 0.218f
C3620 a_6848_6578# a_6427_6578# 0.0104f
C3621 a_3825_7947# vdd 0.135f
C3622 a_4080_3522# a_3823_3712# 0.0467f
C3623 a_8195_6562# a_7802_6064# 0.0192f
C3624 a_11405_1027# a_10888_1271# 0.0467f
C3625 a_13855_7398# vdd 0.133f
C3626 a_7939_4546# a_8877_4302# 0.316f
C3627 a_7804_1652# a_7830_2919# 0.347f
C3628 a_17091_199# a_16895_5026# 0.0424f
C3629 a_17865_4947# a_18116_7146# 0.0192f
C3630 a_6951_194# a_6738_194# 0.448f
C3631 a_8881_6885# a_8877_7062# 0.539f
C3632 a_4079_5728# a_3871_5728# 0.448f
C3633 a_7937_8958# a_8194_8768# 0.0467f
C3634 a_15207_1422# a_15942_1861# 0.155f
C3635 a_6864_5021# a_6750_7102# 0.342f
C3636 a_6750_4902# vdd 0.0342f
C3637 a_13169_8732# a_12961_8732# 0.448f
C3638 a_11725_4866# a_11512_4866# 0.448f
C3639 a_18907_6513# a_19164_6323# 0.0467f
C3640 a_7939_5649# a_8196_5459# 0.0467f
C3641 a_11839_7185# a_11839_4985# 0.176f
C3642 a_2004_153# a_2778_4901# 0.448f
C3643 a_17970_5654# a_17829_6246# 0.133f
C3644 a_16672_5480# a_16880_5480# 0.241f
C3645 a_3142_1006# vdd 0.183f
C3646 a_11823_7645# a_11822_8748# 0.498f
C3647 a_11617_2130# vdd 0.0342f
C3648 a_12035_158# a_11839_4985# 0.0424f
C3649 a_1587_1022# a_856_712# 0.169f
C3650 a_5909_6268# a_6427_6578# 0.11f
C3651 a_11755_8156# a_11839_7185# 0.263f
C3652 a_1808_7180# vdd 0.0369f
C3653 a_14663_138# a_14876_138# 0.448f
C3654 a_17833_6069# a_17829_6246# 0.518f
C3655 a_5492_1307# d0 0.0235f
C3656 d0 a_18910_8542# 0.0138f
C3657 a_16672_5480# vdd 0.0342f
C3658 a_1586_3228# a_855_2918# 0.169f
C3659 a_10149_5980# vdd 0.135f
C3660 a_18910_3758# a_17975_3271# 0.254f
C3661 a_15206_3628# a_15522_3518# 0.0467f
C3662 a_3140_4315# d1 0.0233f
C3663 a_15734_5724# vdd 0.0342f
C3664 a_12916_1201# a_13855_1511# 0.112f
C3665 a_1803_7061# a_1793_5434# 0.206f
C3666 a_13900_9042# a_14108_9042# 0.448f
C3667 a_8878_2096# a_9135_1906# 0.0467f
C3668 a_13173_1011# a_12916_1201# 0.0467f
C3669 a_17834_3863# a_18087_3850# 0.11f
C3670 a_13851_7575# vdd 0.314f
C3671 a_3871_1865# a_4079_1865# 0.448f
C3672 a_17835_1657# a_18228_2155# 0.0192f
C3673 a_120_917# a_648_712# 0.194f
C3674 a_13853_3163# a_13903_2424# 0.011f
C3675 a_6958_4902# a_6537_4902# 0.0104f
C3676 a_16880_5480# a_16879_6583# 0.504f
C3677 a_18911_6336# vdd 0.133f
C3678 a_18087_3850# vdd 0.183f
C3679 a_10147_8643# a_10147_8873# 0.0292f
C3680 a_9134_7975# a_7942_7678# 0.0192f
C3681 a_6851_1063# a_5912_753# 0.206f
C3682 a_12821_8221# a_12807_7118# 0.19f
C3683 a_853_8987# a_1583_8743# 0.195f
C3684 a_857_1266# a_120_917# 0.112f
C3685 a_13857_1883# a_14110_1870# 0.125f
C3686 a_7830_5119# a_6859_4902# 0.409f
C3687 a_6570_1574# d2 0.0235f
C3688 a_16895_5026# a_17865_4947# 0.233f
C3689 a_2932_5418# a_2883_5608# 0.219f
C3690 a_5053_133# vdd 0.114f
C3691 a_16879_6583# vdd 0.0373f
C3692 a_7940_3443# a_7799_4035# 0.133f
C3693 a_2998_8216# a_2790_8216# 0.448f
C3694 a_18913_5787# a_18956_6323# 0.0185f
C3695 a_15941_7930# a_15204_8040# 0.277f
C3696 a_7986_8768# vdd 0.0325f
C3697 a_10885_5129# a_10149_4690# 0.155f
C3698 a_12822_6015# vdd 0.0325f
C3699 a_7940_2340# a_7944_2163# 0.518f
C3700 a_11823_6542# vdd 0.0373f
C3701 a_16600_3785# d2 0.0235f
C3702 a_10886_5683# vdd 0.455f
C3703 a_6847_8784# a_6864_7221# 0.14f
C3704 a_12916_8745# a_13900_9042# 0.292f
C3705 a_16568_7107# a_16895_5026# 0.0104f
C3706 a_9133_9078# a_8876_9268# 0.0467f
C3707 a_14110_4630# a_13902_4630# 0.448f
C3708 a_2885_8740# a_3869_9037# 0.292f
C3709 a_10885_4026# vdd 0.0799f
C3710 a_2778_2701# a_2747_3817# 0.206f
C3711 a_11756_5950# vdd 0.0342f
C3712 a_7937_8958# a_9132_8524# 0.0192f
C3713 a_10464_7889# a_10677_7889# 0.448f
C3714 a_1795_1022# vdd 0.0273f
C3715 a_6641_5475# vdd 0.0342f
C3716 a_12774_3999# a_12809_2706# 0.298f
C3717 a_5704_3513# a_5175_3394# 0.143f
C3718 a_8925_6318# a_8880_6331# 0.154f
C3719 a_7987_7665# a_7832_7154# 0.0267f
C3720 a_8875_8714# vdd 0.314f
C3721 a_10150_3587# a_10150_3358# 0.539f
C3722 a_13854_8501# vdd 0.133f
C3723 a_12913_6716# a_13170_6526# 0.0467f
C3724 a_3825_4084# vdd 0.133f
C3725 a_13851_6472# a_13855_6295# 0.559f
C3726 a_3872_3522# a_3823_3712# 0.218f
C3727 a_13900_6282# vdd 0.0325f
C3728 a_1805_2649# a_1810_2768# 0.586f
C3729 a_8195_6562# a_7987_6562# 0.448f
C3730 a_8877_4302# a_8926_4112# 0.218f
C3731 a_5911_1856# a_6850_2166# 0.302f
C3732 a_15204_7124# a_15204_6937# 0.0625f
C3733 a_2883_4505# a_3822_4815# 0.112f
C3734 a_15521_1861# a_15942_1861# 0.0104f
C3735 a_17972_1242# a_18911_1552# 0.112f
C3736 a_15520_5170# vdd 0.178f
C3737 a_7940_3443# vdd 0.439f
C3738 a_13852_7026# a_12917_6539# 0.254f
C3739 a_2748_1611# a_2744_1788# 0.518f
C3740 a_19165_5220# vdd 0.183f
C3741 a_15941_4067# a_15733_4067# 0.3f
C3742 a_2931_6521# a_2772_7290# 0.0774f
C3743 a_7938_6752# a_7942_6575# 0.518f
C3744 a_16672_4377# vdd 0.0342f
C3745 a_19165_5220# a_18912_5233# 0.125f
C3746 a_7987_7665# a_7797_8447# 0.251f
C3747 a_13850_8678# a_13856_7952# 0.0622f
C3748 a_15736_1312# a_15207_1193# 0.143f
C3749 a_15732_7376# a_15204_6937# 0.011f
C3750 a_3822_5918# a_2883_5608# 0.112f
C3751 a_10676_7335# a_10463_7335# 0.448f
C3752 a_5908_8474# a_5173_8035# 0.155f
C3753 a_16879_6583# a_16812_5991# 0.195f
C3754 a_14110_5733# d0 0.0233f
C3755 a_10149_5564# vdd 0.128f
C3756 a_3826_5741# d0 0.00533f
C3757 a_5701_6268# a_5174_5829# 0.011f
C3758 a_10149_4461# vdd 0.128f
C3759 a_10676_6232# a_10884_6232# 0.3f
C3760 a_17972_1242# vdd 0.439f
C3761 a_7830_5119# a_7834_4942# 0.518f
C3762 a_18116_7146# a_17863_7159# 0.11f
C3763 a_852_8433# vdd 0.0799f
C3764 a_12914_4510# a_13852_4266# 0.316f
C3765 a_2888_3225# a_2933_3212# 0.181f
C3766 a_8057_1639# a_7804_1652# 0.11f
C3767 vdd a_5490_1856# 0.178f
C3768 a_2881_8917# a_3138_8727# 0.0467f
C3769 a_7828_7331# a_7942_6575# 0.0437f
C3770 a_10886_5683# a_10465_5683# 0.0104f
C3771 a_13853_3163# vdd 0.314f
C3772 a_3031_4888# a_2004_153# 0.0192f
C3773 a_3821_5364# vdd 0.314f
C3774 a_3872_762# a_3827_775# 0.154f
C3775 a_8881_6885# vdd 0.145f
C3776 a_4080_3522# a_3872_3522# 0.448f
C3777 a_12821_8221# a_12776_8234# 0.157f
C3778 a_4078_5174# vdd 0.183f
C3779 a_19164_9083# vdd 0.183f
C3780 a_15206_3399# a_15943_3518# 0.426f
C3781 a_18225_8773# a_18017_8773# 0.448f
C3782 a_12920_1024# a_12916_1201# 0.518f
C3783 a_1808_4980# a_1902_4861# 0.214f
C3784 a_11841_2773# vdd 0.038f
C3785 a_10151_1381# a_10151_1568# 0.0622f
C3786 a_12918_5436# a_12914_5613# 0.518f
C3787 a_7877_7141# vdd 0.0325f
C3788 a_18957_5220# a_18913_4684# 0.0185f
C3789 a_17877_8262# a_18085_8262# 0.448f
C3790 a_1803_7061# a_1584_6537# 0.0267f
C3791 a_3821_7021# a_3824_6290# 0.0292f
C3792 a_4077_6277# a_2882_6711# 0.0192f
C3793 a_8877_5405# vdd 0.314f
C3794 a_3823_3712# a_2884_3402# 0.112f
C3795 a_13856_7952# a_14109_7939# 0.11f
C3796 a_12854_4893# a_13062_4893# 0.448f
C3797 a_15205_6021# vdd 0.135f
C3798 a_8879_8537# d0 0.0138f
C3799 a_10887_3477# a_10150_3358# 0.426f
C3800 a_1483_2649# vdd 0.178f
C3801 a_10148_8186# a_10677_7889# 0.0185f
C3802 a_1791_8743# a_1792_7640# 0.498f
C3803 a_6951_194# a_5178_859# 0.0111f
C3804 a_13857_2986# vdd 0.133f
C3805 a_1795_1022# a_856_712# 0.206f
C3806 a_10148_6667# a_10677_6786# 0.143f
C3807 a_12134_158# a_14663_138# 0.0467f
C3808 a_119_3582# a_119_3769# 0.0622f
C3809 a_18227_5464# a_18019_5464# 0.448f
C3810 a_13900_7385# a_13855_7398# 0.154f
C3811 a_3820_9227# vdd 0.311f
C3812 a_10466_717# a_10151_922# 0.0467f
C3813 a_15939_8479# a_15940_9033# 0.498f
C3814 a_13852_4266# a_13856_4089# 0.559f
C3815 a_854_7884# a_853_7330# 0.498f
C3816 a_2791_6010# vdd 0.0325f
C3817 a_16879_6583# a_16458_6583# 0.0104f
C3818 d0 a_15522_3518# 0.0235f
C3819 a_15204_6937# vdd 0.323f
C3820 a_12914_5613# a_13853_5923# 0.112f
C3821 a_12805_2883# a_12779_1616# 0.347f
C3822 a_18913_4684# a_18908_5410# 0.0625f
C3823 a_5173_7119# a_5909_7371# 0.279f
C3824 a_854_7884# a_117_7535# 0.112f
C3825 a_7943_4369# a_8878_4856# 0.254f
C3826 a_2884_2299# a_2888_2122# 0.518f
C3827 a_2933_2109# vdd 0.0325f
C3828 a_13903_767# a_13858_780# 0.154f
C3829 a_17976_1065# a_18909_2101# 0.155f
C3830 a_7804_1652# a_8197_2150# 0.0192f
C3831 a_4077_9037# d0 0.0233f
C3832 a_12912_8922# a_12776_8234# 0.345f
C3833 a_11725_4866# a_11834_4866# 0.117f
C3834 a_10465_5683# a_10149_5564# 0.125f
C3835 a_5702_5165# vdd 0.0342f
C3836 a_3029_7100# a_2821_7100# 0.448f
C3837 a_11836_2654# a_11825_2130# 0.328f
C3838 a_17970_5654# vdd 0.439f
C3839 a_16673_2171# vdd 0.0342f
C3840 a_10677_5129# a_10885_5129# 0.3f
C3841 a_2934_1006# a_3142_1006# 0.448f
C3842 a_6640_7681# vdd 0.0342f
C3843 a_17970_5654# a_18912_5233# 0.426f
C3844 a_10464_6786# d0 0.0235f
C3845 a_19166_4671# d0 0.0233f
C3846 a_8881_5228# d0 0.0138f
C3847 d0 a_3827_2432# 0.00533f
C3848 a_18910_998# a_17972_1242# 0.316f
C3849 a_10462_8438# vdd 0.178f
C3850 a_17833_6069# vdd 0.0273f
C3851 a_6782_3780# vdd 0.0342f
C3852 a_17969_7860# a_18908_8170# 0.112f
C3853 a_18909_3204# a_18913_3027# 0.559f
C3854 a_15206_3815# a_15205_4272# 0.519f
C3855 a_118_5975# a_118_5788# 0.0622f
C3856 a_5175_2520# a_5703_2959# 0.011f
C3857 a_10150_3358# a_10466_3477# 0.125f
C3858 a_10678_4580# a_10149_4690# 0.194f
C3859 a_6429_2166# vdd 0.178f
C3860 a_5909_6268# a_5174_5829# 0.155f
C3861 a_13901_7939# a_12917_7642# 0.292f
C3862 a_15204_6708# a_15204_6937# 0.539f
C3863 a_117_7994# a_433_7884# 0.0467f
C3864 a_5176_1604# vdd 0.135f
C3865 a_10679_3477# a_10150_3358# 0.143f
C3866 a_8882_4679# d0 0.00533f
C3867 a_13851_7575# a_13900_7385# 0.218f
C3868 a_434_1815# a_120_1563# 0.11f
C3869 a_15204_6478# a_15732_6273# 0.194f
C3870 a_3827_3535# vdd 0.135f
C3871 a_1372_4331# d1 0.0235f
C3872 a_119_3582# a_119_3353# 0.539f
C3873 a_10465_2923# a_10150_2671# 0.11f
C3874 a_13857_4643# a_13901_5179# 0.0185f
C3875 a_15522_758# vdd 0.178f
C3876 a_120_1376# a_857_1266# 0.277f
C3877 a_8884_1370# a_8929_1357# 0.151f
C3878 a_5910_5165# a_6428_5475# 0.11f
C3879 a_11822_8748# a_11839_7185# 0.14f
C3880 a_15939_8479# a_15731_8479# 0.3f
C3881 a_2886_6534# a_4078_6831# 0.0192f
C3882 vdd a_12823_3809# 0.0325f
C3883 a_11713_158# a_12134_158# 0.0104f
C3884 a_13853_2060# a_12920_1024# 0.155f
C3885 a_1795_1022# a_1514_1533# 0.11f
C3886 a_3872_762# vdd 0.0325f
C3887 a_9134_4112# a_8877_4302# 0.0467f
C3888 a_8878_2096# a_8929_1357# 0.011f
C3889 d0 a_13857_5746# 0.00533f
C3890 a_13852_4266# a_12919_3230# 0.155f
C3891 a_13856_7952# vdd 0.135f
C3892 a_15203_9143# vdd 0.323f
C3893 a_856_2369# a_1805_2649# 0.276f
C3894 a_11618_1027# a_11405_1027# 0.448f
C3895 a_11514_2654# a_11836_2654# 0.11f
C3896 a_10883_8438# a_11822_8748# 0.302f
C3897 a_2741_8406# vdd 0.0316f
C3898 a_8927_3009# a_7940_3443# 0.283f
C3899 a_119_3582# a_435_3472# 0.0467f
C3900 a_17878_6056# a_18086_6056# 0.448f
C3901 a_15522_758# a_15943_758# 0.0104f
C3902 a_11404_3233# vdd 0.178f
C3903 a_435_2369# a_119_2250# 0.125f
C3904 a_11824_5439# a_11543_5950# 0.11f
C3905 a_16781_7107# vdd 0.0342f
C3906 a_18229_1052# a_17831_1834# 0.0192f
C3907 a_6782_3780# a_6569_3780# 0.448f
C3908 a_11757_3744# a_11841_2773# 0.263f
C3909 a_854_5124# a_1793_5434# 0.206f
C3910 a_14110_2973# d0 0.0233f
C3911 a_10148_7083# a_10463_7335# 0.11f
C3912 a_4078_4071# d0 0.0233f
C3913 a_1803_7061# a_854_6781# 0.28f
C3914 a_7834_2742# a_7799_4035# 0.298f
C3915 a_18226_7670# a_17828_8452# 0.0192f
C3916 a_12803_7295# a_12777_6028# 0.347f
C3917 a_117_6891# a_433_6781# 0.0467f
C3918 a_8878_3199# vdd 0.314f
C3919 a_14108_6282# a_13851_6472# 0.0467f
C3920 a_6848_7681# a_5909_7371# 0.206f
C3921 a_15205_4502# vdd 0.128f
C3922 a_13902_5733# a_13851_6472# 0.011f
C3923 a_7989_3253# a_7940_3443# 0.219f
C3924 a_116_8868# a_116_8638# 0.0292f
C3925 a_1512_5945# a_1725_5945# 0.448f
C3926 a_431_8433# a_644_8433# 0.448f
C3927 a_1586_3228# vdd 0.0342f
C3928 a_16461_1068# vdd 0.178f
C3929 a_18914_2478# vdd 0.145f
C3930 a_7942_6575# a_9134_6872# 0.0192f
C3931 a_11402_7645# a_11823_7645# 0.0104f
C3932 a_13857_4643# vdd 0.146f
C3933 a_15940_7376# a_15941_7930# 0.498f
C3934 a_12918_5436# a_13853_5923# 0.254f
C3935 a_9136_2460# a_8883_2473# 0.11f
C3936 a_7939_5649# vdd 0.439f
C3937 a_13173_1011# d1 0.0233f
C3938 a_10151_1568# a_10150_2025# 0.519f
C3939 a_13029_8221# d2 0.0233f
C3940 a_15523_1312# vdd 0.178f
C3941 a_6539_2690# vdd 0.178f
C3942 a_7939_4546# a_8881_4125# 0.426f
C3943 a_14109_6836# vdd 0.183f
C3944 a_5702_5165# a_5174_4913# 0.14f
C3945 a_2746_6023# a_2999_6010# 0.11f
C3946 a_7987_6562# a_7802_6064# 0.231f
C3947 a_1808_4980# a_1481_7061# 0.0104f
C3948 a_12779_1616# a_13172_2114# 0.0192f
C3949 a_3029_7100# a_2778_4901# 0.0192f
C3950 a_16671_6583# a_15940_6273# 0.169f
C3951 a_15943_2415# vdd 0.454f
C3952 a_17861_5124# a_18118_2734# 0.0192f
C3953 a_2778_2701# a_2774_2878# 0.484f
C3954 a_13853_3163# a_13902_2973# 0.218f
C3955 a_5488_7371# a_5909_7371# 0.0104f
C3956 a_16461_1068# a_15943_758# 0.11f
C3957 a_7834_2742# vdd 0.0269f
C3958 a_12807_7118# a_12772_8411# 0.298f
C3959 a_5487_8474# a_5908_8474# 0.0104f
C3960 a_2823_2688# a_2778_2701# 0.128f
C3961 a_5489_7925# a_5910_7925# 0.0104f
C3962 a_15205_5375# a_15941_5170# 0.255f
C3963 a_13060_7105# a_12852_7105# 0.448f
C3964 a_13859_1334# vdd 0.135f
C3965 a_6859_7102# a_6781_5986# 0.198f
C3966 vout vdd 0.0176f
C3967 d2 a_16599_5991# 0.0235f
C3968 a_17968_8963# a_17832_8275# 0.345f
C3969 a_12774_3999# a_13172_3217# 0.0192f
C3970 a_17830_4040# a_18087_3850# 0.0467f
C3971 d0 a_5491_2410# 0.0235f
C3972 a_5701_9028# a_5172_8909# 0.143f
C3973 a_16881_2171# a_16601_1579# 0.0467f
C3974 a_18226_6567# vdd 0.183f
C3975 a_5174_4726# a_5703_4616# 0.194f
C3976 a_12035_158# a_11713_158# 0.11f
C3977 a_17865_4947# a_17829_6246# 0.181f
C3978 a_10883_8438# a_10148_8186# 0.279f
C3979 a_5175_2520# a_5911_2959# 0.155f
C3980 a_15207_1422# vdd 0.323f
C3981 a_11403_5439# a_10885_5129# 0.11f
C3982 a_16674_1068# vdd 0.0342f
C3983 a_17974_4374# a_18909_4861# 0.254f
C3984 a_5910_6822# vdd 0.454f
C3985 a_13857_2986# a_13902_2973# 0.154f
C3986 a_13173_1011# a_12965_1011# 0.448f
C3987 a_4080_2419# d0 0.0233f
C3988 a_11755_8156# a_11822_8748# 0.195f
C3989 a_15205_4731# a_15205_4502# 0.539f
C3990 a_15206_3628# a_15206_3399# 0.539f
C3991 a_6642_2166# a_5912_2410# 0.195f
C3992 a_10149_4877# vdd 0.144f
C3993 a_1792_7640# vdd 0.0273f
C3994 a_1794_2125# a_1727_1533# 0.195f
C3995 a_6642_2166# a_6861_2690# 0.0267f
C3996 a_17091_199# a_16982_199# 0.117f
C3997 a_12809_4906# vdd 0.0264f
C3998 a_16890_4907# a_15942_4621# 0.0518f
C3999 a_5488_6268# d0 0.0235f
C4000 a_119_2666# a_119_2479# 0.0625f
C4001 a_15941_4067# a_16672_4377# 0.169f
C4002 a_17880_1644# vdd 0.0325f
C4003 a_5173_6703# d0 0.0138f
C4004 a_8879_8537# a_8875_8714# 0.559f
C4005 a_118_4456# d0 0.0138f
C4006 a_10463_8992# a_10884_8992# 0.0104f
C4007 a_1724_8151# a_1511_8151# 0.448f
C4008 a_10677_5129# a_10464_5129# 0.448f
C4009 a_16674_1068# a_15943_758# 0.169f
C4010 a_10676_7335# a_10148_6896# 0.011f
C4011 a_7943_4369# a_7803_3858# 0.206f
C4012 a_13904_1321# vdd 0.0325f
C4013 a_9135_4666# vdd 0.183f
C4014 a_18956_9083# a_17972_8786# 0.292f
C4015 a_5175_2061# a_5911_1856# 0.255f
C4016 a_16897_2814# a_15942_2964# 0.0355f
C4017 a_16895_5026# a_15941_6827# 0.132f
C4018 a_433_4021# a_118_4226# 0.0467f
C4019 a_8883_3576# a_8879_3753# 0.539f
C4020 a_2742_6200# a_2772_7290# 0.14f
C4021 a_6568_5986# a_6781_5986# 0.448f
C4022 a_853_8987# a_1791_8743# 0.133f
C4023 a_8929_1357# a_8880_1547# 0.218f
C4024 a_11834_7066# a_11839_7185# 0.464f
C4025 a_15940_9033# a_16670_8789# 0.195f
C4026 a_8196_4356# d1 0.0233f
C4027 a_13852_5369# a_13902_4630# 0.011f
C4028 a_647_2918# a_119_2479# 0.011f
C4029 a_6783_1574# a_6861_2690# 0.198f
C4030 a_3822_5918# a_3825_5187# 0.0292f
C4031 a_7989_2150# vdd 0.0325f
C4032 a_8881_4125# a_8926_4112# 0.154f
C4033 a_10885_4026# a_10886_4580# 0.498f
C4034 a_18909_3204# a_19166_3014# 0.0467f
C4035 a_5172_8679# vdd 0.312f
C4036 a_7987_7665# a_7942_7678# 0.181f
C4037 a_16989_4907# a_15942_4621# 0.0863f
C4038 a_17970_4551# a_17974_4374# 0.518f
C4039 a_13902_1870# vdd 0.0325f
C4040 a_14109_5179# d0 0.0233f
C4041 a_5175_2520# vdd 0.323f
C4042 a_10147_8873# vdd 0.128f
C4043 a_13853_4820# vdd 0.311f
C4044 a_10148_6437# a_10885_6786# 0.112f
C4045 a_7879_4929# a_7939_5649# 0.0121f
C4046 a_16895_7226# vdd 0.0369f
C4047 a_8056_3845# a_7803_3858# 0.11f
C4048 a_1808_4980# a_2778_4901# 0.233f
C4049 a_10885_7889# vdd 0.455f
C4050 a_12772_8411# a_12776_8234# 0.524f
C4051 a_5704_2410# a_5491_2410# 0.448f
C4052 a_119_2250# a_648_2369# 0.143f
C4053 a_18959_3568# a_18910_3758# 0.218f
C4054 a_3871_2968# a_2884_3402# 0.283f
C4055 a_10150_2671# vdd 0.143f
C4056 a_116_8868# d0 0.0138f
C4057 a_8878_3199# a_8927_3009# 0.218f
C4058 a_13171_4320# a_12963_4320# 0.448f
C4059 a_13854_2614# a_14111_2424# 0.0467f
C4060 a_117_6891# a_117_6662# 0.539f
C4061 a_16671_6583# a_15941_6827# 0.195f
C4062 a_17969_6757# vdd 0.439f
C4063 a_15206_3815# a_15206_3628# 0.0622f
C4064 a_11402_7645# a_11615_7645# 0.448f
C4065 a_3823_2609# a_3826_1878# 0.0292f
C4066 a_15521_1861# vdd 0.178f
C4067 a_12919_2127# a_13854_2614# 0.254f
C4068 a_10678_2923# a_10150_2671# 0.14f
C4069 a_18957_6877# a_18912_6890# 0.151f
C4070 a_119_2250# d0 0.0138f
C4071 a_2743_3994# a_2888_3225# 0.326f
C4072 d5 vdd 0.178f
C4073 a_15206_3169# a_15206_3399# 0.0292f
C4074 a_10149_4461# a_10886_4580# 0.426f
C4075 a_15207_963# a_15207_1193# 0.0292f
C4076 a_5911_4616# a_5910_4062# 0.498f
C4077 a_19164_6323# d0 0.0233f
C4078 a_5705_1307# a_5176_1604# 0.0185f
C4079 a_6639_8784# a_5908_8474# 0.169f
C4080 a_8926_6872# a_7942_6575# 0.292f
C4081 a_14111_3527# a_13854_3717# 0.0467f
C4082 a_11727_2654# vdd 0.0342f
C4083 a_8926_5215# a_9134_5215# 0.448f
C4084 a_5912_2410# a_6861_2690# 0.276f
C4085 d6 a_14663_138# 0.0235f
C4086 a_13900_6282# a_13857_5746# 0.0185f
C4087 a_18227_5464# a_17974_5477# 0.11f
C4088 a_13171_5423# d1 0.0233f
C4089 a_10150_2255# vdd 0.128f
C4090 a_12807_7118# a_12803_7295# 0.606f
C4091 a_12805_5083# a_13062_2693# 0.0192f
C4092 a_118_4872# a_646_5124# 0.14f
C4093 a_1371_6537# a_1584_6537# 0.448f
C4094 a_11404_2130# vdd 0.178f
C4095 a_12920_1024# a_12965_1011# 0.181f
C4096 a_3000_3804# d2 0.0233f
C4097 a_646_5124# a_433_5124# 0.448f
C4098 a_8883_816# a_8880_1547# 0.0292f
C4099 a_15206_2525# a_15735_2415# 0.194f
C4100 a_13851_7575# a_12917_6539# 0.155f
C4101 a_14107_8488# d0 0.0233f
C4102 a_17832_8275# a_17863_7159# 0.206f
C4103 a_18957_4117# a_17970_4551# 0.283f
C4104 a_18906_8719# a_17968_8963# 0.316f
C4105 vdd a_15735_3518# 0.0342f
C4106 a_17091_199# vdd 0.0211f
C4107 a_18906_8719# a_18912_7993# 0.0622f
C4108 a_10148_7999# a_10885_7889# 0.277f
C4109 a_854_5124# a_118_4685# 0.155f
C4110 a_15941_5170# a_15205_4918# 0.279f
C4111 a_7938_7855# a_7832_7154# 0.423f
C4112 a_2821_7100# a_2778_4901# 0.208f
C4113 a_15943_2415# a_16783_2695# 0.0126f
C4114 a_1586_3228# a_1373_3228# 0.448f
C4115 a_4078_4071# a_3825_4084# 0.125f
C4116 a_16811_8197# vdd 0.0342f
C4117 a_15939_8479# a_16670_8789# 0.169f
C4118 a_17835_1657# a_17831_1834# 0.518f
C4119 a_8878_5959# a_7943_5472# 0.254f
C4120 a_10148_7540# a_10463_7335# 0.0467f
C4121 a_5701_9028# a_5488_9028# 0.448f
C4122 a_853_6227# a_1584_6537# 0.169f
C4123 a_12778_3822# vdd 0.0273f
C4124 a_15207_1609# a_15206_2066# 0.519f
C4125 a_15207_1193# d0 0.0138f
C4126 a_15940_7376# a_16879_7686# 0.206f
C4127 a_7830_2919# a_8087_2729# 0.0467f
C4128 a_8877_5405# a_8881_5228# 0.559f
C4129 a_7834_2742# a_7989_3253# 0.0267f
C4130 a_11834_7066# a_11839_4985# 0.594f
C4131 a_6426_8784# vdd 0.178f
C4132 a_4077_9037# a_3820_9227# 0.0467f
C4133 a_4081_1316# a_3828_1329# 0.11f
C4134 a_1370_8743# d1 0.0235f
C4135 a_8877_8165# a_8881_7988# 0.539f
C4136 a_10463_6232# vdd 0.178f
C4137 a_7944_3266# a_8197_3253# 0.11f
C4138 a_5909_7371# a_5701_7371# 0.3f
C4139 a_17828_8452# a_17832_8275# 0.524f
C4140 a_6849_5475# a_6859_7102# 0.206f
C4141 a_17091_199# a_14985_138# 0.294f
C4142 a_15206_3399# d0 0.0138f
C4143 a_116_8868# a_116_9097# 0.539f
C4144 a_13858_3540# a_12919_3230# 0.278f
C4145 a_8882_4679# a_8877_5405# 0.0625f
C4146 a_7938_7855# a_7797_8447# 0.133f
C4147 a_11616_5439# a_10885_5129# 0.169f
C4148 a_2741_8406# a_2790_8216# 0.22f
C4149 a_7830_5119# a_7830_2919# 0.176f
C4150 a_5912_2410# a_6752_2690# 0.0126f
C4151 a_8196_4356# a_7803_3858# 0.0192f
C4152 a_6861_2690# a_6752_2690# 0.117f
C4153 d0 a_10150_3358# 0.0138f
C4154 a_18907_7616# a_19164_7426# 0.0467f
C4155 a_19165_4117# a_18912_4130# 0.125f
C4156 a_2998_8216# a_2776_7113# 0.0192f
C4157 a_434_1815# d0 0.0235f
C4158 a_17968_8963# vdd 0.439f
C4159 a_5053_133# a_7060_194# 0.0224f
C4160 a_1805_2649# a_1586_2125# 0.0267f
C4161 a_17865_4947# vdd 0.0264f
C4162 a_11725_4866# a_11933_4866# 0.337f
C4163 a_10148_7083# a_10148_6896# 0.0625f
C4164 a_18912_7993# vdd 0.135f
C4165 a_3828_1329# a_3871_1865# 0.0185f
C4166 a_433_6781# d0 0.0235f
C4167 a_3139_6521# vdd 0.183f
C4168 a_13853_3163# a_14110_2973# 0.0467f
C4169 a_18021_1052# a_17976_1065# 0.181f
C4170 a_3827_775# a_2885_1196# 0.426f
C4171 a_19164_6323# a_18956_6323# 0.448f
C4172 a_10887_3477# a_10150_3587# 0.277f
C4173 a_1512_5945# a_1792_6537# 0.0467f
C4174 a_3871_1865# a_2884_2299# 0.283f
C4175 a_2887_4328# a_3871_4625# 0.292f
C4176 a_8882_3022# vdd 0.133f
C4177 a_13854_2614# a_13903_2424# 0.218f
C4178 a_18909_4861# vdd 0.311f
C4179 a_14109_4076# d0 0.0233f
C4180 a_18956_7426# a_18912_6890# 0.0185f
C4181 a_16568_7107# vdd 0.178f
C4182 a_18959_2465# a_18909_3204# 0.011f
C4183 a_17973_6580# vdd 0.0951f
C4184 a_9134_4112# a_8881_4125# 0.125f
C4185 a_13851_9232# a_14108_9042# 0.0467f
C4186 a_13899_8488# a_13854_8501# 0.154f
C4187 a_3872_2419# vdd 0.0325f
C4188 a_10883_8438# a_10884_8992# 0.498f
C4189 a_11617_2130# a_11836_2654# 0.0267f
C4190 a_1584_7640# a_853_7330# 0.169f
C4191 a_15204_8227# vdd 0.135f
C4192 a_4079_5728# d0 0.0233f
C4193 a_644_8433# a_116_8638# 0.194f
C4194 a_8876_7611# a_8925_7421# 0.218f
C4195 a_17974_5477# a_19166_5774# 0.0192f
C4196 a_14108_7385# d0 0.0233f
C4197 a_6849_5475# a_6568_5986# 0.11f
C4198 a_10150_2484# a_10150_2671# 0.0625f
C4199 a_3821_4261# a_2883_4505# 0.316f
C4200 a_7938_6752# a_7828_7331# 0.285f
C4201 a_18909_2101# vdd 0.314f
C4202 a_15206_3815# a_15733_4067# 0.14f
C4203 a_7988_4356# a_7939_4546# 0.243f
C4204 a_4079_1865# a_3826_1878# 0.125f
C4205 a_12914_5613# a_12773_6205# 0.133f
C4206 a_13857_2986# a_14110_2973# 0.125f
C4207 a_12805_2883# a_12775_1793# 0.14f
C4208 a_119_3123# a_119_3353# 0.0292f
C4209 a_853_8987# vdd 0.454f
C4210 a_18958_1911# vdd 0.0325f
C4211 a_1371_6537# a_854_6781# 0.0467f
C4212 a_14110_4630# vdd 0.183f
C4213 d0 a_9133_7421# 0.0233f
C4214 a_12916_8745# a_13851_9232# 0.254f
C4215 a_17973_6580# a_19165_6877# 0.0192f
C4216 a_10150_3587# a_10466_3477# 0.0467f
C4217 a_17970_4551# a_17834_3863# 0.345f
C4218 a_646_7884# vdd 0.0342f
C4219 a_15206_3815# d0 0.00888f
C4220 a_7940_2340# vdd 0.439f
C4221 a_8196_5459# a_7798_6241# 0.0192f
C4222 a_10150_3587# a_10679_3477# 0.194f
C4223 a_3001_1598# a_2748_1611# 0.11f
C4224 a_17865_2747# a_18020_3258# 0.0267f
C4225 a_434_2918# d0 0.0235f
C4226 a_13852_5369# a_13856_5192# 0.559f
C4227 a_5175_3623# a_5491_3513# 0.0467f
C4228 a_117_6432# a_854_6781# 0.112f
C4229 a_10150_2484# a_10150_2255# 0.539f
C4230 a_17970_4551# vdd 0.439f
C4231 a_11615_6542# a_11834_7066# 0.0267f
C4232 a_5173_7119# a_5702_6822# 0.0185f
C4233 a_16879_6583# a_16599_5991# 0.0467f
C4234 a_8928_3563# a_7944_3266# 0.292f
C4235 a_18909_2101# a_18915_1375# 0.0622f
C4236 a_18909_5964# a_17974_5477# 0.254f
C4237 a_9888_17# a_5053_133# 0.569f
C4238 a_2889_1019# a_2885_1196# 0.518f
C4239 a_4079_4625# a_3822_4815# 0.0467f
C4240 a_9136_3563# a_8883_3576# 0.11f
C4241 a_853_6227# a_854_6781# 0.498f
C4242 a_8881_7988# d0 0.00533f
C4243 a_10885_5129# a_10149_5334# 0.255f
C4244 a_12914_4510# a_13856_4089# 0.426f
C4245 a_2776_7113# a_2772_7290# 0.606f
C4246 a_16878_8789# a_16879_7686# 0.498f
C4247 a_12915_3407# a_12964_3217# 0.219f
C4248 d3 a_3031_2688# 0.0233f
C4249 a_118_4872# a_433_5124# 0.11f
C4250 a_13854_957# a_14111_767# 0.0467f
C4251 a_15521_4621# a_15942_4621# 0.0104f
C4252 a_18958_1911# a_18915_1375# 0.0185f
C4253 a_18911_6336# a_19164_6323# 0.125f
C4254 a_5910_7925# vdd 0.455f
C4255 a_2792_3804# a_2743_3994# 0.22f
C4256 a_2888_3225# vdd 0.0799f
C4257 d0 a_3824_6290# 0.0138f
C4258 a_10886_2923# a_10465_2923# 0.0104f
C4259 a_8927_1906# a_7940_2340# 0.283f
C4260 a_2778_2701# a_3000_3804# 0.0192f
C4261 a_1694_7061# a_1808_7180# 0.178f
C4262 a_3142_1006# d1 0.0233f
C4263 a_15519_6273# vdd 0.178f
C4264 a_8926_6872# a_8876_7611# 0.011f
C4265 a_12803_7295# a_12962_6526# 0.0774f
C4266 a_10150_2025# a_10887_2374# 0.112f
C4267 a_7939_5649# a_8881_5228# 0.426f
C4268 a_2885_1196# vdd 0.439f
C4269 a_15204_7581# a_15941_7930# 0.112f
C4270 a_9133_9078# a_8880_9091# 0.11f
C4271 a_10887_3477# a_11825_3233# 0.322f
C4272 a_10148_6896# a_10677_6786# 0.194f
C4273 a_1512_5945# d2 0.0235f
C4274 a_119_3582# vdd 0.323f
C4275 a_854_4021# a_1372_4331# 0.11f
C4276 a_1793_4331# a_1585_4331# 0.26f
C4277 a_11824_5439# a_11403_5439# 0.0104f
C4278 a_3869_9037# a_3820_9227# 0.218f
C4279 a_10884_6232# a_10149_5980# 0.279f
C4280 a_13854_2614# vdd 0.311f
C4281 a_6864_7221# vdd 0.0369f
C4282 a_5913_1307# vdd 0.455f
C4283 a_647_1815# vdd 0.0342f
C4284 a_3821_4261# a_3870_4071# 0.218f
C4285 a_117_7765# vdd 0.128f
C4286 a_1481_4861# a_1902_4861# 0.0104f
C4287 a_8879_993# a_9136_803# 0.0467f
C4288 a_10148_6437# vdd 0.312f
C4289 a_13857_4643# a_12918_4333# 0.278f
C4290 a_10465_1820# vdd 0.178f
C4291 a_16879_6583# a_16890_7107# 0.328f
C4292 a_5703_1856# a_5176_1417# 0.011f
C4293 a_12914_5613# a_13171_5423# 0.0467f
C4294 a_18018_6567# vdd 0.0325f
C4295 a_17863_7159# vdd 0.0269f
C4296 a_14108_9042# vdd 0.183f
C4297 a_15206_3169# a_15206_2712# 0.519f
C4298 a_3029_7100# d3 0.0233f
C4299 a_16671_7686# vdd 0.0342f
C4300 a_16673_2171# a_16460_2171# 0.448f
C4301 a_12913_6716# a_13855_6295# 0.426f
C4302 a_10887_3477# a_10466_3477# 0.0104f
C4303 a_4632_133# a_5053_133# 0.0104f
C4304 a_1587_1022# a_1374_1022# 0.448f
C4305 a_2774_5078# a_2743_3994# 0.198f
C4306 a_10887_3477# a_10679_3477# 0.291f
C4307 a_10884_6232# a_11823_6542# 0.302f
C4308 a_3823_952# a_3827_775# 0.559f
C4309 a_3821_8124# vdd 0.311f
C4310 a_18020_2155# a_17971_2345# 0.243f
C4311 a_12918_5436# a_12773_6205# 0.326f
C4312 a_17968_8963# a_18910_8542# 0.426f
C4313 a_14108_7385# a_13855_7398# 0.125f
C4314 a_13854_8501# a_14107_8488# 0.125f
C4315 a_11725_4866# vdd 0.0342f
C4316 a_12809_2706# a_13031_3809# 0.0192f
C4317 a_6427_7681# vdd 0.178f
C4318 a_645_6227# a_118_5788# 0.011f
C4319 a_3821_7021# a_3870_6831# 0.218f
C4320 a_11841_2773# a_11836_2654# 0.586f
C4321 a_7832_7154# vdd 0.0269f
C4322 a_7937_8958# a_8876_9268# 0.112f
C4323 a_2791_6010# a_2742_6200# 0.22f
C4324 a_857_1266# a_436_1266# 0.0104f
C4325 a_9132_8524# a_8924_8524# 0.448f
C4326 a_117_6662# d0 0.0138f
C4327 a_435_2369# a_856_2369# 0.0104f
C4328 a_646_4021# a_119_3769# 0.14f
C4329 a_8882_3022# a_8927_3009# 0.154f
C4330 a_9136_3563# a_8879_3753# 0.0467f
C4331 a_17828_8452# vdd 0.0316f
C4332 a_856_2369# a_1586_2125# 0.195f
C4333 a_19167_2465# vdd 0.183f
C4334 a_15940_7376# a_15204_6937# 0.155f
C4335 a_12916_8745# vdd 0.021f
C4336 a_18088_1644# vdd 0.183f
C4337 a_18955_8529# a_17968_8963# 0.283f
C4338 a_5704_3513# a_5175_3623# 0.194f
C4339 a_16890_4907# a_16895_5026# 0.498f
C4340 a_2745_8229# vdd 0.0273f
C4341 a_18955_8529# a_18912_7993# 0.0185f
C4342 a_10151_1568# a_10680_1271# 0.0185f
C4343 a_3868_8483# vdd 0.0325f
C4344 a_8194_8768# a_7941_8781# 0.11f
C4345 a_17974_4374# a_18908_5410# 0.155f
C4346 a_13851_6472# vdd 0.314f
C4347 a_13899_8488# a_13856_7952# 0.0185f
C4348 d0 a_18912_6890# 0.00533f
C4349 a_10676_7335# vdd 0.0342f
C4350 a_6641_5475# a_6428_5475# 0.448f
C4351 a_1792_6537# a_1725_5945# 0.195f
C4352 a_18227_5464# a_17829_6246# 0.0192f
C4353 a_10149_5793# a_10678_5683# 0.194f
C4354 a_15940_9033# a_15519_9033# 0.0104f
C4355 a_1895_153# a_122_818# 0.0111f
C4356 a_7797_8447# vdd 0.0316f
C4357 a_10679_3477# a_10466_3477# 0.448f
C4358 a_8927_5769# a_7943_5472# 0.292f
C4359 a_3031_4888# a_2778_4901# 0.11f
C4360 a_13851_7575# a_14108_7385# 0.0467f
C4361 a_6951_194# vdd 0.0342f
C4362 a_3822_4815# vdd 0.311f
C4363 a_119_3123# a_855_2918# 0.255f
C4364 a_10885_6786# a_10677_6786# 0.291f
C4365 a_15206_2712# d0 0.00888f
C4366 a_17975_2168# a_18020_2155# 0.181f
C4367 a_12854_4893# a_12035_158# 0.282f
C4368 a_645_6227# a_118_5975# 0.14f
C4369 a_16989_4907# a_16895_5026# 0.214f
C4370 a_5489_6822# vdd 0.178f
C4371 a_9135_4666# a_8882_4679# 0.11f
C4372 a_7803_3858# a_7848_3845# 0.157f
C4373 a_15206_2296# d0 0.0138f
C4374 a_18958_4671# a_18913_4684# 0.151f
C4375 a_5702_4062# a_5910_4062# 0.3f
C4376 a_12917_6539# a_14109_6836# 0.0192f
C4377 a_10679_2374# vdd 0.0342f
C4378 a_7940_3443# a_7879_2729# 0.0126f
C4379 a_9137_1357# a_8929_1357# 0.448f
C4380 a_10676_8992# a_10884_8992# 0.291f
C4381 a_15940_6273# vdd 0.0799f
C4382 a_8195_7665# a_7797_8447# 0.0192f
C4383 a_1808_4980# a_1481_4861# 0.0467f
C4384 a_3820_6467# vdd 0.314f
C4385 a_3868_8483# a_4076_8483# 0.448f
C4386 a_15205_5375# a_15733_5170# 0.194f
C4387 a_122_818# a_2103_153# 0.53f
C4388 a_12803_7295# a_12913_6716# 0.285f
C4389 a_19167_3568# vdd 0.183f
C4390 a_1726_3739# vdd 0.0342f
C4391 a_11512_4866# a_11839_4985# 0.0467f
C4392 a_11826_1027# vdd 0.0273f
C4393 a_17971_3448# a_18958_3014# 0.283f
C4394 a_18914_3581# d0 0.00533f
C4395 a_1803_7061# a_1808_4980# 0.594f
C4396 a_13062_4893# vdd 0.183f
C4397 a_18906_8719# a_18957_7980# 0.011f
C4398 a_5175_3810# a_5910_4062# 0.279f
C4399 a_18956_7426# a_18911_7439# 0.154f
C4400 a_18118_4934# a_17910_4934# 0.448f
C4401 a_2748_1611# a_2888_2122# 0.206f
C4402 a_15203_8914# a_15203_8684# 0.0292f
C4403 a_18086_6056# d2 0.0233f
C4404 a_2748_1611# a_2884_2299# 0.345f
C4405 a_1793_5434# vdd 0.0273f
C4406 a_4954_133# a_5053_133# 3.47f
C4407 a_15734_4621# a_15205_4918# 0.0185f
C4408 a_12807_7118# a_12913_7819# 0.423f
C4409 a_432_8987# d0 0.0235f
C4410 a_16897_2814# vdd 0.038f
C4411 a_2931_6521# a_3139_6521# 0.448f
C4412 a_431_8433# a_116_8638# 0.0467f
C4413 a_12918_4333# a_13853_4820# 0.254f
C4414 a_13853_2060# a_13859_1334# 0.0622f
C4415 a_18914_3581# a_18910_3758# 0.539f
C4416 a_2889_1019# a_2744_1788# 0.326f
C4417 a_856_3472# a_119_3353# 0.426f
C4418 a_7939_5649# a_7060_194# 0.137f
C4419 a_12918_5436# a_13171_5423# 0.11f
C4420 a_6859_4902# vdd 0.0264f
C4421 a_3823_952# vdd 0.314f
C4422 a_7941_1237# a_8880_1547# 0.112f
C4423 a_8876_6508# vdd 0.314f
C4424 a_3824_1506# a_3827_775# 0.0292f
C4425 a_6642_3269# a_5912_3513# 0.219f
C4426 a_18020_2155# a_18228_2155# 0.448f
C4427 a_3139_7624# vdd 0.183f
C4428 a_15943_2415# a_16460_2171# 0.0467f
C4429 a_857_1266# a_649_1266# 0.291f
C4430 a_17880_1644# a_17861_2924# 0.255f
C4431 a_10464_5129# a_10149_5334# 0.0467f
C4432 a_10148_7770# vdd 0.128f
C4433 a_5490_5719# a_5174_5829# 0.0467f
C4434 a_5491_3513# vdd 0.178f
C4435 a_11402_6542# a_11615_6542# 0.448f
C4436 a_18908_7067# a_18912_6890# 0.539f
C4437 a_12919_2127# a_12779_1616# 0.206f
C4438 a_15522_3518# a_15735_3518# 0.448f
C4439 a_117_7994# a_852_8433# 0.155f
C4440 a_17973_7683# a_18912_7993# 0.278f
C4441 a_854_5124# a_1372_5434# 0.11f
C4442 a_8876_9268# a_8880_9091# 0.539f
C4443 a_8194_8768# vdd 0.183f
C4444 a_12824_1603# a_12779_1616# 0.157f
C4445 a_7939_4546# vdd 0.439f
C4446 a_2792_3804# vdd 0.0325f
C4447 a_7938_7855# a_7942_7678# 0.518f
C4448 a_119_2666# a_855_2918# 0.279f
C4449 a_5492_1307# a_5913_1307# 0.0104f
C4450 a_17865_2747# a_17834_3863# 0.206f
C4451 a_120_1376# a_436_1266# 0.0467f
C4452 a_435_3472# a_856_3472# 0.0104f
C4453 a_2744_1788# vdd 0.0316f
C4454 a_11616_5439# a_11824_5439# 0.241f
C4455 a_8055_6051# a_7798_6241# 0.0467f
C4456 a_15942_1861# a_15206_2066# 0.255f
C4457 a_11543_5950# vdd 0.178f
C4458 a_7944_3266# a_8877_4302# 0.155f
C4459 a_18957_7980# vdd 0.0325f
C4460 a_17865_2747# vdd 0.0269f
C4461 a_16813_3785# a_16881_3274# 0.146f
C4462 a_8883_3576# d0 0.00533f
C4463 a_15203_8914# d0 0.0138f
C4464 a_8881_7988# a_8875_8714# 0.0622f
C4465 a_15205_5375# a_15942_5724# 0.112f
C4466 a_15206_3628# a_15943_3518# 0.277f
C4467 a_4078_6831# a_3825_6844# 0.11f
C4468 a_647_2918# a_855_2918# 0.3f
C4469 a_15521_5724# a_15942_5724# 0.0104f
C4470 a_2932_5418# a_2887_5431# 0.181f
C4471 a_13904_1321# a_13853_2060# 0.011f
C4472 a_15206_2525# a_15206_2712# 0.0625f
C4473 a_15943_2415# a_15735_2415# 0.291f
C4474 a_1803_7061# a_1481_7061# 0.11f
C4475 a_9135_5769# vdd 0.183f
C4476 a_10886_2923# vdd 0.1f
C4477 a_2934_1006# a_2885_1196# 0.219f
C4478 a_14985_138# gnd 3.45f  
C4479 a_9888_17# gnd 6.54f  
C4480 vout gnd 0.514f  
C4481 a_9779_17# gnd 0.902f  
C4482 a_9566_17# gnd 1.45f  
C4483 d7 gnd 0.594f  
C4484 a_14876_138# gnd 0.902f  
C4485 a_14663_138# gnd 1.45f  
C4486 d6 gnd 1.19f  
C4487 a_12134_158# gnd 4.59f  
C4488 a_11926_158# gnd 0.902f  
C4489 a_11713_158# gnd 1.45f  
C4490 d5 gnd 2.38f  
C4491 a_16982_199# gnd 0.902f  
C4492 a_16769_199# gnd 1.45f  
C4493 a_4954_133# gnd 3.45f  
C4494 a_5053_133# gnd 7.1f  
C4495 a_4845_133# gnd 0.902f  
C4496 a_4632_133# gnd 1.45f  
C4497 a_2103_153# gnd 4.59f  
C4498 a_1895_153# gnd 0.902f  
C4499 a_1682_153# gnd 1.45f  
C4500 a_6951_194# gnd 0.902f  
C4501 a_6738_194# gnd 1.45f  
C4502 a_18910_998# gnd 2.22f  
C4503 a_15209_864# gnd 6.46f  
C4504 a_15735_758# gnd 0.902f  
C4505 a_15522_758# gnd 1.45f  
C4506 d0 gnd 76.1f  
C4507 a_13854_957# gnd 2.22f  
C4508 a_10153_823# gnd 6.46f  
C4509 a_10679_717# gnd 0.902f  
C4510 a_10466_717# gnd 1.45f  
C4511 a_14111_767# gnd 1.45f  
C4512 a_13903_767# gnd 0.902f  
C4513 a_19167_808# gnd 1.45f  
C4514 a_18959_808# gnd 0.902f  
C4515 a_18914_821# gnd 2.45f  
C4516 a_15207_963# gnd 2.26f  
C4517 a_13858_780# gnd 2.45f  
C4518 a_17972_1242# gnd 2.38f  
C4519 d1 gnd 38f  
C4520 a_18229_1052# gnd 1.45f  
C4521 a_18021_1052# gnd 0.902f  
C4522 a_15943_758# gnd 2.59f  
C4523 a_8879_993# gnd 2.22f  
C4524 a_5178_859# gnd 6.46f  
C4525 a_5704_753# gnd 0.902f  
C4526 a_5491_753# gnd 1.45f  
C4527 a_3823_952# gnd 2.22f  
C4528 a_122_818# gnd 6.46f  
C4529 a_648_712# gnd 0.902f  
C4530 a_435_712# gnd 1.45f  
C4531 a_4080_762# gnd 1.45f  
C4532 a_3872_762# gnd 0.902f  
C4533 a_9136_803# gnd 1.45f  
C4534 a_8928_803# gnd 0.902f  
C4535 a_10151_922# gnd 2.26f  
C4536 a_12916_1201# gnd 2.38f  
C4537 a_13173_1011# gnd 1.45f  
C4538 a_12965_1011# gnd 0.902f  
C4539 a_10887_717# gnd 2.59f  
C4540 a_8883_816# gnd 2.45f  
C4541 a_11618_1027# gnd 0.902f  
C4542 a_11405_1027# gnd 1.45f  
C4543 a_5176_958# gnd 2.26f  
C4544 a_3827_775# gnd 2.45f  
C4545 a_16674_1068# gnd 0.902f  
C4546 a_16461_1068# gnd 1.45f  
C4547 a_15207_1193# gnd 2.45f  
C4548 a_15944_1312# gnd 2.23f  
C4549 a_7941_1237# gnd 2.38f  
C4550 a_8198_1047# gnd 1.45f  
C4551 a_7990_1047# gnd 0.902f  
C4552 a_5912_753# gnd 2.59f  
C4553 a_120_917# gnd 2.26f  
C4554 a_2885_1196# gnd 2.38f  
C4555 a_3142_1006# gnd 1.45f  
C4556 a_2934_1006# gnd 0.902f  
C4557 a_856_712# gnd 2.59f  
C4558 a_1587_1022# gnd 0.902f  
C4559 a_1374_1022# gnd 1.45f  
C4560 a_6643_1063# gnd 0.902f  
C4561 a_6430_1063# gnd 1.45f  
C4562 a_15207_1422# gnd 2.31f  
C4563 a_10151_1152# gnd 2.45f  
C4564 a_10888_1271# gnd 2.23f  
C4565 a_10151_1381# gnd 2.31f  
C4566 a_10680_1271# gnd 0.902f  
C4567 a_10467_1271# gnd 1.45f  
C4568 a_15736_1312# gnd 0.902f  
C4569 a_15523_1312# gnd 1.45f  
C4570 a_17976_1065# gnd 2.59f  
C4571 a_18911_1552# gnd 2.26f  
C4572 a_19168_1362# gnd 1.45f  
C4573 a_18960_1362# gnd 0.902f  
C4574 a_12920_1024# gnd 2.59f  
C4575 a_13855_1511# gnd 2.26f  
C4576 a_14112_1321# gnd 1.45f  
C4577 a_13904_1321# gnd 0.902f  
C4578 a_5176_1188# gnd 2.45f  
C4579 a_5913_1307# gnd 2.23f  
C4580 a_5176_1417# gnd 2.31f  
C4581 a_120_1147# gnd 2.45f  
C4582 a_857_1266# gnd 2.23f  
C4583 a_120_1376# gnd 2.31f  
C4584 a_649_1266# gnd 0.902f  
C4585 a_436_1266# gnd 1.45f  
C4586 a_5705_1307# gnd 0.902f  
C4587 a_5492_1307# gnd 1.45f  
C4588 a_18915_1375# gnd 2.5f  
C4589 a_16882_1068# gnd 1.48f  
C4590 a_7945_1060# gnd 2.59f  
C4591 a_8880_1547# gnd 2.26f  
C4592 a_9137_1357# gnd 1.45f  
C4593 a_8929_1357# gnd 0.902f  
C4594 a_2889_1019# gnd 2.59f  
C4595 a_3824_1506# gnd 2.26f  
C4596 a_4081_1316# gnd 1.45f  
C4597 a_3873_1316# gnd 0.902f  
C4598 a_16814_1579# gnd 0.902f  
C4599 a_16601_1579# gnd 1.45f  
C4600 d2 gnd 19f  
C4601 a_13859_1334# gnd 2.5f  
C4602 a_11826_1027# gnd 1.48f  
C4603 a_11758_1538# gnd 0.902f  
C4604 a_11545_1538# gnd 1.45f  
C4605 a_17831_1834# gnd 1.41f  
C4606 a_18088_1644# gnd 1.45f  
C4607 a_17880_1644# gnd 0.902f  
C4608 a_12775_1793# gnd 1.41f  
C4609 a_13032_1603# gnd 1.45f  
C4610 a_12824_1603# gnd 0.902f  
C4611 a_8884_1370# gnd 2.5f  
C4612 a_6851_1063# gnd 1.48f  
C4613 a_6783_1574# gnd 0.902f  
C4614 a_6570_1574# gnd 1.45f  
C4615 a_3828_1329# gnd 2.5f  
C4616 a_1795_1022# gnd 1.48f  
C4617 a_1727_1533# gnd 0.902f  
C4618 a_1514_1533# gnd 1.45f  
C4619 a_18909_2101# gnd 2.31f  
C4620 a_15207_1609# gnd 2.5f  
C4621 a_7800_1829# gnd 1.41f  
C4622 a_8057_1639# gnd 1.45f  
C4623 a_7849_1639# gnd 0.902f  
C4624 a_2744_1788# gnd 1.41f  
C4625 a_3001_1598# gnd 1.45f  
C4626 a_2793_1598# gnd 0.902f  
C4627 a_15734_1861# gnd 0.902f  
C4628 a_15521_1861# gnd 1.45f  
C4629 a_13853_2060# gnd 2.31f  
C4630 a_10151_1568# gnd 2.5f  
C4631 a_10678_1820# gnd 0.902f  
C4632 a_10465_1820# gnd 1.45f  
C4633 a_14110_1870# gnd 1.45f  
C4634 a_13902_1870# gnd 0.902f  
C4635 a_19166_1911# gnd 1.45f  
C4636 a_18958_1911# gnd 0.902f  
C4637 a_18913_1924# gnd 2.45f  
C4638 a_15206_2066# gnd 2.26f  
C4639 a_13857_1883# gnd 2.45f  
C4640 a_17835_1657# gnd 1.48f  
C4641 a_17971_2345# gnd 2.23f  
C4642 a_18228_2155# gnd 1.45f  
C4643 a_18020_2155# gnd 0.902f  
C4644 a_15942_1861# gnd 2.59f  
C4645 a_16881_2171# gnd 1.41f  
C4646 a_8878_2096# gnd 2.31f  
C4647 a_5176_1604# gnd 2.5f  
C4648 a_5703_1856# gnd 0.902f  
C4649 a_5490_1856# gnd 1.45f  
C4650 a_3822_2055# gnd 2.31f  
C4651 a_120_1563# gnd 2.5f  
C4652 a_647_1815# gnd 0.902f  
C4653 a_434_1815# gnd 1.45f  
C4654 a_4079_1865# gnd 1.45f  
C4655 a_3871_1865# gnd 0.902f  
C4656 a_9135_1906# gnd 1.45f  
C4657 a_8927_1906# gnd 0.902f  
C4658 a_10150_2025# gnd 2.26f  
C4659 a_12779_1616# gnd 1.48f  
C4660 a_12915_2304# gnd 2.23f  
C4661 a_13172_2114# gnd 1.45f  
C4662 a_12964_2114# gnd 0.902f  
C4663 a_10886_1820# gnd 2.59f  
C4664 a_11825_2130# gnd 1.41f  
C4665 a_8882_1919# gnd 2.45f  
C4666 a_11617_2130# gnd 0.902f  
C4667 a_11404_2130# gnd 1.45f  
C4668 a_5175_2061# gnd 2.26f  
C4669 a_3826_1878# gnd 2.45f  
C4670 a_16673_2171# gnd 0.902f  
C4671 a_16460_2171# gnd 1.45f  
C4672 a_15206_2296# gnd 2.45f  
C4673 a_15943_2415# gnd 2.49f  
C4674 a_7804_1652# gnd 1.48f  
C4675 a_7940_2340# gnd 2.23f  
C4676 a_8197_2150# gnd 1.45f  
C4677 a_7989_2150# gnd 0.902f  
C4678 a_5911_1856# gnd 2.59f  
C4679 a_6850_2166# gnd 1.41f  
C4680 a_119_2020# gnd 2.26f  
C4681 a_2748_1611# gnd 1.48f  
C4682 a_2884_2299# gnd 2.23f  
C4683 a_3141_2109# gnd 1.45f  
C4684 a_2933_2109# gnd 0.902f  
C4685 a_855_1815# gnd 2.59f  
C4686 a_1794_2125# gnd 1.41f  
C4687 a_1586_2125# gnd 0.902f  
C4688 a_1373_2125# gnd 1.45f  
C4689 a_6642_2166# gnd 0.902f  
C4690 a_6429_2166# gnd 1.45f  
C4691 a_15206_2525# gnd 2.31f  
C4692 a_10150_2255# gnd 2.45f  
C4693 a_10887_2374# gnd 2.49f  
C4694 a_10150_2484# gnd 2.31f  
C4695 a_10679_2374# gnd 0.902f  
C4696 a_10466_2374# gnd 1.45f  
C4697 a_15735_2415# gnd 0.902f  
C4698 a_15522_2415# gnd 1.45f  
C4699 a_17975_2168# gnd 2.59f  
C4700 a_18910_2655# gnd 2.26f  
C4701 a_19167_2465# gnd 1.45f  
C4702 a_18959_2465# gnd 0.902f  
C4703 a_12919_2127# gnd 2.59f  
C4704 a_13854_2614# gnd 2.26f  
C4705 a_14111_2424# gnd 1.45f  
C4706 a_13903_2424# gnd 0.902f  
C4707 a_5175_2291# gnd 2.45f  
C4708 a_5912_2410# gnd 2.49f  
C4709 a_5175_2520# gnd 2.31f  
C4710 a_119_2250# gnd 2.45f  
C4711 a_856_2369# gnd 2.49f  
C4712 a_119_2479# gnd 2.31f  
C4713 a_648_2369# gnd 0.902f  
C4714 a_435_2369# gnd 1.45f  
C4715 a_5704_2410# gnd 0.902f  
C4716 a_5491_2410# gnd 1.45f  
C4717 a_7944_2163# gnd 2.59f  
C4718 a_8879_2650# gnd 2.26f  
C4719 a_9136_2460# gnd 1.45f  
C4720 a_8928_2460# gnd 0.902f  
C4721 a_2888_2122# gnd 2.59f  
C4722 a_3823_2609# gnd 2.26f  
C4723 a_4080_2419# gnd 1.45f  
C4724 a_3872_2419# gnd 0.902f  
C4725 a_16892_2695# gnd 2.27f  
C4726 a_11836_2654# gnd 2.27f  
C4727 a_18914_2478# gnd 2.5f  
C4728 a_16783_2695# gnd 0.902f  
C4729 a_16570_2695# gnd 1.45f  
C4730 d3 gnd 9.51f  
C4731 a_13858_2437# gnd 2.5f  
C4732 a_17861_2924# gnd 2.04f  
C4733 a_18118_2734# gnd 1.45f  
C4734 a_17910_2734# gnd 0.902f  
C4735 a_11727_2654# gnd 0.902f  
C4736 a_11514_2654# gnd 1.45f  
C4737 a_12805_2883# gnd 2.04f  
C4738 a_13062_2693# gnd 1.45f  
C4739 a_12854_2693# gnd 0.902f  
C4740 a_6861_2690# gnd 2.27f  
C4741 a_1805_2649# gnd 2.27f  
C4742 a_8883_2473# gnd 2.5f  
C4743 a_18909_3204# gnd 2.31f  
C4744 a_15206_2712# gnd 2.5f  
C4745 a_6752_2690# gnd 0.902f  
C4746 a_6539_2690# gnd 1.45f  
C4747 a_3827_2432# gnd 2.5f  
C4748 a_7830_2919# gnd 2.04f  
C4749 a_8087_2729# gnd 1.45f  
C4750 a_7879_2729# gnd 0.902f  
C4751 a_1696_2649# gnd 0.902f  
C4752 a_1483_2649# gnd 1.45f  
C4753 a_2774_2878# gnd 2.04f  
C4754 a_3031_2688# gnd 1.45f  
C4755 a_2823_2688# gnd 0.902f  
C4756 a_15734_2964# gnd 0.902f  
C4757 a_15521_2964# gnd 1.45f  
C4758 a_13853_3163# gnd 2.31f  
C4759 a_10150_2671# gnd 2.5f  
C4760 a_10678_2923# gnd 0.902f  
C4761 a_10465_2923# gnd 1.45f  
C4762 a_14110_2973# gnd 1.45f  
C4763 a_13902_2973# gnd 0.902f  
C4764 a_19166_3014# gnd 1.45f  
C4765 a_18958_3014# gnd 0.902f  
C4766 a_18913_3027# gnd 2.45f  
C4767 a_15206_3169# gnd 2.26f  
C4768 a_13857_2986# gnd 2.45f  
C4769 a_17971_3448# gnd 2.49f  
C4770 a_18228_3258# gnd 1.45f  
C4771 a_18020_3258# gnd 0.902f  
C4772 a_15942_2964# gnd 2.59f  
C4773 a_8878_3199# gnd 2.31f  
C4774 a_5175_2707# gnd 2.5f  
C4775 a_5703_2959# gnd 0.902f  
C4776 a_5490_2959# gnd 1.45f  
C4777 a_3822_3158# gnd 2.31f  
C4778 a_119_2666# gnd 2.5f  
C4779 a_647_2918# gnd 0.902f  
C4780 a_434_2918# gnd 1.45f  
C4781 a_4079_2968# gnd 1.45f  
C4782 a_3871_2968# gnd 0.902f  
C4783 a_9135_3009# gnd 1.45f  
C4784 a_8927_3009# gnd 0.902f  
C4785 a_10150_3128# gnd 2.26f  
C4786 a_12915_3407# gnd 2.49f  
C4787 a_13172_3217# gnd 1.45f  
C4788 a_12964_3217# gnd 0.902f  
C4789 a_10886_2923# gnd 2.59f  
C4790 a_8882_3022# gnd 2.45f  
C4791 a_11617_3233# gnd 0.902f  
C4792 a_11404_3233# gnd 1.45f  
C4793 a_5175_3164# gnd 2.26f  
C4794 a_3826_2981# gnd 2.45f  
C4795 a_16673_3274# gnd 0.902f  
C4796 a_16460_3274# gnd 1.45f  
C4797 a_15206_3399# gnd 2.45f  
C4798 a_15943_3518# gnd 2.23f  
C4799 a_7940_3443# gnd 2.49f  
C4800 a_8197_3253# gnd 1.45f  
C4801 a_7989_3253# gnd 0.902f  
C4802 a_5911_2959# gnd 2.59f  
C4803 a_119_3123# gnd 2.26f  
C4804 a_2884_3402# gnd 2.49f  
C4805 a_3141_3212# gnd 1.45f  
C4806 a_2933_3212# gnd 0.902f  
C4807 a_855_2918# gnd 2.59f  
C4808 a_1586_3228# gnd 0.902f  
C4809 a_1373_3228# gnd 1.45f  
C4810 a_6642_3269# gnd 0.902f  
C4811 a_6429_3269# gnd 1.45f  
C4812 a_15206_3628# gnd 2.31f  
C4813 a_10150_3358# gnd 2.45f  
C4814 a_10887_3477# gnd 2.23f  
C4815 a_10150_3587# gnd 2.31f  
C4816 a_10679_3477# gnd 0.902f  
C4817 a_10466_3477# gnd 1.45f  
C4818 a_15735_3518# gnd 0.902f  
C4819 a_15522_3518# gnd 1.45f  
C4820 a_17975_3271# gnd 2.59f  
C4821 a_18910_3758# gnd 2.26f  
C4822 a_19167_3568# gnd 1.45f  
C4823 a_18959_3568# gnd 0.902f  
C4824 a_12919_3230# gnd 2.59f  
C4825 a_13854_3717# gnd 2.26f  
C4826 a_14111_3527# gnd 1.45f  
C4827 a_13903_3527# gnd 0.902f  
C4828 a_5175_3394# gnd 2.45f  
C4829 a_5912_3513# gnd 2.23f  
C4830 a_5175_3623# gnd 2.31f  
C4831 a_119_3353# gnd 2.45f  
C4832 a_856_3472# gnd 2.23f  
C4833 a_119_3582# gnd 2.31f  
C4834 a_648_3472# gnd 0.902f  
C4835 a_435_3472# gnd 1.45f  
C4836 a_5704_3513# gnd 0.902f  
C4837 a_5491_3513# gnd 1.45f  
C4838 a_18914_3581# gnd 2.5f  
C4839 a_16881_3274# gnd 1.48f  
C4840 a_16897_2814# gnd 2.45f  
C4841 a_7944_3266# gnd 2.59f  
C4842 a_8879_3753# gnd 2.26f  
C4843 a_9136_3563# gnd 1.45f  
C4844 a_8928_3563# gnd 0.902f  
C4845 a_2888_3225# gnd 2.59f  
C4846 a_3823_3712# gnd 2.26f  
C4847 a_4080_3522# gnd 1.45f  
C4848 a_3872_3522# gnd 0.902f  
C4849 a_16813_3785# gnd 0.902f  
C4850 a_16600_3785# gnd 1.45f  
C4851 a_13858_3540# gnd 2.5f  
C4852 a_11825_3233# gnd 1.48f  
C4853 a_11841_2773# gnd 2.45f  
C4854 a_11757_3744# gnd 0.902f  
C4855 a_11544_3744# gnd 1.45f  
C4856 a_17865_2747# gnd 2.33f  
C4857 a_17830_4040# gnd 1.41f  
C4858 a_18087_3850# gnd 1.45f  
C4859 a_17879_3850# gnd 0.902f  
C4860 a_12809_2706# gnd 2.33f  
C4861 a_12774_3999# gnd 1.41f  
C4862 a_13031_3809# gnd 1.45f  
C4863 a_12823_3809# gnd 0.902f  
C4864 a_8883_3576# gnd 2.5f  
C4865 a_6850_3269# gnd 1.48f  
C4866 a_6866_2809# gnd 2.45f  
C4867 a_6782_3780# gnd 0.902f  
C4868 a_6569_3780# gnd 1.45f  
C4869 a_3827_3535# gnd 2.5f  
C4870 a_1794_3228# gnd 1.48f  
C4871 a_1810_2768# gnd 2.45f  
C4872 a_1726_3739# gnd 0.902f  
C4873 a_1513_3739# gnd 1.45f  
C4874 a_18908_4307# gnd 2.31f  
C4875 a_15206_3815# gnd 2.5f  
C4876 a_7834_2742# gnd 2.33f  
C4877 a_7799_4035# gnd 1.41f  
C4878 a_8056_3845# gnd 1.45f  
C4879 a_7848_3845# gnd 0.902f  
C4880 a_2778_2701# gnd 2.33f  
C4881 a_2743_3994# gnd 1.41f  
C4882 a_3000_3804# gnd 1.45f  
C4883 a_2792_3804# gnd 0.902f  
C4884 a_15733_4067# gnd 0.902f  
C4885 a_15520_4067# gnd 1.45f  
C4886 a_13852_4266# gnd 2.31f  
C4887 a_10150_3774# gnd 2.5f  
C4888 a_10677_4026# gnd 0.902f  
C4889 a_10464_4026# gnd 1.45f  
C4890 a_14109_4076# gnd 1.45f  
C4891 a_13901_4076# gnd 0.902f  
C4892 a_19165_4117# gnd 1.45f  
C4893 a_18957_4117# gnd 0.902f  
C4894 a_18912_4130# gnd 2.45f  
C4895 a_15205_4272# gnd 2.26f  
C4896 a_13856_4089# gnd 2.45f  
C4897 a_17834_3863# gnd 1.48f  
C4898 a_17970_4551# gnd 2.23f  
C4899 a_18227_4361# gnd 1.45f  
C4900 a_18019_4361# gnd 0.902f  
C4901 a_15941_4067# gnd 2.59f  
C4902 a_16880_4377# gnd 1.41f  
C4903 a_8877_4302# gnd 2.31f  
C4904 a_5175_3810# gnd 2.5f  
C4905 a_5702_4062# gnd 0.902f  
C4906 a_5489_4062# gnd 1.45f  
C4907 a_3821_4261# gnd 2.31f  
C4908 a_119_3769# gnd 2.5f  
C4909 a_646_4021# gnd 0.902f  
C4910 a_433_4021# gnd 1.45f  
C4911 a_4078_4071# gnd 1.45f  
C4912 a_3870_4071# gnd 0.902f  
C4913 a_9134_4112# gnd 1.45f  
C4914 a_8926_4112# gnd 0.902f  
C4915 a_10149_4231# gnd 2.26f  
C4916 a_12778_3822# gnd 1.48f  
C4917 a_12914_4510# gnd 2.23f  
C4918 a_13171_4320# gnd 1.45f  
C4919 a_12963_4320# gnd 0.902f  
C4920 a_10885_4026# gnd 2.59f  
C4921 a_11824_4336# gnd 1.41f  
C4922 a_8881_4125# gnd 2.45f  
C4923 a_11616_4336# gnd 0.902f  
C4924 a_11403_4336# gnd 1.45f  
C4925 a_5174_4267# gnd 2.26f  
C4926 a_3825_4084# gnd 2.45f  
C4927 a_16672_4377# gnd 0.902f  
C4928 a_16459_4377# gnd 1.45f  
C4929 a_15205_4502# gnd 2.45f  
C4930 a_15942_4621# gnd 2.48f  
C4931 a_7803_3858# gnd 1.48f  
C4932 a_7939_4546# gnd 2.23f  
C4933 a_8196_4356# gnd 1.45f  
C4934 a_7988_4356# gnd 0.902f  
C4935 a_5910_4062# gnd 2.59f  
C4936 a_6849_4372# gnd 1.41f  
C4937 a_118_4226# gnd 2.26f  
C4938 a_2747_3817# gnd 1.48f  
C4939 a_2883_4505# gnd 2.23f  
C4940 a_3140_4315# gnd 1.45f  
C4941 a_2932_4315# gnd 0.902f  
C4942 a_854_4021# gnd 2.59f  
C4943 a_1793_4331# gnd 1.41f  
C4944 a_1585_4331# gnd 0.902f  
C4945 a_1372_4331# gnd 1.45f  
C4946 a_6641_4372# gnd 0.902f  
C4947 a_6428_4372# gnd 1.45f  
C4948 a_15205_4731# gnd 2.31f  
C4949 a_10149_4461# gnd 2.45f  
C4950 a_10886_4580# gnd 2.48f  
C4951 a_10149_4690# gnd 2.31f  
C4952 a_17974_4374# gnd 2.59f  
C4953 a_18909_4861# gnd 2.26f  
C4954 a_15734_4621# gnd 0.902f  
C4955 a_15521_4621# gnd 1.45f  
C4956 a_19166_4671# gnd 1.45f  
C4957 a_18958_4671# gnd 0.902f  
C4958 a_12918_4333# gnd 2.59f  
C4959 a_13853_4820# gnd 2.26f  
C4960 a_10678_4580# gnd 0.902f  
C4961 a_10465_4580# gnd 1.45f  
C4962 a_14110_4630# gnd 1.45f  
C4963 a_13902_4630# gnd 0.902f  
C4964 a_5174_4497# gnd 2.45f  
C4965 a_5911_4616# gnd 2.48f  
C4966 a_5174_4726# gnd 2.31f  
C4967 a_118_4456# gnd 2.45f  
C4968 a_855_4575# gnd 2.48f  
C4969 a_118_4685# gnd 2.31f  
C4970 a_7943_4369# gnd 2.59f  
C4971 a_8878_4856# gnd 2.26f  
C4972 a_5703_4616# gnd 0.902f  
C4973 a_5490_4616# gnd 1.45f  
C4974 a_9135_4666# gnd 1.45f  
C4975 a_8927_4666# gnd 0.902f  
C4976 a_18913_4684# gnd 2.51f  
C4977 a_17091_199# gnd 6.47f  
C4978 a_16890_4907# gnd 3.67f  
C4979 a_16989_4907# gnd 5.48f  
C4980 a_16781_4907# gnd 0.902f  
C4981 a_16568_4907# gnd 1.45f  
C4982 d4 gnd 4.75f  
C4983 a_13857_4643# gnd 2.51f  
C4984 a_17861_5124# gnd 3.32f  
C4985 a_18118_4934# gnd 1.45f  
C4986 a_17910_4934# gnd 0.902f  
C4987 a_12035_158# gnd 6.47f  
C4988 a_11834_4866# gnd 3.67f  
C4989 a_11933_4866# gnd 5.48f  
C4990 a_2887_4328# gnd 2.59f  
C4991 a_3822_4815# gnd 2.26f  
C4992 a_647_4575# gnd 0.902f  
C4993 a_434_4575# gnd 1.45f  
C4994 a_4079_4625# gnd 1.45f  
C4995 a_3871_4625# gnd 0.902f  
C4996 a_11725_4866# gnd 0.902f  
C4997 a_11512_4866# gnd 1.45f  
C4998 a_12805_5083# gnd 3.32f  
C4999 a_13062_4893# gnd 1.45f  
C5000 a_12854_4893# gnd 0.902f  
C5001 a_8882_4679# gnd 2.51f  
C5002 a_18908_5410# gnd 2.31f  
C5003 a_15205_4918# gnd 2.51f  
C5004 a_7060_194# gnd 6.47f  
C5005 a_6859_4902# gnd 3.67f  
C5006 a_6958_4902# gnd 5.48f  
C5007 a_6750_4902# gnd 0.902f  
C5008 a_6537_4902# gnd 1.45f  
C5009 a_3826_4638# gnd 2.51f  
C5010 a_7830_5119# gnd 3.32f  
C5011 a_8087_4929# gnd 1.45f  
C5012 a_7879_4929# gnd 0.902f  
C5013 a_2004_153# gnd 6.47f  
C5014 a_1803_4861# gnd 3.67f  
C5015 a_1902_4861# gnd 5.48f  
C5016 a_1694_4861# gnd 0.902f  
C5017 a_1481_4861# gnd 1.45f  
C5018 a_2774_5078# gnd 3.32f  
C5019 a_3031_4888# gnd 1.45f  
C5020 a_2823_4888# gnd 0.902f  
C5021 a_15733_5170# gnd 0.902f  
C5022 a_15520_5170# gnd 1.45f  
C5023 a_13852_5369# gnd 2.31f  
C5024 a_10149_4877# gnd 2.51f  
C5025 a_10677_5129# gnd 0.902f  
C5026 a_10464_5129# gnd 1.45f  
C5027 a_14109_5179# gnd 1.45f  
C5028 a_13901_5179# gnd 0.902f  
C5029 a_19165_5220# gnd 1.45f  
C5030 a_18957_5220# gnd 0.902f  
C5031 a_18912_5233# gnd 2.45f  
C5032 a_15205_5375# gnd 2.26f  
C5033 a_13856_5192# gnd 2.45f  
C5034 a_17970_5654# gnd 2.48f  
C5035 a_18227_5464# gnd 1.45f  
C5036 a_18019_5464# gnd 0.902f  
C5037 a_15941_5170# gnd 2.59f  
C5038 a_8877_5405# gnd 2.31f  
C5039 a_5174_4913# gnd 2.51f  
C5040 a_5702_5165# gnd 0.902f  
C5041 a_5489_5165# gnd 1.45f  
C5042 a_3821_5364# gnd 2.31f  
C5043 a_118_4872# gnd 2.51f  
C5044 a_646_5124# gnd 0.902f  
C5045 a_433_5124# gnd 1.45f  
C5046 a_4078_5174# gnd 1.45f  
C5047 a_3870_5174# gnd 0.902f  
C5048 a_9134_5215# gnd 1.45f  
C5049 a_8926_5215# gnd 0.902f  
C5050 a_10149_5334# gnd 2.26f  
C5051 a_12914_5613# gnd 2.48f  
C5052 a_13171_5423# gnd 1.45f  
C5053 a_12963_5423# gnd 0.902f  
C5054 a_10885_5129# gnd 2.59f  
C5055 a_8881_5228# gnd 2.45f  
C5056 a_11616_5439# gnd 0.902f  
C5057 a_11403_5439# gnd 1.45f  
C5058 a_5174_5370# gnd 2.26f  
C5059 a_3825_5187# gnd 2.45f  
C5060 a_16672_5480# gnd 0.902f  
C5061 a_16459_5480# gnd 1.45f  
C5062 a_15205_5605# gnd 2.45f  
C5063 a_15942_5724# gnd 2.23f  
C5064 a_7939_5649# gnd 2.48f  
C5065 a_8196_5459# gnd 1.45f  
C5066 a_7988_5459# gnd 0.902f  
C5067 a_5910_5165# gnd 2.59f  
C5068 a_118_5329# gnd 2.26f  
C5069 a_2883_5608# gnd 2.48f  
C5070 a_3140_5418# gnd 1.45f  
C5071 a_2932_5418# gnd 0.902f  
C5072 a_854_5124# gnd 2.59f  
C5073 a_1585_5434# gnd 0.902f  
C5074 a_1372_5434# gnd 1.45f  
C5075 a_6641_5475# gnd 0.902f  
C5076 a_6428_5475# gnd 1.45f  
C5077 a_15205_5834# gnd 2.31f  
C5078 a_10149_5564# gnd 2.45f  
C5079 a_10886_5683# gnd 2.23f  
C5080 a_10149_5793# gnd 2.31f  
C5081 a_10678_5683# gnd 0.902f  
C5082 a_10465_5683# gnd 1.45f  
C5083 a_15734_5724# gnd 0.902f  
C5084 a_15521_5724# gnd 1.45f  
C5085 a_17974_5477# gnd 2.59f  
C5086 a_18909_5964# gnd 2.26f  
C5087 a_19166_5774# gnd 1.45f  
C5088 a_18958_5774# gnd 0.902f  
C5089 a_12918_5436# gnd 2.59f  
C5090 a_13853_5923# gnd 2.26f  
C5091 a_14110_5733# gnd 1.45f  
C5092 a_13902_5733# gnd 0.902f  
C5093 a_5174_5600# gnd 2.45f  
C5094 a_5911_5719# gnd 2.23f  
C5095 a_5174_5829# gnd 2.31f  
C5096 a_118_5559# gnd 2.45f  
C5097 a_855_5678# gnd 2.23f  
C5098 a_118_5788# gnd 2.31f  
C5099 a_647_5678# gnd 0.902f  
C5100 a_434_5678# gnd 1.45f  
C5101 a_5703_5719# gnd 0.902f  
C5102 a_5490_5719# gnd 1.45f  
C5103 a_18913_5787# gnd 2.5f  
C5104 a_16880_5480# gnd 1.48f  
C5105 a_7943_5472# gnd 2.59f  
C5106 a_8878_5959# gnd 2.26f  
C5107 a_9135_5769# gnd 1.45f  
C5108 a_8927_5769# gnd 0.902f  
C5109 a_2887_5431# gnd 2.59f  
C5110 a_3822_5918# gnd 2.26f  
C5111 a_4079_5728# gnd 1.45f  
C5112 a_3871_5728# gnd 0.902f  
C5113 a_16812_5991# gnd 0.902f  
C5114 a_16599_5991# gnd 1.45f  
C5115 a_13857_5746# gnd 2.5f  
C5116 a_11824_5439# gnd 1.48f  
C5117 a_11756_5950# gnd 0.902f  
C5118 a_11543_5950# gnd 1.45f  
C5119 a_17829_6246# gnd 1.41f  
C5120 a_18086_6056# gnd 1.45f  
C5121 a_17878_6056# gnd 0.902f  
C5122 a_12773_6205# gnd 1.41f  
C5123 a_13030_6015# gnd 1.45f  
C5124 a_12822_6015# gnd 0.902f  
C5125 a_8882_5782# gnd 2.5f  
C5126 a_6849_5475# gnd 1.48f  
C5127 a_6781_5986# gnd 0.902f  
C5128 a_6568_5986# gnd 1.45f  
C5129 a_3826_5741# gnd 2.5f  
C5130 a_1793_5434# gnd 1.48f  
C5131 a_1725_5945# gnd 0.902f  
C5132 a_1512_5945# gnd 1.45f  
C5133 a_18907_6513# gnd 2.31f  
C5134 a_15205_6021# gnd 2.5f  
C5135 a_7798_6241# gnd 1.41f  
C5136 a_8055_6051# gnd 1.45f  
C5137 a_7847_6051# gnd 0.902f  
C5138 a_2742_6200# gnd 1.41f  
C5139 a_2999_6010# gnd 1.45f  
C5140 a_2791_6010# gnd 0.902f  
C5141 a_15732_6273# gnd 0.902f  
C5142 a_15519_6273# gnd 1.45f  
C5143 a_13851_6472# gnd 2.31f  
C5144 a_10149_5980# gnd 2.5f  
C5145 a_10676_6232# gnd 0.902f  
C5146 a_10463_6232# gnd 1.45f  
C5147 a_14108_6282# gnd 1.45f  
C5148 a_13900_6282# gnd 0.902f  
C5149 a_19164_6323# gnd 1.45f  
C5150 a_18956_6323# gnd 0.902f  
C5151 a_18911_6336# gnd 2.45f  
C5152 a_15204_6478# gnd 2.26f  
C5153 a_13855_6295# gnd 2.45f  
C5154 a_17833_6069# gnd 1.48f  
C5155 a_17969_6757# gnd 2.23f  
C5156 a_18226_6567# gnd 1.45f  
C5157 a_18018_6567# gnd 0.902f  
C5158 a_15940_6273# gnd 2.59f  
C5159 a_16879_6583# gnd 1.41f  
C5160 a_8876_6508# gnd 2.31f  
C5161 a_5174_6016# gnd 2.5f  
C5162 a_5701_6268# gnd 0.902f  
C5163 a_5488_6268# gnd 1.45f  
C5164 a_3820_6467# gnd 2.31f  
C5165 a_118_5975# gnd 2.5f  
C5166 a_645_6227# gnd 0.902f  
C5167 a_432_6227# gnd 1.45f  
C5168 a_4077_6277# gnd 1.45f  
C5169 a_3869_6277# gnd 0.902f  
C5170 a_9133_6318# gnd 1.45f  
C5171 a_8925_6318# gnd 0.902f  
C5172 a_10148_6437# gnd 2.26f  
C5173 a_12777_6028# gnd 1.48f  
C5174 a_12913_6716# gnd 2.23f  
C5175 a_13170_6526# gnd 1.45f  
C5176 a_12962_6526# gnd 0.902f  
C5177 a_10884_6232# gnd 2.59f  
C5178 a_11823_6542# gnd 1.41f  
C5179 a_8880_6331# gnd 2.45f  
C5180 a_11615_6542# gnd 0.902f  
C5181 a_11402_6542# gnd 1.45f  
C5182 a_5173_6473# gnd 2.26f  
C5183 a_3824_6290# gnd 2.45f  
C5184 a_16671_6583# gnd 0.902f  
C5185 a_16458_6583# gnd 1.45f  
C5186 a_15204_6708# gnd 2.45f  
C5187 a_15941_6827# gnd 2.49f  
C5188 a_7802_6064# gnd 1.48f  
C5189 a_7938_6752# gnd 2.23f  
C5190 a_8195_6562# gnd 1.45f  
C5191 a_7987_6562# gnd 0.902f  
C5192 a_5909_6268# gnd 2.59f  
C5193 a_6848_6578# gnd 1.41f  
C5194 a_117_6432# gnd 2.26f  
C5195 a_2746_6023# gnd 1.48f  
C5196 a_2882_6711# gnd 2.23f  
C5197 a_3139_6521# gnd 1.45f  
C5198 a_2931_6521# gnd 0.902f  
C5199 a_853_6227# gnd 2.59f  
C5200 a_1792_6537# gnd 1.41f  
C5201 a_1584_6537# gnd 0.902f  
C5202 a_1371_6537# gnd 1.45f  
C5203 a_6640_6578# gnd 0.902f  
C5204 a_6427_6578# gnd 1.45f  
C5205 a_15204_6937# gnd 2.31f  
C5206 a_10148_6667# gnd 2.45f  
C5207 a_10885_6786# gnd 2.49f  
C5208 a_10148_6896# gnd 2.31f  
C5209 a_10677_6786# gnd 0.902f  
C5210 a_10464_6786# gnd 1.45f  
C5211 a_15733_6827# gnd 0.902f  
C5212 a_15520_6827# gnd 1.45f  
C5213 a_17973_6580# gnd 2.59f  
C5214 a_18908_7067# gnd 2.26f  
C5215 a_19165_6877# gnd 1.45f  
C5216 a_18957_6877# gnd 0.902f  
C5217 a_12917_6539# gnd 2.59f  
C5218 a_13852_7026# gnd 2.26f  
C5219 a_14109_6836# gnd 1.45f  
C5220 a_13901_6836# gnd 0.902f  
C5221 a_5173_6703# gnd 2.45f  
C5222 a_5910_6822# gnd 2.49f  
C5223 a_5173_6932# gnd 2.31f  
C5224 a_117_6662# gnd 2.45f  
C5225 a_854_6781# gnd 2.49f  
C5226 a_117_6891# gnd 2.31f  
C5227 a_646_6781# gnd 0.902f  
C5228 a_433_6781# gnd 1.45f  
C5229 a_5702_6822# gnd 0.902f  
C5230 a_5489_6822# gnd 1.45f  
C5231 a_7942_6575# gnd 2.59f  
C5232 a_8877_7062# gnd 2.26f  
C5233 a_9134_6872# gnd 1.45f  
C5234 a_8926_6872# gnd 0.902f  
C5235 a_2886_6534# gnd 2.59f  
C5236 a_3821_7021# gnd 2.26f  
C5237 a_4078_6831# gnd 1.45f  
C5238 a_3870_6831# gnd 0.902f  
C5239 a_16890_7107# gnd 2.33f  
C5240 a_16895_5026# gnd 3.32f  
C5241 a_11834_7066# gnd 2.33f  
C5242 a_11839_4985# gnd 3.32f  
C5243 a_18912_6890# gnd 2.5f  
C5244 a_17865_4947# gnd 3.67f  
C5245 a_16781_7107# gnd 0.902f  
C5246 a_16568_7107# gnd 1.45f  
C5247 a_13856_6849# gnd 2.5f  
C5248 a_17859_7336# gnd 2.45f  
C5249 a_18116_7146# gnd 1.45f  
C5250 a_17908_7146# gnd 0.902f  
C5251 a_12809_4906# gnd 3.67f  
C5252 a_11725_7066# gnd 0.902f  
C5253 a_11512_7066# gnd 1.45f  
C5254 a_12803_7295# gnd 2.45f  
C5255 a_13060_7105# gnd 1.45f  
C5256 a_12852_7105# gnd 0.902f  
C5257 a_6859_7102# gnd 2.33f  
C5258 a_6864_5021# gnd 3.32f  
C5259 a_1803_7061# gnd 2.33f  
C5260 a_1808_4980# gnd 3.32f  
C5261 a_8881_6885# gnd 2.5f  
C5262 a_18907_7616# gnd 2.31f  
C5263 a_15204_7124# gnd 2.5f  
C5264 a_7834_4942# gnd 3.67f  
C5265 a_6750_7102# gnd 0.902f  
C5266 a_6537_7102# gnd 1.45f  
C5267 a_3825_6844# gnd 2.5f  
C5268 a_7828_7331# gnd 2.45f  
C5269 a_8085_7141# gnd 1.45f  
C5270 a_7877_7141# gnd 0.902f  
C5271 a_2778_4901# gnd 3.67f  
C5272 a_1694_7061# gnd 0.902f  
C5273 a_1481_7061# gnd 1.45f  
C5274 a_2772_7290# gnd 2.45f  
C5275 a_3029_7100# gnd 1.45f  
C5276 a_2821_7100# gnd 0.902f  
C5277 a_15732_7376# gnd 0.902f  
C5278 a_15519_7376# gnd 1.45f  
C5279 a_13851_7575# gnd 2.31f  
C5280 a_10148_7083# gnd 2.5f  
C5281 a_10676_7335# gnd 0.902f  
C5282 a_10463_7335# gnd 1.45f  
C5283 a_14108_7385# gnd 1.45f  
C5284 a_13900_7385# gnd 0.902f  
C5285 a_19164_7426# gnd 1.45f  
C5286 a_18956_7426# gnd 0.902f  
C5287 a_18911_7439# gnd 2.45f  
C5288 a_15204_7581# gnd 2.26f  
C5289 a_13855_7398# gnd 2.45f  
C5290 a_17969_7860# gnd 2.49f  
C5291 a_18226_7670# gnd 1.45f  
C5292 a_18018_7670# gnd 0.902f  
C5293 a_15940_7376# gnd 2.59f  
C5294 a_8876_7611# gnd 2.31f  
C5295 a_5173_7119# gnd 2.5f  
C5296 a_5701_7371# gnd 0.902f  
C5297 a_5488_7371# gnd 1.45f  
C5298 a_3820_7570# gnd 2.31f  
C5299 a_117_7078# gnd 2.5f  
C5300 a_645_7330# gnd 0.902f  
C5301 a_432_7330# gnd 1.45f  
C5302 a_4077_7380# gnd 1.45f  
C5303 a_3869_7380# gnd 0.902f  
C5304 a_9133_7421# gnd 1.45f  
C5305 a_8925_7421# gnd 0.902f  
C5306 a_10148_7540# gnd 2.26f  
C5307 a_12913_7819# gnd 2.49f  
C5308 a_13170_7629# gnd 1.45f  
C5309 a_12962_7629# gnd 0.902f  
C5310 a_10884_7335# gnd 2.59f  
C5311 a_8880_7434# gnd 2.45f  
C5312 a_11615_7645# gnd 0.902f  
C5313 a_11402_7645# gnd 1.45f  
C5314 a_5173_7576# gnd 2.26f  
C5315 a_3824_7393# gnd 2.45f  
C5316 a_16671_7686# gnd 0.902f  
C5317 a_16458_7686# gnd 1.45f  
C5318 a_15204_7811# gnd 2.45f  
C5319 a_15941_7930# gnd 2.23f  
C5320 a_7938_7855# gnd 2.49f  
C5321 a_8195_7665# gnd 1.45f  
C5322 a_7987_7665# gnd 0.902f  
C5323 a_5909_7371# gnd 2.59f  
C5324 a_117_7535# gnd 2.26f  
C5325 a_2882_7814# gnd 2.49f  
C5326 a_3139_7624# gnd 1.45f  
C5327 a_2931_7624# gnd 0.902f  
C5328 a_853_7330# gnd 2.59f  
C5329 a_1584_7640# gnd 0.902f  
C5330 a_1371_7640# gnd 1.45f  
C5331 a_6640_7681# gnd 0.902f  
C5332 a_6427_7681# gnd 1.45f  
C5333 a_15204_8040# gnd 2.31f  
C5334 a_10148_7770# gnd 2.45f  
C5335 a_10885_7889# gnd 2.23f  
C5336 a_10148_7999# gnd 2.31f  
C5337 a_10677_7889# gnd 0.902f  
C5338 a_10464_7889# gnd 1.45f  
C5339 a_15733_7930# gnd 0.902f  
C5340 a_15520_7930# gnd 1.45f  
C5341 a_17973_7683# gnd 2.59f  
C5342 a_18908_8170# gnd 2.26f  
C5343 a_19165_7980# gnd 1.45f  
C5344 a_18957_7980# gnd 0.902f  
C5345 a_12917_7642# gnd 2.59f  
C5346 a_13852_8129# gnd 2.26f  
C5347 a_14109_7939# gnd 1.45f  
C5348 a_13901_7939# gnd 0.902f  
C5349 a_5173_7806# gnd 2.45f  
C5350 a_5910_7925# gnd 2.23f  
C5351 a_5173_8035# gnd 2.31f  
C5352 a_117_7765# gnd 2.45f  
C5353 a_854_7884# gnd 2.23f  
C5354 a_117_7994# gnd 2.31f  
C5355 a_646_7884# gnd 0.902f  
C5356 a_433_7884# gnd 1.45f  
C5357 a_5702_7925# gnd 0.902f  
C5358 a_5489_7925# gnd 1.45f  
C5359 a_18912_7993# gnd 2.5f  
C5360 a_16879_7686# gnd 1.48f  
C5361 a_16895_7226# gnd 2.04f  
C5362 a_7942_7678# gnd 2.59f  
C5363 a_8877_8165# gnd 2.26f  
C5364 a_9134_7975# gnd 1.45f  
C5365 a_8926_7975# gnd 0.902f  
C5366 a_2886_7637# gnd 2.59f  
C5367 a_3821_8124# gnd 2.26f  
C5368 a_4078_7934# gnd 1.45f  
C5369 a_3870_7934# gnd 0.902f  
C5370 a_16811_8197# gnd 0.902f  
C5371 a_16598_8197# gnd 1.45f  
C5372 a_13856_7952# gnd 2.5f  
C5373 a_11823_7645# gnd 1.48f  
C5374 a_11839_7185# gnd 2.04f  
C5375 a_11755_8156# gnd 0.902f  
C5376 a_11542_8156# gnd 1.45f  
C5377 a_17863_7159# gnd 2.27f  
C5378 a_17828_8452# gnd 1.41f  
C5379 a_18085_8262# gnd 1.45f  
C5380 a_17877_8262# gnd 0.902f  
C5381 a_12807_7118# gnd 2.27f  
C5382 a_12772_8411# gnd 1.41f  
C5383 a_13029_8221# gnd 1.45f  
C5384 a_12821_8221# gnd 0.902f  
C5385 a_8881_7988# gnd 2.5f  
C5386 a_6848_7681# gnd 1.48f  
C5387 a_6864_7221# gnd 2.04f  
C5388 a_6780_8192# gnd 0.902f  
C5389 a_6567_8192# gnd 1.45f  
C5390 a_3825_7947# gnd 2.5f  
C5391 a_1792_7640# gnd 1.48f  
C5392 a_1808_7180# gnd 2.04f  
C5393 a_1724_8151# gnd 0.902f  
C5394 a_1511_8151# gnd 1.45f  
C5395 a_18906_8719# gnd 2.31f  
C5396 a_15204_8227# gnd 2.5f  
C5397 a_7832_7154# gnd 2.27f  
C5398 a_7797_8447# gnd 1.41f  
C5399 a_8054_8257# gnd 1.45f  
C5400 a_7846_8257# gnd 0.902f  
C5401 a_2776_7113# gnd 2.27f  
C5402 a_2741_8406# gnd 1.41f  
C5403 a_2998_8216# gnd 1.45f  
C5404 a_2790_8216# gnd 0.902f  
C5405 a_15731_8479# gnd 0.902f  
C5406 a_15518_8479# gnd 1.45f  
C5407 a_13850_8678# gnd 2.31f  
C5408 a_10148_8186# gnd 2.5f  
C5409 a_10675_8438# gnd 0.902f  
C5410 a_10462_8438# gnd 1.45f  
C5411 a_14107_8488# gnd 1.45f  
C5412 a_13899_8488# gnd 0.902f  
C5413 a_19163_8529# gnd 1.45f  
C5414 a_18955_8529# gnd 0.902f  
C5415 a_18910_8542# gnd 2.45f  
C5416 a_15203_8684# gnd 2.26f  
C5417 a_13854_8501# gnd 2.45f  
C5418 a_17832_8275# gnd 1.48f  
C5419 a_17968_8963# gnd 2.23f  
C5420 a_18225_8773# gnd 1.45f  
C5421 a_18017_8773# gnd 0.902f  
C5422 a_15939_8479# gnd 2.59f  
C5423 a_16878_8789# gnd 1.41f  
C5424 a_8875_8714# gnd 2.31f  
C5425 a_5173_8222# gnd 2.5f  
C5426 a_5700_8474# gnd 0.902f  
C5427 a_5487_8474# gnd 1.45f  
C5428 a_3819_8673# gnd 2.31f  
C5429 a_117_8181# gnd 2.5f  
C5430 a_644_8433# gnd 0.902f  
C5431 a_431_8433# gnd 1.45f  
C5432 a_4076_8483# gnd 1.45f  
C5433 a_3868_8483# gnd 0.902f  
C5434 a_9132_8524# gnd 1.45f  
C5435 a_8924_8524# gnd 0.902f  
C5436 a_10147_8643# gnd 2.26f  
C5437 a_12776_8234# gnd 1.48f  
C5438 a_12912_8922# gnd 2.23f  
C5439 a_13169_8732# gnd 1.45f  
C5440 a_12961_8732# gnd 0.902f  
C5441 a_10883_8438# gnd 2.59f  
C5442 a_11822_8748# gnd 1.41f  
C5443 a_8879_8537# gnd 2.45f  
C5444 a_11614_8748# gnd 0.902f  
C5445 a_11401_8748# gnd 1.45f  
C5446 a_5172_8679# gnd 2.26f  
C5447 a_3823_8496# gnd 2.45f  
C5448 a_16670_8789# gnd 0.902f  
C5449 a_16457_8789# gnd 1.45f  
C5450 a_15203_8914# gnd 2.45f  
C5451 a_15940_9033# gnd 2.38f  
C5452 a_7801_8270# gnd 1.48f  
C5453 a_7937_8958# gnd 2.23f  
C5454 a_8194_8768# gnd 1.45f  
C5455 a_7986_8768# gnd 0.902f  
C5456 a_5908_8474# gnd 2.59f  
C5457 a_6847_8784# gnd 1.41f  
C5458 a_116_8638# gnd 2.26f  
C5459 a_2745_8229# gnd 1.48f  
C5460 a_2881_8917# gnd 2.23f  
C5461 a_3138_8727# gnd 1.45f  
C5462 a_2930_8727# gnd 0.902f  
C5463 a_852_8433# gnd 2.59f  
C5464 a_1791_8743# gnd 1.41f  
C5465 a_1583_8743# gnd 0.902f  
C5466 a_1370_8743# gnd 1.45f  
C5467 a_6639_8784# gnd 0.902f  
C5468 a_6426_8784# gnd 1.45f  
C5469 a_15203_9143# gnd 2.22f  
C5470 a_10147_8873# gnd 2.45f  
C5471 a_10884_8992# gnd 2.38f  
C5472 a_10147_9102# gnd 2.22f  
C5473 a_10676_8992# gnd 0.902f  
C5474 a_10463_8992# gnd 1.45f  
C5475 a_15732_9033# gnd 0.902f  
C5476 a_15519_9033# gnd 1.45f  
C5477 a_17972_8786# gnd 2.87f  
C5478 a_18907_9273# gnd 2.79f  
C5479 a_19164_9083# gnd 1.56f  
C5480 a_18956_9083# gnd 1.05f  
C5481 a_12916_8745# gnd 2.59f  
C5482 a_13851_9232# gnd 2.26f  
C5483 a_14108_9042# gnd 1.45f  
C5484 a_13900_9042# gnd 0.902f  
C5485 a_5172_8909# gnd 2.45f  
C5486 a_5909_9028# gnd 2.38f  
C5487 a_5172_9138# gnd 2.22f  
C5488 a_116_8868# gnd 2.45f  
C5489 a_853_8987# gnd 2.38f  
C5490 a_116_9097# gnd 2.22f  
C5491 a_645_8987# gnd 0.902f  
C5492 a_432_8987# gnd 1.45f  
C5493 a_5701_9028# gnd 0.902f  
C5494 a_5488_9028# gnd 1.45f  
C5495 a_13855_9055# gnd 3.01f  
C5496 a_8880_9091# gnd 2.83f  
C5497 a_7941_8781# gnd 2.59f  
C5498 a_8876_9268# gnd 2.26f  
C5499 a_9133_9078# gnd 1.45f  
C5500 a_8925_9078# gnd 0.902f  
C5501 a_2885_8740# gnd 2.59f  
C5502 a_3820_9227# gnd 2.26f  
C5503 a_4077_9037# gnd 1.45f  
C5504 a_3869_9037# gnd 0.902f  
C5505 vref gnd 0.154f  
C5506 a_3824_9050# gnd 3.01f  
C5507 vdd gnd 0.578p  

Vdd vdd 0 dc 3.3
Vin1 vref 0 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5us 10us)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10us 20us)
Vd2 d2 0 pulse(0 1.8 0ns 0.1ns 0.1ns 20us 40us)
Vd3 d3 0 pulse(0 1.8 0ns 0.1ns 0.1ns 40us 80us)
Vd4 d4 0 pulse(0 1.8 0ns 0.1ns 0.1ns 80us 160us)
Vd5 d5 0 pulse(0 1.8 0ns 0.1ns 0.1ns 160us 320us)
Vd6 d6 0 pulse(0 1.8 0ns 0.1ns 0.1ns 320us 640us)
Vd7 d7 0 pulse(0 1.8 0ns 0.1ns 0.1ns 640us 1280us)

*.tran 0.1us 1280us
*.control
*run
*plot V(vout) 
*.endc
*.end

*.tran 0.001us 20us
*.tran 10us 1280us
.tran 10us 1280us


* Control Statements 
.control
run
print allv > plot_data_v.txt
print alli > plot_data_i.txt

print v(vout) > output_v.txt

plot vout
.endc
.end