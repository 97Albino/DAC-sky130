** sch_path: /home/97ms/uci/ip/dac5v/1.schematics/2bit_dac.sch

.include sw.spice

.subckt 2bit_dac vdd vss vrefh vrefl d0 d1 vout
XR1 net3 vrefh vss sky130_fd_pr__res_high_po_0p35 L=1.09 mult=1
XR2 net4 net3 vss sky130_fd_pr__res_high_po_0p35 L=1.09 mult=1
XR3 net5 net4 vss sky130_fd_pr__res_high_po_0p35 L=1.09 mult=1
XR4 vrefl net5 vss sky130_fd_pr__res_high_po_0p35 L=1.09 mult=1
X1 vdd vss d0 net3 net4 net2 sw
X2 vdd vss d0 net5 vrefl net1 sw
X3 vdd vss d1 net2 net1 vout sw
.ends
