magic
tech sky130B
magscale 1 2
timestamp 1687966408
<< locali >>
rect 0 700 1650 720
rect 0 660 70 700
rect 1580 660 1650 700
rect 0 568 1650 660
rect 0 70 70 568
rect 1580 70 1650 568
rect 0 0 1650 70
rect 0 -270 1650 -200
rect 0 -634 70 -270
rect 1586 -634 1650 -270
rect 0 -726 1650 -634
rect 0 -766 70 -726
rect 1580 -766 1650 -726
rect 0 -786 1650 -766
<< viali >>
rect 70 660 1580 700
rect 70 -766 1580 -726
<< metal1 >>
rect 0 700 1650 720
rect 0 660 70 700
rect 1580 660 1650 700
rect 0 568 1650 660
rect 70 420 150 568
rect 70 218 190 420
rect 224 178 272 460
rect 456 420 516 568
rect 302 218 402 420
rect 456 218 576 420
rect 200 -60 292 132
rect 0 -140 292 -60
rect 200 -332 292 -140
rect 332 -60 402 218
rect 608 178 656 460
rect 688 408 788 420
rect 688 230 710 408
rect 770 230 788 408
rect 688 218 788 230
rect 862 408 962 420
rect 862 230 880 408
rect 940 230 962 408
rect 862 218 962 230
rect 994 178 1042 460
rect 1074 218 1348 420
rect 586 -60 678 132
rect 972 -60 1064 132
rect 332 -140 1064 -60
rect 70 -494 190 -410
rect 70 -634 150 -494
rect 222 -526 270 -378
rect 332 -410 402 -140
rect 586 -332 678 -140
rect 972 -332 1064 -140
rect 302 -494 402 -410
rect 456 -494 576 -410
rect 456 -634 536 -494
rect 608 -526 656 -378
rect 688 -422 788 -410
rect 688 -482 710 -422
rect 770 -482 788 -422
rect 688 -494 788 -482
rect 862 -422 962 -410
rect 862 -482 880 -422
rect 940 -482 962 -422
rect 862 -494 962 -482
rect 994 -526 1042 -378
rect 1170 -410 1252 218
rect 1380 178 1428 460
rect 1460 400 1720 420
rect 1460 240 1640 400
rect 1700 240 1720 400
rect 1460 218 1720 240
rect 1358 -70 1450 132
rect 1358 -130 1374 -70
rect 1434 -130 1450 -70
rect 1358 -332 1450 -130
rect 1074 -494 1348 -410
rect 1380 -526 1428 -378
rect 1460 -422 1580 -410
rect 1460 -482 1510 -422
rect 1570 -482 1580 -422
rect 1460 -494 1580 -482
rect 0 -726 1650 -634
rect 0 -766 70 -726
rect 1580 -766 1650 -726
rect 0 -786 1650 -766
<< via1 >>
rect 710 230 770 408
rect 880 230 940 408
rect 710 -482 770 -422
rect 880 -482 940 -422
rect 1640 240 1700 400
rect 1374 -130 1434 -70
rect 1510 -482 1570 -422
<< metal2 >>
rect 870 520 1580 600
rect 700 408 780 420
rect 700 230 710 408
rect 770 230 780 408
rect 700 -60 780 230
rect 870 408 950 520
rect 870 230 880 408
rect 940 230 950 408
rect 870 220 950 230
rect 700 -70 1450 -60
rect 700 -130 1374 -70
rect 1434 -130 1450 -70
rect 700 -140 1450 -130
rect 700 -422 780 -140
rect 700 -482 710 -422
rect 770 -482 780 -422
rect 700 -492 780 -482
rect 870 -422 950 -412
rect 870 -482 880 -422
rect 940 -482 950 -422
rect 870 -586 950 -482
rect 1500 -422 1580 520
rect 1500 -482 1510 -422
rect 1570 -482 1580 -422
rect 1500 -494 1580 -482
rect 1630 400 1710 410
rect 1630 240 1640 400
rect 1700 240 1710 400
rect 1630 -586 1710 240
rect 870 -666 1710 -586
use sky130_fd_pr__pfet_01v8_XPYSY6  XM1
timestamp 1687761602
transform 1 0 246 0 1 319
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_XPYSY6  XM2
timestamp 1687761602
transform 1 0 632 0 1 319
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_XPYSY6  XM3
timestamp 1687761602
transform 1 0 1018 0 1 319
box -246 -319 246 319
use sky130_fd_pr__pfet_01v8_XPYSY6  XM4
timestamp 1687761602
transform 1 0 1404 0 1 319
box -246 -319 246 319
use sky130_fd_pr__nfet_01v8_ZFH27D  XM5
timestamp 1687760742
transform 1 0 246 0 1 -452
box -246 -252 246 252
use sky130_fd_pr__nfet_01v8_ZFH27D  XM6
timestamp 1687760742
transform 1 0 632 0 1 -452
box -246 -252 246 252
use sky130_fd_pr__nfet_01v8_ZFH27D  XM7
timestamp 1687760742
transform 1 0 1018 0 1 -452
box -246 -252 246 252
use sky130_fd_pr__nfet_01v8_ZFH27D  XM8
timestamp 1687760742
transform 1 0 1404 0 1 -452
box -246 -252 246 252
<< labels >>
flabel metal1 20 660 60 700 0 FreeSans 128 0 0 0 vdd
port 0 nsew
flabel metal1 20 -766 60 -726 0 FreeSans 128 0 0 0 vss
port 1 nsew
flabel metal1 0 -120 40 -80 0 FreeSans 128 0 0 0 din
port 2 nsew
flabel metal1 862 380 902 420 0 FreeSans 128 0 0 0 vin1
port 3 nsew
flabel metal1 862 -494 902 -454 0 FreeSans 128 0 0 0 vin2
port 4 nsew
flabel metal1 1180 -120 1220 -80 0 FreeSans 128 0 0 0 vout
port 5 nsew
<< end >>
