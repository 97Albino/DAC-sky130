magic
tech sky130B
magscale 1 2
timestamp 1687795939
<< pwell >>
rect -201 -707 201 707
<< psubdiff >>
rect -165 637 -69 671
rect 69 637 165 671
rect -165 575 -131 637
rect 131 575 165 637
rect -165 -637 -131 -575
rect 131 -637 165 -575
rect -165 -671 -69 -637
rect 69 -671 165 -637
<< psubdiffcont >>
rect -69 637 69 671
rect -165 -575 -131 575
rect 131 -575 165 575
rect -69 -671 69 -637
<< xpolycontact >>
rect -35 109 35 541
rect -35 -541 35 -109
<< ppolyres >>
rect -35 -109 35 109
<< locali >>
rect -165 637 -69 671
rect 69 637 165 671
rect -165 575 -131 637
rect 131 575 165 637
rect -165 -637 -131 -575
rect 131 -637 165 -575
rect -165 -671 -69 -637
rect 69 -671 165 -637
<< viali >>
rect -19 126 19 523
rect -19 -523 19 -126
<< metal1 >>
rect -25 523 25 535
rect -25 126 -19 523
rect 19 126 25 523
rect -25 114 25 126
rect -25 -126 25 -114
rect -25 -523 -19 -126
rect 19 -523 25 -126
rect -25 -535 25 -523
<< res0p35 >>
rect -37 -111 37 111
<< properties >>
string FIXED_BBOX -148 -654 148 654
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 1.09 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.109k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
