MACRO SW
  ORIGIN 0 0 ;
  FOREIGN SW 0 0 ;
  SIZE 5.16 BY 30.24 ;
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
      LAYER M2 ;
        RECT 2.84 6.58 4.04 6.86 ;
      LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
      LAYER M2 ;
        RECT 2.84 14.14 4.04 14.42 ;
      LAYER M2 ;
        RECT 2.84 15.82 4.04 16.1 ;
      LAYER M2 ;
        RECT 1.12 29.26 2.32 29.54 ;
      LAYER M2 ;
        RECT 3.28 0.7 3.6 0.98 ;
      LAYER M3 ;
        RECT 3.3 0.84 3.58 6.72 ;
      LAYER M2 ;
        RECT 3.28 6.58 3.6 6.86 ;
      LAYER M3 ;
        RECT 3.3 6.72 3.58 8.4 ;
      LAYER M2 ;
        RECT 3.28 8.26 3.6 8.54 ;
      LAYER M3 ;
        RECT 3.3 8.4 3.58 14.28 ;
      LAYER M2 ;
        RECT 3.28 14.14 3.6 14.42 ;
      LAYER M3 ;
        RECT 3.3 14.28 3.58 15.96 ;
      LAYER M2 ;
        RECT 3.28 15.82 3.6 16.1 ;
      LAYER M2 ;
        RECT 2.85 15.82 3.17 16.1 ;
      LAYER M1 ;
        RECT 2.885 15.96 3.135 28.98 ;
      LAYER M2 ;
        RECT 2.15 28.84 3.01 29.12 ;
      LAYER M1 ;
        RECT 2.025 28.98 2.275 29.4 ;
      LAYER M2 ;
        RECT 1.99 29.26 2.31 29.54 ;
    END
  END VDD
  PIN DIGITAL_INPUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
      LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
      LAYER M2 ;
        RECT 2.15 0.28 3.01 0.56 ;
    END
  END DIGITAL_INPUT
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 17.92 2.32 18.2 ;
      LAYER M2 ;
        RECT 2.84 17.92 4.04 18.2 ;
      LAYER M2 ;
        RECT 2.15 17.92 3.01 18.2 ;
      LAYER M2 ;
        RECT 1.12 27.16 2.32 27.44 ;
      LAYER M2 ;
        RECT 2.84 27.16 4.04 27.44 ;
      LAYER M2 ;
        RECT 2.15 27.16 3.01 27.44 ;
      LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
      LAYER M3 ;
        RECT 2.01 18.06 2.29 27.3 ;
      LAYER M2 ;
        RECT 1.99 27.16 2.31 27.44 ;
    END
  END VOUT
  PIN VIN2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.69 21.7 1.89 21.98 ;
      LAYER M2 ;
        RECT 0.69 23.38 1.89 23.66 ;
      LAYER M2 ;
        RECT 1.13 21.7 1.45 21.98 ;
      LAYER M3 ;
        RECT 1.15 21.84 1.43 23.52 ;
      LAYER M2 ;
        RECT 1.13 23.38 1.45 23.66 ;
    END
  END VIN2
  PIN VIN1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.27 21.7 4.47 21.98 ;
      LAYER M2 ;
        RECT 3.27 23.38 4.47 23.66 ;
      LAYER M2 ;
        RECT 3.71 21.7 4.03 21.98 ;
      LAYER M3 ;
        RECT 3.73 21.84 4.01 23.52 ;
      LAYER M2 ;
        RECT 3.71 23.38 4.03 23.66 ;
    END
  END VIN1
  OBS 
  LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
  LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
  LAYER M2 ;
        RECT 2.15 4.48 3.01 4.76 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 2.15 7.84 3.01 8.12 ;
  LAYER M2 ;
        RECT 1.12 22.12 2.32 22.4 ;
  LAYER M2 ;
        RECT 2.84 22.12 4.04 22.4 ;
  LAYER M2 ;
        RECT 2.15 22.12 3.01 22.4 ;
  LAYER M2 ;
        RECT 2.42 4.48 2.74 4.76 ;
  LAYER M1 ;
        RECT 2.455 4.62 2.705 7.98 ;
  LAYER M2 ;
        RECT 2.42 7.84 2.74 8.12 ;
  LAYER M1 ;
        RECT 2.455 7.98 2.705 22.26 ;
  LAYER M2 ;
        RECT 2.42 22.12 2.74 22.4 ;
  LAYER M1 ;
        RECT 2.455 4.535 2.705 4.705 ;
  LAYER M2 ;
        RECT 2.41 4.48 2.75 4.76 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 8.065 ;
  LAYER M2 ;
        RECT 2.41 7.84 2.75 8.12 ;
  LAYER M1 ;
        RECT 2.455 4.535 2.705 4.705 ;
  LAYER M2 ;
        RECT 2.41 4.48 2.75 4.76 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 8.065 ;
  LAYER M2 ;
        RECT 2.41 7.84 2.75 8.12 ;
  LAYER M1 ;
        RECT 2.455 4.535 2.705 4.705 ;
  LAYER M2 ;
        RECT 2.41 4.48 2.75 4.76 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 8.065 ;
  LAYER M2 ;
        RECT 2.41 7.84 2.75 8.12 ;
  LAYER M1 ;
        RECT 2.455 22.175 2.705 22.345 ;
  LAYER M2 ;
        RECT 2.41 22.12 2.75 22.4 ;
  LAYER M1 ;
        RECT 2.455 4.535 2.705 4.705 ;
  LAYER M2 ;
        RECT 2.41 4.48 2.75 4.76 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 8.065 ;
  LAYER M2 ;
        RECT 2.41 7.84 2.75 8.12 ;
  LAYER M1 ;
        RECT 2.455 22.175 2.705 22.345 ;
  LAYER M2 ;
        RECT 2.41 22.12 2.75 22.4 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 1.12 14.14 2.32 14.42 ;
  LAYER M2 ;
        RECT 1.12 15.82 2.32 16.1 ;
  LAYER M2 ;
        RECT 2.84 29.26 4.04 29.54 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.84 1.86 6.72 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.72 1.86 8.4 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.4 1.86 14.28 ;
  LAYER M2 ;
        RECT 1.56 14.14 1.88 14.42 ;
  LAYER M3 ;
        RECT 1.58 14.28 1.86 15.96 ;
  LAYER M2 ;
        RECT 1.56 15.82 1.88 16.1 ;
  LAYER M2 ;
        RECT 1.99 15.82 2.31 16.1 ;
  LAYER M1 ;
        RECT 2.025 15.96 2.275 28.56 ;
  LAYER M2 ;
        RECT 2.15 28.42 3.01 28.7 ;
  LAYER M3 ;
        RECT 2.87 28.56 3.15 29.4 ;
  LAYER M2 ;
        RECT 2.85 29.26 3.17 29.54 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 14.14 1.88 14.42 ;
  LAYER M3 ;
        RECT 1.58 14.12 1.86 14.44 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 14.14 1.88 14.42 ;
  LAYER M3 ;
        RECT 1.58 14.12 1.86 14.44 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 14.14 1.88 14.42 ;
  LAYER M3 ;
        RECT 1.58 14.12 1.86 14.44 ;
  LAYER M2 ;
        RECT 1.56 15.82 1.88 16.1 ;
  LAYER M3 ;
        RECT 1.58 15.8 1.86 16.12 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 14.14 1.88 14.42 ;
  LAYER M3 ;
        RECT 1.58 14.12 1.86 14.44 ;
  LAYER M2 ;
        RECT 1.56 15.82 1.88 16.1 ;
  LAYER M3 ;
        RECT 1.58 15.8 1.86 16.12 ;
  LAYER M1 ;
        RECT 2.025 15.875 2.275 16.045 ;
  LAYER M2 ;
        RECT 1.98 15.82 2.32 16.1 ;
  LAYER M1 ;
        RECT 2.025 28.475 2.275 28.645 ;
  LAYER M2 ;
        RECT 1.98 28.42 2.32 28.7 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 14.14 1.88 14.42 ;
  LAYER M3 ;
        RECT 1.58 14.12 1.86 14.44 ;
  LAYER M2 ;
        RECT 1.56 15.82 1.88 16.1 ;
  LAYER M3 ;
        RECT 1.58 15.8 1.86 16.12 ;
  LAYER M2 ;
        RECT 2.85 28.42 3.17 28.7 ;
  LAYER M3 ;
        RECT 2.87 28.4 3.15 28.72 ;
  LAYER M2 ;
        RECT 2.85 29.26 3.17 29.54 ;
  LAYER M3 ;
        RECT 2.87 29.24 3.15 29.56 ;
  LAYER M1 ;
        RECT 2.025 15.875 2.275 16.045 ;
  LAYER M2 ;
        RECT 1.98 15.82 2.32 16.1 ;
  LAYER M1 ;
        RECT 2.025 28.475 2.275 28.645 ;
  LAYER M2 ;
        RECT 1.98 28.42 2.32 28.7 ;
  LAYER M2 ;
        RECT 1.56 0.7 1.88 0.98 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 1 ;
  LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
  LAYER M3 ;
        RECT 1.58 6.56 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 14.14 1.88 14.42 ;
  LAYER M3 ;
        RECT 1.58 14.12 1.86 14.44 ;
  LAYER M2 ;
        RECT 1.56 15.82 1.88 16.1 ;
  LAYER M3 ;
        RECT 1.58 15.8 1.86 16.12 ;
  LAYER M2 ;
        RECT 2.85 28.42 3.17 28.7 ;
  LAYER M3 ;
        RECT 2.87 28.4 3.15 28.72 ;
  LAYER M2 ;
        RECT 2.85 29.26 3.17 29.54 ;
  LAYER M3 ;
        RECT 2.87 29.24 3.15 29.56 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M2 ;
        RECT 2.15 12.04 3.01 12.32 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M2 ;
        RECT 2.84 22.96 4.04 23.24 ;
  LAYER M2 ;
        RECT 2.15 22.96 3.01 23.24 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.18 2.72 23.1 ;
  LAYER M2 ;
        RECT 2.42 22.96 2.74 23.24 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 22.96 2.74 23.24 ;
  LAYER M3 ;
        RECT 2.44 22.94 2.72 23.26 ;
  LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
  LAYER M3 ;
        RECT 2.44 12.02 2.72 12.34 ;
  LAYER M2 ;
        RECT 2.42 22.96 2.74 23.24 ;
  LAYER M3 ;
        RECT 2.44 22.94 2.72 23.26 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 3.865 ;
  LAYER M1 ;
        RECT 3.745 4.115 3.995 5.125 ;
  LAYER M1 ;
        RECT 3.745 6.215 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 3.865 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 3.865 ;
  LAYER M2 ;
        RECT 2.84 6.58 4.04 6.86 ;
  LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
  LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 3.865 ;
  LAYER M1 ;
        RECT 1.165 4.115 1.415 5.125 ;
  LAYER M1 ;
        RECT 1.165 6.215 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.595 0.335 1.845 3.865 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
  LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 2.84 14.14 4.04 14.42 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 1.12 14.14 2.32 14.42 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M1 ;
        RECT 3.745 18.815 3.995 22.345 ;
  LAYER M1 ;
        RECT 3.745 17.555 3.995 18.565 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 16.465 ;
  LAYER M1 ;
        RECT 3.315 18.815 3.565 22.345 ;
  LAYER M1 ;
        RECT 4.175 18.815 4.425 22.345 ;
  LAYER M2 ;
        RECT 2.84 15.82 4.04 16.1 ;
  LAYER M2 ;
        RECT 2.84 22.12 4.04 22.4 ;
  LAYER M2 ;
        RECT 2.84 17.92 4.04 18.2 ;
  LAYER M2 ;
        RECT 3.27 21.7 4.47 21.98 ;
  LAYER M1 ;
        RECT 1.165 18.815 1.415 22.345 ;
  LAYER M1 ;
        RECT 1.165 17.555 1.415 18.565 ;
  LAYER M1 ;
        RECT 1.165 15.455 1.415 16.465 ;
  LAYER M1 ;
        RECT 1.595 18.815 1.845 22.345 ;
  LAYER M1 ;
        RECT 0.735 18.815 0.985 22.345 ;
  LAYER M2 ;
        RECT 1.12 15.82 2.32 16.1 ;
  LAYER M2 ;
        RECT 1.12 22.12 2.32 22.4 ;
  LAYER M2 ;
        RECT 1.12 17.92 2.32 18.2 ;
  LAYER M2 ;
        RECT 0.69 21.7 1.89 21.98 ;
  LAYER M1 ;
        RECT 1.165 23.015 1.415 26.545 ;
  LAYER M1 ;
        RECT 1.165 26.795 1.415 27.805 ;
  LAYER M1 ;
        RECT 1.165 28.895 1.415 29.905 ;
  LAYER M1 ;
        RECT 1.595 23.015 1.845 26.545 ;
  LAYER M1 ;
        RECT 0.735 23.015 0.985 26.545 ;
  LAYER M2 ;
        RECT 1.12 29.26 2.32 29.54 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M2 ;
        RECT 1.12 27.16 2.32 27.44 ;
  LAYER M2 ;
        RECT 0.69 23.38 1.89 23.66 ;
  LAYER M1 ;
        RECT 3.745 23.015 3.995 26.545 ;
  LAYER M1 ;
        RECT 3.745 26.795 3.995 27.805 ;
  LAYER M1 ;
        RECT 3.745 28.895 3.995 29.905 ;
  LAYER M1 ;
        RECT 3.315 23.015 3.565 26.545 ;
  LAYER M1 ;
        RECT 4.175 23.015 4.425 26.545 ;
  LAYER M2 ;
        RECT 2.84 29.26 4.04 29.54 ;
  LAYER M2 ;
        RECT 2.84 22.96 4.04 23.24 ;
  LAYER M2 ;
        RECT 2.84 27.16 4.04 27.44 ;
  LAYER M2 ;
        RECT 3.27 23.38 4.47 23.66 ;
  END 
END SW
