magic
tech sky130B
magscale 1 2
timestamp 1688567721
<< metal1 >>
rect 6760 34894 21920 34910
rect 6760 34834 6770 34894
rect 6830 34834 21850 34894
rect 21910 34834 21920 34894
rect 6760 34820 21920 34834
rect 7630 34716 21280 34730
rect 7630 34656 7640 34716
rect 7700 34714 21280 34716
rect 7700 34656 21210 34714
rect 7630 34654 21210 34656
rect 21270 34654 21280 34714
rect 7630 34640 21280 34654
rect 7220 34540 21650 34550
rect 7220 34470 7230 34540
rect 7300 34538 21650 34540
rect 7300 34470 21570 34538
rect 21638 34470 21650 34538
rect 7220 34460 21650 34470
rect 280 33720 480 33920
rect 3590 33884 3690 33984
rect 13874 33570 14806 34002
rect 28206 33706 28406 33906
rect 1920 33162 1960 33202
rect 3442 32508 3542 32608
rect 4100 32236 4180 32316
rect 4400 30290 4480 30370
rect 4400 26518 4480 26598
rect 4400 18894 4480 18974
rect 6760 18902 6770 18962
rect 6830 18902 6840 18962
rect 21840 18902 21850 18962
rect 21910 18902 21920 18962
rect 13660 2666 15020 2746
rect 9860 2530 24580 2540
rect 9860 2470 9870 2530
rect 9930 2470 24510 2530
rect 24570 2470 24580 2530
rect 9860 2460 24580 2470
rect 5120 2310 19660 2320
rect 5120 2308 19590 2310
rect 5120 2248 5130 2308
rect 5190 2250 19590 2308
rect 19650 2250 19660 2310
rect 5190 2248 19660 2250
rect 5120 2240 19660 2248
rect 7000 1954 19054 2106
rect 6496 1680 6506 1740
rect 6566 1680 6576 1740
rect 5120 1316 5430 1326
rect 5120 1256 5130 1316
rect 5190 1256 5430 1316
rect 5120 1246 5430 1256
rect 13400 1246 13480 1326
rect 19580 1316 19990 1326
rect 14570 1200 14650 1280
rect 19580 1256 19590 1316
rect 19650 1256 19990 1316
rect 19580 1246 19990 1256
rect 21160 1100 21170 1160
rect 21230 1100 21240 1160
rect 7612 600 19990 752
<< via1 >>
rect 6770 34834 6830 34894
rect 21850 34834 21910 34894
rect 7640 34656 7700 34716
rect 21210 34654 21270 34714
rect 7230 34470 7300 34540
rect 21570 34470 21638 34538
rect 9870 2470 9930 2530
rect 24510 2470 24570 2530
rect 5130 2248 5190 2308
rect 19590 2250 19650 2310
rect 6506 1680 6566 1740
rect 5130 1256 5190 1316
rect 19590 1256 19650 1316
rect 21170 1100 21230 1160
<< metal2 >>
rect 6760 34894 6840 34910
rect 6760 34834 6770 34894
rect 6830 34834 6840 34894
rect 6760 18962 6840 34834
rect 21840 34894 21920 34910
rect 21840 34834 21850 34894
rect 21910 34834 21920 34894
rect 7630 34716 7710 34730
rect 7630 34656 7640 34716
rect 7700 34656 7710 34716
rect 7220 34540 7310 34550
rect 7220 34470 7230 34540
rect 7300 34470 7310 34540
rect 7220 30364 7310 34470
rect 7220 30296 7230 30364
rect 7298 30296 7310 30364
rect 7220 30286 7310 30296
rect 7630 26554 7710 34656
rect 21200 34714 21280 34730
rect 21200 34654 21210 34714
rect 21270 34654 21280 34714
rect 21200 26512 21280 34654
rect 21560 34538 21650 34550
rect 21560 34470 21570 34538
rect 21638 34470 21650 34538
rect 21560 30364 21650 34470
rect 21560 30296 21572 30364
rect 21640 30296 21650 30364
rect 21560 30286 21650 30296
rect 6760 18902 6770 18962
rect 6830 18902 6840 18962
rect 6760 18892 6840 18902
rect 21840 18962 21920 34834
rect 21840 18902 21850 18962
rect 21910 18902 21920 18962
rect 21840 18892 21920 18902
rect 9860 2530 9940 4426
rect 9860 2470 9870 2530
rect 9930 2470 9940 2530
rect 9860 2460 9940 2470
rect 24500 2530 24580 4506
rect 24500 2470 24510 2530
rect 24570 2470 24580 2530
rect 24500 2460 24580 2470
rect 5120 2308 5200 2320
rect 5120 2248 5130 2308
rect 5190 2248 5200 2308
rect 5120 1316 5200 2248
rect 19580 2310 19660 2320
rect 19580 2250 19590 2310
rect 19650 2250 19660 2310
rect 7750 1906 14270 1986
rect 6500 1740 6730 1750
rect 6500 1680 6506 1740
rect 6566 1680 6660 1740
rect 6720 1680 6730 1740
rect 6500 1670 6730 1680
rect 7750 1740 7830 1906
rect 7750 1680 7760 1740
rect 7820 1680 7830 1740
rect 7750 1670 7830 1680
rect 5120 1256 5130 1316
rect 5190 1256 5200 1316
rect 5120 1246 5200 1256
rect 19580 1316 19660 2250
rect 19580 1256 19590 1316
rect 19650 1256 19660 1316
rect 19580 1246 19660 1256
rect 20370 1160 20590 1170
rect 20370 1100 20520 1160
rect 20580 1100 20590 1160
rect 20370 1090 20590 1100
rect 20950 1160 21240 1170
rect 20950 1100 20960 1160
rect 21020 1100 21170 1160
rect 21230 1100 21240 1160
rect 20950 1090 21240 1100
rect 20370 800 20450 1090
rect 15110 720 20450 800
<< via2 >>
rect 7230 30296 7298 30364
rect 21572 30296 21640 30364
rect 6770 18902 6830 18962
rect 21850 18902 21910 18962
rect 6660 1680 6720 1740
rect 7760 1680 7820 1740
rect 20520 1100 20580 1160
rect 20960 1100 21020 1160
<< metal3 >>
rect 7220 30364 7310 30374
rect 7220 30296 7230 30364
rect 7298 30296 7310 30364
rect 7220 30286 7310 30296
rect 21560 30364 21654 30374
rect 21560 30296 21572 30364
rect 21640 30296 21654 30364
rect 21560 30286 21654 30296
rect 6760 18962 6840 18976
rect 6760 18902 6770 18962
rect 6830 18902 6840 18962
rect 6760 18892 6840 18902
rect 21840 18962 21920 18967
rect 21840 18902 21850 18962
rect 21910 18902 21920 18962
rect 21840 18897 21920 18902
rect 6646 1740 7830 1750
rect 6646 1680 6660 1740
rect 6720 1680 7760 1740
rect 7820 1680 7830 1740
rect 6646 1670 7830 1680
rect 20510 1160 21030 1170
rect 20510 1100 20520 1160
rect 20580 1100 20960 1160
rect 21020 1100 21030 1160
rect 20510 1090 21030 1100
use 6bit_dac  X1
timestamp 1688392753
transform 1 0 0 0 1 3306
box 0 -2706 14040 31000
use 6bit_dac  X2
timestamp 1688392753
transform 1 0 14640 0 1 3306
box 0 -2706 14040 31000
use sw  X3
timestamp 1687966408
transform 1 0 13400 0 1 1386
box 0 -786 1720 720
<< labels >>
flabel metal1 280 33720 480 33920 0 FreeSans 256 0 0 0 vrefh
port 2 nsew
flabel metal1 28206 33706 28406 33906 0 FreeSans 256 0 0 0 vrefl
port 3 nsew
flabel metal1 3590 33884 3690 33984 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 3442 32508 3542 32608 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 4100 32236 4180 32316 0 FreeSans 256 0 0 0 d1
port 5 nsew
flabel metal1 4400 30290 4480 30370 0 FreeSans 256 0 0 0 d2
port 6 nsew
flabel metal1 4400 26518 4480 26598 0 FreeSans 256 0 0 0 d3
port 7 nsew
flabel metal1 4400 18894 4480 18974 0 FreeSans 256 0 0 0 d4
port 8 nsew
flabel metal1 5350 1246 5430 1326 0 FreeSans 256 0 0 0 d5
port 9 nsew
flabel metal1 13400 1246 13480 1326 0 FreeSans 256 0 0 0 d6
port 10 nsew
flabel metal1 14570 1200 14650 1280 0 FreeSans 256 0 0 0 vout
port 11 nsew
flabel metal1 1920 33162 1960 33202 0 FreeSans 256 0 0 0 d0
port 4 nsew
<< end >>
