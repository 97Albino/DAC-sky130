* SPICE3 file created from 8bit_dac.ext - technology: sky130B

.subckt sky130_fd_pr__res_high_po_0p35_2NY7PZ a_n35_109# a_n165_n671# a_n35_n541#
X0 a_n35_n541# a_n35_109# a_n165_n671# sky130_fd_pr__res_high_po_0p35 l=1.09
C0 a_n35_109# a_n35_n541# 0.0153f
C1 a_n35_n541# a_n165_n671# 0.583f
C2 a_n35_109# a_n165_n671# 0.583f
.ends

.subckt sky130_fd_pr__pfet_01v8_XPYSY6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
+ VSUBS
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 w_n246_n319# a_50_n100# 0.0852f
C1 w_n246_n319# a_n108_n100# 0.0852f
C2 a_n50_n197# w_n246_n319# 0.119f
C3 a_n108_n100# a_50_n100# 0.0906f
C4 a_n50_n197# a_50_n100# 0.0163f
C5 a_n50_n197# a_n108_n100# 0.0163f
C6 a_50_n100# VSUBS 0.0558f
C7 a_n108_n100# VSUBS 0.0558f
C8 a_n50_n197# VSUBS 0.179f
C9 w_n246_n319# VSUBS 1.41f
.ends

.subckt sky130_fd_pr__nfet_01v8_ZFH27D a_50_n42# a_n210_n216# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n210_n216# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
C0 a_n50_n130# a_50_n42# 0.00909f
C1 a_n108_n42# a_50_n42# 0.0391f
C2 a_n50_n130# a_n108_n42# 0.00909f
C3 a_50_n42# a_n210_n216# 0.0801f
C4 a_n108_n42# a_n210_n216# 0.0801f
C5 a_n50_n130# a_n210_n216# 0.439f
.ends

.subckt sw vin1 vin2 vout vdd din m1_688_n494# vss m1_994_178#
XXM1 vdd din m1_994_178# vdd vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM2 vdd m1_994_178# m1_688_n494# vdd vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM3 vdd m1_994_178# vout vin1 vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM4 vdd m1_688_n494# vin2 vout vss sky130_fd_pr__pfet_01v8_XPYSY6
XXM5 m1_994_178# vss vss din sky130_fd_pr__nfet_01v8_ZFH27D
XXM6 m1_688_n494# vss vss m1_994_178# sky130_fd_pr__nfet_01v8_ZFH27D
XXM7 vout vss vin2 m1_994_178# sky130_fd_pr__nfet_01v8_ZFH27D
XXM8 vin1 vss vout m1_688_n494# sky130_fd_pr__nfet_01v8_ZFH27D
C0 m1_688_n494# vin1 0.382f
C1 m1_994_178# din 0.477f
C2 vin2 m1_994_178# 0.0836f
C3 vout vin1 -0.0258f
C4 vdd m1_994_178# 0.619f
C5 vin2 din 4.93e-19
C6 vdd din 0.31f
C7 vdd vin2 0.147f
C8 m1_994_178# m1_688_n494# 0.393f
C9 m1_994_178# vout 0.323f
C10 m1_688_n494# din 0.00777f
C11 m1_994_178# vin1 0.154f
C12 vin2 m1_688_n494# 0.247f
C13 vdd m1_688_n494# 0.182f
C14 vin2 vout -0.0571f
C15 vdd vout 0.192f
C16 vin1 din 5.3e-19
C17 vin2 vin1 0.514f
C18 vdd vin1 0.259f
C19 m1_688_n494# vout 0.374f
C20 din vss 0.855f
C21 vin1 vss 0.327f
C22 vout vss 0.355f
C23 m1_688_n494# vss 1.01f
C24 m1_994_178# vss 1.62f
C25 vin2 vss 0.759f
C26 vdd vss 4.95f
.ends

.subckt x2bit_dac X1/vin2 X3/vin2 vout vrefl X2/m1_994_178# d0 X2/m1_688_n494# X3/m1_688_n494#
+ X1/m1_688_n494# X1/m1_994_178# vdd vrefh X1/vin1 X2/vin1 d1 vss X3/vin1 X3/m1_994_178#
XXR1 vrefh vss X1/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XXR2 X1/vin2 vss X1/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XXR3 X1/vin2 vss X2/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XXR4 vrefl vss X2/vin1 sky130_fd_pr__res_high_po_0p35_2NY7PZ
XX1 X1/vin1 X1/vin2 X3/vin1 vdd d0 X1/m1_688_n494# vss X1/m1_994_178# sw
XX2 X2/vin1 vrefl X3/vin2 vdd d0 X2/m1_688_n494# vss X2/m1_994_178# sw
XX3 X3/vin1 X3/vin2 vout vdd d1 X3/m1_688_n494# vss X3/m1_994_178# sw
C0 X2/vin1 d1 7.58e-19
C1 X1/vin2 X3/m1_688_n494# 0.00743f
C2 X2/m1_688_n494# X2/vin1 0.0109f
C3 vrefh d0 1.28e-19
C4 X1/m1_688_n494# X3/vin1 0.121f
C5 vrefh X1/vin1 0.0879f
C6 X1/vin2 vrefl 0.0763f
C7 X1/vin2 vdd 0.167f
C8 X2/m1_688_n494# X3/m1_688_n494# 4.77e-21
C9 X3/vin2 X2/vin1 0.133f
C10 X1/m1_688_n494# d0 0.0316f
C11 X1/m1_994_178# X2/vin1 1.78e-19
C12 X1/m1_688_n494# X3/m1_994_178# 1.06e-19
C13 X1/m1_688_n494# X1/vin1 0.0288f
C14 vrefl d1 7.29e-21
C15 vout d1 -2.03e-24
C16 vdd d1 0.0712f
C17 vrefl X2/m1_688_n494# 0.0375f
C18 X3/vin2 X3/m1_688_n494# 0.0138f
C19 vdd X2/m1_688_n494# 0.0636f
C20 X3/vin1 d0 4.36e-19
C21 X3/vin1 X3/m1_994_178# 0.0297f
C22 X1/vin2 vrefh 0.0964f
C23 X3/vin1 X1/vin1 0.102f
C24 X2/m1_994_178# d0 0.0126f
C25 vrefl X3/vin2 0.111f
C26 X2/vin1 X3/m1_688_n494# 0.00351f
C27 vdd X3/vin2 0.118f
C28 X1/vin1 d0 0.0483f
C29 X1/vin2 X1/m1_688_n494# 0.0102f
C30 vdd X1/m1_994_178# 6.99e-19
C31 vrefl X2/vin1 0.067f
C32 vdd X2/vin1 0.234f
C33 X1/m1_688_n494# d1 2.7e-19
C34 X1/vin2 X3/vin1 0.157f
C35 X1/m1_688_n494# X2/m1_688_n494# 0.00198f
C36 X1/vin2 d0 0.177f
C37 X1/vin2 X3/m1_994_178# 0.00113f
C38 X1/vin2 X2/m1_994_178# 1.78e-19
C39 vdd X3/m1_688_n494# -0.00126f
C40 X3/vin1 d1 0.0273f
C41 X1/vin2 X1/vin1 0.167f
C42 X1/m1_688_n494# X3/vin2 7.84e-19
C43 X3/vin1 X2/m1_688_n494# 0.00207f
C44 X1/m1_994_178# X1/m1_688_n494# -5.68e-32
C45 X2/m1_688_n494# d0 0.0412f
C46 X2/m1_994_178# d1 2.92e-22
C47 X3/m1_994_178# X2/m1_688_n494# 1.15e-20
C48 vdd vrefl 0.186f
C49 X1/vin1 d1 1.51e-19
C50 X1/m1_688_n494# X2/vin1 8.88e-20
C51 X3/vin1 X3/vin2 0.0734f
C52 X1/m1_994_178# X3/vin1 0.00578f
C53 X3/vin2 d0 4.34e-19
C54 X3/m1_994_178# X3/vin2 0.0079f
C55 X1/m1_994_178# d0 0.00943f
C56 X2/m1_994_178# X3/vin2 0.00558f
C57 X1/m1_994_178# X2/m1_994_178# 0.00396f
C58 X1/m1_688_n494# X3/m1_688_n494# 4.2e-20
C59 X1/vin1 X3/vin2 2.23e-19
C60 X3/vin1 X2/vin1 0.00117f
C61 vdd vrefh 9.92e-19
C62 X1/m1_994_178# X1/vin1 0.025f
C63 X1/vin2 d1 0.00147f
C64 X2/vin1 d0 0.199f
C65 X1/vin2 X2/m1_688_n494# 8.88e-20
C66 X3/m1_994_178# X2/vin1 5.34e-19
C67 X2/m1_994_178# X2/vin1 0.0261f
C68 X3/vin1 X3/m1_688_n494# 0.0365f
C69 X1/vin1 X2/vin1 0.0689f
C70 vdd X1/m1_688_n494# 0.0775f
C71 X2/m1_688_n494# d1 0.00148f
C72 X3/m1_994_178# X3/m1_688_n494# 2.84e-32
C73 X1/vin2 X3/vin2 8.93e-19
C74 X1/vin2 X1/m1_994_178# 0.0269f
C75 X3/vin1 vrefl 0.00118f
C76 X3/vin1 vout 8.02e-19
C77 vdd X3/vin1 0.313f
C78 vrefl d0 0.0255f
C79 X3/vin2 d1 0.012f
C80 vdd d0 0.152f
C81 X1/vin2 X2/vin1 0.227f
C82 X2/m1_688_n494# X3/vin2 0.168f
C83 X1/m1_994_178# d1 2.25e-20
C84 vrefl X2/m1_994_178# 0.0258f
C85 vdd X2/m1_994_178# 6.68e-20
C86 vdd X1/vin1 0.252f
C87 d1 vss 0.545f
C88 vout vss 0.2f
C89 X3/m1_688_n494# vss 0.858f
C90 X3/m1_994_178# vss 1.15f
C91 vdd vss 15.8f
C92 d0 vss 1.67f
C93 X2/vin1 vss 1.77f
C94 X3/vin2 vss 1.43f
C95 X2/m1_688_n494# vss 0.858f
C96 X2/m1_994_178# vss 1.15f
C97 vrefl vss 3f
C98 X1/vin1 vss 2.28f
C99 X3/vin1 vss 0.845f
C100 X1/m1_688_n494# vss 0.853f
C101 X1/m1_994_178# vss 1.15f
C102 X1/vin2 vss 2.16f
C103 vrefh vss 1.34f
.ends

.subckt x3bit_dac d1 d2 X2/X1/m1_994_178# X1/X2/m1_688_n494# X2/X1/vin1 X2/X1/m1_688_n494#
+ X2/X2/vin1 X1/X3/vin2 X1/X3/vin1 X1/vout X2/X2/m1_994_178# sw_0/m1_994_178# X1/X1/m1_994_178#
+ sw_0/m1_688_n494# X1/X2/vin1 vdd X2/X3/vin2 X2/X3/vin1 X2/X2/m1_688_n494# X1/X3/m1_994_178#
+ X1/X1/m1_688_n494# X1/X3/m1_688_n494# vrefl X2/X3/m1_688_n494# vout d0 X1/X1/vin1
+ X1/X1/vin2 vrefh X2/vrefh vss X2/vout X1/X2/m1_994_178# X2/X3/m1_994_178# X2/X1/vin2
XX1 X1/X1/vin2 X1/X3/vin2 X1/vout X2/vrefh X1/X2/m1_994_178# d0 X1/X2/m1_688_n494#
+ X1/X3/m1_688_n494# X1/X1/m1_688_n494# X1/X1/m1_994_178# vdd vrefh X1/X1/vin1 X1/X2/vin1
+ d1 vss X1/X3/vin1 X1/X3/m1_994_178# x2bit_dac
XX2 X2/X1/vin2 X2/X3/vin2 X2/vout vrefl X2/X2/m1_994_178# d0 X2/X2/m1_688_n494# X2/X3/m1_688_n494#
+ X2/X1/m1_688_n494# X2/X1/m1_994_178# vdd X2/vrefh X2/X1/vin1 X2/X2/vin1 d1 vss X2/X3/vin1
+ X2/X3/m1_994_178# x2bit_dac
Xsw_0 X1/vout X2/vout vout vdd d2 sw_0/m1_688_n494# vss sw_0/m1_994_178# sw
C0 X2/X3/m1_688_n494# d1 0.0412f
C1 X2/X3/m1_994_178# d2 3.33e-19
C2 X1/X3/m1_994_178# vdd 6.99e-19
C3 vdd X2/X3/vin2 -0.00176f
C4 X1/X3/vin2 X1/vout 0.27f
C5 X2/X1/vin2 X2/X3/vin1 -0.00988f
C6 X1/X2/vin1 d1 0.0136f
C7 X2/X1/m1_688_n494# vdd -0.00178f
C8 X1/vout X2/vout 3.21e-19
C9 X1/X3/vin2 d1 0.141f
C10 X1/X2/vin1 d0 0.0624f
C11 sw_0/m1_994_178# X1/X3/m1_688_n494# 3.14e-19
C12 X1/X2/m1_994_178# vdd 5.52e-19
C13 X1/X3/m1_994_178# X1/vout 0.0106f
C14 X2/X1/vin2 d2 7.2e-20
C15 X2/vout d1 0.033f
C16 sw_0/m1_994_178# vdd 7.35e-19
C17 X1/X3/vin1 vdd 0.0299f
C18 sw_0/m1_688_n494# X2/X3/vin1 0.00874f
C19 X1/X3/m1_994_178# d1 0.00943f
C20 X2/X3/vin2 d1 9.56e-19
C21 X1/X3/m1_688_n494# vout 1.52e-19
C22 X2/X1/vin2 X2/X1/vin1 -0.0277f
C23 X1/X2/m1_994_178# X2/X1/m1_994_178# 0.00396f
C24 X2/X3/vin1 vdd -0.0214f
C25 X2/X1/m1_688_n494# d1 7.06e-20
C26 sw_0/m1_994_178# X1/vout 7.31e-20
C27 X1/X3/vin1 X1/vout 0.00864f
C28 X2/vrefh X1/X2/vin1 -0.033f
C29 X2/X1/m1_688_n494# d0 0.028f
C30 X2/vrefh X1/X3/vin2 -0.0182f
C31 vdd d2 0.0019f
C32 sw_0/m1_994_178# d1 0.00705f
C33 X1/X3/vin1 d1 0.00177f
C34 X2/X1/vin2 X2/X3/m1_994_178# -0.00113f
C35 X2/X2/vin1 d0 2.3e-20
C36 X2/X1/vin1 vdd -0.00426f
C37 X2/X3/vin1 d1 0.12f
C38 vrefh d0 1.38e-20
C39 X2/vrefh X2/X1/m1_688_n494# 8.22e-20
C40 d1 d2 0.0105f
C41 sw_0/m1_688_n494# X2/X3/m1_994_178# 3.31e-19
C42 X2/X1/m1_994_178# X2/X1/vin1 -1.07e-19
C43 X2/X3/m1_994_178# vdd 5.31e-20
C44 X2/X1/vin1 d1 0.0116f
C45 X2/X1/vin1 d0 0.219f
C46 vrefl d0 1.55e-19
C47 X2/vrefh X2/X3/vin1 2.33e-19
C48 X2/X3/m1_688_n494# X2/vout 0.0187f
C49 X1/X3/vin2 X1/X2/vin1 -0.00316f
C50 X2/X1/vin2 vdd -0.0121f
C51 X2/vrefh d2 6.65e-20
C52 X2/X3/m1_994_178# d1 0.0126f
C53 X1/X2/vin1 X1/X3/m1_994_178# -5.34e-19
C54 X1/X3/m1_688_n494# sw_0/m1_688_n494# 4.19e-20
C55 X2/vrefh X2/X1/vin1 0.164f
C56 X1/X3/vin2 X1/X3/m1_994_178# -3.03e-19
C57 sw_0/m1_688_n494# vdd 4.24e-19
C58 sw_0/m1_994_178# X2/X3/m1_688_n494# 3.38e-19
C59 X1/X3/m1_688_n494# vdd 0.0893f
C60 X2/X3/vin2 X2/vout 0.00734f
C61 X1/X3/vin2 X2/X1/m1_688_n494# 8.07e-19
C62 X2/X1/vin2 d1 0.0971f
C63 X1/X2/m1_688_n494# X2/X1/m1_688_n494# 0.00198f
C64 X2/X1/vin2 d0 0.0754f
C65 X2/X3/vin1 X2/X3/m1_688_n494# -0.00752f
C66 X2/X3/m1_688_n494# vout 9.7e-20
C67 sw_0/m1_994_178# X1/X3/vin2 0.00546f
C68 X1/vout sw_0/m1_688_n494# 1.18e-19
C69 X1/X3/vin1 X1/X3/vin2 -0.00351f
C70 X1/X3/m1_688_n494# X1/vout 0.0222f
C71 sw_0/m1_994_178# X1/X2/m1_688_n494# 2.95e-20
C72 sw_0/m1_994_178# X2/vout 1.78e-19
C73 X1/vout vdd 0.0747f
C74 sw_0/m1_688_n494# d1 0.0467f
C75 X1/X1/vin2 d0 0.0233f
C76 X1/X3/m1_688_n494# d1 0.0316f
C77 X1/X3/vin2 X2/X3/vin1 1.22e-19
C78 sw_0/m1_994_178# X1/X3/m1_994_178# 6.1e-19
C79 vdd d1 0.48f
C80 X1/X2/vin1 d2 6e-20
C81 X2/X3/vin1 X2/vout 0.221f
C82 X2/vrefh X2/X1/vin2 0.00388f
C83 vdd d0 0.0538f
C84 X1/X3/vin2 d2 0.00417f
C85 sw_0/m1_994_178# X2/X1/m1_688_n494# 2.68e-20
C86 X2/X3/vin1 X2/X3/vin2 -2.38e-19
C87 X1/X2/m1_688_n494# d2 4.64e-19
C88 X1/vout d1 0.0238f
C89 X2/vrefh X1/X1/vin2 -2.85e-19
C90 X1/X3/vin2 X2/X1/vin1 5.19e-19
C91 X1/X3/m1_994_178# d2 3.09e-19
C92 X1/X2/m1_688_n494# X2/X1/vin1 8.22e-20
C93 X2/X1/m1_994_178# d0 0.0069f
C94 sw_0/m1_994_178# X2/X3/vin1 0.00329f
C95 X2/X1/m1_688_n494# d2 6.36e-19
C96 X2/vrefh vdd 0.0108f
C97 X2/X1/m1_688_n494# X2/X1/vin1 -0.00247f
C98 X2/X1/vin2 X2/X3/m1_688_n494# -0.00743f
C99 X1/X2/m1_994_178# X2/X1/vin1 1.64e-19
C100 X2/vrefh X2/X1/m1_994_178# 1.64e-19
C101 X2/X3/m1_994_178# X2/vout 0.011f
C102 X2/X3/vin1 d2 0.00216f
C103 X2/vrefh d1 0.0738f
C104 X2/X1/vin2 X1/X3/vin2 3.94e-19
C105 X2/vrefh d0 0.818f
C106 sw_0/m1_688_n494# X2/X3/m1_688_n494# 5.55e-20
C107 vdd X2/X3/m1_688_n494# -0.00442f
C108 sw_0/m1_994_178# X2/X3/m1_994_178# 6.71e-19
C109 X2/X1/vin1 d2 9.24e-20
C110 X1/X2/vin1 X1/X3/m1_688_n494# -0.00351f
C111 X1/X3/vin2 sw_0/m1_688_n494# 0.00815f
C112 X1/X3/vin2 X1/X3/m1_688_n494# -0.00934f
C113 X1/X2/vin1 vdd -5.68e-32
C114 X1/X3/vin2 vdd 0.228f
C115 sw_0/m1_688_n494# X2/vout 1.76e-19
C116 X2/X3/vin1 X2/X3/m1_994_178# 2.84e-32
C117 X1/X2/m1_688_n494# vdd 6.35e-19
C118 X1/X3/m1_994_178# sw_0/m1_688_n494# 2.86e-19
C119 sw_0/m1_688_n494# X2/X3/vin2 3.85e-19
C120 X1/X3/m1_994_178# X1/X3/m1_688_n494# -2.84e-32
C121 vdd X2/vout 0.105f
C122 d2 vss 0.62f
C123 vout vss 0.2f
C124 sw_0/m1_688_n494# vss 0.859f
C125 sw_0/m1_994_178# vss 1.15f
C126 d1 vss 1.95f
C127 X2/vout vss 0.945f
C128 X2/X3/m1_688_n494# vss 0.949f
C129 X2/X3/m1_994_178# vss 1.15f
C130 vdd vss 35.7f
C131 d0 vss 3.81f
C132 X2/X2/vin1 vss 1.46f
C133 X2/X3/vin2 vss 1.4f
C134 X2/X2/m1_688_n494# vss 0.858f
C135 X2/X2/m1_994_178# vss 1.15f
C136 vrefl vss 2.39f
C137 X2/X1/vin1 vss 1.92f
C138 X2/X3/vin1 vss 0.868f
C139 X2/X1/m1_688_n494# vss 0.858f
C140 X2/X1/m1_994_178# vss 1.15f
C141 X2/X1/vin2 vss 1.73f
C142 X1/vout vss 0.698f
C143 X1/X3/m1_688_n494# vss 0.856f
C144 X1/X3/m1_994_178# vss 1.15f
C145 X1/X2/vin1 vss 1.46f
C146 X1/X3/vin2 vss 1.2f
C147 X1/X2/m1_688_n494# vss 0.858f
C148 X1/X2/m1_994_178# vss 1.15f
C149 X2/vrefh vss 3.29f
C150 X1/X1/vin1 vss 1.91f
C151 X1/X3/vin1 vss 0.813f
C152 X1/X1/m1_688_n494# vss 0.858f
C153 X1/X1/m1_994_178# vss 1.15f
C154 X1/X1/vin2 vss 1.73f
C155 vrefh vss 1.11f
.ends

.subckt x4bit_dac vrefh d3 X2/X2/X1/m1_688_n494# X2/X1/X2/vin1 X2/X1/X1/vin2 X2/X2/vrefh
+ X1/X1/X3/vin1 X1/X1/X3/vin2 X2/X2/X1/vin2 X1/X1/vout vrefl X1/X1/X3/m1_994_178#
+ d1 X1/X2/X3/vin2 X3/vin2 X1/X1/X3/m1_688_n494# X1/X2/X3/vin1 X3/m1_994_178# vout
+ X1/sw_0/m1_994_178# X1/X2/X1/vin1 X2/X1/X3/vin1 X2/X2/X3/vin2 X1/X2/X2/vin1 X2/sw_0/m1_688_n494#
+ X2/X2/X3/vin1 X2/X2/X2/m1_994_178# X1/X1/X2/m1_994_178# X1/X2/X3/m1_994_178# X2/X2/vout
+ X3/vin1 X2/X2/X2/m1_688_n494# X2/X2/X1/m1_994_178# X2/sw_0/m1_994_178# X2/X1/X3/m1_688_n494#
+ X2/X2/X1/vin1 X2/X1/vout X1/X2/vout X1/X1/X1/vin1 X2/X2/X2/vin1 X1/X1/X1/vin2 X3/m1_688_n494#
+ vdd X2/X1/X3/vin2 X1/X1/X2/vin1 X1/sw_0/m1_688_n494# X1/X2/vrefh X2/X2/X3/m1_994_178#
+ d0 X2/X1/X3/m1_994_178# X2/X2/X3/m1_688_n494# X1/X2/X3/m1_688_n494# X1/X1/X1/m1_994_178#
+ d2 vss X2/vrefh X1/X1/X2/m1_688_n494# X1/X1/X1/m1_688_n494# X2/X1/X1/vin1 X1/X2/X1/vin2
XX1 d1 d2 X1/X2/X1/m1_994_178# X1/X1/X2/m1_688_n494# X1/X2/X1/vin1 X1/X2/X1/m1_688_n494#
+ X1/X2/X2/vin1 X1/X1/X3/vin2 X1/X1/X3/vin1 X1/X1/vout X1/X2/X2/m1_994_178# X1/sw_0/m1_994_178#
+ X1/X1/X1/m1_994_178# X1/sw_0/m1_688_n494# X1/X1/X2/vin1 vdd X1/X2/X3/vin2 X1/X2/X3/vin1
+ X1/X2/X2/m1_688_n494# X1/X1/X3/m1_994_178# X1/X1/X1/m1_688_n494# X1/X1/X3/m1_688_n494#
+ X2/vrefh X1/X2/X3/m1_688_n494# X3/vin1 d0 X1/X1/X1/vin1 X1/X1/X1/vin2 vrefh X1/X2/vrefh
+ vss X1/X2/vout X1/X1/X2/m1_994_178# X1/X2/X3/m1_994_178# X1/X2/X1/vin2 x3bit_dac
XX2 d1 d2 X2/X2/X1/m1_994_178# X2/X1/X2/m1_688_n494# X2/X2/X1/vin1 X2/X2/X1/m1_688_n494#
+ X2/X2/X2/vin1 X2/X1/X3/vin2 X2/X1/X3/vin1 X2/X1/vout X2/X2/X2/m1_994_178# X2/sw_0/m1_994_178#
+ X2/X1/X1/m1_994_178# X2/sw_0/m1_688_n494# X2/X1/X2/vin1 vdd X2/X2/X3/vin2 X2/X2/X3/vin1
+ X2/X2/X2/m1_688_n494# X2/X1/X3/m1_994_178# X2/X1/X1/m1_688_n494# X2/X1/X3/m1_688_n494#
+ vrefl X2/X2/X3/m1_688_n494# X3/vin2 d0 X2/X1/X1/vin1 X2/X1/X1/vin2 X2/vrefh X2/X2/vrefh
+ vss X2/X2/vout X2/X1/X2/m1_994_178# X2/X2/X3/m1_994_178# X2/X2/X1/vin2 x3bit_dac
XX3 X3/vin1 X3/vin2 vout vdd d3 X3/m1_688_n494# vss X3/m1_994_178# sw
C0 X1/X2/X3/m1_688_n494# X3/vin1 8.57e-19
C1 d1 vdd 0.519f
C2 X1/X2/X2/vin1 d3 8.68e-20
C3 X1/X2/X3/vin2 d3 3.9e-19
C4 X1/X2/X2/m1_994_178# X2/X1/X1/m1_994_178# 0.00396f
C5 X1/X2/X3/m1_994_178# vdd 6.13e-19
C6 X1/X2/X2/m1_688_n494# d3 1.89e-19
C7 X1/X1/vout X1/X2/vout -0.00707f
C8 X1/X2/X2/m1_994_178# d2 0.00533f
C9 X1/sw_0/m1_688_n494# X1/sw_0/m1_994_178# -8.53e-32
C10 X2/vrefh X2/X1/X1/m1_688_n494# 8.22e-20
C11 X2/X1/X1/vin2 d3 3.99e-21
C12 X3/m1_994_178# d2 0.00703f
C13 X1/sw_0/m1_994_178# d1 -9.18e-19
C14 X2/X1/X3/vin1 vdd -0.0496f
C15 vdd d0 0.0538f
C16 X2/X1/X2/m1_688_n494# d2 0.00618f
C17 X1/X1/X3/vin2 vdd -0.00143f
C18 X1/X2/vout d2 7.51e-19
C19 X1/X2/X1/vin2 d1 -0.0945f
C20 d1 X3/m1_688_n494# 0.0363f
C21 X2/X1/X3/m1_994_178# X3/m1_994_178# 6.2e-19
C22 X3/vin1 X3/m1_994_178# -2.84e-32
C23 X2/vrefh d1 0.00744f
C24 X1/X2/vout X3/vin1 0.325f
C25 X2/X2/vout d2 4.55e-20
C26 X2/X2/vrefh X2/X1/X3/vin2 -0.00423f
C27 X1/X2/X3/m1_994_178# X3/m1_688_n494# 3.08e-19
C28 X1/X2/X1/vin2 d0 0.0233f
C29 X2/X2/vrefh d2 0.168f
C30 X2/X1/X3/vin1 X3/m1_688_n494# 0.00837f
C31 d1 X2/X1/X1/m1_688_n494# 1.25e-19
C32 X2/vrefh X2/X1/X3/vin1 2.33e-19
C33 X2/X2/X3/vin1 d2 0.0524f
C34 X2/vrefh d0 0.818f
C35 X2/X1/vout X2/sw_0/m1_994_178# -0.00141f
C36 X2/X1/X1/vin1 vdd -0.00426f
C37 X2/X1/X3/vin2 d2 0.167f
C38 X1/X1/vout d2 8.47e-20
C39 X2/X2/vout X3/vin2 0.0142f
C40 X2/X1/X1/m1_994_178# d2 0.00272f
C41 X1/sw_0/m1_688_n494# d1 -0.00449f
C42 d1 vout 0.00166f
C43 X1/X1/vout X3/vin1 0.0265f
C44 X2/X1/X1/m1_688_n494# d0 0.028f
C45 X1/X2/X3/m1_994_178# d1 0.00692f
C46 X2/X2/X3/vin1 X3/vin2 1.42e-20
C47 X2/X1/X3/m1_994_178# d2 7.31e-20
C48 X3/vin1 d2 0.00136f
C49 X1/X2/X2/vin1 vdd -0.00217f
C50 X2/X1/X3/vin2 X3/vin2 0.0533f
C51 d1 X2/X1/X3/vin1 0.122f
C52 X2/vrefh X2/X1/X1/vin1 0.164f
C53 X1/X2/X3/vin2 vdd 0.0265f
C54 X2/sw_0/m1_688_n494# d2 0.0108f
C55 X1/X1/X3/vin2 d1 -7.83e-19
C56 X2/X1/X1/vin2 X2/X1/X3/m1_688_n494# -0.00743f
C57 X2/X1/X2/vin1 d2 0.0318f
C58 X1/X2/X2/m1_688_n494# vdd 0.00105f
C59 X3/vin2 d2 0.00193f
C60 d1 X2/sw_0/m1_994_178# -9.18e-19
C61 X1/X2/X1/vin1 d2 0.0114f
C62 X2/X1/X1/vin2 vdd -0.0393f
C63 X3/vin1 X3/vin2 0.0399f
C64 X1/X2/X3/vin1 X1/X2/vout -0.00915f
C65 X2/X1/X1/m1_688_n494# X2/X1/X1/vin1 -0.00247f
C66 X1/X2/X3/m1_688_n494# vdd -0.00137f
C67 d2 d3 0.00639f
C68 X2/sw_0/m1_688_n494# X3/vin2 0.0239f
C69 X2/vrefh X1/X2/X2/vin1 -0.033f
C70 X1/X2/X3/vin2 X3/m1_688_n494# 0.00846f
C71 X2/vrefh X1/X2/X3/vin2 -0.0225f
C72 d1 X2/X1/X1/vin1 0.0116f
C73 X2/X2/X3/m1_994_178# d2 2.71e-19
C74 X2/X1/X3/m1_994_178# d3 3.17e-19
C75 X3/vin1 d3 1.11e-34
C76 X2/vrefh X2/X1/X1/vin2 0.00388f
C77 X2/X1/X3/m1_688_n494# X3/m1_994_178# 3.21e-19
C78 X1/X2/X2/m1_994_178# vdd 5.58e-19
C79 X1/X2/X3/m1_688_n494# X3/m1_688_n494# 4.41e-20
C80 vdd X3/m1_994_178# 0.00418f
C81 X2/X1/X1/vin1 d0 0.219f
C82 X1/X2/X2/m1_688_n494# X2/X1/X1/m1_688_n494# 0.00198f
C83 X1/X2/vout vdd -0.00265f
C84 X1/X2/X2/vin1 d1 -6.55e-19
C85 X1/X2/X3/vin1 d2 0.153f
C86 X1/X2/X3/vin2 d1 0.126f
C87 X1/X2/X2/vin1 X1/X2/X3/m1_994_178# -5.34e-19
C88 vdd X2/X2/vout -4.16e-19
C89 X1/X2/X2/m1_688_n494# d1 3.02e-20
C90 X1/sw_0/m1_994_178# X1/X2/vout -1.42e-32
C91 d1 X2/X1/X1/vin2 -0.00107f
C92 X1/X2/X3/vin1 X3/vin1 0.0174f
C93 X2/X1/vout X3/m1_994_178# 1.64e-19
C94 X1/X2/X1/m1_688_n494# d2 0.00416f
C95 X1/X2/X2/vin1 d0 0.0624f
C96 X2/X2/vrefh vdd -0.0152f
C97 X3/m1_994_178# X3/m1_688_n494# -1.71e-31
C98 X1/X2/X3/m1_688_n494# vout 1.64e-19
C99 X2/X2/X3/vin1 vdd -0.00249f
C100 X1/X2/X3/m1_688_n494# d1 0.026f
C101 X2/X1/X3/vin2 vdd -0.0369f
C102 X2/X1/vout X2/X2/vout -4.3e-19
C103 X2/X1/X1/vin2 X2/X1/X3/vin1 -0.0141f
C104 X1/X2/X3/m1_994_178# X1/X2/X3/m1_688_n494# 5.68e-32
C105 X2/X1/X1/vin2 d0 0.0754f
C106 vdd d2 2.08f
C107 X2/X1/X1/m1_688_n494# X3/m1_994_178# 5.36e-21
C108 X2/X1/X3/m1_994_178# X2/X1/X3/m1_688_n494# 5.68e-32
C109 X1/X1/vout X1/sw_0/m1_994_178# -0.00129f
C110 X2/X1/X3/m1_994_178# vdd 5.01e-20
C111 X3/vin1 vdd 0.101f
C112 X2/X1/X3/vin2 X2/X1/vout -0.0165f
C113 X2/X1/X3/m1_688_n494# X3/vin2 8.57e-19
C114 d1 X3/m1_994_178# 0.0135f
C115 X1/sw_0/m1_688_n494# X1/X2/vout -0.00889f
C116 X2/X1/X3/vin2 X3/m1_688_n494# 3.49e-19
C117 X1/sw_0/m1_994_178# d2 0.0176f
C118 X2/sw_0/m1_688_n494# vdd -7.94e-19
C119 X1/X2/X2/m1_688_n494# X2/X1/X1/vin1 8.22e-20
C120 X2/X1/X2/vin1 vdd -0.00219f
C121 X1/X2/X1/vin2 d2 0.226f
C122 X1/X2/X3/m1_994_178# X3/m1_994_178# 6.48e-19
C123 vdd X3/vin2 0.696f
C124 X2/X1/vout d2 0.00121f
C125 X2/vrefh X2/X1/X1/m1_994_178# 1.64e-19
C126 X2/X1/X1/vin2 X2/X1/X1/vin1 -0.0277f
C127 d2 X3/m1_688_n494# 0.00112f
C128 X1/sw_0/m1_994_178# X3/vin1 0.014f
C129 X2/vrefh d2 0.158f
C130 X2/X1/X3/vin1 X3/m1_994_178# 0.00298f
C131 X2/X1/X3/m1_994_178# X3/m1_688_n494# 2.97e-19
C132 vdd d3 0.0106f
C133 X1/X2/X3/vin2 X1/X2/X2/vin1 -0.00316f
C134 X2/X2/vrefh d1 -0.0615f
C135 X2/X1/vout X2/sw_0/m1_688_n494# -0.00792f
C136 X2/X1/X1/m1_994_178# X2/X1/X1/m1_688_n494# 1.14e-31
C137 d1 X2/X2/X3/vin1 -5.52e-19
C138 X2/X1/vout X3/vin2 0.295f
C139 X2/X1/X1/m1_688_n494# d2 0.00328f
C140 X1/X1/vout X1/sw_0/m1_688_n494# -0.00463f
C141 d1 X2/X1/X3/vin2 -0.00276f
C142 X1/sw_0/m1_688_n494# d2 0.0105f
C143 d2 vout 1.57e-20
C144 X1/X2/X2/m1_994_178# X2/X1/X1/vin1 1.64e-19
C145 X2/X2/vrefh d0 1.55e-19
C146 X1/X2/X2/vin1 X1/X2/X3/m1_688_n494# -0.00351f
C147 d1 d2 1.31f
C148 X2/vrefh d3 6.65e-20
C149 X1/X2/X3/m1_994_178# d2 2.71e-19
C150 X1/sw_0/m1_688_n494# X3/vin1 0.0362f
C151 d1 X2/X1/X3/m1_994_178# 0.0101f
C152 d1 X3/vin1 0.00179f
C153 X2/X1/X1/m1_994_178# d0 0.0069f
C154 X1/X2/X3/vin1 vdd -0.0352f
C155 d1 X2/sw_0/m1_688_n494# -0.00449f
C156 X2/X1/X3/vin1 d2 0.104f
C157 d0 d2 4.31e-19
C158 X1/X1/X3/vin2 d2 0.0586f
C159 d1 X2/X1/X2/vin1 -0.0143f
C160 d1 X3/vin2 0.00807f
C161 X2/X1/X1/m1_688_n494# d3 0.00112f
C162 X2/sw_0/m1_994_178# d2 0.0197f
C163 X1/X2/X3/vin2 X3/m1_994_178# 0.00143f
C164 X1/X2/X3/vin2 X1/X2/vout -0.00497f
C165 X1/X2/X1/m1_994_178# d2 0.00351f
C166 X1/X2/X1/vin2 X1/X2/X3/vin1 -0.00423f
C167 X1/X2/X2/m1_688_n494# X3/m1_994_178# 4.72e-20
C168 d1 d3 0.0143f
C169 X2/X1/X2/m1_994_178# d2 0.00464f
C170 X2/X1/X2/vin1 d0 2.3e-20
C171 X2/X1/X3/vin1 X3/vin2 0.0321f
C172 X2/X1/X3/m1_688_n494# vdd -0.00348f
C173 X2/X1/X1/m1_994_178# X2/X1/X1/vin1 -1.07e-19
C174 X1/X1/X3/m1_994_178# d2 7.31e-20
C175 X1/X2/X3/m1_994_178# d3 3.25e-19
C176 X2/sw_0/m1_994_178# X3/vin2 0.0147f
C177 X2/X1/X1/vin1 d2 0.0105f
C178 X1/X2/X3/m1_688_n494# X3/m1_994_178# 3.3e-19
C179 X2/X1/X3/vin1 d3 0.00192f
C180 X1/X2/vrefh d0 1.38e-20
C181 X2/X1/X3/m1_688_n494# X3/m1_688_n494# 5.25e-20
C182 X1/X2/X1/vin2 vdd -0.0262f
C183 X1/X2/X2/vin1 d2 0.0329f
C184 X2/X1/vout vdd -0.00524f
C185 X1/X2/X3/vin1 d1 -0.00179f
C186 vdd X3/m1_688_n494# 0.0122f
C187 X1/X2/X3/vin2 d2 0.0902f
C188 X2/vrefh vdd 0.00674f
C189 X1/X2/X2/m1_688_n494# d2 0.00792f
C190 X1/X2/vout X3/m1_994_178# 7.93e-20
C191 X2/X1/X1/vin1 d3 6.34e-20
C192 X2/X1/X1/vin2 d2 0.231f
C193 X1/X2/X3/vin2 X3/vin1 0.0565f
C194 X2/X1/X1/m1_688_n494# vdd -0.00178f
C195 X2/X1/X1/vin2 X2/X1/X3/m1_994_178# -0.00113f
C196 X2/X1/X3/m1_688_n494# vout 7.93e-20
C197 X1/X2/X1/vin2 X2/vrefh -2.85e-19
C198 d1 X2/X1/X3/m1_688_n494# 0.0355f
C199 d3 vss 0.621f
C200 vout vss 0.2f
C201 X3/m1_688_n494# vss 0.86f
C202 X3/m1_994_178# vss 1.15f
C203 d2 vss 2.17f
C204 X3/vin2 vss 1.83f
C205 X2/sw_0/m1_688_n494# vss 0.858f
C206 X2/sw_0/m1_994_178# vss 1.15f
C207 X2/X2/vout vss 0.868f
C208 X2/X2/X3/m1_688_n494# vss 0.858f
C209 X2/X2/X3/m1_994_178# vss 1.15f
C210 vdd vss 73.9f
C211 d0 vss 8.26f
C212 X2/X2/X2/vin1 vss 1.46f
C213 X2/X2/X3/vin2 vss 1.23f
C214 X2/X2/X2/m1_688_n494# vss 0.858f
C215 X2/X2/X2/m1_994_178# vss 1.15f
C216 vrefl vss 2.39f
C217 X2/X2/X1/vin1 vss 1.91f
C218 X2/X2/X3/vin1 vss 0.814f
C219 X2/X2/X1/m1_688_n494# vss 0.858f
C220 X2/X2/X1/m1_994_178# vss 1.15f
C221 X2/X2/X1/vin2 vss 1.73f
C222 X2/X1/vout vss 0.606f
C223 X2/X1/X3/m1_688_n494# vss 0.858f
C224 X2/X1/X3/m1_994_178# vss 1.15f
C225 X2/X1/X2/vin1 vss 1.46f
C226 X2/X1/X3/vin2 vss 1.23f
C227 X2/X1/X2/m1_688_n494# vss 0.858f
C228 X2/X1/X2/m1_994_178# vss 1.15f
C229 X2/X2/vrefh vss 3.27f
C230 X2/X1/X1/vin1 vss 1.92f
C231 X2/X1/X3/vin1 vss 0.839f
C232 X2/X1/X1/m1_688_n494# vss 0.858f
C233 X2/X1/X1/m1_994_178# vss 1.15f
C234 X2/X1/X1/vin2 vss 1.73f
C235 X3/vin1 vss 2.22f
C236 X1/sw_0/m1_688_n494# vss 0.857f
C237 X1/sw_0/m1_994_178# vss 1.15f
C238 d1 vss 3.57f
C239 X1/X2/vout vss 0.85f
C240 X1/X2/X3/m1_688_n494# vss 0.856f
C241 X1/X2/X3/m1_994_178# vss 1.15f
C242 X1/X2/X2/vin1 vss 1.46f
C243 X1/X2/X3/vin2 vss 1.21f
C244 X1/X2/X2/m1_688_n494# vss 0.858f
C245 X1/X2/X2/m1_994_178# vss 1.15f
C246 X2/vrefh vss 3.29f
C247 X1/X2/X1/vin1 vss 1.91f
C248 X1/X2/X3/vin1 vss 0.811f
C249 X1/X2/X1/m1_688_n494# vss 0.858f
C250 X1/X2/X1/m1_994_178# vss 1.15f
C251 X1/X2/X1/vin2 vss 1.73f
C252 X1/X1/vout vss 0.607f
C253 X1/X1/X3/m1_688_n494# vss 0.858f
C254 X1/X1/X3/m1_994_178# vss 1.15f
C255 X1/X1/X2/vin1 vss 1.46f
C256 X1/X1/X3/vin2 vss 1.23f
C257 X1/X1/X2/m1_688_n494# vss 0.858f
C258 X1/X1/X2/m1_994_178# vss 1.15f
C259 X1/X2/vrefh vss 3.27f
C260 X1/X1/X1/vin1 vss 1.91f
C261 X1/X1/X3/vin1 vss 0.816f
C262 X1/X1/X1/m1_688_n494# vss 0.858f
C263 X1/X1/X1/m1_994_178# vss 1.15f
C264 X1/X1/X1/vin2 vss 1.73f
C265 vrefh vss 1.11f
.ends

.subckt x5bit_dac d4 vout X1/X1/X2/X2/vin1 X1/X2/X1/X1/vin2 X2/X2/X2/vout X1/X2/X2/X1/vin1
+ X1/X2/X2/X2/vin1 X2/X1/X2/X1/vin1 X1/X1/X1/X3/vin2 X2/X1/X2/X2/vin1 X1/X1/X1/X3/vin1
+ X1/X1/X1/X3/m1_994_178# X2/X1/X2/X1/vin2 X1/X2/X1/X1/vin1 X1/X1/X1/vout X2/X2/X2/X1/vin1
+ X2/X3/m1_688_n494# X1/X2/X1/X2/vin1 X1/X2/X2/X1/vin2 X2/X1/X1/X1/vin1 X2/X2/sw_0/m1_994_178#
+ X2/X1/X1/X2/vin1 vrefh X1/X2/X1/X3/m1_688_n494# X1/X1/X2/X3/vin2 X1/X1/X1/X3/m1_688_n494#
+ X1/X1/X2/X3/vin1 X2/X1/X2/vrefh X2/X2/X1/X1/vin1 X1/X2/X2/X3/vin2 X2/X1/X1/X3/m1_688_n494#
+ X2/X2/sw_0/m1_688_n494# X2/X2/X1/X2/vin1 X1/X3/m1_688_n494# X1/X1/X2/vrefh X1/X2/X1/vout
+ X1/X2/X2/X3/vin1 X1/X1/X1/X1/vin2 X2/X2/X1/X1/vin2 X2/X1/X1/X3/vin1 X1/X1/X1/X1/m1_994_178#
+ X1/X1/X1/X1/vin1 X1/X3/vin1 X1/X1/X2/vout X2/X2/X2/X2/vin1 X1/X2/X2/X3/m1_994_178#
+ X2/X1/X1/vout X1/X1/sw_0/m1_994_178# X2/X2/X1/X3/vin2 X2/X2/X1/vout X1/X1/sw_0/m1_688_n494#
+ X2/X1/X2/X3/m1_688_n494# X2/X2/X1/X3/vin1 X2/X2/X2/X2/m1_688_n494# X2/X3/vin2 X2/X2/X1/X3/m1_994_178#
+ X2/X3/vin1 X2/X1/X1/X3/vin2 X2/X1/X1/X3/m1_994_178# X2/X2/vrefh X1/X1/X1/X1/m1_688_n494#
+ X1/X2/X2/vrefh X1/X3/vin2 X2/X2/X2/vrefh X3/vin1 X2/X2/X2/X2/m1_994_178# X1/X2/sw_0/m1_688_n494#
+ X2/X2/X1/X3/m1_688_n494# X1/X1/X2/X3/m1_994_178# X3/m1_688_n494# X1/X1/X2/X1/vin2
+ X2/X2/X2/X1/vin2 X2/X1/X2/vout X1/X2/vrefh X2/X2/X2/X3/m1_994_178# X1/X1/X2/X1/vin1
+ X2/X2/X2/X3/m1_688_n494# vdd X1/X2/X2/vout X2/X1/X1/X1/vin2 X1/X2/X2/X3/m1_688_n494#
+ d3 X1/X1/X2/X3/m1_688_n494# d1 X2/X2/X2/X3/vin2 d2 X1/X1/X1/X2/vin1 X2/X1/sw_0/m1_688_n494#
+ d0 vss X3/m1_994_178# X2/vrefh X2/X2/X2/X3/vin1 X3/vin2 vrefl
XX1 vrefh d3 X1/X2/X2/X1/m1_688_n494# X1/X2/X1/X2/vin1 X1/X2/X1/X1/vin2 X1/X2/X2/vrefh
+ X1/X1/X1/X3/vin1 X1/X1/X1/X3/vin2 X1/X2/X2/X1/vin2 X1/X1/X1/vout X2/vrefh X1/X1/X1/X3/m1_994_178#
+ d1 X1/X1/X2/X3/vin2 X1/X3/vin2 X1/X1/X1/X3/m1_688_n494# X1/X1/X2/X3/vin1 X1/X3/m1_994_178#
+ X3/vin1 X1/X1/sw_0/m1_994_178# X1/X1/X2/X1/vin1 X1/X2/X1/X3/vin1 X1/X2/X2/X3/vin2
+ X1/X1/X2/X2/vin1 X1/X2/sw_0/m1_688_n494# X1/X2/X2/X3/vin1 X1/X2/X2/X2/m1_994_178#
+ X1/X1/X1/X2/m1_994_178# X1/X1/X2/X3/m1_994_178# X1/X2/X2/vout X1/X3/vin1 X1/X2/X2/X2/m1_688_n494#
+ X1/X2/X2/X1/m1_994_178# X1/X2/sw_0/m1_994_178# X1/X2/X1/X3/m1_688_n494# X1/X2/X2/X1/vin1
+ X1/X2/X1/vout X1/X1/X2/vout X1/X1/X1/X1/vin1 X1/X2/X2/X2/vin1 X1/X1/X1/X1/vin2 X1/X3/m1_688_n494#
+ vdd X1/X2/X1/X3/vin2 X1/X1/X1/X2/vin1 X1/X1/sw_0/m1_688_n494# X1/X1/X2/vrefh X1/X2/X2/X3/m1_994_178#
+ d0 X1/X2/X1/X3/m1_994_178# X1/X2/X2/X3/m1_688_n494# X1/X1/X2/X3/m1_688_n494# X1/X1/X1/X1/m1_994_178#
+ d2 vss X1/X2/vrefh X1/X1/X1/X2/m1_688_n494# X1/X1/X1/X1/m1_688_n494# X1/X2/X1/X1/vin1
+ X1/X1/X2/X1/vin2 x4bit_dac
XX2 X2/vrefh d3 X2/X2/X2/X1/m1_688_n494# X2/X2/X1/X2/vin1 X2/X2/X1/X1/vin2 X2/X2/X2/vrefh
+ X2/X1/X1/X3/vin1 X2/X1/X1/X3/vin2 X2/X2/X2/X1/vin2 X2/X1/X1/vout vrefl X2/X1/X1/X3/m1_994_178#
+ d1 X2/X1/X2/X3/vin2 X2/X3/vin2 X2/X1/X1/X3/m1_688_n494# X2/X1/X2/X3/vin1 X2/X3/m1_994_178#
+ X3/vin2 X2/X1/sw_0/m1_994_178# X2/X1/X2/X1/vin1 X2/X2/X1/X3/vin1 X2/X2/X2/X3/vin2
+ X2/X1/X2/X2/vin1 X2/X2/sw_0/m1_688_n494# X2/X2/X2/X3/vin1 X2/X2/X2/X2/m1_994_178#
+ X2/X1/X1/X2/m1_994_178# X2/X1/X2/X3/m1_994_178# X2/X2/X2/vout X2/X3/vin1 X2/X2/X2/X2/m1_688_n494#
+ X2/X2/X2/X1/m1_994_178# X2/X2/sw_0/m1_994_178# X2/X2/X1/X3/m1_688_n494# X2/X2/X2/X1/vin1
+ X2/X2/X1/vout X2/X1/X2/vout X2/X1/X1/X1/vin1 X2/X2/X2/X2/vin1 X2/X1/X1/X1/vin2 X2/X3/m1_688_n494#
+ vdd X2/X2/X1/X3/vin2 X2/X1/X1/X2/vin1 X2/X1/sw_0/m1_688_n494# X2/X1/X2/vrefh X2/X2/X2/X3/m1_994_178#
+ d0 X2/X2/X1/X3/m1_994_178# X2/X2/X2/X3/m1_688_n494# X2/X1/X2/X3/m1_688_n494# X2/X1/X1/X1/m1_994_178#
+ d2 vss X2/X2/vrefh X2/X1/X1/X2/m1_688_n494# X2/X1/X1/X1/m1_688_n494# X2/X2/X1/X1/vin1
+ X2/X1/X2/X1/vin2 x4bit_dac
XX3 X3/vin1 X3/vin2 vout vdd d4 X3/m1_688_n494# vss X3/m1_994_178# sw
C0 X2/X1/X1/vout X3/vin2 0.0524f
C1 X1/X2/X1/X3/vin1 X3/vin1 0.0131f
C2 vdd X3/m1_688_n494# 7.42e-19
C3 X1/X2/X2/X1/m1_994_178# d2 0.00274f
C4 X1/X2/sw_0/m1_688_n494# d3 5.8e-19
C5 X1/X2/X1/vout d3 0.00226f
C6 vdd X2/X1/X1/X3/m1_994_178# 5.01e-20
C7 d2 d4 0.0103f
C8 X2/X1/X1/X2/vin1 d2 0.0309f
C9 X1/X2/X2/vrefh d0 1.38e-20
C10 X1/X2/X2/X1/vin2 d2 0.231f
C11 X2/X1/X2/X3/m1_688_n494# d3 0.00106f
C12 X2/X3/vin1 X2/X3/m1_994_178# -7.49e-19
C13 vdd d3 1.03f
C14 X2/X1/X1/X3/vin2 d2 0.106f
C15 X2/X1/X1/X3/vin1 X3/m1_994_178# 0.00298f
C16 X2/X1/X1/X1/vin2 d4 3.99e-21
C17 X2/X1/X1/X3/vin1 d2 0.104f
C18 X1/X3/m1_688_n494# X3/vin1 0.109f
C19 X1/X2/X2/X2/vin1 d0 0.0624f
C20 X2/X1/X2/vrefh X2/X1/X1/X3/vin2 -0.00423f
C21 vdd X2/X1/X1/X3/m1_688_n494# -0.00348f
C22 X2/X1/X1/X1/vin2 X2/X1/X1/X3/vin1 -0.0141f
C23 X2/X1/X1/X3/m1_994_178# d4 3.17e-19
C24 X1/X1/X2/X3/vin2 vdd -2.84e-32
C25 X1/X1/X2/X3/vin1 d3 2.1e-19
C26 X2/X3/m1_994_178# d2 -0.00133f
C27 X2/X1/X1/X3/vin2 X3/m1_688_n494# 3.49e-19
C28 X1/X3/vin1 X1/X3/m1_994_178# -0.0012f
C29 vdd X1/X2/X2/X3/m1_688_n494# -1.82e-19
C30 X1/X3/m1_688_n494# d2 -4.03e-19
C31 X2/vrefh vdd -0.00501f
C32 X2/X1/X2/vout d3 0.0232f
C33 X2/X3/vin1 X2/X3/vin2 -0.00203f
C34 X2/X3/m1_688_n494# X3/vin2 0.0523f
C35 X2/X1/X1/X3/vin1 X3/m1_688_n494# 0.00837f
C36 X1/X2/X1/X3/vin1 d3 0.0176f
C37 X1/X2/X2/X3/m1_994_178# X1/X2/X2/X2/vin1 -5.34e-19
C38 vdd X1/X2/X2/X2/m1_688_n494# 6.24e-19
C39 X2/X1/X2/X3/vin2 d3 0.0114f
C40 X2/X1/X1/X1/vin1 d2 0.0116f
C41 d1 vdd 0.355f
C42 X2/X3/vin1 d2 3.74e-20
C43 X2/vrefh X2/X1/X1/X1/m1_688_n494# 8.22e-20
C44 X2/X1/X2/X3/vin1 d3 2.1e-19
C45 vdd X2/X1/X1/vout -6.12e-19
C46 X1/X2/X2/X2/m1_688_n494# X2/X1/X1/X1/m1_688_n494# 0.00198f
C47 X2/X1/X1/X1/vin2 X2/X1/X1/X1/vin1 -0.0277f
C48 X1/X2/X2/X2/m1_994_178# X2/X1/X1/X1/m1_994_178# 0.00396f
C49 X3/vin1 d2 6.26e-19
C50 X1/X3/vin1 X1/X3/vin2 -0.00783f
C51 vdd X1/X2/X2/vout 0.165f
C52 d1 X2/X1/X1/X1/m1_688_n494# 1.25e-19
C53 X2/vrefh d4 6.65e-20
C54 X2/X2/X1/X3/vin2 d3 7.71e-19
C55 X2/X3/m1_994_178# d3 0.119f
C56 d2 X3/m1_994_178# 0.0123f
C57 X1/X3/m1_688_n494# d3 0.273f
C58 X1/X2/X2/X1/vin2 X2/vrefh -2.85e-19
C59 X1/X2/X2/X2/m1_688_n494# d4 1.89e-19
C60 vdd X1/X2/X2/X3/vin2 0.0508f
C61 X2/X1/X1/X1/m1_994_178# X2/X1/X1/X1/m1_688_n494# -2.84e-32
C62 X1/X2/X2/X3/vin1 vdd -0.0314f
C63 d1 d4 0.0105f
C64 X2/vrefh X2/X1/X1/X3/vin1 2.33e-19
C65 d1 X2/X1/X1/X2/vin1 -0.0143f
C66 X2/X1/X1/X2/m1_994_178# d2 0.00414f
C67 d1 X1/X2/X2/X1/vin2 -0.0983f
C68 X2/X1/X1/X1/vin2 d2 0.231f
C69 X1/X2/X2/X3/vin2 X2/X1/X1/X1/m1_688_n494# 8.07e-19
C70 X2/X2/X1/X3/m1_994_178# d3 0.00146f
C71 X2/X3/vin1 d3 0.374f
C72 d1 X2/X1/X1/X3/vin2 -0.00197f
C73 X2/X1/X2/vrefh d2 0.177f
C74 d1 X2/X1/X1/X3/vin1 0.117f
C75 X2/X1/X1/X3/m1_994_178# X3/m1_994_178# 6.2e-19
C76 d2 X3/m1_688_n494# 0.00172f
C77 X2/X3/vin2 d3 0.152f
C78 X3/vin1 d3 0.673f
C79 X1/X2/X2/X3/vin2 d4 0.00458f
C80 vdd X1/X2/X2/X2/vin1 -0.00217f
C81 vdd X2/X3/m1_688_n494# -0.00177f
C82 X3/m1_994_178# d3 7.7e-20
C83 X1/X2/sw_0/m1_994_178# vdd 1.48e-19
C84 d1 X2/X3/m1_994_178# -9.18e-19
C85 d1 X1/X3/m1_688_n494# -0.00449f
C86 X2/vrefh X2/X1/X1/X1/vin1 0.164f
C87 X1/X2/X2/X1/vin2 X1/X2/X2/X3/vin1 -0.00423f
C88 X2/X1/X2/X3/m1_994_178# d3 7.52e-19
C89 d2 d3 0.0129f
C90 X2/X1/X1/X1/vin2 X2/X1/X1/X3/m1_994_178# -0.00113f
C91 vdd X1/X3/vin2 0.0287f
C92 X1/X2/X1/X3/vin1 X1/X3/m1_994_178# -4.64e-19
C93 X1/X2/X2/X3/vin2 X2/X1/X1/X3/vin1 1.22e-19
C94 X1/X2/X2/X2/m1_688_n494# X2/X1/X1/X1/vin1 8.22e-20
C95 vdd X2/X2/X1/X3/vin1 -0.00133f
C96 vdd d0 0.0538f
C97 X2/X1/X1/X3/m1_688_n494# X3/m1_994_178# 3.21e-19
C98 X1/X2/X2/X3/m1_688_n494# X3/vin1 5.31e-19
C99 X2/X1/X1/X3/m1_994_178# X3/m1_688_n494# 2.97e-19
C100 X2/X1/sw_0/m1_688_n494# d2 7.88e-19
C101 d1 X2/X1/X1/X1/vin1 0.0109f
C102 d2 vout 5.3e-20
C103 d1 X2/X3/vin1 -2.22e-34
C104 X1/X2/X2/X3/m1_688_n494# X3/m1_994_178# 3.3e-19
C105 X1/X2/X2/X2/vin1 d4 8.68e-20
C106 X2/X1/X2/X3/m1_688_n494# X3/vin2 4.38e-19
C107 X2/X1/X1/X1/m1_994_178# X2/X1/X1/X1/vin1 -1.07e-19
C108 d3 X3/m1_688_n494# 0.0466f
C109 vdd X3/vin2 0.121f
C110 X2/X1/X1/X1/m1_688_n494# d0 0.028f
C111 X1/X2/X2/X2/m1_688_n494# X3/m1_994_178# 4.72e-20
C112 X2/X1/X1/X1/vin2 X2/X1/X1/X3/m1_688_n494# -0.00743f
C113 X1/X2/X2/X3/m1_994_178# vdd 6.13e-19
C114 X1/X2/X1/X3/m1_994_178# d3 0.00146f
C115 X2/vrefh d2 0.173f
C116 d1 X3/vin1 0.0079f
C117 X1/X2/X2/X2/m1_688_n494# d2 0.00583f
C118 X1/X3/m1_994_178# X1/X3/m1_688_n494# -0.00446f
C119 d1 X3/m1_994_178# 0.00705f
C120 X1/X2/X2/X3/vin2 X2/X1/X1/X1/vin1 5.19e-19
C121 X2/vrefh X2/X1/X1/X1/vin2 0.00388f
C122 X2/X1/X1/X3/m1_688_n494# X3/m1_688_n494# 5.25e-20
C123 X2/X1/X1/vout X3/m1_994_178# 1.64e-19
C124 X1/X2/X2/X1/m1_688_n494# d2 0.0033f
C125 X2/X1/X1/X2/vin1 d0 2.3e-20
C126 d1 d2 0.981f
C127 X1/X2/X2/X1/vin2 d0 0.0233f
C128 X1/X2/X2/vout X3/vin1 0.2f
C129 X2/X1/X1/X3/m1_994_178# X2/X1/X1/X3/m1_688_n494# -1.14e-31
C130 X2/X1/X1/vout d2 0.00107f
C131 X1/X1/X2/X3/m1_994_178# d3 7.52e-19
C132 X1/X2/X2/X3/m1_688_n494# X3/m1_688_n494# 4.41e-20
C133 X1/X2/X2/vout X3/m1_994_178# 7.93e-20
C134 X1/X2/X2/X3/vin2 X3/vin1 0.139f
C135 X2/X1/sw_0/m1_688_n494# d3 0.0466f
C136 X2/X1/X1/X1/m1_994_178# d2 0.00256f
C137 X2/X1/X2/vout X3/vin2 0.197f
C138 d1 X2/X1/X1/X1/vin2 -0.00132f
C139 X2/X3/m1_994_178# X2/X3/m1_688_n494# -0.00446f
C140 X2/X1/X1/X3/m1_688_n494# d3 3.07e-19
C141 X1/X2/X2/vout d2 6.28e-19
C142 X1/X2/X2/X3/vin2 X3/m1_994_178# 0.00601f
C143 d1 X2/X1/X2/vrefh -0.0667f
C144 X1/X2/X2/X3/m1_994_178# d4 3.25e-19
C145 X1/X2/X2/X3/vin1 X3/vin1 0.0131f
C146 X2/X1/X2/X3/vin2 X3/vin2 0.102f
C147 X1/X2/X1/X3/vin2 X3/vin1 0.0903f
C148 X1/X1/X2/X3/vin2 d3 0.0207f
C149 X2/X1/X1/X3/vin2 X3/vin2 0.0943f
C150 X1/X2/X2/X3/m1_688_n494# d3 3.07e-19
C151 X1/X2/X2/X3/vin2 d2 0.113f
C152 X1/X3/m1_994_178# X3/vin1 0.00755f
C153 X1/X3/vin2 X1/X3/m1_688_n494# -0.0217f
C154 X2/X2/X1/X3/m1_688_n494# d3 0.00148f
C155 d1 X3/m1_688_n494# 0.0467f
C156 X2/X2/X1/X3/vin1 X2/X3/m1_994_178# -4.64e-19
C157 X2/X1/X2/X3/vin1 X3/vin2 0.0131f
C158 X2/X1/X1/X3/vin1 X3/vin2 0.0425f
C159 X2/X1/X1/X3/m1_688_n494# vout 7.93e-20
C160 d1 X2/X1/X1/X3/m1_994_178# 0.0101f
C161 X1/X2/X2/X3/vin1 d2 0.0988f
C162 X1/X1/X2/X3/m1_688_n494# d3 7.51e-19
C163 X2/X3/vin1 X2/X3/m1_688_n494# -0.0187f
C164 X1/X1/X2/vout d3 6.06e-19
C165 X1/X2/X2/X3/vin2 X2/X1/X1/X1/vin2 3.94e-19
C166 X1/X3/m1_994_178# d2 -0.00133f
C167 X1/X2/sw_0/m1_688_n494# vdd 0.0909f
C168 X1/X2/X1/vout vdd 0.0297f
C169 X1/X2/X2/X3/m1_688_n494# vout 1.64e-19
C170 d1 d3 0.0179f
C171 X2/X3/m1_994_178# X3/vin2 0.00595f
C172 X2/X3/vin2 X2/X3/m1_688_n494# -2.84e-32
C173 X2/X1/X1/vout d3 0.00883f
C174 X2/X1/X1/X1/vin1 d0 0.219f
C175 X1/X2/X2/X3/vin2 X3/m1_688_n494# 0.00846f
C176 X1/X2/X2/X2/m1_994_178# vdd 5.58e-19
C177 X1/X2/X2/vout d3 8.47e-19
C178 X1/X2/X2/X2/vin1 d2 0.0314f
C179 X1/X3/vin2 X3/vin1 0.346f
C180 X2/X2/X1/vout d3 0.00146f
C181 d1 X2/X1/X1/X3/m1_688_n494# 0.0355f
C182 d2 X2/X3/m1_688_n494# -4.03e-19
C183 X1/X3/vin1 X1/X3/m1_688_n494# -0.00636f
C184 X1/X2/sw_0/m1_994_178# d2 0.00443f
C185 X1/X2/X2/X1/vin1 d2 0.0106f
C186 X2/X3/vin1 X3/vin2 0.345f
C187 d1 X1/X2/X2/X3/m1_688_n494# 0.026f
C188 vdd X2/X1/X1/X1/m1_688_n494# -0.00178f
C189 d1 X2/vrefh 0.00964f
C190 X1/X3/vin2 d2 1.57e-20
C191 X1/X2/X1/X3/vin2 d3 2.81e-19
C192 d0 d2 3.82e-19
C193 X1/X3/m1_994_178# d3 0.119f
C194 X2/X3/vin2 X3/vin2 0.097f
C195 X3/vin1 X3/vin2 0.0453f
C196 X2/vrefh X2/X1/X1/X1/m1_994_178# 1.64e-19
C197 vdd d4 0.00182f
C198 X1/X2/X1/X3/vin1 vdd -0.00133f
C199 vdd X2/X1/X1/X2/vin1 -0.00219f
C200 X1/X2/X2/X1/vin2 vdd -0.0272f
C201 X2/X1/X1/X1/vin2 d0 0.0754f
C202 X1/X2/X2/X3/m1_994_178# X3/m1_994_178# 6.48e-19
C203 vdd X2/X1/X1/X3/vin2 -0.034f
C204 X2/X1/X2/vrefh d0 1.55e-19
C205 d2 X3/vin2 4.24e-19
C206 X2/vrefh X1/X2/X2/X3/vin2 -0.0225f
C207 X1/X3/vin1 X3/vin1 0.095f
C208 X2/X1/X1/X1/m1_688_n494# d4 0.00112f
C209 X2/X3/m1_688_n494# d3 0.28f
C210 vdd X2/X1/X1/X3/vin1 -0.0496f
C211 X2/X1/sw_0/m1_994_178# d2 0.00659f
C212 X1/X1/X2/X3/vin2 X1/X3/m1_994_178# -6.6e-19
C213 X1/X2/X1/X3/m1_688_n494# X3/vin1 4.49e-19
C214 d1 X1/X2/X2/X3/vin2 0.138f
C215 X1/X3/vin2 d3 0.385f
C216 X2/X2/X1/X3/vin1 d3 0.0176f
C217 d1 X1/X2/X2/X3/vin1 -0.00124f
C218 X1/X2/X2/X3/m1_994_178# X3/m1_688_n494# 3.08e-19
C219 d1 X1/X3/m1_994_178# -9.18e-19
C220 X1/X2/X2/X2/vin1 X1/X2/X2/X3/m1_688_n494# -0.00351f
C221 X2/vrefh X1/X2/X2/X2/vin1 -0.033f
C222 X2/X1/X1/X3/vin1 d4 0.00192f
C223 X3/vin2 d3 0.474f
C224 vdd X2/X1/X1/X1/vin1 -0.00437f
C225 X1/X2/X2/X2/m1_994_178# X2/X1/X1/X1/vin1 1.64e-19
C226 vdd X2/X3/vin1 -0.00261f
C227 X1/X2/X1/vout X3/vin1 0.038f
C228 X1/X2/sw_0/m1_688_n494# X3/vin1 7.98e-19
C229 X2/X1/sw_0/m1_994_178# d3 7.7e-20
C230 d1 X1/X2/X2/X2/vin1 -6.55e-19
C231 d1 X2/X3/m1_688_n494# -0.00465f
C232 X2/vrefh d0 0.818f
C233 X2/X1/sw_0/m1_688_n494# X3/vin2 0.00292f
C234 X1/X3/vin1 d3 0.0863f
C235 X2/X1/X1/X1/m1_688_n494# X2/X1/X1/X1/vin1 -0.00247f
C236 vdd X3/vin1 0.56f
C237 X2/X1/X1/X3/m1_688_n494# X3/vin2 5.21e-19
C238 X1/X2/sw_0/m1_688_n494# d2 5.29e-19
C239 vdd X3/m1_994_178# 6.63e-19
C240 X1/X2/X1/X3/m1_688_n494# d3 0.00179f
C241 vdd d2 1.8f
C242 X1/X2/X2/X3/m1_994_178# X1/X2/X2/X3/m1_688_n494# 1.42e-32
C243 X1/X2/X2/X3/vin2 X1/X2/X2/X2/vin1 -0.00316f
C244 X1/X2/X2/X2/m1_994_178# d2 0.00441f
C245 X2/X1/X1/X1/vin1 d4 6.34e-20
C246 X1/X2/X2/vout X1/X3/vin2 -2.1e-19
C247 X2/X1/X1/X1/m1_994_178# d0 0.0069f
C248 X2/X1/X1/X2/m1_688_n494# d2 0.00543f
C249 X2/X1/X1/X1/m1_688_n494# X3/m1_994_178# 5.36e-21
C250 vdd X2/X1/X1/X1/vin2 -0.0393f
C251 d1 X3/vin2 0.0113f
C252 X2/X1/X2/vrefh vdd -0.0165f
C253 X2/X1/X1/X1/m1_688_n494# d2 0.00309f
C254 d1 X1/X2/X2/X3/m1_994_178# 0.00692f
C255 d4 vss 0.621f
C256 vout vss 0.2f
C257 X3/m1_688_n494# vss 0.86f
C258 X3/m1_994_178# vss 1.15f
C259 d3 vss 3.6f
C260 X3/vin2 vss 1.91f
C261 X2/X3/m1_688_n494# vss 0.858f
C262 X2/X3/m1_994_178# vss 1.15f
C263 d2 vss 4.48f
C264 X2/X3/vin2 vss 1.75f
C265 X2/X2/sw_0/m1_688_n494# vss 0.858f
C266 X2/X2/sw_0/m1_994_178# vss 1.15f
C267 X2/X2/X2/vout vss 0.868f
C268 X2/X2/X2/X3/m1_688_n494# vss 0.858f
C269 X2/X2/X2/X3/m1_994_178# vss 1.15f
C270 d0 vss 17.2f
C271 X2/X2/X2/X2/vin1 vss 1.46f
C272 X2/X2/X2/X3/vin2 vss 1.23f
C273 X2/X2/X2/X2/m1_688_n494# vss 0.858f
C274 X2/X2/X2/X2/m1_994_178# vss 1.15f
C275 vrefl vss 2.39f
C276 X2/X2/X2/X1/vin1 vss 1.91f
C277 X2/X2/X2/X3/vin1 vss 0.816f
C278 X2/X2/X2/X1/m1_688_n494# vss 0.858f
C279 X2/X2/X2/X1/m1_994_178# vss 1.15f
C280 X2/X2/X2/X1/vin2 vss 1.73f
C281 X2/X2/X1/vout vss 0.607f
C282 X2/X2/X1/X3/m1_688_n494# vss 0.858f
C283 X2/X2/X1/X3/m1_994_178# vss 1.15f
C284 X2/X2/X1/X2/vin1 vss 1.46f
C285 X2/X2/X1/X3/vin2 vss 1.23f
C286 X2/X2/X1/X2/m1_688_n494# vss 0.858f
C287 X2/X2/X1/X2/m1_994_178# vss 1.15f
C288 X2/X2/X2/vrefh vss 3.27f
C289 X2/X2/X1/X1/vin1 vss 1.91f
C290 X2/X2/X1/X3/vin1 vss 0.816f
C291 X2/X2/X1/X1/m1_688_n494# vss 0.858f
C292 X2/X2/X1/X1/m1_994_178# vss 1.15f
C293 X2/X2/X1/X1/vin2 vss 1.73f
C294 X2/X3/vin1 vss 1.49f
C295 X2/X1/sw_0/m1_688_n494# vss 0.858f
C296 X2/X1/sw_0/m1_994_178# vss 1.15f
C297 X2/X1/X2/vout vss 0.868f
C298 X2/X1/X2/X3/m1_688_n494# vss 0.858f
C299 X2/X1/X2/X3/m1_994_178# vss 1.15f
C300 X2/X1/X2/X2/vin1 vss 1.46f
C301 X2/X1/X2/X3/vin2 vss 1.23f
C302 X2/X1/X2/X2/m1_688_n494# vss 0.858f
C303 X2/X1/X2/X2/m1_994_178# vss 1.15f
C304 X2/X2/vrefh vss 3.27f
C305 X2/X1/X2/X1/vin1 vss 1.91f
C306 X2/X1/X2/X3/vin1 vss 0.816f
C307 X2/X1/X2/X1/m1_688_n494# vss 0.858f
C308 X2/X1/X2/X1/m1_994_178# vss 1.15f
C309 X2/X1/X2/X1/vin2 vss 1.73f
C310 X2/X1/X1/vout vss 0.607f
C311 X2/X1/X1/X3/m1_688_n494# vss 0.858f
C312 X2/X1/X1/X3/m1_994_178# vss 1.15f
C313 X2/X1/X1/X2/vin1 vss 1.46f
C314 X2/X1/X1/X3/vin2 vss 1.23f
C315 X2/X1/X1/X2/m1_688_n494# vss 0.858f
C316 X2/X1/X1/X2/m1_994_178# vss 1.15f
C317 X2/X1/X2/vrefh vss 3.27f
C318 X2/X1/X1/X1/vin1 vss 1.92f
C319 X2/X1/X1/X3/vin1 vss 0.839f
C320 X2/X1/X1/X1/m1_688_n494# vss 0.858f
C321 X2/X1/X1/X1/m1_994_178# vss 1.15f
C322 X2/X1/X1/X1/vin2 vss 1.73f
C323 X3/vin1 vss 1.68f
C324 X1/X3/m1_688_n494# vss 0.856f
C325 X1/X3/m1_994_178# vss 1.15f
C326 X1/X3/vin2 vss 1.75f
C327 X1/X2/sw_0/m1_688_n494# vss 0.858f
C328 X1/X2/sw_0/m1_994_178# vss 1.15f
C329 X1/X2/X2/vout vss 0.868f
C330 X1/X2/X2/X3/m1_688_n494# vss 0.856f
C331 X1/X2/X2/X3/m1_994_178# vss 1.15f
C332 vdd vss 0.152p
C333 X1/X2/X2/X2/vin1 vss 1.46f
C334 X1/X2/X2/X3/vin2 vss 1.21f
C335 X1/X2/X2/X2/m1_688_n494# vss 0.858f
C336 X1/X2/X2/X2/m1_994_178# vss 1.15f
C337 X2/vrefh vss 3.29f
C338 X1/X2/X2/X1/vin1 vss 1.91f
C339 X1/X2/X2/X3/vin1 vss 0.813f
C340 X1/X2/X2/X1/m1_688_n494# vss 0.858f
C341 X1/X2/X2/X1/m1_994_178# vss 1.15f
C342 X1/X2/X2/X1/vin2 vss 1.73f
C343 X1/X2/X1/vout vss 0.607f
C344 X1/X2/X1/X3/m1_688_n494# vss 0.858f
C345 X1/X2/X1/X3/m1_994_178# vss 1.15f
C346 X1/X2/X1/X2/vin1 vss 1.46f
C347 X1/X2/X1/X3/vin2 vss 1.23f
C348 X1/X2/X1/X2/m1_688_n494# vss 0.858f
C349 X1/X2/X1/X2/m1_994_178# vss 1.15f
C350 X1/X2/X2/vrefh vss 3.27f
C351 X1/X2/X1/X1/vin1 vss 1.91f
C352 X1/X2/X1/X3/vin1 vss 0.816f
C353 X1/X2/X1/X1/m1_688_n494# vss 0.858f
C354 X1/X2/X1/X1/m1_994_178# vss 1.15f
C355 X1/X2/X1/X1/vin2 vss 1.73f
C356 X1/X3/vin1 vss 1.49f
C357 X1/X1/sw_0/m1_688_n494# vss 0.858f
C358 X1/X1/sw_0/m1_994_178# vss 1.15f
C359 d1 vss 6.92f
C360 X1/X1/X2/vout vss 0.868f
C361 X1/X1/X2/X3/m1_688_n494# vss 0.858f
C362 X1/X1/X2/X3/m1_994_178# vss 1.15f
C363 X1/X1/X2/X2/vin1 vss 1.46f
C364 X1/X1/X2/X3/vin2 vss 1.23f
C365 X1/X1/X2/X2/m1_688_n494# vss 0.858f
C366 X1/X1/X2/X2/m1_994_178# vss 1.15f
C367 X1/X2/vrefh vss 3.27f
C368 X1/X1/X2/X1/vin1 vss 1.91f
C369 X1/X1/X2/X3/vin1 vss 0.816f
C370 X1/X1/X2/X1/m1_688_n494# vss 0.858f
C371 X1/X1/X2/X1/m1_994_178# vss 1.15f
C372 X1/X1/X2/X1/vin2 vss 1.73f
C373 X1/X1/X1/vout vss 0.607f
C374 X1/X1/X1/X3/m1_688_n494# vss 0.858f
C375 X1/X1/X1/X3/m1_994_178# vss 1.15f
C376 X1/X1/X1/X2/vin1 vss 1.46f
C377 X1/X1/X1/X3/vin2 vss 1.23f
C378 X1/X1/X1/X2/m1_688_n494# vss 0.858f
C379 X1/X1/X1/X2/m1_994_178# vss 1.15f
C380 X1/X1/X2/vrefh vss 3.27f
C381 X1/X1/X1/X1/vin1 vss 1.91f
C382 X1/X1/X1/X3/vin1 vss 0.816f
C383 X1/X1/X1/X1/m1_688_n494# vss 0.858f
C384 X1/X1/X1/X1/m1_994_178# vss 1.15f
C385 X1/X1/X1/X1/vin2 vss 1.73f
C386 vrefh vss 1.11f
.ends

.subckt x6bit_dac vrefh d5 vout X1/X1/X1/X1/X3/vin1 X2/X2/X1/sw_0/m1_688_n494# X2/X2/X1/X2/vout
+ X2/X1/X1/X2/X2/vin1 X3/vin1 X1/X1/X2/X1/X1/vin1 X1/X2/X2/X2/X1/vin2 X1/X1/X2/X1/X2/vin1
+ X1/X2/X1/X1/X1/vin1 X1/X2/X2/X2/X2/m1_688_n494# X1/X2/X2/X2/X1/vin1 X1/X2/vrefh
+ X2/X1/X2/X2/X1/vin1 X1/X1/X1/X2/vrefh X1/X2/X1/X1/X1/vin2 X1/X2/X1/X1/X2/vin1 X1/X2/X1/X2/vrefh
+ X2/X1/X2/X2/X2/vin1 X2/X2/X1/X2/X1/vin1 X2/X1/X1/X2/X1/vin2 X2/X2/X1/X2/X2/vin1
+ X1/X1/X1/X2/X3/vin2 X1/X2/X2/X1/X1/vin1 X1/X1/X2/X1/X1/vin2 X1/X1/X1/X2/X3/vin1
+ X2/X2/X1/X1/X3/m1_688_n494# X1/X2/X2/X1/X2/vin1 X2/X1/X1/X1/X2/vin1 X1/X1/X2/X1/X3/m1_688_n494#
+ X2/X2/X1/X1/X1/vin2 X2/X2/X2/X1/X3/vin2 X2/X2/X2/X2/X3/vin1 X2/X1/X2/X1/X1/vin1
+ X2/X1/X1/X1/X1/m1_994_178# X3/vin2 d4 X2/X1/X1/X1/X1/m1_688_n494# X1/X1/X3/m1_688_n494#
+ X2/X1/X2/X1/X2/vin1 X2/X2/X2/X2/X2/vin1 X2/X2/X1/X1/X1/vin1 X1/X2/X1/X1/X3/vin1
+ X2/X3/m1_688_n494# X1/X1/X3/vin1 X1/X1/X1/X2/X3/m1_994_178# X1/X2/X1/X2/X1/vin2
+ X2/X2/X1/X2/X3/m1_688_n494# X1/X1/X1/X2/X3/m1_688_n494# X2/X2/X1/X1/X2/vin1 X1/X2/X2/X2/X2/vin1
+ X2/X1/X2/X1/X1/vin2 X1/X1/X2/X2/vrefh X2/X2/X2/X1/X3/m1_994_178# X1/X2/X2/X2/vrefh
+ X2/X2/X2/X1/X3/m1_688_n494# X2/X2/X2/sw_0/m1_994_178# X2/X2/X1/X2/vrefh X1/X3/vin2
+ X2/X2/X2/sw_0/m1_688_n494# X1/X1/X1/X1/X1/m1_994_178# X2/X2/X2/X1/X1/vin1 X1/X1/X2/vrefh
+ X1/X1/X2/X1/vout X1/X1/X2/X2/X1/vin2 X2/X1/X2/vrefh X2/X2/X2/X1/X2/vin1 X1/X1/X1/X2/vout
+ X2/X2/X1/X2/X1/vin2 X2/X2/X2/X2/X3/m1_994_178# d1 X2/X2/X2/X2/X3/m1_688_n494# X2/X2/X2/X1/X3/vin1
+ X2/X1/X1/X1/X3/vin1 X3/m1_994_178# X1/X1/X1/X1/X3/m1_994_178# X1/X1/X1/X1/X1/vin2
+ X1/X1/X1/X1/X3/m1_688_n494# X2/X2/X2/X2/vout X1/X1/X3/vin2 X2/X2/X2/X2/X1/vin2 X1/X1/X2/sw_0/m1_688_n494#
+ X2/X1/X2/X2/X1/vin2 X2/X1/X2/X2/vrefh X2/X2/X2/X2/X1/vin1 X1/X1/X1/X2/X1/vin1 X2/X2/X2/X2/vrefh
+ X2/X2/X3/vin1 X2/X2/X1/X1/vout X1/X3/vin1 X1/X1/X1/X1/X1/m1_688_n494# X2/X3/vin2
+ X1/X2/X2/X1/X1/vin2 X1/X1/X1/X2/X2/vin1 X2/X2/X2/X2/X2/m1_994_178# X2/X3/vin1 X2/X2/X2/X2/X2/m1_688_n494#
+ X2/X2/X3/vin2 X1/X2/X2/vrefh X1/X2/X2/X2/X2/m1_994_178# X1/X1/X2/X2/vout X2/X2/X2/vrefh
+ d3 X1/X1/X1/X1/vout X1/X1/X2/X2/X1/vin1 X1/X3/m1_688_n494# X2/X2/vrefh X3/m1_688_n494#
+ X1/X1/X1/X1/X1/vin1 X1/X1/X1/X2/X1/vin2 X1/X1/X2/X2/X2/vin1 X1/X1/X2/X2/X3/m1_688_n494#
+ vdd X1/X2/X1/X2/X1/vin1 d2 X2/X2/X2/X1/X1/vin2 X2/X2/X2/X2/X3/vin2 X2/X2/X3/m1_688_n494#
+ X1/X1/X1/X1/X2/vin1 X1/X2/X1/X2/X2/vin1 X1/X1/X1/sw_0/m1_688_n494# X2/X1/X1/X1/X1/vin2
+ X2/X2/X2/X1/vout X1/X1/X1/X1/X3/vin2 X2/vrefh d0 vrefl vss X2/X1/X1/X2/X1/vin1 X2/X1/X1/X2/vrefh
+ X2/X1/X1/X1/X1/vin1
XX1 d4 X3/vin1 X1/X1/X1/X2/X2/vin1 X1/X1/X2/X1/X1/vin2 X1/X2/X2/X2/vout X1/X1/X2/X2/X1/vin1
+ X1/X1/X2/X2/X2/vin1 X1/X2/X1/X2/X1/vin1 X1/X1/X1/X1/X3/vin2 X1/X2/X1/X2/X2/vin1
+ X1/X1/X1/X1/X3/vin1 X1/X1/X1/X1/X3/m1_994_178# X1/X2/X1/X2/X1/vin2 X1/X1/X2/X1/X1/vin1
+ X1/X1/X1/X1/vout X1/X2/X2/X2/X1/vin1 X1/X2/X3/m1_688_n494# X1/X1/X2/X1/X2/vin1 X1/X1/X2/X2/X1/vin2
+ X1/X2/X1/X1/X1/vin1 X1/X2/X2/sw_0/m1_994_178# X1/X2/X1/X1/X2/vin1 vrefh X1/X1/X2/X1/X3/m1_688_n494#
+ X1/X1/X1/X2/X3/vin2 X1/X1/X1/X1/X3/m1_688_n494# X1/X1/X1/X2/X3/vin1 X1/X2/X1/X2/vrefh
+ X1/X2/X2/X1/X1/vin1 X1/X1/X2/X2/X3/vin2 X1/X2/X1/X1/X3/m1_688_n494# X1/X2/X2/sw_0/m1_688_n494#
+ X1/X2/X2/X1/X2/vin1 X1/X1/X3/m1_688_n494# X1/X1/X1/X2/vrefh X1/X1/X2/X1/vout X1/X1/X2/X2/X3/vin1
+ X1/X1/X1/X1/X1/vin2 X1/X2/X2/X1/X1/vin2 X1/X2/X1/X1/X3/vin1 X1/X1/X1/X1/X1/m1_994_178#
+ X1/X1/X1/X1/X1/vin1 X1/X1/X3/vin1 X1/X1/X1/X2/vout X1/X2/X2/X2/X2/vin1 X1/X1/X2/X2/X3/m1_994_178#
+ X1/X2/X1/X1/vout X1/X1/X1/sw_0/m1_994_178# X1/X2/X2/X1/X3/vin2 X1/X2/X2/X1/vout
+ X1/X1/X1/sw_0/m1_688_n494# X1/X2/X1/X2/X3/m1_688_n494# X1/X2/X2/X1/X3/vin1 X1/X2/X2/X2/X2/m1_688_n494#
+ X1/X2/X3/vin2 X1/X2/X2/X1/X3/m1_994_178# X1/X2/X3/vin1 X1/X2/X1/X1/X3/vin2 X1/X2/X1/X1/X3/m1_994_178#
+ X1/X2/X2/vrefh X1/X1/X1/X1/X1/m1_688_n494# X1/X1/X2/X2/vrefh X1/X1/X3/vin2 X1/X2/X2/X2/vrefh
+ X1/X3/vin1 X1/X2/X2/X2/X2/m1_994_178# X1/X1/X2/sw_0/m1_688_n494# X1/X2/X2/X1/X3/m1_688_n494#
+ X1/X1/X1/X2/X3/m1_994_178# X1/X3/m1_688_n494# X1/X1/X1/X2/X1/vin2 X1/X2/X2/X2/X1/vin2
+ X1/X2/X1/X2/vout X1/X1/X2/vrefh X1/X2/X2/X2/X3/m1_994_178# X1/X1/X1/X2/X1/vin1 X1/X2/X2/X2/X3/m1_688_n494#
+ vdd X1/X1/X2/X2/vout X1/X2/X1/X1/X1/vin2 X1/X1/X2/X2/X3/m1_688_n494# d3 X1/X1/X1/X2/X3/m1_688_n494#
+ d1 X1/X2/X2/X2/X3/vin2 d2 X1/X1/X1/X1/X2/vin1 X1/X2/X1/sw_0/m1_688_n494# d0 vss
+ X1/X3/m1_994_178# X1/X2/vrefh X1/X2/X2/X2/X3/vin1 X1/X3/vin2 X2/vrefh x5bit_dac
XX2 d4 X3/vin2 X2/X1/X1/X2/X2/vin1 X2/X1/X2/X1/X1/vin2 X2/X2/X2/X2/vout X2/X1/X2/X2/X1/vin1
+ X2/X1/X2/X2/X2/vin1 X2/X2/X1/X2/X1/vin1 X2/X1/X1/X1/X3/vin2 X2/X2/X1/X2/X2/vin1
+ X2/X1/X1/X1/X3/vin1 X2/X1/X1/X1/X3/m1_994_178# X2/X2/X1/X2/X1/vin2 X2/X1/X2/X1/X1/vin1
+ X2/X1/X1/X1/vout X2/X2/X2/X2/X1/vin1 X2/X2/X3/m1_688_n494# X2/X1/X2/X1/X2/vin1 X2/X1/X2/X2/X1/vin2
+ X2/X2/X1/X1/X1/vin1 X2/X2/X2/sw_0/m1_994_178# X2/X2/X1/X1/X2/vin1 X2/vrefh X2/X1/X2/X1/X3/m1_688_n494#
+ X2/X1/X1/X2/X3/vin2 X2/X1/X1/X1/X3/m1_688_n494# X2/X1/X1/X2/X3/vin1 X2/X2/X1/X2/vrefh
+ X2/X2/X2/X1/X1/vin1 X2/X1/X2/X2/X3/vin2 X2/X2/X1/X1/X3/m1_688_n494# X2/X2/X2/sw_0/m1_688_n494#
+ X2/X2/X2/X1/X2/vin1 X2/X1/X3/m1_688_n494# X2/X1/X1/X2/vrefh X2/X1/X2/X1/vout X2/X1/X2/X2/X3/vin1
+ X2/X1/X1/X1/X1/vin2 X2/X2/X2/X1/X1/vin2 X2/X2/X1/X1/X3/vin1 X2/X1/X1/X1/X1/m1_994_178#
+ X2/X1/X1/X1/X1/vin1 X2/X1/X3/vin1 X2/X1/X1/X2/vout X2/X2/X2/X2/X2/vin1 X2/X1/X2/X2/X3/m1_994_178#
+ X2/X2/X1/X1/vout X2/X1/X1/sw_0/m1_994_178# X2/X2/X2/X1/X3/vin2 X2/X2/X2/X1/vout
+ X2/X1/X1/sw_0/m1_688_n494# X2/X2/X1/X2/X3/m1_688_n494# X2/X2/X2/X1/X3/vin1 X2/X2/X2/X2/X2/m1_688_n494#
+ X2/X2/X3/vin2 X2/X2/X2/X1/X3/m1_994_178# X2/X2/X3/vin1 X2/X2/X1/X1/X3/vin2 X2/X2/X1/X1/X3/m1_994_178#
+ X2/X2/X2/vrefh X2/X1/X1/X1/X1/m1_688_n494# X2/X1/X2/X2/vrefh X2/X1/X3/vin2 X2/X2/X2/X2/vrefh
+ X2/X3/vin1 X2/X2/X2/X2/X2/m1_994_178# X2/X1/X2/sw_0/m1_688_n494# X2/X2/X2/X1/X3/m1_688_n494#
+ X2/X1/X1/X2/X3/m1_994_178# X2/X3/m1_688_n494# X2/X1/X1/X2/X1/vin2 X2/X2/X2/X2/X1/vin2
+ X2/X2/X1/X2/vout X2/X1/X2/vrefh X2/X2/X2/X2/X3/m1_994_178# X2/X1/X1/X2/X1/vin1 X2/X2/X2/X2/X3/m1_688_n494#
+ vdd X2/X1/X2/X2/vout X2/X2/X1/X1/X1/vin2 X2/X1/X2/X2/X3/m1_688_n494# d3 X2/X1/X1/X2/X3/m1_688_n494#
+ d1 X2/X2/X2/X2/X3/vin2 d2 X2/X1/X1/X1/X2/vin1 X2/X2/X1/sw_0/m1_688_n494# d0 vss
+ X2/X3/m1_994_178# X2/X2/vrefh X2/X2/X2/X2/X3/vin1 X2/X3/vin2 vrefl x5bit_dac
XX3 X3/vin1 X3/vin2 vout vdd d5 X3/m1_688_n494# vss X3/m1_994_178# sw
C0 X1/X2/X2/X1/vout X3/vin1 0.0215f
C1 X1/X1/X1/X1/X3/vin2 d2 0.00327f
C2 d1 X1/X3/m1_688_n494# -0.00429f
C3 X2/vrefh X1/X2/X2/X2/X2/vin1 -0.033f
C4 d3 d4 0.135f
C5 X1/X1/X3/vin1 d2 0.0581f
C6 d3 X2/X3/vin1 0.00305f
C7 d2 X2/X2/X2/X1/X3/m1_688_n494# 0.00123f
C8 X2/vrefh X3/vin1 0.178f
C9 X1/X1/X1/sw_0/m1_994_178# d2 0.0861f
C10 vdd X1/X2/X2/X2/X3/m1_994_178# 2.74e-19
C11 X1/X2/X2/X1/X3/vin2 X3/vin1 0.049f
C12 X2/X1/X1/X1/X1/vin2 X2/X1/X1/X1/X3/vin1 -0.00988f
C13 X1/X2/X2/X1/X3/vin1 d2 3.6e-20
C14 vdd X1/X1/X1/X2/vout -8.37e-19
C15 X2/X2/X2/sw_0/m1_688_n494# X2/X2/X2/X2/vout -1.42e-32
C16 vdd X1/X3/vin2 3.59e-19
C17 X1/X1/X1/X2/X3/vin2 d2 6.41e-19
C18 X3/vin1 X2/X1/X2/X2/X3/m1_688_n494# 8.66e-20
C19 X2/X3/m1_688_n494# X3/vin2 0.0515f
C20 vdd X2/X2/X2/X2/X3/m1_994_178# 2.74e-19
C21 X2/X2/X2/X2/vout X2/X2/X3/vin2 -2.26e-19
C22 d2 X2/X1/X1/X2/vout 0.105f
C23 X1/X3/vin1 X1/X3/m1_688_n494# -0.00223f
C24 X1/X2/X2/X2/X3/m1_688_n494# d2 0.00202f
C25 X1/X2/X1/X2/X3/m1_688_n494# X3/vin1 2.12e-19
C26 X1/X2/X2/X1/vout d2 0.0891f
C27 X1/X2/X2/X1/X3/m1_994_178# d2 0.00129f
C28 X1/X2/X1/X1/X3/m1_994_178# d4 0.00144f
C29 d3 X2/X2/X1/sw_0/m1_688_n494# 8.75e-19
C30 d2 X2/X1/X1/X2/X3/vin2 4.29e-19
C31 X1/X2/X2/X2/vout X3/vin1 0.0857f
C32 d1 X1/X2/X2/X2/X2/vin1 0.0136f
C33 X2/X1/X2/X1/vout X3/vin2 3.2e-19
C34 d3 X2/X2/X1/X1/X3/m1_688_n494# 1.6e-19
C35 d1 X3/vin1 0.046f
C36 vdd d4 0.163f
C37 vdd X2/X3/vin1 -0.00202f
C38 X1/X2/X2/X1/X3/vin2 d2 0.00316f
C39 X2/X2/X2/X2/X3/vin1 X2/X2/X3/vin2 -1.42e-20
C40 X1/X2/X2/X2/X3/vin2 X1/X2/X2/X2/X2/vin1 -0.00316f
C41 d0 X2/X1/X1/X1/X2/vin1 2.3e-20
C42 X2/X3/m1_994_178# X2/X3/m1_688_n494# -0.00318f
C43 d2 X2/X2/X2/X1/vout 0.113f
C44 X1/X2/X2/X2/X3/vin2 X3/vin1 0.049f
C45 d2 X2/X1/X1/X2/X3/vin1 0.0022f
C46 X2/vrefh X3/m1_994_178# 7.23e-19
C47 X1/X3/m1_688_n494# X3/vin1 0.0703f
C48 X2/X1/X1/X1/X1/vin2 X2/X1/X1/X1/X1/vin1 -0.0277f
C49 X1/X2/X2/X2/vout X1/X2/X3/vin2 -2.26e-19
C50 X1/X1/X3/vin1 d3 1.13e-19
C51 d0 X2/X1/X1/X1/X1/vin1 0.22f
C52 X1/X2/X1/X1/X3/m1_688_n494# d4 0.00142f
C53 X1/X1/X1/X1/vout X1/X1/X1/sw_0/m1_688_n494# -1.15e-19
C54 X1/X2/X1/sw_0/m1_688_n494# X3/vin2 2.04e-19
C55 X1/X2/X2/X2/X1/vin2 X2/vrefh -2.85e-19
C56 X3/vin1 X2/X1/X3/vin1 0.00304f
C57 d0 d5 1.37e-19
C58 d1 X1/X3/m1_994_178# -8.86e-19
C59 X1/X2/X3/m1_688_n494# X3/vin2 3.68e-19
C60 X1/X2/X3/vin1 d3 0.00118f
C61 X1/X1/X1/X1/vout d2 0.0897f
C62 X1/X3/vin1 X3/vin1 0.0837f
C63 X1/X2/X2/X2/vout d2 0.11f
C64 X1/X2/X1/X1/X3/vin2 X3/vin1 8.36e-19
C65 X2/X1/X1/X1/X1/m1_994_178# X2/X1/X1/X1/X1/m1_688_n494# -2.84e-32
C66 X1/X3/m1_994_178# X1/X3/m1_688_n494# -0.00605f
C67 X1/X1/X2/X2/X3/vin1 d4 2.08e-19
C68 d1 d2 0.0186f
C69 X1/X2/X3/vin2 X2/X1/X3/vin1 0.0604f
C70 vdd X3/m1_688_n494# -5.68e-32
C71 X1/X2/X1/X2/vout X3/vin1 3.08e-19
C72 X1/X2/X2/X2/X3/vin2 d2 8.42e-19
C73 X1/X3/vin1 X2/X3/vin2 0.273f
C74 d2 X1/X3/m1_688_n494# -3.96e-19
C75 X2/X2/X2/sw_0/m1_688_n494# X2/X2/X3/vin2 -0.00108f
C76 X2/X3/m1_994_178# X3/vin2 0.00629f
C77 d0 X3/vin2 0.0421f
C78 X1/X2/X2/X2/vrefh d0 1.38e-20
C79 vdd X1/X1/X1/X1/X3/vin2 1.47e-19
C80 vdd X1/X1/X2/X2/X3/vin2 -7.11e-33
C81 d4 X2/X3/m1_688_n494# 0.273f
C82 X2/X1/X3/m1_688_n494# X3/vin2 6.66e-19
C83 X1/X3/vin1 X1/X3/m1_994_178# -7.49e-19
C84 X2/X3/vin1 X2/X3/m1_688_n494# -0.0172f
C85 vdd X1/X1/X3/vin1 -0.00158f
C86 X2/X2/X1/X1/X3/vin1 X2/X3/m1_994_178# -4.21e-19
C87 X1/X2/X1/X1/X3/vin1 X1/X3/m1_994_178# -6.53e-19
C88 d2 X2/X1/X3/vin1 0.0605f
C89 X1/X2/X2/X2/X2/m1_994_178# d0 9.39e-20
C90 X2/vrefh X2/X1/X1/X1/X1/m1_688_n494# 4.89e-19
C91 d3 X2/X1/X2/X2/X3/m1_688_n494# 1.6e-19
C92 d0 X2/X1/X1/X1/X1/vin2 0.0754f
C93 X1/X2/X3/vin2 X3/vin1 0.0816f
C94 X1/X3/vin2 X3/vin2 3.82e-19
C95 X2/X1/X1/X1/vout X2/X1/X1/X2/vout -3.21e-19
C96 vdd X2/X1/X1/X2/vout -8.37e-19
C97 X1/X2/X1/X2/X3/m1_688_n494# d3 1.6e-19
C98 X1/X3/m1_994_178# X3/vin1 0.0057f
C99 vdd X1/X2/X2/X2/X3/m1_688_n494# -0.00154f
C100 d1 X2/X1/X1/X1/X3/m1_688_n494# 0.0358f
C101 d2 X2/X2/X2/X1/X3/vin1 6.75e-20
C102 d2 X3/vin1 0.1f
C103 X3/vin1 X2/X1/X2/sw_0/m1_688_n494# 2.24e-19
C104 vdd X2/vrefh 0.281f
C105 vdd X1/X1/X2/X2/vout 2.22e-34
C106 X2/X2/X1/X1/X3/vin2 d4 6.94e-19
C107 d2 X2/X2/X2/sw_0/m1_994_178# 0.105f
C108 d2 X2/X1/X1/X2/X3/m1_994_178# 0.00227f
C109 d4 X3/vin2 0.288f
C110 X3/vin1 X2/X1/X3/vin2 6.26e-19
C111 X2/X3/vin1 X3/vin2 1.05f
C112 d3 X1/X3/m1_688_n494# 3.43e-19
C113 vdd X2/X2/X2/X1/vout -2.57e-19
C114 d1 X2/X1/X1/X1/X3/m1_994_178# 0.0106f
C115 d1 X2/X1/X1/X1/X1/m1_688_n494# 6.3e-19
C116 d4 X2/X2/X1/X1/X3/vin1 0.0174f
C117 X1/X2/X3/vin2 d2 0.0481f
C118 X1/X2/X1/X1/vout d4 0.00145f
C119 X1/X1/X3/m1_688_n494# d3 0.00305f
C120 X1/X1/X2/X2/X3/m1_688_n494# d4 7.27e-19
C121 d3 X2/X1/X3/vin1 1.13e-19
C122 X1/X1/X1/X1/X3/vin1 d2 1.69e-19
C123 d2 X1/X3/m1_994_178# -0.00126f
C124 d3 X2/X2/X3/m1_688_n494# 0.00211f
C125 X1/X3/vin1 d3 0.0384f
C126 X1/X1/X1/sw_0/m1_688_n494# d2 0.236f
C127 d4 X2/X3/m1_994_178# 0.129f
C128 X2/X3/vin1 X2/X3/m1_994_178# -7.85e-19
C129 X2/X1/X1/X1/X1/m1_994_178# X2/X1/X1/X1/X1/vin1 -1.07e-19
C130 vdd X1/X2/X2/X2/vout -8.37e-19
C131 d1 X2/X1/X1/X1/vout 1.44e-19
C132 X1/X3/vin1 X1/X1/X3/vin2 7.11e-33
C133 vdd d1 1.13f
C134 X2/X1/X1/X2/X3/m1_688_n494# X3/vin2 2.33e-19
C135 X1/X2/X1/X2/vout d3 7.11e-33
C136 X3/vin1 X2/X1/X1/sw_0/m1_688_n494# 6.45e-19
C137 X1/X2/X2/sw_0/m1_688_n494# X3/vin2 5.84e-19
C138 X3/vin1 X2/X1/X1/X1/X3/m1_688_n494# 8.66e-20
C139 vdd X1/X2/X2/X2/X3/vin2 0.0139f
C140 d1 X2/X1/X1/X1/X3/vin2 0.00117f
C141 X2/X2/X2/X1/vout X2/X2/X2/X2/vout -3.21e-19
C142 X3/vin2 X3/m1_688_n494# 0.00463f
C143 d3 X3/vin1 0.834f
C144 X1/X3/vin2 d4 0.0958f
C145 X1/X3/vin2 X2/X3/vin1 1.22e-19
C146 d0 X2/X1/X1/X2/vrefh 1.55e-19
C147 d1 X2/X1/X1/X1/X3/vin1 0.127f
C148 X2/X1/X1/X1/vout X2/X1/X3/vin1 -2.19e-19
C149 vdd X2/X1/X3/vin1 -0.00158f
C150 X2/vrefh X2/X1/X1/X1/X1/vin1 0.0393f
C151 X1/X3/vin1 vdd 5.96e-19
C152 X1/X2/X3/vin2 d3 0.00302f
C153 d3 X2/X3/vin2 0.0437f
C154 X1/X1/X1/X2/X3/vin1 d2 0.00271f
C155 X1/X1/X1/X1/X3/m1_994_178# d2 0.00129f
C156 vdd X1/X2/X1/X1/X3/vin1 -0.00133f
C157 d0 X3/m1_688_n494# 3.19e-19
C158 X2/vrefh d5 3.62e-19
C159 X1/X2/X3/vin1 X3/vin2 4.41e-19
C160 vdd X2/X1/X2/X2/X3/vin2 -1.42e-32
C161 X1/X1/X3/vin1 X2/X2/X3/vin2 0.0604f
C162 d2 X2/X1/X1/sw_0/m1_688_n494# 0.254f
C163 X1/X1/X3/vin2 X2/X3/vin2 7.46e-20
C164 d4 X2/X3/vin1 0.0859f
C165 d2 X2/X1/X1/X1/X3/m1_688_n494# 0.00123f
C166 X2/X1/X1/X2/vout X3/vin2 0.0898f
C167 d1 X1/X2/X2/X2/X3/vin1 0.00168f
C168 d3 X2/X1/X2/sw_0/m1_688_n494# 3.43e-19
C169 X3/vin1 X2/X1/X1/X1/vout 5.53e-20
C170 vdd X1/X2/X2/X2/X2/vin1 -8.53e-32
C171 X1/X2/X2/X1/vout X3/vin2 4.93e-20
C172 X3/vin2 vout 9.83e-25
C173 d0 X2/X1/X1/X1/X1/m1_994_178# 0.00699f
C174 d1 X2/X3/m1_688_n494# -0.00429f
C175 vdd X3/vin1 0.147f
C176 X1/X1/X2/X1/X3/m1_688_n494# d3 1.6e-19
C177 X2/X1/X1/X2/X3/vin2 X3/vin2 0.0523f
C178 d3 X2/X1/X3/vin2 0.00178f
C179 X2/vrefh X3/vin2 0.15f
C180 d2 X2/X1/X1/X1/X3/m1_994_178# 0.00213f
C181 d4 X2/X2/X1/X1/X3/m1_994_178# 0.0013f
C182 X2/X1/X1/X2/X3/vin1 X3/vin2 0.00836f
C183 vdd X1/X2/X3/vin2 -2.37e-19
C184 vdd X2/X3/vin2 4.3e-19
C185 X1/X2/X1/X1/X3/m1_688_n494# X3/vin1 2.12e-19
C186 X1/X2/X2/X2/X2/m1_994_178# X2/vrefh 9.79e-19
C187 X2/X1/X2/X2/X3/m1_688_n494# X3/vin2 2.33e-19
C188 X2/X2/X2/X1/vout X2/X2/X2/sw_0/m1_688_n494# -1.15e-19
C189 d0 vout -1e-23
C190 X1/X1/X1/X1/X3/vin1 vdd 0.00759f
C191 d4 X2/X2/X1/X1/X3/m1_688_n494# 0.0013f
C192 X2/vrefh X2/X1/X1/X1/X1/vin2 -3.82e-19
C193 X3/vin1 X2/X1/X2/X1/X3/m1_688_n494# 8.66e-20
C194 d2 X2/X2/X2/X2/X3/m1_688_n494# 0.00138f
C195 X2/vrefh d0 4.64f
C196 X1/X2/X2/X2/X2/m1_688_n494# d0 4.7e-20
C197 X1/X2/X2/X2/X3/m1_994_178# X1/X2/X2/X2/X3/m1_688_n494# 5.68e-32
C198 d2 X2/X1/X1/X1/vout 0.114f
C199 vdd d2 0.427f
C200 X1/X1/X2/X2/X3/vin2 d4 0.0219f
C201 d2 X2/X1/X1/sw_0/m1_994_178# 0.106f
C202 X1/X2/X2/X2/vout X3/vin2 1.5e-19
C203 d1 X3/vin2 0.0461f
C204 d2 X2/X1/X1/X1/X3/vin2 0.00536f
C205 X1/X2/X2/X2/X3/vin1 X3/vin1 0.00789f
C206 X3/vin1 X2/X3/m1_688_n494# 5.87e-20
C207 X1/X3/m1_688_n494# X3/vin2 6.58e-20
C208 X2/X1/X1/X1/X3/m1_994_178# X2/X1/X1/X1/X3/m1_688_n494# -1.14e-31
C209 d2 X2/X1/X1/X1/X3/vin1 3e-19
C210 X1/X1/X3/vin2 d3 0.00413f
C211 X1/X1/X2/X2/X3/m1_994_178# d4 7.44e-19
C212 X1/X2/X2/X2/X3/vin1 X1/X2/X3/vin2 -1.42e-20
C213 d1 X2/X1/X1/X1/X1/vin2 0.0778f
C214 X2/X1/X2/X2/vout X3/vin2 3.38e-19
C215 X2/X1/X3/vin1 X3/vin2 0.0361f
C216 d3 X2/X2/X1/X2/X3/m1_688_n494# 1.6e-19
C217 d1 X2/X3/m1_994_178# -6.71e-19
C218 X1/X1/X1/X2/X3/m1_994_178# d2 0.00333f
C219 d4 X2/X2/X1/X1/vout 0.00132f
C220 X1/X3/vin1 X3/vin2 7.53e-21
C221 X1/X1/X1/X1/X3/m1_994_178# vdd 3.24e-19
C222 d2 X2/X2/X2/X2/vout 0.107f
C223 X2/X1/X1/X1/vout X2/X1/X1/sw_0/m1_688_n494# -1.15e-19
C224 X2/X1/X2/X2/X3/vin2 X3/vin2 0.0011f
C225 X1/X1/X1/X1/vout X1/X1/X1/X2/vout -3.21e-19
C226 X1/X1/X2/X2/vout d4 6.02e-19
C227 d1 X1/X2/X2/X2/X3/m1_994_178# 0.00733f
C228 X1/X2/X2/X2/X3/vin1 d2 0.00319f
C229 vdd X2/X1/X1/X1/X3/m1_688_n494# -0.00334f
C230 d2 X2/X2/X2/X2/X3/vin2 5.81e-19
C231 X1/X1/X1/X1/X3/m1_688_n494# d2 7.51e-19
C232 X1/X3/vin1 X2/X2/X3/vin2 0.00719f
C233 d2 X2/X3/m1_688_n494# -2.59e-19
C234 vdd d3 0.0118f
C235 X1/X2/X1/sw_0/m1_688_n494# X3/vin1 3.28e-19
C236 d4 X2/X1/X2/X2/X3/m1_688_n494# 8.66e-19
C237 X2/X1/X3/vin1 X2/X1/X3/m1_688_n494# 2.84e-32
C238 d2 X2/X2/X2/X2/X3/vin1 0.00254f
C239 X3/vin1 X3/vin2 2.73f
C240 X1/X1/X3/vin2 vdd -8.88e-34
C241 X1/X2/X3/m1_688_n494# X3/vin1 6.09e-19
C242 X1/X3/vin2 X1/X3/m1_688_n494# -0.03f
C243 vdd X2/X1/X1/X1/X3/m1_994_178# 3.24e-19
C244 X2/X1/X2/X2/X3/vin2 X2/X3/m1_994_178# -8.37e-19
C245 d2 X2/X2/X2/X1/X3/vin2 0.00524f
C246 vdd X2/X1/X1/X1/X1/m1_688_n494# -0.00178f
C247 X1/X2/X2/X1/vout X1/X2/X2/sw_0/m1_688_n494# -1.15e-19
C248 X1/X2/X1/X1/vout X3/vin1 2.91e-19
C249 X1/X2/X1/X1/X3/m1_688_n494# d3 1.6e-19
C250 d3 X2/X2/X1/X2/vout 3.55e-33
C251 X1/X2/X3/vin2 X3/vin2 0.00254f
C252 X2/X3/vin2 X3/vin2 0.0982f
C253 X1/X1/X2/sw_0/m1_688_n494# d3 3.43e-19
C254 d3 X2/X1/X2/X1/X3/m1_688_n494# 1.6e-19
C255 X1/X2/X3/vin2 X1/X2/X3/m1_688_n494# 2.84e-32
C256 d1 d4 0.0167f
C257 X1/X3/vin1 X1/X3/vin2 -0.00705f
C258 X1/X2/X2/X2/X2/vin1 d0 0.0624f
C259 X2/vrefh X3/m1_688_n494# 7.3e-19
C260 d0 X3/vin1 0.0436f
C261 vdd X2/X2/X2/X2/X3/m1_688_n494# 1.37e-19
C262 X1/X3/m1_688_n494# d4 0.249f
C263 vdd X2/X1/X1/X1/vout -2.57e-19
C264 X3/vin1 X2/X1/X3/m1_688_n494# 3.93e-19
C265 X1/X2/X2/X2/X3/m1_994_178# X1/X2/X2/X2/X2/vin1 -5.34e-19
C266 d2 X2/X2/X2/X1/X3/m1_994_178# 0.00213f
C267 d2 X3/vin2 0.1f
C268 X2/X1/X2/sw_0/m1_688_n494# X3/vin2 3.67e-19
C269 vdd X2/X1/X1/X1/X3/vin2 -0.00178f
C270 X2/vrefh X2/X1/X1/X1/X1/m1_994_178# 9.79e-19
C271 d4 X2/X1/X2/X2/vout 6.95e-19
C272 X2/X1/X3/vin2 X3/vin2 0.039f
C273 d2 X2/X2/X2/sw_0/m1_688_n494# 0.254f
C274 d3 X2/X3/m1_688_n494# 3.43e-19
C275 X1/X3/vin2 X3/vin1 0.964f
C276 X1/X3/vin1 d4 0.0842f
C277 X1/X2/X1/X1/X3/vin2 d4 4.77e-19
C278 X1/X2/X1/X1/X3/vin1 d4 0.0186f
C279 X1/X2/X2/sw_0/m1_688_n494# X1/X2/X2/X2/vout -1.69e-19
C280 vdd X2/X1/X1/X1/X3/vin1 -0.0131f
C281 d2 X2/X2/X3/vin2 0.0665f
C282 d4 X2/X1/X2/X2/X3/vin2 0.0218f
C283 d2 X2/X3/m1_994_178# -0.00102f
C284 d4 X2/X1/X2/X2/X3/vin1 2.52e-19
C285 X1/X1/X1/X1/vout X1/X1/X3/vin1 -2.19e-19
C286 X1/X2/X2/sw_0/m1_994_178# d2 0.0861f
C287 X2/X1/X1/X1/X1/m1_688_n494# X2/X1/X1/X1/X1/vin1 -0.00247f
C288 vdd X2/X2/X2/X2/vout -8.37e-19
C289 d0 X3/m1_994_178# 2.73e-19
C290 X1/X1/X1/X2/vout X1/X1/X1/sw_0/m1_688_n494# -1.69e-19
C291 X1/X3/m1_994_178# X1/X3/vin2 -1.42e-32
C292 X1/X2/X2/X2/X3/m1_994_178# d2 0.00333f
C293 X3/vin1 d4 0.286f
C294 X2/vrefh X1/X2/X2/X2/X2/m1_688_n494# 4.89e-19
C295 X3/vin1 X2/X3/vin1 3.45e-19
C296 X2/X1/X1/sw_0/m1_688_n494# X3/vin2 0.00111f
C297 X1/X1/X1/X2/vout d2 0.11f
C298 X2/X1/X1/X1/X3/m1_688_n494# X3/vin2 2.33e-19
C299 vdd X2/X2/X2/X2/X3/vin2 0.0273f
C300 X1/X1/X1/X1/X3/m1_688_n494# vdd 1.62e-19
C301 vdd X2/X3/m1_688_n494# -0.00177f
C302 X1/X2/X2/X2/X1/vin2 d0 0.0233f
C303 X1/X2/X1/sw_0/m1_688_n494# d3 3.43e-19
C304 d2 X2/X2/X2/X2/X3/m1_994_178# 0.00233f
C305 d3 X2/X2/X3/vin1 0.00118f
C306 d3 X3/vin2 0.77f
C307 d4 X2/X3/vin2 0.0986f
C308 X1/X3/vin2 X2/X1/X3/vin2 7.46e-20
C309 X1/X2/X3/vin2 X2/X3/vin1 7.46e-20
C310 X2/X3/vin1 X2/X3/vin2 -2.4e-19
C311 X1/X2/X3/m1_688_n494# d3 0.00211f
C312 vdd X2/X1/X1/X1/X1/vin1 -0.00426f
C313 X1/X3/m1_994_178# d4 0.128f
C314 X1/X2/X2/X1/vout X1/X2/X2/X2/vout -3.21e-19
C315 vdd X2/X2/X2/X1/X3/vin2 -1.62e-19
C316 d1 X1/X2/X2/X2/X3/m1_688_n494# 0.0262f
C317 X1/X2/X1/X1/vout d3 3.55e-33
C318 X1/X1/X2/X2/X3/m1_688_n494# d3 1.6e-19
C319 X1/X1/X1/X2/X3/m1_688_n494# d2 0.00202f
C320 X2/X1/X1/X1/X1/vin2 X2/X1/X1/X1/X3/m1_688_n494# -0.00743f
C321 d3 X2/X2/X3/vin2 0.00583f
C322 X3/vin1 X2/X1/X1/X2/X3/m1_688_n494# 8.66e-20
C323 d2 d4 0.0119f
C324 X1/X2/X2/sw_0/m1_688_n494# X3/vin1 9.8e-19
C325 d1 X2/vrefh 0.062f
C326 X1/X2/X2/X1/X3/m1_688_n494# X3/vin1 2.12e-19
C327 X2/X1/X3/vin2 X2/X3/vin1 -1.42e-32
C328 X2/vrefh X1/X2/X2/X2/X3/vin2 -0.0116f
C329 d3 X2/X1/X3/m1_688_n494# 0.00305f
C330 X2/X1/X1/X1/X1/vin2 X2/X1/X1/X1/X3/m1_994_178# -0.00113f
C331 X1/X2/X2/sw_0/m1_688_n494# X1/X2/X3/vin2 -0.00108f
C332 X2/X1/X1/X1/vout X3/vin2 0.033f
C333 d0 X2/X1/X1/X1/X1/m1_688_n494# 0.0281f
C334 vdd X3/vin2 0.157f
C335 X1/X3/vin2 d3 0.00989f
C336 X2/X1/X1/X1/X3/vin2 X3/vin2 0.0523f
C337 X1/X2/X2/X1/X3/vin1 X3/vin1 0.00789f
C338 vdd X2/X2/X1/X1/X3/vin1 -0.00133f
C339 vdd X2/X2/X2/sw_0/m1_688_n494# -1.42e-32
C340 X1/X2/X3/vin1 X3/vin1 7.18e-19
C341 d2 X2/X1/X1/X2/X3/m1_688_n494# 0.00138f
C342 d1 X1/X2/X2/X2/vout 5.72e-20
C343 X1/X2/X2/sw_0/m1_688_n494# d2 0.236f
C344 vdd X2/X2/X3/vin2 -4.43e-19
C345 X2/X1/X1/X1/X3/vin1 X3/vin2 0.00836f
C346 X1/X1/X2/X2/X3/vin2 X1/X3/m1_994_178# -9.61e-19
C347 X1/X2/X2/X1/X3/m1_688_n494# d2 7.51e-19
C348 X1/X2/X2/X2/X2/vin1 X1/X2/X2/X2/X3/m1_688_n494# -0.00351f
C349 vdd X2/X1/X1/X1/X1/vin2 -0.0121f
C350 X3/vin1 X2/X1/X1/X2/vout 1.71e-19
C351 d4 X2/X1/X2/X2/X3/m1_994_178# 8.64e-19
C352 X1/X2/X2/X2/X3/m1_688_n494# X3/vin1 2.12e-19
C353 X1/X1/X3/vin1 X1/X1/X1/sw_0/m1_688_n494# -0.00197f
C354 vdd d0 0.311f
C355 d1 X1/X2/X2/X2/X3/vin2 0.201f
C356 X2/X1/X2/X1/X3/m1_688_n494# X3/vin2 2.33e-19
C357 d5 vss 0.613f
C358 vout vss 0.2f
C359 X3/m1_688_n494# vss 0.861f
C360 X3/m1_994_178# vss 1.15f
C361 X3/vin2 vss 1.98f
C362 X2/X3/m1_688_n494# vss 0.858f
C363 X2/X3/m1_994_178# vss 1.15f
C364 X2/X3/vin2 vss 1.85f
C365 X2/X2/X3/m1_688_n494# vss 0.858f
C366 X2/X2/X3/m1_994_178# vss 1.15f
C367 X2/X2/X3/vin2 vss 1.75f
C368 X2/X2/X2/sw_0/m1_688_n494# vss 0.858f
C369 X2/X2/X2/sw_0/m1_994_178# vss 1.15f
C370 X2/X2/X2/X2/vout vss 0.868f
C371 X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C372 X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C373 X2/X2/X2/X2/X2/vin1 vss 1.46f
C374 X2/X2/X2/X2/X3/vin2 vss 1.23f
C375 X2/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C376 X2/X2/X2/X2/X2/m1_994_178# vss 1.15f
C377 vrefl vss 2.39f
C378 X2/X2/X2/X2/X1/vin1 vss 1.91f
C379 X2/X2/X2/X2/X3/vin1 vss 0.816f
C380 X2/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C381 X2/X2/X2/X2/X1/m1_994_178# vss 1.15f
C382 X2/X2/X2/X2/X1/vin2 vss 1.73f
C383 X2/X2/X2/X1/vout vss 0.607f
C384 X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C385 X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C386 X2/X2/X2/X1/X2/vin1 vss 1.46f
C387 X2/X2/X2/X1/X3/vin2 vss 1.23f
C388 X2/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C389 X2/X2/X2/X1/X2/m1_994_178# vss 1.15f
C390 X2/X2/X2/X2/vrefh vss 3.27f
C391 X2/X2/X2/X1/X1/vin1 vss 1.91f
C392 X2/X2/X2/X1/X3/vin1 vss 0.816f
C393 X2/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C394 X2/X2/X2/X1/X1/m1_994_178# vss 1.15f
C395 X2/X2/X2/X1/X1/vin2 vss 1.73f
C396 X2/X2/X3/vin1 vss 1.49f
C397 X2/X2/X1/sw_0/m1_688_n494# vss 0.858f
C398 X2/X2/X1/sw_0/m1_994_178# vss 1.15f
C399 X2/X2/X1/X2/vout vss 0.868f
C400 X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C401 X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C402 X2/X2/X1/X2/X2/vin1 vss 1.46f
C403 X2/X2/X1/X2/X3/vin2 vss 1.23f
C404 X2/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C405 X2/X2/X1/X2/X2/m1_994_178# vss 1.15f
C406 X2/X2/X2/vrefh vss 3.27f
C407 X2/X2/X1/X2/X1/vin1 vss 1.91f
C408 X2/X2/X1/X2/X3/vin1 vss 0.816f
C409 X2/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C410 X2/X2/X1/X2/X1/m1_994_178# vss 1.15f
C411 X2/X2/X1/X2/X1/vin2 vss 1.73f
C412 X2/X2/X1/X1/vout vss 0.607f
C413 X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C414 X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C415 X2/X2/X1/X1/X2/vin1 vss 1.46f
C416 X2/X2/X1/X1/X3/vin2 vss 1.23f
C417 X2/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C418 X2/X2/X1/X1/X2/m1_994_178# vss 1.15f
C419 X2/X2/X1/X2/vrefh vss 3.27f
C420 X2/X2/X1/X1/X1/vin1 vss 1.91f
C421 X2/X2/X1/X1/X3/vin1 vss 0.816f
C422 X2/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C423 X2/X2/X1/X1/X1/m1_994_178# vss 1.15f
C424 X2/X2/X1/X1/X1/vin2 vss 1.73f
C425 X2/X3/vin1 vss 1.6f
C426 X2/X1/X3/m1_688_n494# vss 0.858f
C427 X2/X1/X3/m1_994_178# vss 1.15f
C428 X2/X1/X3/vin2 vss 1.75f
C429 X2/X1/X2/sw_0/m1_688_n494# vss 0.858f
C430 X2/X1/X2/sw_0/m1_994_178# vss 1.15f
C431 X2/X1/X2/X2/vout vss 0.868f
C432 X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C433 X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C434 X2/X1/X2/X2/X2/vin1 vss 1.46f
C435 X2/X1/X2/X2/X3/vin2 vss 1.23f
C436 X2/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C437 X2/X1/X2/X2/X2/m1_994_178# vss 1.15f
C438 X2/X2/vrefh vss 3.27f
C439 X2/X1/X2/X2/X1/vin1 vss 1.91f
C440 X2/X1/X2/X2/X3/vin1 vss 0.816f
C441 X2/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C442 X2/X1/X2/X2/X1/m1_994_178# vss 1.15f
C443 X2/X1/X2/X2/X1/vin2 vss 1.73f
C444 X2/X1/X2/X1/vout vss 0.607f
C445 X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C446 X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C447 X2/X1/X2/X1/X2/vin1 vss 1.46f
C448 X2/X1/X2/X1/X3/vin2 vss 1.23f
C449 X2/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C450 X2/X1/X2/X1/X2/m1_994_178# vss 1.15f
C451 X2/X1/X2/X2/vrefh vss 3.27f
C452 X2/X1/X2/X1/X1/vin1 vss 1.91f
C453 X2/X1/X2/X1/X3/vin1 vss 0.816f
C454 X2/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C455 X2/X1/X2/X1/X1/m1_994_178# vss 1.15f
C456 X2/X1/X2/X1/X1/vin2 vss 1.73f
C457 X2/X1/X3/vin1 vss 1.49f
C458 X2/X1/X1/sw_0/m1_688_n494# vss 0.858f
C459 X2/X1/X1/sw_0/m1_994_178# vss 1.15f
C460 X2/X1/X1/X2/vout vss 0.868f
C461 X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C462 X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C463 X2/X1/X1/X2/X2/vin1 vss 1.46f
C464 X2/X1/X1/X2/X3/vin2 vss 1.23f
C465 X2/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C466 X2/X1/X1/X2/X2/m1_994_178# vss 1.15f
C467 X2/X1/X2/vrefh vss 3.27f
C468 X2/X1/X1/X2/X1/vin1 vss 1.91f
C469 X2/X1/X1/X2/X3/vin1 vss 0.816f
C470 X2/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C471 X2/X1/X1/X2/X1/m1_994_178# vss 1.15f
C472 X2/X1/X1/X2/X1/vin2 vss 1.73f
C473 X2/X1/X1/X1/vout vss 0.607f
C474 X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C475 X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C476 X2/X1/X1/X1/X2/vin1 vss 1.46f
C477 X2/X1/X1/X1/X3/vin2 vss 1.23f
C478 X2/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C479 X2/X1/X1/X1/X2/m1_994_178# vss 1.15f
C480 X2/X1/X1/X2/vrefh vss 3.27f
C481 X2/X1/X1/X1/X1/vin1 vss 1.94f
C482 X2/X1/X1/X1/X3/vin1 vss 0.823f
C483 X2/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C484 X2/X1/X1/X1/X1/m1_994_178# vss 1.15f
C485 X2/X1/X1/X1/X1/vin2 vss 1.74f
C486 d4 vss 2.04f
C487 X3/vin1 vss 1.24f
C488 X1/X3/m1_688_n494# vss 0.857f
C489 X1/X3/m1_994_178# vss 1.15f
C490 d3 vss 7.57f
C491 X1/X3/vin2 vss 1.85f
C492 X1/X2/X3/m1_688_n494# vss 0.858f
C493 X1/X2/X3/m1_994_178# vss 1.15f
C494 d2 vss 11.5f
C495 X1/X2/X3/vin2 vss 1.75f
C496 X1/X2/X2/sw_0/m1_688_n494# vss 0.858f
C497 X1/X2/X2/sw_0/m1_994_178# vss 1.15f
C498 X1/X2/X2/X2/vout vss 0.868f
C499 X1/X2/X2/X2/X3/m1_688_n494# vss 0.856f
C500 X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C501 d0 vss 37f
C502 X1/X2/X2/X2/X2/vin1 vss 1.46f
C503 X1/X2/X2/X2/X3/vin2 vss 1.21f
C504 X1/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C505 X1/X2/X2/X2/X2/m1_994_178# vss 1.15f
C506 X2/vrefh vss 8.33f
C507 X1/X2/X2/X2/X1/vin1 vss 1.91f
C508 X1/X2/X2/X2/X3/vin1 vss 0.813f
C509 X1/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C510 X1/X2/X2/X2/X1/m1_994_178# vss 1.15f
C511 X1/X2/X2/X2/X1/vin2 vss 1.73f
C512 X1/X2/X2/X1/vout vss 0.607f
C513 X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C514 X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C515 X1/X2/X2/X1/X2/vin1 vss 1.46f
C516 X1/X2/X2/X1/X3/vin2 vss 1.23f
C517 X1/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C518 X1/X2/X2/X1/X2/m1_994_178# vss 1.15f
C519 X1/X2/X2/X2/vrefh vss 3.27f
C520 X1/X2/X2/X1/X1/vin1 vss 1.91f
C521 X1/X2/X2/X1/X3/vin1 vss 0.816f
C522 X1/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C523 X1/X2/X2/X1/X1/m1_994_178# vss 1.15f
C524 X1/X2/X2/X1/X1/vin2 vss 1.73f
C525 X1/X2/X3/vin1 vss 1.49f
C526 X1/X2/X1/sw_0/m1_688_n494# vss 0.858f
C527 X1/X2/X1/sw_0/m1_994_178# vss 1.15f
C528 X1/X2/X1/X2/vout vss 0.868f
C529 X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C530 X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C531 X1/X2/X1/X2/X2/vin1 vss 1.46f
C532 X1/X2/X1/X2/X3/vin2 vss 1.23f
C533 X1/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C534 X1/X2/X1/X2/X2/m1_994_178# vss 1.15f
C535 X1/X2/X2/vrefh vss 3.27f
C536 X1/X2/X1/X2/X1/vin1 vss 1.91f
C537 X1/X2/X1/X2/X3/vin1 vss 0.816f
C538 X1/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C539 X1/X2/X1/X2/X1/m1_994_178# vss 1.15f
C540 X1/X2/X1/X2/X1/vin2 vss 1.73f
C541 X1/X2/X1/X1/vout vss 0.607f
C542 X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C543 X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C544 X1/X2/X1/X1/X2/vin1 vss 1.46f
C545 X1/X2/X1/X1/X3/vin2 vss 1.23f
C546 X1/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C547 X1/X2/X1/X1/X2/m1_994_178# vss 1.15f
C548 X1/X2/X1/X2/vrefh vss 3.27f
C549 X1/X2/X1/X1/X1/vin1 vss 1.91f
C550 X1/X2/X1/X1/X3/vin1 vss 0.816f
C551 X1/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C552 X1/X2/X1/X1/X1/m1_994_178# vss 1.15f
C553 X1/X2/X1/X1/X1/vin2 vss 1.73f
C554 X1/X3/vin1 vss 1.6f
C555 X1/X1/X3/m1_688_n494# vss 0.858f
C556 X1/X1/X3/m1_994_178# vss 1.15f
C557 X1/X1/X3/vin2 vss 1.75f
C558 X1/X1/X2/sw_0/m1_688_n494# vss 0.858f
C559 X1/X1/X2/sw_0/m1_994_178# vss 1.15f
C560 X1/X1/X2/X2/vout vss 0.868f
C561 X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C562 X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C563 vdd vss 0.311p
C564 X1/X1/X2/X2/X2/vin1 vss 1.46f
C565 X1/X1/X2/X2/X3/vin2 vss 1.23f
C566 X1/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C567 X1/X1/X2/X2/X2/m1_994_178# vss 1.15f
C568 X1/X2/vrefh vss 3.27f
C569 X1/X1/X2/X2/X1/vin1 vss 1.91f
C570 X1/X1/X2/X2/X3/vin1 vss 0.816f
C571 X1/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C572 X1/X1/X2/X2/X1/m1_994_178# vss 1.15f
C573 X1/X1/X2/X2/X1/vin2 vss 1.73f
C574 X1/X1/X2/X1/vout vss 0.607f
C575 X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C576 X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C577 X1/X1/X2/X1/X2/vin1 vss 1.46f
C578 X1/X1/X2/X1/X3/vin2 vss 1.23f
C579 X1/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C580 X1/X1/X2/X1/X2/m1_994_178# vss 1.15f
C581 X1/X1/X2/X2/vrefh vss 3.27f
C582 X1/X1/X2/X1/X1/vin1 vss 1.91f
C583 X1/X1/X2/X1/X3/vin1 vss 0.816f
C584 X1/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C585 X1/X1/X2/X1/X1/m1_994_178# vss 1.15f
C586 X1/X1/X2/X1/X1/vin2 vss 1.73f
C587 X1/X1/X3/vin1 vss 1.49f
C588 X1/X1/X1/sw_0/m1_688_n494# vss 0.858f
C589 X1/X1/X1/sw_0/m1_994_178# vss 1.15f
C590 d1 vss 15.2f
C591 X1/X1/X1/X2/vout vss 0.868f
C592 X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C593 X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C594 X1/X1/X1/X2/X2/vin1 vss 1.46f
C595 X1/X1/X1/X2/X3/vin2 vss 1.23f
C596 X1/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C597 X1/X1/X1/X2/X2/m1_994_178# vss 1.15f
C598 X1/X1/X2/vrefh vss 3.27f
C599 X1/X1/X1/X2/X1/vin1 vss 1.91f
C600 X1/X1/X1/X2/X3/vin1 vss 0.816f
C601 X1/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C602 X1/X1/X1/X2/X1/m1_994_178# vss 1.15f
C603 X1/X1/X1/X2/X1/vin2 vss 1.73f
C604 X1/X1/X1/X1/vout vss 0.607f
C605 X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C606 X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C607 X1/X1/X1/X1/X2/vin1 vss 1.46f
C608 X1/X1/X1/X1/X3/vin2 vss 1.23f
C609 X1/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C610 X1/X1/X1/X1/X2/m1_994_178# vss 1.15f
C611 X1/X1/X1/X2/vrefh vss 3.27f
C612 X1/X1/X1/X1/X1/vin1 vss 1.96f
C613 X1/X1/X1/X1/X3/vin1 vss 0.823f
C614 X1/X1/X1/X1/X1/m1_688_n494# vss 0.859f
C615 X1/X1/X1/X1/X1/m1_994_178# vss 1.15f
C616 X1/X1/X1/X1/X1/vin2 vss 1.74f
C617 vrefh vss 1.11f
.ends

.subckt x7bit_dac d2 d4 d6 vout X2/X2/X1/X2/X1/X1/vin1 X1/X1/X2/X1/X2/vrefh X2/X2/X1/X2/X1/X2/vin1
+ X3/vin1 X1/X2/X2/X2/X2/X3/vin2 X2/X2/X2/X1/X1/X1/vin1 X1/X1/X1/X1/X2/X1/vin1 X2/X2/X1/X1/X1/X1/m1_994_178#
+ X2/X2/X2/X1/X1/X2/vin1 X2/X2/X1/X1/X1/X1/m1_688_n494# X1/X1/X1/X2/X1/X1/vin2 X1/X1/X1/X1/X2/X2/vin1
+ X2/X2/X1/X1/X2/X1/vin2 X2/X2/X1/X2/X2/vrefh X2/X2/X2/X2/X1/X1/vin1 X2/X2/X2/X2/X2/vrefh
+ X1/X1/X1/X1/X1/X1/m1_688_n494# X2/X3/m1_688_n494# X1/X1/X1/X2/X2/X1/vin1 X2/X2/X2/X2/X2/X1/vin2
+ X2/X2/X2/X2/X1/X2/vin1 X1/X1/X1/X1/X1/X1/vin1 X1/X1/X1/X2/X2/X2/vin1 X1/X1/X2/X1/X2/X1/vin2
+ X1/X1/X2/X1/X2/X1/vin1 X2/X2/X2/X2/X2/X1/vin1 X1/X1/X1/X2/X2/vrefh X1/X1/X2/X1/X2/X2/vin1
+ X1/X1/X2/X2/X2/vrefh X3/vin2 X2/X2/X2/X1/X1/X1/vin2 X2/X2/vrefh X1/X3/m1_994_178#
+ X1/X1/X1/X2/X2/X1/vin2 X1/X1/X1/X2/X1/X1/vin1 X1/X1/X2/X2/X2/X1/vin1 X1/X1/X1/X1/X1/X3/m1_994_178#
+ X2/X2/X1/X2/vrefh X1/X1/X1/X1/X1/X3/m1_688_n494# X1/X1/X2/X2/vrefh X1/X1/X1/X2/X1/X2/vin1
+ X1/X1/X2/X2/X2/X2/vin1 X1/X1/X2/X1/X1/X1/vin1 X1/X1/X1/X1/X1/X2/vin1 X2/X2/X1/X2/X1/X1/vin2
+ X1/X1/X1/X1/X1/X1/vin2 X1/X1/X2/X1/X1/X2/vin1 X1/X3/vin2 X2/X2/X2/X2/X2/X2/m1_994_178#
+ X1/X3/vin1 X2/X2/X2/X2/X2/X2/m1_688_n494# X1/X2/X2/X2/X2/X2/m1_994_178# vrefl X1/X2/X2/X2/X2/X2/m1_688_n494#
+ X2/X2/X2/X2/X2/X2/vin1 d1 X1/X1/X2/X2/X1/X1/vin1 X1/X1/X2/X2/X1/X1/vin2 X1/X3/m1_688_n494#
+ X2/X2/X2/X1/X2/X1/vin2 X3/m1_994_178# X1/X1/X2/X2/X1/X2/vin1 X2/X2/X1/X1/X2/X1/vin1
+ X2/X2/X1/X1/X2/X2/vin1 X2/X2/X2/X2/vrefh X2/X2/X1/X2/X2/X1/vin2 X1/X1/X1/X1/X2/X1/vin2
+ X2/X3/vin2 X1/X1/X1/X1/X1/X3/vin1 X1/X2/X2/X2/X2/X2/vin1 X2/X3/vin1 X2/X2/X1/X2/X2/X1/vin1
+ X2/X2/X2/vrefh X2/X2/X1/X1/X1/X1/vin2 X2/X2/X2/X1/X2/X1/vin1 X2/X2/X1/X2/X2/X2/vin1
+ X2/X2/X1/X1/X1/X1/vin1 X2/X2/X2/X2/X2/X3/vin2 X2/X2/X1/X1/X2/vrefh X1/X1/X2/X2/X2/X1/vin2
+ X1/X1/X2/X2/X2/X2/m1_994_178# X3/m1_688_n494# X1/X1/X2/X2/X2/X2/m1_688_n494# d5
+ X2/X2/X2/X1/X2/vrefh X2/X2/X2/X1/X2/X2/vin1 X2/X2/X1/X1/X1/X2/vin1 vdd X2/X1/X1/X1/X1/X1/vin2
+ d3 X1/X1/X1/X1/X1/X1/m1_994_178# vrefh X2/X3/m1_994_178# X2/X1/X1/X1/X1/X1/vin1
+ X2/X2/X2/X2/X1/X1/vin2 X1/X2/vrefh X2/vrefh vss X1/X1/X2/vrefh X1/X1/X1/X1/X2/vrefh
+ d0 X1/X1/X1/X2/vrefh X1/X1/X2/X1/X1/X1/vin2
XX1 vrefh d5 X3/vin1 X1/X1/X1/X1/X1/X3/vin1 X1/X2/X2/X1/sw_0/m1_688_n494# X1/X2/X2/X1/X2/vout
+ X1/X2/X1/X1/X2/X2/vin1 X1/X3/vin1 X1/X1/X1/X2/X1/X1/vin1 X1/X1/X2/X2/X2/X1/vin2
+ X1/X1/X1/X2/X1/X2/vin1 X1/X1/X2/X1/X1/X1/vin1 X1/X1/X2/X2/X2/X2/m1_688_n494# X1/X1/X2/X2/X2/X1/vin1
+ X1/X1/X2/vrefh X1/X2/X1/X2/X2/X1/vin1 X1/X1/X1/X1/X2/vrefh X1/X1/X2/X1/X1/X1/vin2
+ X1/X1/X2/X1/X1/X2/vin1 X1/X1/X2/X1/X2/vrefh X1/X2/X1/X2/X2/X2/vin1 X1/X2/X2/X1/X2/X1/vin1
+ X1/X2/X1/X1/X2/X1/vin2 X1/X2/X2/X1/X2/X2/vin1 X1/X1/X1/X1/X2/X3/vin2 X1/X1/X2/X2/X1/X1/vin1
+ X1/X1/X1/X2/X1/X1/vin2 X1/X1/X1/X1/X2/X3/vin1 X1/X2/X2/X1/X1/X3/m1_688_n494# X1/X1/X2/X2/X1/X2/vin1
+ X1/X2/X1/X1/X1/X2/vin1 X1/X1/X1/X2/X1/X3/m1_688_n494# X1/X2/X2/X1/X1/X1/vin2 X1/X2/X2/X2/X1/X3/vin2
+ X1/X2/X2/X2/X2/X3/vin1 X1/X2/X1/X2/X1/X1/vin1 X1/X2/X1/X1/X1/X1/m1_994_178# X1/X3/vin2
+ d4 X1/X2/X1/X1/X1/X1/m1_688_n494# X1/X1/X1/X3/m1_688_n494# X1/X2/X1/X2/X1/X2/vin1
+ X1/X2/X2/X2/X2/X2/vin1 X1/X2/X2/X1/X1/X1/vin1 X1/X1/X2/X1/X1/X3/vin1 X1/X2/X3/m1_688_n494#
+ X1/X1/X1/X3/vin1 X1/X1/X1/X1/X2/X3/m1_994_178# X1/X1/X2/X1/X2/X1/vin2 X1/X2/X2/X1/X2/X3/m1_688_n494#
+ X1/X1/X1/X1/X2/X3/m1_688_n494# X1/X2/X2/X1/X1/X2/vin1 X1/X1/X2/X2/X2/X2/vin1 X1/X2/X1/X2/X1/X1/vin2
+ X1/X1/X1/X2/X2/vrefh X1/X2/X2/X2/X1/X3/m1_994_178# X1/X1/X2/X2/X2/vrefh X1/X2/X2/X2/X1/X3/m1_688_n494#
+ X1/X2/X2/X2/sw_0/m1_994_178# X1/X2/X2/X1/X2/vrefh X1/X1/X3/vin2 X1/X2/X2/X2/sw_0/m1_688_n494#
+ X1/X1/X1/X1/X1/X1/m1_994_178# X1/X2/X2/X2/X1/X1/vin1 X1/X1/X1/X2/vrefh X1/X1/X1/X2/X1/vout
+ X1/X1/X1/X2/X2/X1/vin2 X1/X2/X1/X2/vrefh X1/X2/X2/X2/X1/X2/vin1 X1/X1/X1/X1/X2/vout
+ X1/X2/X2/X1/X2/X1/vin2 X1/X2/X2/X2/X2/X3/m1_994_178# d1 X1/X2/X2/X2/X2/X3/m1_688_n494#
+ X1/X2/X2/X2/X1/X3/vin1 X1/X2/X1/X1/X1/X3/vin1 X1/X3/m1_994_178# X1/X1/X1/X1/X1/X3/m1_994_178#
+ X1/X1/X1/X1/X1/X1/vin2 X1/X1/X1/X1/X1/X3/m1_688_n494# X1/X2/X2/X2/X2/vout X1/X1/X1/X3/vin2
+ X1/X2/X2/X2/X2/X1/vin2 X1/X1/X1/X2/sw_0/m1_688_n494# X1/X2/X1/X2/X2/X1/vin2 X1/X2/X1/X2/X2/vrefh
+ X1/X2/X2/X2/X2/X1/vin1 X1/X1/X1/X1/X2/X1/vin1 X1/X2/X2/X2/X2/vrefh X1/X2/X2/X3/vin1
+ X1/X2/X2/X1/X1/vout X1/X1/X3/vin1 X1/X1/X1/X1/X1/X1/m1_688_n494# X1/X2/X3/vin2 X1/X1/X2/X2/X1/X1/vin2
+ X1/X1/X1/X1/X2/X2/vin1 X1/X2/X2/X2/X2/X2/m1_994_178# X1/X2/X3/vin1 X1/X2/X2/X2/X2/X2/m1_688_n494#
+ X1/X2/X2/X3/vin2 X1/X1/X2/X2/vrefh X1/X1/X2/X2/X2/X2/m1_994_178# X1/X1/X1/X2/X2/vout
+ X1/X2/X2/X2/vrefh d3 X1/X1/X1/X1/X1/vout X1/X1/X1/X2/X2/X1/vin1 X1/X1/X3/m1_688_n494#
+ X1/X2/X2/vrefh X1/X3/m1_688_n494# X1/X1/X1/X1/X1/X1/vin1 X1/X1/X1/X1/X2/X1/vin2
+ X1/X1/X1/X2/X2/X2/vin1 X1/X1/X1/X2/X2/X3/m1_688_n494# vdd X1/X1/X2/X1/X2/X1/vin1
+ d2 X1/X2/X2/X2/X1/X1/vin2 X1/X2/X2/X2/X2/X3/vin2 X1/X2/X2/X3/m1_688_n494# X1/X1/X1/X1/X1/X2/vin1
+ X1/X1/X2/X1/X2/X2/vin1 X1/X1/X1/X1/sw_0/m1_688_n494# X1/X2/X1/X1/X1/X1/vin2 X1/X2/X2/X2/X1/vout
+ X1/X1/X1/X1/X1/X3/vin2 X1/X2/vrefh d0 X2/vrefh vss X1/X2/X1/X1/X2/X1/vin1 X1/X2/X1/X1/X2/vrefh
+ X1/X2/X1/X1/X1/X1/vin1 x6bit_dac
XX2 X2/vrefh d5 X3/vin2 X2/X1/X1/X1/X1/X3/vin1 X2/X2/X2/X1/sw_0/m1_688_n494# X2/X2/X2/X1/X2/vout
+ X2/X2/X1/X1/X2/X2/vin1 X2/X3/vin1 X2/X1/X1/X2/X1/X1/vin1 X2/X1/X2/X2/X2/X1/vin2
+ X2/X1/X1/X2/X1/X2/vin1 X2/X1/X2/X1/X1/X1/vin1 X2/X1/X2/X2/X2/X2/m1_688_n494# X2/X1/X2/X2/X2/X1/vin1
+ X2/X1/X2/vrefh X2/X2/X1/X2/X2/X1/vin1 X2/X1/X1/X1/X2/vrefh X2/X1/X2/X1/X1/X1/vin2
+ X2/X1/X2/X1/X1/X2/vin1 X2/X1/X2/X1/X2/vrefh X2/X2/X1/X2/X2/X2/vin1 X2/X2/X2/X1/X2/X1/vin1
+ X2/X2/X1/X1/X2/X1/vin2 X2/X2/X2/X1/X2/X2/vin1 X2/X1/X1/X1/X2/X3/vin2 X2/X1/X2/X2/X1/X1/vin1
+ X2/X1/X1/X2/X1/X1/vin2 X2/X1/X1/X1/X2/X3/vin1 X2/X2/X2/X1/X1/X3/m1_688_n494# X2/X1/X2/X2/X1/X2/vin1
+ X2/X2/X1/X1/X1/X2/vin1 X2/X1/X1/X2/X1/X3/m1_688_n494# X2/X2/X2/X1/X1/X1/vin2 X2/X2/X2/X2/X1/X3/vin2
+ X2/X2/X2/X2/X2/X3/vin1 X2/X2/X1/X2/X1/X1/vin1 X2/X2/X1/X1/X1/X1/m1_994_178# X2/X3/vin2
+ d4 X2/X2/X1/X1/X1/X1/m1_688_n494# X2/X1/X1/X3/m1_688_n494# X2/X2/X1/X2/X1/X2/vin1
+ X2/X2/X2/X2/X2/X2/vin1 X2/X2/X2/X1/X1/X1/vin1 X2/X1/X2/X1/X1/X3/vin1 X2/X2/X3/m1_688_n494#
+ X2/X1/X1/X3/vin1 X2/X1/X1/X1/X2/X3/m1_994_178# X2/X1/X2/X1/X2/X1/vin2 X2/X2/X2/X1/X2/X3/m1_688_n494#
+ X2/X1/X1/X1/X2/X3/m1_688_n494# X2/X2/X2/X1/X1/X2/vin1 X2/X1/X2/X2/X2/X2/vin1 X2/X2/X1/X2/X1/X1/vin2
+ X2/X1/X1/X2/X2/vrefh X2/X2/X2/X2/X1/X3/m1_994_178# X2/X1/X2/X2/X2/vrefh X2/X2/X2/X2/X1/X3/m1_688_n494#
+ X2/X2/X2/X2/sw_0/m1_994_178# X2/X2/X2/X1/X2/vrefh X2/X1/X3/vin2 X2/X2/X2/X2/sw_0/m1_688_n494#
+ X2/X1/X1/X1/X1/X1/m1_994_178# X2/X2/X2/X2/X1/X1/vin1 X2/X1/X1/X2/vrefh X2/X1/X1/X2/X1/vout
+ X2/X1/X1/X2/X2/X1/vin2 X2/X2/X1/X2/vrefh X2/X2/X2/X2/X1/X2/vin1 X2/X1/X1/X1/X2/vout
+ X2/X2/X2/X1/X2/X1/vin2 X2/X2/X2/X2/X2/X3/m1_994_178# d1 X2/X2/X2/X2/X2/X3/m1_688_n494#
+ X2/X2/X2/X2/X1/X3/vin1 X2/X2/X1/X1/X1/X3/vin1 X2/X3/m1_994_178# X2/X1/X1/X1/X1/X3/m1_994_178#
+ X2/X1/X1/X1/X1/X1/vin2 X2/X1/X1/X1/X1/X3/m1_688_n494# X2/X2/X2/X2/X2/vout X2/X1/X1/X3/vin2
+ X2/X2/X2/X2/X2/X1/vin2 X2/X1/X1/X2/sw_0/m1_688_n494# X2/X2/X1/X2/X2/X1/vin2 X2/X2/X1/X2/X2/vrefh
+ X2/X2/X2/X2/X2/X1/vin1 X2/X1/X1/X1/X2/X1/vin1 X2/X2/X2/X2/X2/vrefh X2/X2/X2/X3/vin1
+ X2/X2/X2/X1/X1/vout X2/X1/X3/vin1 X2/X1/X1/X1/X1/X1/m1_688_n494# X2/X2/X3/vin2 X2/X1/X2/X2/X1/X1/vin2
+ X2/X1/X1/X1/X2/X2/vin1 X2/X2/X2/X2/X2/X2/m1_994_178# X2/X2/X3/vin1 X2/X2/X2/X2/X2/X2/m1_688_n494#
+ X2/X2/X2/X3/vin2 X2/X1/X2/X2/vrefh X2/X1/X2/X2/X2/X2/m1_994_178# X2/X1/X1/X2/X2/vout
+ X2/X2/X2/X2/vrefh d3 X2/X1/X1/X1/X1/vout X2/X1/X1/X2/X2/X1/vin1 X2/X1/X3/m1_688_n494#
+ X2/X2/X2/vrefh X2/X3/m1_688_n494# X2/X1/X1/X1/X1/X1/vin1 X2/X1/X1/X1/X2/X1/vin2
+ X2/X1/X1/X2/X2/X2/vin1 X2/X1/X1/X2/X2/X3/m1_688_n494# vdd X2/X1/X2/X1/X2/X1/vin1
+ d2 X2/X2/X2/X2/X1/X1/vin2 X2/X2/X2/X2/X2/X3/vin2 X2/X2/X2/X3/m1_688_n494# X2/X1/X1/X1/X1/X2/vin1
+ X2/X1/X2/X1/X2/X2/vin1 X2/X1/X1/X1/sw_0/m1_688_n494# X2/X2/X1/X1/X1/X1/vin2 X2/X2/X2/X2/X1/vout
+ X2/X1/X1/X1/X1/X3/vin2 X2/X2/vrefh d0 vrefl vss X2/X2/X1/X1/X2/X1/vin1 X2/X2/X1/X1/X2/vrefh
+ X2/X2/X1/X1/X1/X1/vin1 x6bit_dac
XX3 X3/vin1 X3/vin2 vout vdd d6 X3/m1_688_n494# vss X3/m1_994_178# sw
C0 d4 X2/X1/X1/X3/m1_688_n494# 3.47e-19
C1 d2 X1/X1/X1/X1/X2/vout -0.00114f
C2 d2 X2/vrefh 0.168f
C3 d1 X3/vin1 0.0299f
C4 d3 X2/X1/X1/X1/X2/vout 0.125f
C5 X1/X2/X1/X2/X1/X2/vin1 X2/X1/X2/X1/X2/X1/vin2 0.00232f
C6 d1 X1/X2/X1/X1/X1/X3/vin1 0.00275f
C7 d1 X2/X3/vin1 0.0441f
C8 d3 X2/X2/X2/X3/vin1 3.57e-20
C9 d3 X1/X1/X3/vin1 -0.0356f
C10 X1/X2/X2/X2/X1/X2/vin1 X2/X1/X1/X1/X2/X1/vin2 0.00232f
C11 X1/X2/X2/X2/X2/X1/vin2 X2/X1/X1/X1/X1/X2/vin1 0.00232f
C12 X1/X3/vin2 X3/vin1 0.165f
C13 d3 X2/X1/X1/X1/X2/X3/vin2 0.0775f
C14 d3 X1/X2/X2/X3/m1_688_n494# 0.00146f
C15 d4 X2/X2/X2/X2/X2/vout 0.0955f
C16 X1/X2/X1/X2/vrefh X2/X1/X2/X2/X1/X1/vin2 0.0128f
C17 X1/X2/vrefh d1 0.195f
C18 d2 X1/X2/X2/X2/X2/X3/m1_688_n494# 2.8e-19
C19 X2/X3/m1_994_178# X2/X3/m1_688_n494# -0.0124f
C20 X2/vrefh X2/X1/X1/X1/X1/X1/vin1 0.0048f
C21 X1/X2/X1/X2/vrefh d0 0.00385f
C22 vdd X3/vin1 1.07f
C23 d3 X2/X1/X1/X1/X2/X3/vin1 0.0103f
C24 X1/X2/X1/X1/X1/X3/vin1 vdd -5.98e-19
C25 vdd X2/X3/vin1 -0.00138f
C26 d4 X2/X2/X2/X2/X2/X3/vin2 0.0533f
C27 d3 X2/X2/X2/X2/sw_0/m1_688_n494# 2.73e-19
C28 d3 X2/X1/X1/X1/X1/X3/vin2 0.0678f
C29 d2 X1/X2/X2/X2/X2/X2/m1_688_n494# 1.95e-19
C30 d4 X2/X2/X3/m1_688_n494# 1.8e-19
C31 d3 X2/X1/X1/X1/X1/X3/vin1 0.0103f
C32 d3 X1/X2/X2/X2/X1/X3/vin1 0.0137f
C33 d4 X2/X2/X2/X2/X2/X3/vin1 0.00851f
C34 d2 X2/X1/X1/X1/X1/X3/m1_688_n494# 2.32e-19
C35 X1/X2/vrefh vdd 0.003f
C36 d4 X2/X1/X3/vin1 0.425f
C37 d0 d2 3.9e-19
C38 X1/X2/X2/X2/X2/X1/vin1 X2/X1/X1/X1/X2/vrefh 0.00437f
C39 d0 X3/vin2 0.00479f
C40 X2/X2/vrefh X3/vin2 4.75e-20
C41 d3 d2 5.76f
C42 d4 X2/X2/X2/X1/X2/X3/m1_688_n494# 2.4e-19
C43 X1/X3/m1_688_n494# d5 0.0322f
C44 X2/X3/vin2 d5 -4.93e-19
C45 d3 X1/X2/X3/vin2 -0.00604f
C46 d4 X1/X2/X2/X2/X2/X2/m1_994_178# 1.8e-19
C47 X1/X2/X1/X1/X2/X2/vin1 X2/X1/X2/X2/X1/X1/vin2 0.00232f
C48 d2 X1/X2/X2/X2/X2/vout -0.00473f
C49 X2/X3/m1_994_178# X3/vin2 0.161f
C50 X2/X1/X3/vin1 X2/X2/X2/X3/vin2 -0.00712f
C51 d0 X1/X2/X2/vrefh 0.00385f
C52 d3 X2/X1/X1/X1/sw_0/m1_688_n494# 0.00177f
C53 d1 X2/X3/m1_688_n494# 5.18e-19
C54 X1/X1/X1/X1/X2/X3/vin1 d4 0.00851f
C55 X1/X3/vin1 d5 0.057f
C56 d2 X1/X2/X2/X2/X2/X3/vin2 0.00369f
C57 d0 d6 2.49e-19
C58 X1/X2/X1/X1/X2/vrefh X2/X1/X2/X2/X2/vrefh 0.117f
C59 d4 X2/X3/vin2 0.0087f
C60 d3 X2/X1/X1/X3/vin1 0.0658f
C61 X1/X2/X2/X1/X2/X1/vin1 X2/X1/X1/X2/X2/vrefh 0.00437f
C62 X1/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X2/X1/vin1 0.00437f
C63 d3 X2/X2/X2/X2/X1/vout 3.57e-20
C64 X2/vrefh X2/X1/X1/X1/X1/X1/vin2 0.0128f
C65 d4 X2/X1/X3/m1_688_n494# 1.04e-19
C66 d3 X2/X1/X1/X1/X1/X1/vin1 0.00492f
C67 d2 X2/X1/X1/X1/X1/vout 1.23e-19
C68 X1/X2/X2/X1/X1/X1/vin2 X2/X1/X1/X2/X2/X2/vin1 0.00232f
C69 X1/X2/X2/X1/X2/vrefh X2/X1/X1/X2/X2/X1/vin1 0.00437f
C70 d2 X1/X2/X2/X2/X2/X3/vin1 1.78e-33
C71 X1/X1/X3/vin1 X1/X2/X2/X3/vin2 -0.00712f
C72 X1/X3/vin1 d4 0.00102f
C73 d3 X2/X1/X1/X3/vin2 0.0441f
C74 d4 X2/X2/X2/X3/vin2 0.0939f
C75 d0 X2/X1/X2/X2/X2/vrefh 0.00385f
C76 d3 X1/X1/X3/vin2 -0.00208f
C77 X1/X3/vin1 X1/X3/m1_688_n494# -0.0204f
C78 d2 X2/X1/X1/X1/X1/X1/m1_994_178# 3.9e-19
C79 d4 X2/X2/X2/X1/X2/vout 3.47e-19
C80 X1/X1/X1/X3/vin2 d4 0.0401f
C81 X3/vin1 d5 0.0932f
C82 X2/X3/vin1 d5 0.00714f
C83 d1 X2/X2/X1/X1/X1/X1/m1_688_n494# 1.57e-19
C84 d1 d2 1.48e-20
C85 d1 X3/vin2 0.00146f
C86 X1/X2/vrefh d5 9.61e-19
C87 d2 X1/X2/X2/X2/X1/X3/m1_994_178# -7.81e-36
C88 X1/X2/X1/X2/X1/X1/vin2 X2/X1/X2/X1/X2/X2/vin1 0.00232f
C89 X1/X3/m1_688_n494# X3/vin1 0.0615f
C90 d2 X1/X2/X2/X2/sw_0/m1_688_n494# 1.51e-19
C91 d3 X2/X2/X2/X3/m1_688_n494# 1.23e-19
C92 d4 X1/X2/X2/X2/X1/vout 4.78e-20
C93 d2 vdd 0.159f
C94 d2 X2/X2/X2/X2/X2/X3/m1_688_n494# 1.89e-19
C95 d3 X2/X1/X1/X1/X1/X1/vin2 1.14e-19
C96 vdd X1/X2/X3/vin2 -7.09e-20
C97 d2 X1/X2/X2/X3/vin2 -7.11e-33
C98 vdd X3/vin2 0.0704f
C99 X1/X3/vin1 X3/vin1 0.169f
C100 d1 d6 2.34e-19
C101 d3 X1/X1/X1/X1/X2/vout 7.64e-20
C102 d3 X2/vrefh 0.00665f
C103 X1/X2/X2/X1/X2/X2/vin1 X2/X1/X1/X2/X1/X1/vin2 0.00232f
C104 vdd X2/X1/X1/X3/vin1 -2.84e-32
C105 d1 X2/X2/X1/X1/X1/X3/vin1 0.00275f
C106 X1/X1/X1/X2/X1/X3/m1_688_n494# d4 2.4e-19
C107 X1/X2/X1/X1/X2/vrefh X2/X1/X2/X2/X2/X1/vin2 0.0128f
C108 d0 X1/X2/X1/X1/X2/vrefh 0.00385f
C109 d4 X2/X1/X1/X1/X1/X1/m1_688_n494# 8.99e-20
C110 d3 X1/X2/X2/X2/X2/X3/m1_688_n494# 4.75e-19
C111 d4 X2/X1/X1/X1/X2/vout 1.45e-19
C112 d2 X1/X2/X2/X2/X2/X3/m1_994_178# 2.78e-35
C113 X2/X3/m1_688_n494# d5 0.0242f
C114 vdd X2/X2/X1/X1/X1/X3/vin1 -5.98e-19
C115 d3 X2/X2/X3/vin2 -0.0367f
C116 d4 X2/X2/X2/X3/vin1 8.41e-19
C117 d0 X3/m1_994_178# 2.73e-19
C118 X1/X1/X3/vin1 d4 0.917f
C119 d3 X1/X2/X2/X2/X2/X2/m1_688_n494# 1.28e-19
C120 d2 X2/X2/X2/X2/X2/vout -0.0013f
C121 d0 X2/X1/X2/X1/X2/vrefh 0.00385f
C122 X1/X2/X2/X1/X2/X1/vin2 X2/X1/X1/X2/X1/X2/vin1 0.00232f
C123 d0 X2/X2/vrefh 0.0562f
C124 X1/X2/X1/X1/X1/X1/vin2 X2/X2/vrefh 0.0128f
C125 X1/X2/vrefh X3/vin1 0.0451f
C126 d3 X2/X1/X1/X1/X1/X3/m1_688_n494# 3.23e-19
C127 d4 X1/X2/X2/X3/m1_688_n494# 3.58e-19
C128 d0 X1/X2/X1/X2/X2/vrefh 0.00385f
C129 X1/X2/X2/X1/X1/X2/vin1 X2/X1/X1/X2/X2/X1/vin2 0.00232f
C130 X1/X2/X1/X2/X2/vrefh X2/X1/X2/X1/X2/vrefh 0.117f
C131 d3 d0 2.56e-19
C132 X1/X2/X2/X2/X1/X1/vin1 X2/X1/X1/X2/vrefh 0.00437f
C133 d0 X1/X2/X2/X1/X2/vrefh 0.00385f
C134 X1/X2/X1/X2/X2/vrefh X2/X1/X2/X1/X2/X1/vin2 0.0128f
C135 X1/X1/X3/m1_688_n494# d4 1.99e-19
C136 d1 X2/X2/X1/X1/X1/X1/vin1 0.00581f
C137 X1/X2/X2/X2/X2/X2/vin1 X2/X1/X1/X1/X1/X1/vin2 0.00232f
C138 X2/X3/vin2 X2/X3/m1_688_n494# -0.0288f
C139 d4 X2/X2/X2/X2/sw_0/m1_688_n494# 0.00116f
C140 d0 X1/X2/X2/X2/X2/vrefh 0.00385f
C141 d4 X2/X2/X2/X2/X1/X3/m1_688_n494# 2.4e-19
C142 d3 X1/X2/X2/X2/X2/vout 0.222f
C143 X1/X2/X1/X1/X1/X1/vin1 X2/X2/vrefh 0.00437f
C144 d0 X3/m1_688_n494# 1.37e-19
C145 X1/X1/X1/X1/X1/X3/vin1 d4 0.00851f
C146 X3/vin2 d5 0.0456f
C147 X2/X2/vrefh X3/m1_688_n494# 2.22e-19
C148 vdd X2/vrefh 1.11e-34
C149 d3 X1/X2/X2/X2/X2/X3/vin2 0.109f
C150 d2 X1/X2/X2/X2/X2/X2/m1_994_178# 3.9e-19
C151 d3 X2/X1/X3/vin2 -5.8e-19
C152 d4 X1/X2/X2/X1/sw_0/m1_688_n494# 1.54e-19
C153 d2 d4 1.65f
C154 d0 X1/X2/X2/X2/vrefh 0.00385f
C155 d3 X2/X1/X1/X1/X1/vout 0.0408f
C156 d4 X1/X2/X3/vin2 0.436f
C157 X1/X1/X1/X2/X2/X3/m1_688_n494# d4 2.4e-19
C158 d3 X1/X2/X2/X2/X2/X3/vin1 0.0137f
C159 d4 X2/X1/X1/X1/sw_0/m1_688_n494# 5.68e-19
C160 d3 X1/X2/X2/X2/X1/X3/vin2 0.0944f
C161 X1/X2/X1/X1/X2/X1/vin2 X2/X1/X2/X2/X2/vrefh 0.0128f
C162 X2/X3/vin2 X3/vin2 0.0745f
C163 d5 d6 4.95e-19
C164 d1 X3/m1_994_178# 4.67e-19
C165 d1 d0 3.77f
C166 X1/X3/m1_994_178# d5 0.0065f
C167 X2/X3/vin1 X2/X3/m1_688_n494# -0.00513f
C168 d4 X2/X1/X1/X3/vin1 0.00246f
C169 X1/X2/X2/X2/X1/X1/vin2 X2/X1/X1/X2/vrefh 0.0128f
C170 d4 X2/X2/X2/X2/X1/vout 0.0233f
C171 d3 X2/X1/X1/X1/X1/X1/m1_994_178# 2.56e-19
C172 d1 X1/X2/X1/X1/X1/X1/vin2 0.0193f
C173 d1 X2/X2/vrefh 0.196f
C174 d1 X2/X2/X1/X1/X1/X1/vin2 0.0193f
C175 d4 X2/X1/X1/X1/X1/X1/vin1 0.00332f
C176 vdd X2/X2/X3/vin2 -7.09e-20
C177 d4 X2/X1/X1/X2/sw_0/m1_688_n494# 1.99e-19
C178 d0 X1/X3/vin2 -0.0053f
C179 X1/X1/X1/X1/X2/X3/m1_688_n494# d4 2.4e-19
C180 d4 X2/X2/X2/X2/X1/X3/vin2 0.0533f
C181 d1 X2/X3/m1_994_178# 4.67e-19
C182 d4 X2/X1/X1/X3/vin2 0.00419f
C183 d0 vdd -0.324f
C184 X1/X1/X3/vin2 d4 0.0377f
C185 X1/X2/X1/X2/X2/X1/vin2 X2/X1/X2/X1/X1/X2/vin1 0.00232f
C186 d3 X1/X2/X2/X3/vin1 4.39e-19
C187 d4 X2/X2/X2/X2/X1/X3/vin1 0.00851f
C188 vdd X2/X2/vrefh 0.00159f
C189 X2/X1/X1/X3/vin1 X2/X2/X2/X3/vin2 -2.1e-20
C190 d1 X1/X2/X1/X1/X1/X1/vin1 0.0129f
C191 d3 X1/X2/X2/X2/sw_0/m1_688_n494# 0.00329f
C192 d3 vdd 0.244f
C193 d1 X3/m1_688_n494# 2.34e-19
C194 d1 X2/X1/X2/X2/X2/X2/m1_688_n494# 1.39e-20
C195 d4 X2/X2/X2/X1/sw_0/m1_688_n494# 2.94e-19
C196 X1/X3/vin1 X1/X3/m1_994_178# -7.13e-19
C197 d3 X1/X2/X2/X3/vin2 0.258f
C198 X1/X1/X1/X3/m1_688_n494# d4 6.91e-19
C199 X1/X1/X1/X3/vin1 d3 0.00108f
C200 d4 X2/X2/X2/X1/X1/X3/m1_688_n494# 2.4e-19
C201 X2/X3/vin1 X3/vin2 0.0157f
C202 d2 X1/X2/X2/X2/X1/vout 1.32e-19
C203 d1 X1/X2/X1/X1/X1/X1/m1_994_178# 2.78e-20
C204 X1/X2/X1/X1/X2/vrefh X2/X1/X2/X2/X2/X1/vin1 0.00437f
C205 X1/X1/X1/X1/X2/X3/vin2 d4 0.0533f
C206 d0 X2/X1/X1/X2/vrefh 0.00385f
C207 vdd X3/m1_688_n494# -0.00407f
C208 X1/X2/X1/X2/X2/X1/vin1 X2/X1/X2/X1/X2/vrefh 0.00437f
C209 d4 X2/X2/X2/X3/m1_688_n494# 7.15e-19
C210 X1/X1/X1/X1/sw_0/m1_688_n494# d4 0.00116f
C211 X1/X2/X1/X1/X1/X1/vin2 X2/X1/X2/X2/X2/X2/vin1 0.00232f
C212 d4 X2/X1/X1/X1/X1/X1/vin2 8.21e-20
C213 d3 X2/X1/X1/X3/m1_688_n494# 7.75e-19
C214 vdd X2/X1/X1/X1/X1/vout -5.68e-32
C215 X1/X2/X1/X2/X1/X1/vin2 X2/X1/X2/X2/vrefh 0.0128f
C216 X1/X2/X2/vrefh X2/X1/X2/vrefh 0.117f
C217 X1/X2/X1/X2/X2/vrefh X2/X1/X2/X1/X2/X1/vin1 0.00437f
C218 X3/vin1 d6 0.0158f
C219 X1/X2/X1/X2/X2/X1/vin1 X1/X2/X1/X2/X2/vrefh 7.11e-33
C220 X1/X2/X1/X1/X1/X2/vin1 X2/X1/X2/X2/X2/X1/vin2 0.00232f
C221 X1/X3/m1_994_178# X3/vin1 0.00582f
C222 X1/X2/X1/X2/vrefh X2/X1/X2/X2/vrefh 0.117f
C223 X1/X1/X1/X1/X2/vout d4 0.0921f
C224 d4 X2/vrefh 0.00449f
C225 X1/X1/X1/X1/X1/vout d4 0.0336f
C226 X2/X1/X3/vin1 X2/X2/X3/vin2 -0.273f
C227 X1/X2/X1/X2/X2/X2/vin1 X2/X1/X2/X1/X1/X1/vin2 0.00232f
C228 d2 X2/X1/X1/X1/X1/X1/m1_688_n494# 1.95e-19
C229 d3 X2/X2/X2/X2/X2/vout 1.05e-19
C230 d0 X2/X1/X1/X2/X2/vrefh 0.00385f
C231 X1/X2/vrefh d6 4.63e-19
C232 d4 X2/X2/X2/X1/X1/vout 3.29e-19
C233 d2 X2/X1/X1/X1/X2/vout -0.00196f
C234 d1 vdd 0.521f
C235 X1/X2/X2/X1/X2/vrefh X2/X1/X1/X2/X2/vrefh 0.117f
C236 X1/X1/X3/vin1 X1/X2/X3/vin2 -0.273f
C237 vdd X1/X3/vin2 0.0771f
C238 X3/m1_994_178# d5 9.9e-19
C239 d0 d5 0.529f
C240 d4 X2/X2/X3/vin2 0.928f
C241 d4 X1/X2/X2/X2/X2/X2/m1_688_n494# 8.99e-20
C242 d3 X2/X1/X3/vin1 -0.00902f
C243 X2/X2/vrefh d5 9.61e-19
C244 X1/X2/X2/X2/vrefh X2/X1/X1/X2/vrefh 0.117f
C245 X1/X1/X1/X1/X1/X3/vin2 d4 0.0533f
C246 X1/X2/X1/X1/X2/X1/vin1 X2/X1/X2/X2/X2/vrefh 0.00437f
C247 X2/X3/m1_688_n494# X3/vin2 0.285f
C248 d2 X2/X2/X2/X2/sw_0/m1_688_n494# 1.78e-19
C249 X2/X3/m1_994_178# d5 0.00347f
C250 X1/X1/X1/X3/vin1 vdd 1.42e-32
C251 d0 d4 1.8e-19
C252 X1/X1/X1/X1/X1/X3/m1_688_n494# d4 2.4e-19
C253 X1/X1/X1/X3/vin1 X1/X2/X2/X3/vin2 -2.1e-20
C254 d2 X2/X1/X1/X1/X1/X3/vin1 0.00301f
C255 d3 X1/X2/X2/X2/X2/X2/m1_994_178# 2.56e-19
C256 d0 X2/X3/vin2 -0.00805f
C257 d3 d4 6.48f
C258 d2 X1/X2/X2/X2/sw_0/m1_994_178# 1.14e-31
C259 d4 X1/X2/X2/X2/X2/vout 1.45e-19
C260 d5 X3/m1_688_n494# 4.95e-19
C261 d3 X2/X3/vin2 -6.81e-19
C262 X2/X3/m1_994_178# X2/X3/vin2 -0.0015f
C263 d0 X1/X3/vin1 -8.92e-19
C264 X1/X2/X2/X1/X1/X1/vin1 X2/X1/X2/vrefh 0.00437f
C265 X1/X2/X2/X2/X2/X1/vin2 X2/X1/X1/X1/X2/vrefh 0.0128f
C266 d2 X2/X1/X1/X1/X1/X3/m1_994_178# 2.97e-20
C267 d4 X1/X2/X2/X2/X2/X3/vin2 1.57e-19
C268 d4 X2/X1/X3/vin2 0.0236f
C269 d4 X1/X2/X3/m1_688_n494# 9.46e-20
C270 d3 X1/X2/X2/X2/X1/X3/m1_688_n494# 4.75e-19
C271 d3 X2/X2/X2/X3/vin2 -0.00156f
C272 d2 X2/X1/X1/X1/sw_0/m1_688_n494# 6.21e-20
C273 d4 X2/X1/X1/X1/X1/vout 4.78e-20
C274 X1/X2/X2/X2/vrefh X2/X1/X1/X2/X1/X1/vin1 0.00437f
C275 d2 X2/X1/X1/X3/vin1 1.11e-34
C276 d2 X2/X2/X2/X2/X1/vout 7.09e-20
C277 X1/X2/X1/X2/X2/X1/vin2 X2/X1/X2/X1/X2/vrefh 0.0128f
C278 X1/X1/X1/X3/vin2 d3 -0.00232f
C279 d2 X2/X1/X1/X1/X1/X1/vin1 0.0337f
C280 d1 d5 2.27f
C281 X3/vin1 X3/m1_994_178# 0.0255f
C282 d0 X3/vin1 0.0254f
C283 X1/X1/X1/X2/X1/vout d4 3.29e-19
C284 d4 X2/X1/X1/X1/X1/X1/m1_994_178# 1.8e-19
C285 X3/vin1 X2/X2/vrefh 0.00136f
C286 d0 X2/X3/vin1 -0.00364f
C287 X1/X2/X2/vrefh X2/X1/X2/X1/X1/X1/vin1 0.00437f
C288 d0 X2/X1/X2/vrefh 0.00385f
C289 X1/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X2/X1/vin2 0.0128f
C290 d2 X2/X2/X2/X2/X1/X3/vin2 1.39e-35
C291 d4 X2/X2/X3/vin1 4.44e-34
C292 d4 X1/X1/X1/X2/sw_0/m1_688_n494# 3.79e-19
C293 X1/X3/vin2 d5 0.0373f
C294 d4 X1/X1/X1/X2/X2/vout 3.47e-19
C295 vdd X2/X1/X3/vin1 -2.84e-32
C296 X1/X2/X2/X1/X2/vrefh X2/X1/X1/X2/X2/X1/vin2 0.0128f
C297 X1/X2/vrefh d0 0.0571f
C298 X2/X3/vin1 X2/X3/m1_994_178# -4.6e-19
C299 X1/X2/X2/X1/X2/X1/vin2 X2/X1/X1/X2/X2/vrefh 0.0128f
C300 d1 X1/X2/X1/X1/X1/X1/m1_688_n494# 1.71e-19
C301 X1/X2/vrefh X2/X2/vrefh 0.0959f
C302 vdd d5 3.93f
C303 d3 X2/X1/X1/X1/X2/X3/m1_688_n494# 3.23e-19
C304 d1 X2/X3/vin2 0.0431f
C305 d4 X1/X2/X2/X3/vin1 3.38e-19
C306 d3 X1/X2/X2/X2/X1/vout 0.0406f
C307 d0 X2/X1/X1/X1/X2/vrefh 0.00385f
C308 X1/X2/X1/X2/vrefh X2/X1/X2/X2/X1/X1/vin1 0.00437f
C309 X1/X2/X2/X1/X1/X1/vin2 X2/X1/X2/vrefh 0.0128f
C310 d2 X2/X1/X1/X1/X2/X3/m1_994_178# -1.73e-36
C311 d4 X1/X2/X2/X2/sw_0/m1_688_n494# 5.68e-19
C312 X3/vin1 X3/m1_688_n494# 0.035f
C313 vdd d4 0.204f
C314 d4 X2/X2/X2/X2/X2/X3/m1_688_n494# 2.4e-19
C315 d4 X1/X2/X2/X3/vin2 0.0175f
C316 X1/X1/X1/X3/vin1 d4 0.0378f
C317 X1/X2/X2/X2/vrefh X2/X1/X1/X2/X1/X1/vin2 0.0128f
C318 vdd X1/X3/m1_688_n494# -0.00196f
C319 X1/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X2/vrefh 0.117f
C320 X1/X3/vin1 X1/X3/vin2 -2.18e-19
C321 d2 X1/X1/X1/X1/sw_0/m1_688_n494# 8.29e-20
C322 X1/X2/X2/X2/X1/X1/vin2 X2/X1/X1/X1/X2/X2/vin1 0.00232f
C323 d2 X2/X1/X1/X1/X1/X1/vin2 1.68e-19
C324 X1/X1/X2/X1/X1/X3/vin1 d4 1.78e-33
C325 d0 X2/X1/X2/X2/vrefh 0.00385f
C326 X1/X2/X1/X1/X2/X1/vin2 X2/X1/X2/X2/X1/X2/vin1 0.00232f
C327 X1/X2/X2/vrefh X2/X1/X2/X1/X1/X1/vin2 0.0128f
C328 d3 X2/X1/X1/X1/X1/X1/m1_688_n494# 1.28e-19
C329 X1/X2/X1/X2/X1/X1/vin1 X2/X1/X2/X2/vrefh 0.00437f
C330 d1 X2/X1/X2/X2/X2/X2/m1_994_178# 2.78e-20
C331 vdd X1/X3/vin1 0.00162f
C332 d6 vss 0.613f
C333 vout vss 0.2f
C334 X3/m1_688_n494# vss 0.858f
C335 X3/m1_994_178# vss 1.15f
C336 d5 vss 2.57f
C337 X3/vin2 vss 3.08f
C338 X2/X3/m1_688_n494# vss 0.847f
C339 X2/X3/m1_994_178# vss 1.15f
C340 X2/X3/vin2 vss 1.26f
C341 X2/X2/X3/m1_688_n494# vss 0.858f
C342 X2/X2/X3/m1_994_178# vss 1.15f
C343 X2/X2/X3/vin2 vss 1.85f
C344 X2/X2/X2/X3/m1_688_n494# vss 0.858f
C345 X2/X2/X2/X3/m1_994_178# vss 1.15f
C346 X2/X2/X2/X3/vin2 vss 1.75f
C347 X2/X2/X2/X2/sw_0/m1_688_n494# vss 0.858f
C348 X2/X2/X2/X2/sw_0/m1_994_178# vss 1.15f
C349 X2/X2/X2/X2/X2/vout vss 0.868f
C350 X2/X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C351 X2/X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C352 X2/X2/X2/X2/X2/X2/vin1 vss 1.46f
C353 X2/X2/X2/X2/X2/X3/vin2 vss 1.23f
C354 X2/X2/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C355 X2/X2/X2/X2/X2/X2/m1_994_178# vss 1.15f
C356 vrefl vss 2.39f
C357 X2/X2/X2/X2/X2/X1/vin1 vss 1.91f
C358 X2/X2/X2/X2/X2/X3/vin1 vss 0.816f
C359 X2/X2/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C360 X2/X2/X2/X2/X2/X1/m1_994_178# vss 1.15f
C361 X2/X2/X2/X2/X2/X1/vin2 vss 1.73f
C362 X2/X2/X2/X2/X1/vout vss 0.607f
C363 X2/X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C364 X2/X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C365 X2/X2/X2/X2/X1/X2/vin1 vss 1.46f
C366 X2/X2/X2/X2/X1/X3/vin2 vss 1.23f
C367 X2/X2/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C368 X2/X2/X2/X2/X1/X2/m1_994_178# vss 1.15f
C369 X2/X2/X2/X2/X2/vrefh vss 3.27f
C370 X2/X2/X2/X2/X1/X1/vin1 vss 1.91f
C371 X2/X2/X2/X2/X1/X3/vin1 vss 0.816f
C372 X2/X2/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C373 X2/X2/X2/X2/X1/X1/m1_994_178# vss 1.15f
C374 X2/X2/X2/X2/X1/X1/vin2 vss 1.73f
C375 X2/X2/X2/X3/vin1 vss 1.49f
C376 X2/X2/X2/X1/sw_0/m1_688_n494# vss 0.858f
C377 X2/X2/X2/X1/sw_0/m1_994_178# vss 1.15f
C378 X2/X2/X2/X1/X2/vout vss 0.868f
C379 X2/X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C380 X2/X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C381 X2/X2/X2/X1/X2/X2/vin1 vss 1.46f
C382 X2/X2/X2/X1/X2/X3/vin2 vss 1.23f
C383 X2/X2/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C384 X2/X2/X2/X1/X2/X2/m1_994_178# vss 1.15f
C385 X2/X2/X2/X2/vrefh vss 3.27f
C386 X2/X2/X2/X1/X2/X1/vin1 vss 1.91f
C387 X2/X2/X2/X1/X2/X3/vin1 vss 0.816f
C388 X2/X2/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C389 X2/X2/X2/X1/X2/X1/m1_994_178# vss 1.15f
C390 X2/X2/X2/X1/X2/X1/vin2 vss 1.73f
C391 X2/X2/X2/X1/X1/vout vss 0.607f
C392 X2/X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C393 X2/X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C394 X2/X2/X2/X1/X1/X2/vin1 vss 1.46f
C395 X2/X2/X2/X1/X1/X3/vin2 vss 1.23f
C396 X2/X2/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C397 X2/X2/X2/X1/X1/X2/m1_994_178# vss 1.15f
C398 X2/X2/X2/X1/X2/vrefh vss 3.27f
C399 X2/X2/X2/X1/X1/X1/vin1 vss 1.91f
C400 X2/X2/X2/X1/X1/X3/vin1 vss 0.816f
C401 X2/X2/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C402 X2/X2/X2/X1/X1/X1/m1_994_178# vss 1.15f
C403 X2/X2/X2/X1/X1/X1/vin2 vss 1.73f
C404 X2/X2/X3/vin1 vss 1.6f
C405 X2/X2/X1/X3/m1_688_n494# vss 0.858f
C406 X2/X2/X1/X3/m1_994_178# vss 1.15f
C407 X2/X2/X1/X3/vin2 vss 1.75f
C408 X2/X2/X1/X2/sw_0/m1_688_n494# vss 0.858f
C409 X2/X2/X1/X2/sw_0/m1_994_178# vss 1.15f
C410 X2/X2/X1/X2/X2/vout vss 0.868f
C411 X2/X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C412 X2/X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C413 X2/X2/X1/X2/X2/X2/vin1 vss 1.46f
C414 X2/X2/X1/X2/X2/X3/vin2 vss 1.23f
C415 X2/X2/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C416 X2/X2/X1/X2/X2/X2/m1_994_178# vss 1.15f
C417 X2/X2/X2/vrefh vss 3.27f
C418 X2/X2/X1/X2/X2/X1/vin1 vss 1.91f
C419 X2/X2/X1/X2/X2/X3/vin1 vss 0.816f
C420 X2/X2/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C421 X2/X2/X1/X2/X2/X1/m1_994_178# vss 1.15f
C422 X2/X2/X1/X2/X2/X1/vin2 vss 1.73f
C423 X2/X2/X1/X2/X1/vout vss 0.607f
C424 X2/X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C425 X2/X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C426 X2/X2/X1/X2/X1/X2/vin1 vss 1.46f
C427 X2/X2/X1/X2/X1/X3/vin2 vss 1.23f
C428 X2/X2/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C429 X2/X2/X1/X2/X1/X2/m1_994_178# vss 1.15f
C430 X2/X2/X1/X2/X2/vrefh vss 3.27f
C431 X2/X2/X1/X2/X1/X1/vin1 vss 1.91f
C432 X2/X2/X1/X2/X1/X3/vin1 vss 0.816f
C433 X2/X2/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C434 X2/X2/X1/X2/X1/X1/m1_994_178# vss 1.15f
C435 X2/X2/X1/X2/X1/X1/vin2 vss 1.73f
C436 X2/X2/X1/X3/vin1 vss 1.49f
C437 X2/X2/X1/X1/sw_0/m1_688_n494# vss 0.858f
C438 X2/X2/X1/X1/sw_0/m1_994_178# vss 1.15f
C439 X2/X2/X1/X1/X2/vout vss 0.868f
C440 X2/X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C441 X2/X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C442 X2/X2/X1/X1/X2/X2/vin1 vss 1.46f
C443 X2/X2/X1/X1/X2/X3/vin2 vss 1.23f
C444 X2/X2/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C445 X2/X2/X1/X1/X2/X2/m1_994_178# vss 1.15f
C446 X2/X2/X1/X2/vrefh vss 3.27f
C447 X2/X2/X1/X1/X2/X1/vin1 vss 1.91f
C448 X2/X2/X1/X1/X2/X3/vin1 vss 0.816f
C449 X2/X2/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C450 X2/X2/X1/X1/X2/X1/m1_994_178# vss 1.15f
C451 X2/X2/X1/X1/X2/X1/vin2 vss 1.73f
C452 X2/X2/X1/X1/X1/vout vss 0.607f
C453 X2/X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C454 X2/X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C455 X2/X2/X1/X1/X1/X2/vin1 vss 1.46f
C456 X2/X2/X1/X1/X1/X3/vin2 vss 1.23f
C457 X2/X2/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C458 X2/X2/X1/X1/X1/X2/m1_994_178# vss 1.15f
C459 X2/X2/X1/X1/X2/vrefh vss 3.27f
C460 X2/X2/X1/X1/X1/X1/vin1 vss 1.91f
C461 X2/X2/X1/X1/X1/X3/vin1 vss 0.816f
C462 X2/X2/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C463 X2/X2/X1/X1/X1/X1/m1_994_178# vss 1.15f
C464 X2/X2/X1/X1/X1/X1/vin2 vss 1.73f
C465 X2/X3/vin1 vss 1.12f
C466 X2/X1/X3/m1_688_n494# vss 0.858f
C467 X2/X1/X3/m1_994_178# vss 1.15f
C468 X2/X1/X3/vin2 vss 1.85f
C469 X2/X1/X2/X3/m1_688_n494# vss 0.858f
C470 X2/X1/X2/X3/m1_994_178# vss 1.15f
C471 X2/X1/X2/X3/vin2 vss 1.75f
C472 X2/X1/X2/X2/sw_0/m1_688_n494# vss 0.858f
C473 X2/X1/X2/X2/sw_0/m1_994_178# vss 1.15f
C474 X2/X1/X2/X2/X2/vout vss 0.868f
C475 X2/X1/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C476 X2/X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C477 X2/X1/X2/X2/X2/X2/vin1 vss 1.46f
C478 X2/X1/X2/X2/X2/X3/vin2 vss 1.23f
C479 X2/X1/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C480 X2/X1/X2/X2/X2/X2/m1_994_178# vss 1.15f
C481 X2/X2/vrefh vss 6.36f
C482 X2/X1/X2/X2/X2/X1/vin1 vss 1.91f
C483 X2/X1/X2/X2/X2/X3/vin1 vss 0.816f
C484 X2/X1/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C485 X2/X1/X2/X2/X2/X1/m1_994_178# vss 1.15f
C486 X2/X1/X2/X2/X2/X1/vin2 vss 1.74f
C487 X2/X1/X2/X2/X1/vout vss 0.607f
C488 X2/X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C489 X2/X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C490 X2/X1/X2/X2/X1/X2/vin1 vss 1.46f
C491 X2/X1/X2/X2/X1/X3/vin2 vss 1.23f
C492 X2/X1/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C493 X2/X1/X2/X2/X1/X2/m1_994_178# vss 1.15f
C494 X2/X1/X2/X2/X2/vrefh vss 3.27f
C495 X2/X1/X2/X2/X1/X1/vin1 vss 1.91f
C496 X2/X1/X2/X2/X1/X3/vin1 vss 0.816f
C497 X2/X1/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C498 X2/X1/X2/X2/X1/X1/m1_994_178# vss 1.15f
C499 X2/X1/X2/X2/X1/X1/vin2 vss 1.74f
C500 X2/X1/X2/X3/vin1 vss 1.49f
C501 X2/X1/X2/X1/sw_0/m1_688_n494# vss 0.858f
C502 X2/X1/X2/X1/sw_0/m1_994_178# vss 1.15f
C503 X2/X1/X2/X1/X2/vout vss 0.868f
C504 X2/X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C505 X2/X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C506 X2/X1/X2/X1/X2/X2/vin1 vss 1.46f
C507 X2/X1/X2/X1/X2/X3/vin2 vss 1.23f
C508 X2/X1/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C509 X2/X1/X2/X1/X2/X2/m1_994_178# vss 1.15f
C510 X2/X1/X2/X2/vrefh vss 3.27f
C511 X2/X1/X2/X1/X2/X1/vin1 vss 1.91f
C512 X2/X1/X2/X1/X2/X3/vin1 vss 0.816f
C513 X2/X1/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C514 X2/X1/X2/X1/X2/X1/m1_994_178# vss 1.15f
C515 X2/X1/X2/X1/X2/X1/vin2 vss 1.74f
C516 X2/X1/X2/X1/X1/vout vss 0.607f
C517 X2/X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C518 X2/X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C519 X2/X1/X2/X1/X1/X2/vin1 vss 1.46f
C520 X2/X1/X2/X1/X1/X3/vin2 vss 1.23f
C521 X2/X1/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C522 X2/X1/X2/X1/X1/X2/m1_994_178# vss 1.15f
C523 X2/X1/X2/X1/X2/vrefh vss 3.27f
C524 X2/X1/X2/X1/X1/X1/vin1 vss 1.91f
C525 X2/X1/X2/X1/X1/X3/vin1 vss 0.816f
C526 X2/X1/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C527 X2/X1/X2/X1/X1/X1/m1_994_178# vss 1.15f
C528 X2/X1/X2/X1/X1/X1/vin2 vss 1.74f
C529 X2/X1/X3/vin1 vss 1.6f
C530 X2/X1/X1/X3/m1_688_n494# vss 0.858f
C531 X2/X1/X1/X3/m1_994_178# vss 1.15f
C532 X2/X1/X1/X3/vin2 vss 1.75f
C533 X2/X1/X1/X2/sw_0/m1_688_n494# vss 0.858f
C534 X2/X1/X1/X2/sw_0/m1_994_178# vss 1.15f
C535 X2/X1/X1/X2/X2/vout vss 0.868f
C536 X2/X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C537 X2/X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C538 X2/X1/X1/X2/X2/X2/vin1 vss 1.46f
C539 X2/X1/X1/X2/X2/X3/vin2 vss 1.23f
C540 X2/X1/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C541 X2/X1/X1/X2/X2/X2/m1_994_178# vss 1.15f
C542 X2/X1/X2/vrefh vss 3.27f
C543 X2/X1/X1/X2/X2/X1/vin1 vss 1.91f
C544 X2/X1/X1/X2/X2/X3/vin1 vss 0.816f
C545 X2/X1/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C546 X2/X1/X1/X2/X2/X1/m1_994_178# vss 1.15f
C547 X2/X1/X1/X2/X2/X1/vin2 vss 1.74f
C548 X2/X1/X1/X2/X1/vout vss 0.607f
C549 X2/X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C550 X2/X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C551 X2/X1/X1/X2/X1/X2/vin1 vss 1.46f
C552 X2/X1/X1/X2/X1/X3/vin2 vss 1.23f
C553 X2/X1/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C554 X2/X1/X1/X2/X1/X2/m1_994_178# vss 1.15f
C555 X2/X1/X1/X2/X2/vrefh vss 3.27f
C556 X2/X1/X1/X2/X1/X1/vin1 vss 1.91f
C557 X2/X1/X1/X2/X1/X3/vin1 vss 0.816f
C558 X2/X1/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C559 X2/X1/X1/X2/X1/X1/m1_994_178# vss 1.15f
C560 X2/X1/X1/X2/X1/X1/vin2 vss 1.74f
C561 X2/X1/X1/X3/vin1 vss 1.49f
C562 X2/X1/X1/X1/sw_0/m1_688_n494# vss 0.858f
C563 X2/X1/X1/X1/sw_0/m1_994_178# vss 1.15f
C564 X2/X1/X1/X1/X2/vout vss 0.868f
C565 X2/X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C566 X2/X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C567 X2/X1/X1/X1/X2/X2/vin1 vss 1.46f
C568 X2/X1/X1/X1/X2/X3/vin2 vss 1.23f
C569 X2/X1/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C570 X2/X1/X1/X1/X2/X2/m1_994_178# vss 1.15f
C571 X2/X1/X1/X2/vrefh vss 3.27f
C572 X2/X1/X1/X1/X2/X1/vin1 vss 1.91f
C573 X2/X1/X1/X1/X2/X3/vin1 vss 0.816f
C574 X2/X1/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C575 X2/X1/X1/X1/X2/X1/m1_994_178# vss 1.15f
C576 X2/X1/X1/X1/X2/X1/vin2 vss 1.74f
C577 X2/X1/X1/X1/X1/vout vss 0.607f
C578 X2/X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C579 X2/X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C580 X2/X1/X1/X1/X1/X2/vin1 vss 1.46f
C581 X2/X1/X1/X1/X1/X3/vin2 vss 1.23f
C582 X2/X1/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C583 X2/X1/X1/X1/X1/X2/m1_994_178# vss 1.15f
C584 X2/X1/X1/X1/X2/vrefh vss 3.27f
C585 X2/X1/X1/X1/X1/X1/vin1 vss 1.91f
C586 X2/X1/X1/X1/X1/X3/vin1 vss 0.816f
C587 X2/X1/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C588 X2/X1/X1/X1/X1/X1/m1_994_178# vss 1.15f
C589 X2/X1/X1/X1/X1/X1/vin2 vss 1.74f
C590 X3/vin1 vss 1.6f
C591 X1/X3/m1_688_n494# vss 0.858f
C592 X1/X3/m1_994_178# vss 1.15f
C593 X1/X3/vin2 vss 1.27f
C594 X1/X2/X3/m1_688_n494# vss 0.858f
C595 X1/X2/X3/m1_994_178# vss 1.15f
C596 X1/X2/X3/vin2 vss 1.85f
C597 X1/X2/X2/X3/m1_688_n494# vss 0.858f
C598 X1/X2/X2/X3/m1_994_178# vss 1.15f
C599 X1/X2/X2/X3/vin2 vss 1.75f
C600 X1/X2/X2/X2/sw_0/m1_688_n494# vss 0.858f
C601 X1/X2/X2/X2/sw_0/m1_994_178# vss 1.15f
C602 X1/X2/X2/X2/X2/vout vss 0.868f
C603 X1/X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C604 X1/X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C605 X1/X2/X2/X2/X2/X2/vin1 vss 1.46f
C606 X1/X2/X2/X2/X2/X3/vin2 vss 1.23f
C607 X1/X2/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C608 X1/X2/X2/X2/X2/X2/m1_994_178# vss 1.15f
C609 X2/vrefh vss 3.66f
C610 X1/X2/X2/X2/X2/X1/vin1 vss 1.91f
C611 X1/X2/X2/X2/X2/X3/vin1 vss 0.816f
C612 X1/X2/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C613 X1/X2/X2/X2/X2/X1/m1_994_178# vss 1.15f
C614 X1/X2/X2/X2/X2/X1/vin2 vss 1.74f
C615 X1/X2/X2/X2/X1/vout vss 0.607f
C616 X1/X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C617 X1/X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C618 X1/X2/X2/X2/X1/X2/vin1 vss 1.46f
C619 X1/X2/X2/X2/X1/X3/vin2 vss 1.23f
C620 X1/X2/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C621 X1/X2/X2/X2/X1/X2/m1_994_178# vss 1.15f
C622 X1/X2/X2/X2/X2/vrefh vss 3.27f
C623 X1/X2/X2/X2/X1/X1/vin1 vss 1.91f
C624 X1/X2/X2/X2/X1/X3/vin1 vss 0.816f
C625 X1/X2/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C626 X1/X2/X2/X2/X1/X1/m1_994_178# vss 1.15f
C627 X1/X2/X2/X2/X1/X1/vin2 vss 1.74f
C628 X1/X2/X2/X3/vin1 vss 1.49f
C629 X1/X2/X2/X1/sw_0/m1_688_n494# vss 0.858f
C630 X1/X2/X2/X1/sw_0/m1_994_178# vss 1.15f
C631 X1/X2/X2/X1/X2/vout vss 0.868f
C632 X1/X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C633 X1/X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C634 X1/X2/X2/X1/X2/X2/vin1 vss 1.46f
C635 X1/X2/X2/X1/X2/X3/vin2 vss 1.23f
C636 X1/X2/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C637 X1/X2/X2/X1/X2/X2/m1_994_178# vss 1.15f
C638 X1/X2/X2/X2/vrefh vss 3.27f
C639 X1/X2/X2/X1/X2/X1/vin1 vss 1.91f
C640 X1/X2/X2/X1/X2/X3/vin1 vss 0.816f
C641 X1/X2/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C642 X1/X2/X2/X1/X2/X1/m1_994_178# vss 1.15f
C643 X1/X2/X2/X1/X2/X1/vin2 vss 1.74f
C644 X1/X2/X2/X1/X1/vout vss 0.607f
C645 X1/X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C646 X1/X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C647 X1/X2/X2/X1/X1/X2/vin1 vss 1.46f
C648 X1/X2/X2/X1/X1/X3/vin2 vss 1.23f
C649 X1/X2/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C650 X1/X2/X2/X1/X1/X2/m1_994_178# vss 1.15f
C651 X1/X2/X2/X1/X2/vrefh vss 3.27f
C652 X1/X2/X2/X1/X1/X1/vin1 vss 1.91f
C653 X1/X2/X2/X1/X1/X3/vin1 vss 0.816f
C654 X1/X2/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C655 X1/X2/X2/X1/X1/X1/m1_994_178# vss 1.15f
C656 X1/X2/X2/X1/X1/X1/vin2 vss 1.74f
C657 X1/X2/X3/vin1 vss 1.6f
C658 X1/X2/X1/X3/m1_688_n494# vss 0.858f
C659 X1/X2/X1/X3/m1_994_178# vss 1.15f
C660 X1/X2/X1/X3/vin2 vss 1.75f
C661 X1/X2/X1/X2/sw_0/m1_688_n494# vss 0.858f
C662 X1/X2/X1/X2/sw_0/m1_994_178# vss 1.15f
C663 X1/X2/X1/X2/X2/vout vss 0.868f
C664 X1/X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C665 X1/X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C666 X1/X2/X1/X2/X2/X2/vin1 vss 1.46f
C667 X1/X2/X1/X2/X2/X3/vin2 vss 1.23f
C668 X1/X2/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C669 X1/X2/X1/X2/X2/X2/m1_994_178# vss 1.15f
C670 X1/X2/X2/vrefh vss 3.27f
C671 X1/X2/X1/X2/X2/X1/vin1 vss 1.91f
C672 X1/X2/X1/X2/X2/X3/vin1 vss 0.816f
C673 X1/X2/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C674 X1/X2/X1/X2/X2/X1/m1_994_178# vss 1.15f
C675 X1/X2/X1/X2/X2/X1/vin2 vss 1.74f
C676 X1/X2/X1/X2/X1/vout vss 0.607f
C677 X1/X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C678 X1/X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C679 X1/X2/X1/X2/X1/X2/vin1 vss 1.46f
C680 X1/X2/X1/X2/X1/X3/vin2 vss 1.23f
C681 X1/X2/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C682 X1/X2/X1/X2/X1/X2/m1_994_178# vss 1.15f
C683 X1/X2/X1/X2/X2/vrefh vss 3.27f
C684 X1/X2/X1/X2/X1/X1/vin1 vss 1.91f
C685 X1/X2/X1/X2/X1/X3/vin1 vss 0.816f
C686 X1/X2/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C687 X1/X2/X1/X2/X1/X1/m1_994_178# vss 1.15f
C688 X1/X2/X1/X2/X1/X1/vin2 vss 1.74f
C689 X1/X2/X1/X3/vin1 vss 1.49f
C690 X1/X2/X1/X1/sw_0/m1_688_n494# vss 0.858f
C691 X1/X2/X1/X1/sw_0/m1_994_178# vss 1.15f
C692 X1/X2/X1/X1/X2/vout vss 0.868f
C693 X1/X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C694 X1/X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C695 X1/X2/X1/X1/X2/X2/vin1 vss 1.46f
C696 X1/X2/X1/X1/X2/X3/vin2 vss 1.23f
C697 X1/X2/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C698 X1/X2/X1/X1/X2/X2/m1_994_178# vss 1.15f
C699 X1/X2/X1/X2/vrefh vss 3.27f
C700 X1/X2/X1/X1/X2/X1/vin1 vss 1.91f
C701 X1/X2/X1/X1/X2/X3/vin1 vss 0.816f
C702 X1/X2/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C703 X1/X2/X1/X1/X2/X1/m1_994_178# vss 1.15f
C704 X1/X2/X1/X1/X2/X1/vin2 vss 1.74f
C705 X1/X2/X1/X1/X1/vout vss 0.607f
C706 X1/X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C707 X1/X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C708 X1/X2/X1/X1/X1/X2/vin1 vss 1.46f
C709 X1/X2/X1/X1/X1/X3/vin2 vss 1.23f
C710 X1/X2/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C711 X1/X2/X1/X1/X1/X2/m1_994_178# vss 1.15f
C712 X1/X2/X1/X1/X2/vrefh vss 3.27f
C713 X1/X2/X1/X1/X1/X1/vin1 vss 1.91f
C714 X1/X2/X1/X1/X1/X3/vin1 vss 0.816f
C715 X1/X2/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C716 X1/X2/X1/X1/X1/X1/m1_994_178# vss 1.15f
C717 X1/X2/X1/X1/X1/X1/vin2 vss 1.74f
C718 d4 vss 4.6f
C719 X1/X3/vin1 vss 1.12f
C720 X1/X1/X3/m1_688_n494# vss 0.858f
C721 X1/X1/X3/m1_994_178# vss 1.15f
C722 d3 vss 16.7f
C723 X1/X1/X3/vin2 vss 1.85f
C724 X1/X1/X2/X3/m1_688_n494# vss 0.858f
C725 X1/X1/X2/X3/m1_994_178# vss 1.15f
C726 d2 vss 24.8f
C727 X1/X1/X2/X3/vin2 vss 1.75f
C728 X1/X1/X2/X2/sw_0/m1_688_n494# vss 0.858f
C729 X1/X1/X2/X2/sw_0/m1_994_178# vss 1.15f
C730 X1/X1/X2/X2/X2/vout vss 0.868f
C731 X1/X1/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C732 X1/X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C733 d0 vss 72.9f
C734 X1/X1/X2/X2/X2/X2/vin1 vss 1.46f
C735 X1/X1/X2/X2/X2/X3/vin2 vss 1.23f
C736 X1/X1/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C737 X1/X1/X2/X2/X2/X2/m1_994_178# vss 1.15f
C738 X1/X2/vrefh vss 6.35f
C739 X1/X1/X2/X2/X2/X1/vin1 vss 1.91f
C740 X1/X1/X2/X2/X2/X3/vin1 vss 0.816f
C741 X1/X1/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C742 X1/X1/X2/X2/X2/X1/m1_994_178# vss 1.15f
C743 X1/X1/X2/X2/X2/X1/vin2 vss 1.73f
C744 X1/X1/X2/X2/X1/vout vss 0.607f
C745 X1/X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C746 X1/X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C747 X1/X1/X2/X2/X1/X2/vin1 vss 1.46f
C748 X1/X1/X2/X2/X1/X3/vin2 vss 1.23f
C749 X1/X1/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C750 X1/X1/X2/X2/X1/X2/m1_994_178# vss 1.15f
C751 X1/X1/X2/X2/X2/vrefh vss 3.27f
C752 X1/X1/X2/X2/X1/X1/vin1 vss 1.91f
C753 X1/X1/X2/X2/X1/X3/vin1 vss 0.816f
C754 X1/X1/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C755 X1/X1/X2/X2/X1/X1/m1_994_178# vss 1.15f
C756 X1/X1/X2/X2/X1/X1/vin2 vss 1.73f
C757 X1/X1/X2/X3/vin1 vss 1.49f
C758 X1/X1/X2/X1/sw_0/m1_688_n494# vss 0.858f
C759 X1/X1/X2/X1/sw_0/m1_994_178# vss 1.15f
C760 X1/X1/X2/X1/X2/vout vss 0.868f
C761 X1/X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C762 X1/X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C763 X1/X1/X2/X1/X2/X2/vin1 vss 1.46f
C764 X1/X1/X2/X1/X2/X3/vin2 vss 1.23f
C765 X1/X1/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C766 X1/X1/X2/X1/X2/X2/m1_994_178# vss 1.15f
C767 X1/X1/X2/X2/vrefh vss 3.27f
C768 X1/X1/X2/X1/X2/X1/vin1 vss 1.91f
C769 X1/X1/X2/X1/X2/X3/vin1 vss 0.816f
C770 X1/X1/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C771 X1/X1/X2/X1/X2/X1/m1_994_178# vss 1.15f
C772 X1/X1/X2/X1/X2/X1/vin2 vss 1.73f
C773 X1/X1/X2/X1/X1/vout vss 0.607f
C774 X1/X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C775 X1/X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C776 X1/X1/X2/X1/X1/X2/vin1 vss 1.46f
C777 X1/X1/X2/X1/X1/X3/vin2 vss 1.23f
C778 X1/X1/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C779 X1/X1/X2/X1/X1/X2/m1_994_178# vss 1.15f
C780 X1/X1/X2/X1/X2/vrefh vss 3.27f
C781 X1/X1/X2/X1/X1/X1/vin1 vss 1.91f
C782 X1/X1/X2/X1/X1/X3/vin1 vss 0.816f
C783 X1/X1/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C784 X1/X1/X2/X1/X1/X1/m1_994_178# vss 1.15f
C785 X1/X1/X2/X1/X1/X1/vin2 vss 1.73f
C786 X1/X1/X3/vin1 vss 1.6f
C787 X1/X1/X1/X3/m1_688_n494# vss 0.858f
C788 X1/X1/X1/X3/m1_994_178# vss 1.15f
C789 X1/X1/X1/X3/vin2 vss 1.75f
C790 X1/X1/X1/X2/sw_0/m1_688_n494# vss 0.858f
C791 X1/X1/X1/X2/sw_0/m1_994_178# vss 1.15f
C792 X1/X1/X1/X2/X2/vout vss 0.868f
C793 X1/X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C794 X1/X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C795 vdd vss 0.621p
C796 X1/X1/X1/X2/X2/X2/vin1 vss 1.46f
C797 X1/X1/X1/X2/X2/X3/vin2 vss 1.23f
C798 X1/X1/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C799 X1/X1/X1/X2/X2/X2/m1_994_178# vss 1.15f
C800 X1/X1/X2/vrefh vss 3.27f
C801 X1/X1/X1/X2/X2/X1/vin1 vss 1.91f
C802 X1/X1/X1/X2/X2/X3/vin1 vss 0.816f
C803 X1/X1/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C804 X1/X1/X1/X2/X2/X1/m1_994_178# vss 1.15f
C805 X1/X1/X1/X2/X2/X1/vin2 vss 1.73f
C806 X1/X1/X1/X2/X1/vout vss 0.607f
C807 X1/X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C808 X1/X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C809 X1/X1/X1/X2/X1/X2/vin1 vss 1.46f
C810 X1/X1/X1/X2/X1/X3/vin2 vss 1.23f
C811 X1/X1/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C812 X1/X1/X1/X2/X1/X2/m1_994_178# vss 1.15f
C813 X1/X1/X1/X2/X2/vrefh vss 3.27f
C814 X1/X1/X1/X2/X1/X1/vin1 vss 1.91f
C815 X1/X1/X1/X2/X1/X3/vin1 vss 0.816f
C816 X1/X1/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C817 X1/X1/X1/X2/X1/X1/m1_994_178# vss 1.15f
C818 X1/X1/X1/X2/X1/X1/vin2 vss 1.73f
C819 X1/X1/X1/X3/vin1 vss 1.49f
C820 X1/X1/X1/X1/sw_0/m1_688_n494# vss 0.858f
C821 X1/X1/X1/X1/sw_0/m1_994_178# vss 1.15f
C822 d1 vss 31.6f
C823 X1/X1/X1/X1/X2/vout vss 0.868f
C824 X1/X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C825 X1/X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C826 X1/X1/X1/X1/X2/X2/vin1 vss 1.46f
C827 X1/X1/X1/X1/X2/X3/vin2 vss 1.23f
C828 X1/X1/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C829 X1/X1/X1/X1/X2/X2/m1_994_178# vss 1.15f
C830 X1/X1/X1/X2/vrefh vss 3.27f
C831 X1/X1/X1/X1/X2/X1/vin1 vss 1.91f
C832 X1/X1/X1/X1/X2/X3/vin1 vss 0.816f
C833 X1/X1/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C834 X1/X1/X1/X1/X2/X1/m1_994_178# vss 1.15f
C835 X1/X1/X1/X1/X2/X1/vin2 vss 1.73f
C836 X1/X1/X1/X1/X1/vout vss 0.607f
C837 X1/X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C838 X1/X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C839 X1/X1/X1/X1/X1/X2/vin1 vss 1.46f
C840 X1/X1/X1/X1/X1/X3/vin2 vss 1.23f
C841 X1/X1/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C842 X1/X1/X1/X1/X1/X2/m1_994_178# vss 1.15f
C843 X1/X1/X1/X1/X2/vrefh vss 3.27f
C844 X1/X1/X1/X1/X1/X1/vin1 vss 1.91f
C845 X1/X1/X1/X1/X1/X3/vin1 vss 0.816f
C846 X1/X1/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C847 X1/X1/X1/X1/X1/X1/m1_994_178# vss 1.15f
C848 X1/X1/X1/X1/X1/X1/vin2 vss 1.73f
C849 vrefh vss 1.11f
.ends

.subckt x8bit_dac vrefh vrefl d0 d1 d2 d3 d4 d5 d6 d7 vout vss vdd
XX1 d2 d4 d6 X3/vin1 X1/X2/X2/X1/X2/X1/X1/vin1 X1/X1/X1/X2/X1/X2/vrefh X1/X2/X2/X1/X2/X1/X2/vin1
+ X1/X3/vin1 X1/X1/X2/X2/X2/X2/X3/vin2 X1/X2/X2/X2/X1/X1/X1/vin1 X1/X1/X1/X1/X1/X2/X1/vin1
+ X1/X2/X2/X1/X1/X1/X1/m1_994_178# X1/X2/X2/X2/X1/X1/X2/vin1 X1/X2/X2/X1/X1/X1/X1/m1_688_n494#
+ X1/X1/X1/X1/X2/X1/X1/vin2 X1/X1/X1/X1/X1/X2/X2/vin1 X1/X2/X2/X1/X1/X2/X1/vin2 X1/X2/X2/X1/X2/X2/vrefh
+ X1/X2/X2/X2/X2/X1/X1/vin1 X1/X2/X2/X2/X2/X2/vrefh X1/X1/X1/X1/X1/X1/X1/m1_688_n494#
+ X1/X2/X3/m1_688_n494# X1/X1/X1/X1/X2/X2/X1/vin1 X1/X2/X2/X2/X2/X2/X1/vin2 X1/X2/X2/X2/X2/X1/X2/vin1
+ X1/X1/X1/X1/X1/X1/X1/vin1 X1/X1/X1/X1/X2/X2/X2/vin1 X1/X1/X1/X2/X1/X2/X1/vin2 X1/X1/X1/X2/X1/X2/X1/vin1
+ X1/X2/X2/X2/X2/X2/X1/vin1 X1/X1/X1/X1/X2/X2/vrefh X1/X1/X1/X2/X1/X2/X2/vin1 X1/X1/X1/X2/X2/X2/vrefh
+ X1/X3/vin2 X1/X2/X2/X2/X1/X1/X1/vin2 X1/X2/X2/vrefh X1/X1/X3/m1_994_178# X1/X1/X1/X1/X2/X2/X1/vin2
+ X1/X1/X1/X1/X2/X1/X1/vin1 X1/X1/X1/X2/X2/X2/X1/vin1 X1/X1/X1/X1/X1/X1/X3/m1_994_178#
+ X1/X2/X2/X1/X2/vrefh X1/X1/X1/X1/X1/X1/X3/m1_688_n494# X1/X1/X1/X2/X2/vrefh X1/X1/X1/X1/X2/X1/X2/vin1
+ X1/X1/X1/X2/X2/X2/X2/vin1 X1/X1/X1/X2/X1/X1/X1/vin1 X1/X1/X1/X1/X1/X1/X2/vin1 X1/X2/X2/X1/X2/X1/X1/vin2
+ X1/X1/X1/X1/X1/X1/X1/vin2 X1/X1/X1/X2/X1/X1/X2/vin1 X1/X1/X3/vin2 X1/X2/X2/X2/X2/X2/X2/m1_994_178#
+ X1/X1/X3/vin1 X1/X2/X2/X2/X2/X2/X2/m1_688_n494# X1/X1/X2/X2/X2/X2/X2/m1_994_178#
+ X2/vrefh X1/X1/X2/X2/X2/X2/X2/m1_688_n494# X1/X2/X2/X2/X2/X2/X2/vin1 d1 X1/X1/X1/X2/X2/X1/X1/vin1
+ X1/X1/X1/X2/X2/X1/X1/vin2 X1/X1/X3/m1_688_n494# X1/X2/X2/X2/X1/X2/X1/vin2 X1/X3/m1_994_178#
+ X1/X1/X1/X2/X2/X1/X2/vin1 X1/X2/X2/X1/X1/X2/X1/vin1 X1/X2/X2/X1/X1/X2/X2/vin1 X1/X2/X2/X2/X2/vrefh
+ X1/X2/X2/X1/X2/X2/X1/vin2 X1/X1/X1/X1/X1/X2/X1/vin2 X1/X2/X3/vin2 X1/X1/X1/X1/X1/X1/X3/vin1
+ X1/X1/X2/X2/X2/X2/X2/vin1 X1/X2/X3/vin1 X1/X2/X2/X1/X2/X2/X1/vin1 X1/X2/X2/X2/vrefh
+ X1/X2/X2/X1/X1/X1/X1/vin2 X1/X2/X2/X2/X1/X2/X1/vin1 X1/X2/X2/X1/X2/X2/X2/vin1 X1/X2/X2/X1/X1/X1/X1/vin1
+ X1/X2/X2/X2/X2/X2/X3/vin2 X1/X2/X2/X1/X1/X2/vrefh X1/X1/X1/X2/X2/X2/X1/vin2 X1/X1/X1/X2/X2/X2/X2/m1_994_178#
+ X1/X3/m1_688_n494# X1/X1/X1/X2/X2/X2/X2/m1_688_n494# d5 X1/X2/X2/X2/X1/X2/vrefh
+ X1/X2/X2/X2/X1/X2/X2/vin1 X1/X2/X2/X1/X1/X1/X2/vin1 vdd X1/X2/X1/X1/X1/X1/X1/vin2
+ d3 X1/X1/X1/X1/X1/X1/X1/m1_994_178# vrefh X1/X2/X3/m1_994_178# X1/X2/X1/X1/X1/X1/X1/vin1
+ X1/X2/X2/X2/X2/X1/X1/vin2 X1/X1/X2/vrefh X1/X2/vrefh vss X1/X1/X1/X2/vrefh X1/X1/X1/X1/X1/X2/vrefh
+ d0 X1/X1/X1/X1/X2/vrefh X1/X1/X1/X2/X1/X1/X1/vin2 x7bit_dac
XX2 d2 d4 d6 X3/vin2 X2/X2/X2/X1/X2/X1/X1/vin1 X2/X1/X1/X2/X1/X2/vrefh X2/X2/X2/X1/X2/X1/X2/vin1
+ X2/X3/vin1 X2/X1/X2/X2/X2/X2/X3/vin2 X2/X2/X2/X2/X1/X1/X1/vin1 X2/X1/X1/X1/X1/X2/X1/vin1
+ X2/X2/X2/X1/X1/X1/X1/m1_994_178# X2/X2/X2/X2/X1/X1/X2/vin1 X2/X2/X2/X1/X1/X1/X1/m1_688_n494#
+ X2/X1/X1/X1/X2/X1/X1/vin2 X2/X1/X1/X1/X1/X2/X2/vin1 X2/X2/X2/X1/X1/X2/X1/vin2 X2/X2/X2/X1/X2/X2/vrefh
+ X2/X2/X2/X2/X2/X1/X1/vin1 X2/X2/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X1/X1/X1/m1_688_n494#
+ X2/X2/X3/m1_688_n494# X2/X1/X1/X1/X2/X2/X1/vin1 X2/X2/X2/X2/X2/X2/X1/vin2 X2/X2/X2/X2/X2/X1/X2/vin1
+ X2/X1/X1/X1/X1/X1/X1/vin1 X2/X1/X1/X1/X2/X2/X2/vin1 X2/X1/X1/X2/X1/X2/X1/vin2 X2/X1/X1/X2/X1/X2/X1/vin1
+ X2/X2/X2/X2/X2/X2/X1/vin1 X2/X1/X1/X1/X2/X2/vrefh X2/X1/X1/X2/X1/X2/X2/vin1 X2/X1/X1/X2/X2/X2/vrefh
+ X2/X3/vin2 X2/X2/X2/X2/X1/X1/X1/vin2 X2/X2/X2/vrefh X2/X1/X3/m1_994_178# X2/X1/X1/X1/X2/X2/X1/vin2
+ X2/X1/X1/X1/X2/X1/X1/vin1 X2/X1/X1/X2/X2/X2/X1/vin1 X2/X1/X1/X1/X1/X1/X3/m1_994_178#
+ X2/X2/X2/X1/X2/vrefh X2/X1/X1/X1/X1/X1/X3/m1_688_n494# X2/X1/X1/X2/X2/vrefh X2/X1/X1/X1/X2/X1/X2/vin1
+ X2/X1/X1/X2/X2/X2/X2/vin1 X2/X1/X1/X2/X1/X1/X1/vin1 X2/X1/X1/X1/X1/X1/X2/vin1 X2/X2/X2/X1/X2/X1/X1/vin2
+ X2/X1/X1/X1/X1/X1/X1/vin2 X2/X1/X1/X2/X1/X1/X2/vin1 X2/X1/X3/vin2 X2/X2/X2/X2/X2/X2/X2/m1_994_178#
+ X2/X1/X3/vin1 X2/X2/X2/X2/X2/X2/X2/m1_688_n494# X2/X1/X2/X2/X2/X2/X2/m1_994_178#
+ vrefl X2/X1/X2/X2/X2/X2/X2/m1_688_n494# X2/X2/X2/X2/X2/X2/X2/vin1 d1 X2/X1/X1/X2/X2/X1/X1/vin1
+ X2/X1/X1/X2/X2/X1/X1/vin2 X2/X1/X3/m1_688_n494# X2/X2/X2/X2/X1/X2/X1/vin2 X2/X3/m1_994_178#
+ X2/X1/X1/X2/X2/X1/X2/vin1 X2/X2/X2/X1/X1/X2/X1/vin1 X2/X2/X2/X1/X1/X2/X2/vin1 X2/X2/X2/X2/X2/vrefh
+ X2/X2/X2/X1/X2/X2/X1/vin2 X2/X1/X1/X1/X1/X2/X1/vin2 X2/X2/X3/vin2 X2/X1/X1/X1/X1/X1/X3/vin1
+ X2/X1/X2/X2/X2/X2/X2/vin1 X2/X2/X3/vin1 X2/X2/X2/X1/X2/X2/X1/vin1 X2/X2/X2/X2/vrefh
+ X2/X2/X2/X1/X1/X1/X1/vin2 X2/X2/X2/X2/X1/X2/X1/vin1 X2/X2/X2/X1/X2/X2/X2/vin1 X2/X2/X2/X1/X1/X1/X1/vin1
+ X2/X2/X2/X2/X2/X2/X3/vin2 X2/X2/X2/X1/X1/X2/vrefh X2/X1/X1/X2/X2/X2/X1/vin2 X2/X1/X1/X2/X2/X2/X2/m1_994_178#
+ X2/X3/m1_688_n494# X2/X1/X1/X2/X2/X2/X2/m1_688_n494# d5 X2/X2/X2/X2/X1/X2/vrefh
+ X2/X2/X2/X2/X1/X2/X2/vin1 X2/X2/X2/X1/X1/X1/X2/vin1 vdd X2/X2/X1/X1/X1/X1/X1/vin2
+ d3 X2/X1/X1/X1/X1/X1/X1/m1_994_178# X2/vrefh X2/X2/X3/m1_994_178# X2/X2/X1/X1/X1/X1/X1/vin1
+ X2/X2/X2/X2/X2/X1/X1/vin2 X2/X1/X2/vrefh X2/X2/vrefh vss X2/X1/X1/X2/vrefh X2/X1/X1/X1/X1/X2/vrefh
+ d0 X2/X1/X1/X1/X2/vrefh X2/X1/X1/X2/X1/X1/X1/vin2 x7bit_dac
XX3 X3/vin1 X3/vin2 vout vdd d7 X3/m1_688_n494# vss X3/m1_994_178# sw
X0 X1/X2/X1/X1/X2/X1/X1/m1_994_178# d0.t73 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X1 X2/X1/X1/X2/X1/X2/X3/m1_994_178# d1.t75 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X2 X1/X2/X1/X2/X2/X2/X2/m1_994_178# d0.t95 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X3 X2/X2/X2/X1/X2/X1/X2/m1_994_178# d0.t235 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X4 X1/X2/X2/X1/X2/X2/X2/m1_994_178# d0.t111 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X5 X1/X1/X3/m1_994_178# d5.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X6 X1/X1/X2/X2/X2/X1/X1/m1_994_178# d0.t57 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X7 X2/X2/X1/X1/X1/X2/X3/m1_994_178# d1.t99 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X8 X2/X2/X2/X2/X2/X2/X1/m1_994_178# d0.t253 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X9 X1/X2/X1/X1/X2/X2/X2/m1_994_178# d0.t79 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X10 X2/X2/X1/X1/X2/X2/X3/m1_994_178# d1.t103 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X11 X2/X1/X2/X3/m1_994_178# d4.t11 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X12 X1/X1/X2/X1/X1/sw_0/m1_994_178# d2.t9 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X13 X2/X2/X2/X1/X1/X1/X1/m1_994_178# d0.t225 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X14 X1/X1/X2/X2/X2/X2/X3/m1_994_178# d1.t31 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X15 X2/X2/X2/X1/X1/sw_0/m1_994_178# d2.t57 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X16 X2/X1/X1/X1/X2/X2/X1/m1_994_178# d0.t141 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X17 X1/X1/X1/X2/X1/X1/X1/m1_994_178# d0.t17 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X18 X2/X1/X1/X1/X2/X1/X3/m1_994_178# d1.t69 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X19 X2/X2/X1/X2/X1/X2/X2/m1_994_178# d0.t215 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X20 X2/X1/X1/X1/X1/X1/X1/m1_994_178# d0.t129 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X21 X1/X2/X1/X2/X1/X2/X3/m1_994_178# d1.t43 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X22 X1/X2/X2/X2/X2/X1/X2/m1_994_178# d0.t123 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X23 X1/X1/X1/X1/X1/X2/X1/m1_994_178# d0.t5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X24 X2/X1/X1/X2/X2/X1/X2/m1_994_178# d0.t155 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X25 X2/X1/X2/X1/X1/X1/X3/m1_994_178# d1.t81 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X26 X2/X1/X2/X1/X1/X1/X1/m1_994_178# d0.t161 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X27 X2/X2/X3/m1_994_178# d5.t7 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X28 X2/X1/X1/X2/X1/X1/X2/m1_994_178# d0.t147 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X29 X1/X2/X2/X2/X1/X1/X1/m1_994_178# d0.t113 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X30 X2/X2/X2/X1/X2/X2/X3/m1_994_178# d1.t119 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X31 X1/X1/X2/X1/X2/sw_0/m1_994_178# d2.t11 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X32 X1/X1/X2/X1/X1/X2/X3/m1_994_178# d1.t19 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X33 X1/X2/X1/X3/m1_994_178# d4.t5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X34 X2/X2/X2/X1/X1/X2/X3/m1_994_178# d1.t115 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X35 X1/X2/X1/X2/X3/m1_994_178# d3.t11 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X36 X1/X2/X1/X2/X2/X1/X1/m1_994_178# d0.t89 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X37 X2/X1/X2/X1/X2/X1/X1/m1_994_178# d0.t169 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X38 X2/X2/X1/X2/X2/X1/X2/m1_994_178# d0.t219 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X39 X2/X2/X2/X2/X1/X2/X2/m1_994_178# d0.t247 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X40 X1/X1/X1/X1/X2/sw_0/m1_994_178# d2.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X41 X1/X2/X2/X2/X1/sw_0/m1_994_178# d2.t29 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X42 X2/X1/X1/X3/m1_994_178# d4.t9 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X43 X1/X2/X1/X1/X2/X2/X1/m1_994_178# d0.t77 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X44 X2/X1/X1/X2/X3/m1_994_178# d3.t19 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X45 X2/X2/X2/X1/X1/X2/X2/m1_994_178# d0.t231 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X46 X2/X2/X1/X1/X2/X1/X2/m1_994_178# d0.t203 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X47 X1/X2/X2/X1/X2/X1/X2/m1_994_178# d0.t107 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X48 X1/X2/X2/X1/X1/X1/X1/m1_994_178# d0.t97 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X49 X1/X2/X1/X1/X2/X1/X3/m1_994_178# d1.t37 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X50 X1/X2/X2/X2/X3/m1_994_178# d3.t15 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X51 X1/X2/X1/X1/X1/X1/X1/m1_994_178# d0.t65 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X52 X2/X1/X1/X2/X2/X2/X2/m1_994_178# d0.t159 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X53 X2/X2/X1/X1/X3/m1_994_178# d3.t25 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X54 X1/X2/X2/X2/X2/X2/X1/m1_994_178# d0.t125 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X55 X1/X2/X1/X2/X1/X1/X2/m1_994_178# d0.t83 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X56 X1/X1/X1/X1/X1/X1/X2/m1_994_178# d0.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X57 X2/X2/X2/X2/X2/X1/X3/m1_994_178# d1.t125 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X58 X1/X1/X2/X2/X1/X1/X2/m1_994_178# d0.t51 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X59 X1/X2/X1/X2/X2/X1/X3/m1_994_178# d1.t45 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X60 X2/X1/X2/X1/X2/X2/X3/m1_994_178# d1.t87 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X61 X2/X1/X2/X2/X1/X2/X1/m1_994_178# d0.t181 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X62 X2/X1/X1/X1/X1/X2/X3/m1_994_178# d1.t67 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X63 X2/X2/X1/X1/X1/sw_0/m1_994_178# d2.t49 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X64 X2/X1/X1/X1/X2/X2/X3/m1_994_178# d1.t71 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X65 X1/X2/X2/X3/m1_994_178# d4.t7 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X66 X1/X1/X1/X2/X1/X1/X3/m1_994_178# d1.t9 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X67 X1/X2/X2/X1/X1/X2/X3/m1_994_178# d1.t51 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X68 X2/X2/X1/X2/X2/X2/X2/m1_994_178# d0.t223 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X69 X2/X1/X3/m1_994_178# d5.t5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X70 X1/X1/X2/X1/X2/X2/X1/m1_994_178# d0.t45 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X71 X2/X1/X2/X1/X2/X2/X2/m1_994_178# d0.t175 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X72 X2/X1/X1/X2/X1/X2/X2/m1_994_178# d0.t151 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X73 X2/X2/X2/X1/X3/m1_994_178# d3.t29 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X74 X1/X1/X2/X2/X1/X1/X3/m1_994_178# d1.t25 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X75 X2/X2/X2/X1/X2/X1/X3/m1_994_178# d1.t117 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X76 X1/X2/X2/X1/X2/X2/X3/m1_994_178# d1.t55 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X77 X1/X1/X1/X2/X2/X1/X2/m1_994_178# d0.t27 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X78 X1/X1/X2/X1/X1/X1/X3/m1_994_178# d1.t17 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X79 X2/X2/X2/X1/X1/X1/X3/m1_994_178# d1.t113 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X80 X2/X1/X2/X2/X2/X1/X3/m1_994_178# d1.t93 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X81 X2/X2/X1/X2/X1/sw_0/m1_994_178# d2.t53 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X82 X1/X2/X2/X2/X1/X2/X2/m1_994_178# d0.t119 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X83 X1/X1/X1/X1/X2/X1/X1/m1_994_178# d0.t9 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X84 X1/X2/X1/X2/X2/X2/X3/m1_994_178# d1.t47 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X85 X2/X2/X1/X1/X1/X2/X2/m1_994_178# d0.t199 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X86 X1/X2/X1/X1/X1/X2/X3/m1_994_178# d1.t35 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X87 X1/X2/X2/X1/X1/X2/X2/m1_994_178# d0.t103 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X88 X2/X1/X1/X2/X2/X1/X1/m1_994_178# d0.t153 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X89 X1/X2/X1/X1/X2/X2/X3/m1_994_178# d1.t39 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X90 X2/X2/X2/X2/X2/X2/X2/m1_994_178# d0.t255 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X91 X1/X2/X1/X2/X2/X2/X1/m1_994_178# d0.t93 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X92 X2/X1/X1/X1/X2/X1/X2/m1_994_178# d0.t139 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X93 X2/X1/X2/X2/X2/X1/X2/m1_994_178# d0.t187 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X94 X1/X1/X1/X1/X2/X2/X2/m1_994_178# d0.t15 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X95 X1/X1/X2/X2/X1/sw_0/m1_994_178# d2.t13 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X96 X2/X2/X2/X2/X2/sw_0/m1_994_178# d2.t63 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X97 X1/X2/X1/X2/X1/X2/X2/m1_994_178# d0.t87 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X98 X1/X2/X1/X1/X3/m1_994_178# d3.t9 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X99 X1/X2/X2/X2/X2/X1/X3/m1_994_178# d1.t61 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X100 X2/X3/m1_994_178# d6.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X101 X2/X1/X2/X1/X3/m1_994_178# d3.t21 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X102 X2/X1/X2/X1/X2/X1/X3/m1_994_178# d1.t85 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X103 X2/X2/X1/X2/X1/X2/X1/m1_994_178# d0.t213 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X104 X2/X2/X1/X2/X2/X1/X1/m1_994_178# d0.t217 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X105 X2/X2/X2/X2/X2/X1/X1/m1_994_178# d0.t249 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X106 X2/X1/X2/X2/X1/X1/X1/m1_994_178# d0.t177 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X107 X1/X1/X1/X2/X2/X2/X2/m1_994_178# d0.t31 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X108 X2/X2/X1/X1/X1/X1/X3/m1_994_178# d1.t97 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X109 X1/X1/X2/X2/X3/m1_994_178# d3.t7 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X110 X2/X1/X1/X1/X3/m1_994_178# d3.t17 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X111 X1/X2/X1/X1/X1/sw_0/m1_994_178# d2.t17 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X112 X1/X1/X1/X2/X1/X2/X3/m1_994_178# d1.t11 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X113 X1/X1/X2/X1/X1/X1/X2/m1_994_178# d0.t35 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X114 X1/X2/X2/X1/X1/X1/X3/m1_994_178# d1.t49 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X115 X2/X1/X1/X2/X2/X1/X3/m1_994_178# d1.t77 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X116 X2/X1/X1/X1/X1/sw_0/m1_994_178# d2.t33 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X117 X1/X1/X2/X1/X2/X1/X1/m1_994_178# d0.t41 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X118 X2/X2/X2/X2/X1/X2/X3/m1_994_178# d1.t123 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X119 X2/X1/X2/X1/X2/X1/X2/m1_994_178# d0.t171 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X120 X1/X2/X2/X1/X2/X1/X3/m1_994_178# d1.t53 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X121 X1/X2/X1/X1/X2/X1/X2/m1_994_178# d0.t75 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X122 X1/X1/X2/X3/m1_994_178# d4.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X123 X2/X2/X1/X2/X2/X1/X3/m1_994_178# d1.t109 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X124 X2/X1/X2/X2/X2/sw_0/m1_994_178# d2.t47 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X125 X1/X2/X1/X2/X1/sw_0/m1_994_178# d2.t21 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X126 X2/X1/X2/X2/X2/X2/X1/m1_994_178# d0.t189 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X127 X1/X1/X1/X1/X2/X2/X1/m1_994_178# d0.t13 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X128 X1/X1/X1/X1/X2/X1/X3/m1_994_178# d1.t5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X129 X2/X1/X1/X2/X1/sw_0/m1_994_178# d2.t37 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X130 X1/X2/X2/X2/X2/X2/X2/m1_994_178# d0.t127 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X131 X1/X1/X1/X1/X1/X1/X1/m1_994_178# d0.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X132 X1/X1/X2/X2/X1/X2/X1/m1_994_178# d0.t53 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X133 X2/X1/X1/X1/X1/X2/X2/m1_994_178# d0.t135 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X134 X2/X1/X1/X2/X2/X2/X3/m1_994_178# d1.t79 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X135 X2/X1/X2/X2/X1/X2/X3/m1_994_178# d1.t91 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X136 X1/X1/X1/X2/X1/X1/X2/m1_994_178# d0.t19 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X137 X1/X1/X1/X2/X2/X1/X1/m1_994_178# d0.t25 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X138 X2/X2/X1/X2/X1/X1/X1/m1_994_178# d0.t209 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X139 X3/m1_994_178# d7.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X140 X1/X2/X2/X2/X2/X1/X1/m1_994_178# d0.t121 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X141 X2/X1/X1/X2/X2/X2/X1/m1_994_178# d0.t157 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X142 X1/X1/X2/X1/X2/X2/X2/m1_994_178# d0.t47 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X143 X2/X2/X1/X1/X1/X2/X1/m1_994_178# d0.t197 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X144 X1/X1/X1/X3/m1_994_178# d4.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X145 X2/X2/X1/X2/X2/X2/X3/m1_994_178# d1.t111 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X146 X2/X2/X2/X2/X1/X1/X2/m1_994_178# d0.t243 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X147 X1/X2/X2/X1/X3/m1_994_178# d3.t13 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X148 X2/X1/X1/X2/X1/X2/X1/m1_994_178# d0.t149 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X149 X1/X1/X1/X2/X3/m1_994_178# d3.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X150 X2/X1/X2/X2/X1/X2/X2/m1_994_178# d0.t183 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X151 X2/X1/X1/X1/X1/X1/X3/m1_994_178# d1.t65 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X152 X2/X1/X1/X2/X2/sw_0/m1_994_178# d2.t39 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X153 X1/X2/X2/X2/X1/X2/X3/m1_994_178# d1.t59 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X154 X2/X1/X2/X1/X1/X2/X2/m1_994_178# d0.t167 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X155 X2/X2/X1/X2/X2/X2/X1/m1_994_178# d0.t221 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X156 X1/X2/X1/X1/X1/X2/X2/m1_994_178# d0.t71 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X157 X1/X1/X1/X2/X2/X1/X3/m1_994_178# d1.t13 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X158 X2/X2/X2/X1/X1/X1/X2/m1_994_178# d0.t227 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X159 X2/X2/X1/X1/X2/sw_0/m1_994_178# d2.t51 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X160 X2/X2/X2/X1/X2/X2/X1/m1_994_178# d0.t237 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X161 X2/X2/X2/X2/X2/X2/X3/m1_994_178# d1.t127 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X162 X1/X1/X2/X1/X2/X2/X3/m1_994_178# d1.t23 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X163 X2/X2/X1/X2/X2/sw_0/m1_994_178# d2.t55 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X164 X1/X1/X1/X1/X1/X2/X3/m1_994_178# d1.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X165 X1/X1/X2/X2/X2/X1/X2/m1_994_178# d0.t59 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X166 X1/X1/X1/X1/X2/X2/X3/m1_994_178# d1.t7 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X167 X2/X1/X2/X1/X1/X1/X2/m1_994_178# d0.t163 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X168 X1/X2/X2/X2/X2/sw_0/m1_994_178# d2.t31 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X169 X1/X2/X1/X2/X1/X2/X1/m1_994_178# d0.t85 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X170 X1/X1/X2/X2/X1/X1/X1/m1_994_178# d0.t49 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X171 X2/X2/X1/X1/X1/X1/X2/m1_994_178# d0.t195 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X172 X1/X2/X1/X1/X1/X1/X3/m1_994_178# d1.t33 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X173 X2/X2/X2/X1/X2/sw_0/m1_994_178# d2.t59 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X174 X1/X1/X1/X2/X1/X2/X2/m1_994_178# d0.t23 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X175 X1/X1/X2/X1/X1/X2/X1/m1_994_178# d0.t37 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X176 X1/X1/X1/X2/X2/X2/X3/m1_994_178# d1.t15 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X177 X2/X2/X1/X2/X1/X1/X3/m1_994_178# d1.t105 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X178 X2/X1/X2/X2/X2/X2/X3/m1_994_178# d1.t95 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X179 X1/X1/X2/X2/X2/X1/X3/m1_994_178# d1.t29 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X180 X1/X1/X2/X1/X2/X1/X2/m1_994_178# d0.t43 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X181 X2/X1/X1/X2/X1/X1/X1/m1_994_178# d0.t145 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X182 X1/X2/X2/X1/X1/X1/X2/m1_994_178# d0.t99 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X183 X1/X2/X2/X2/X1/X1/X2/m1_994_178# d0.t115 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X184 X1/X1/X1/X2/X2/X2/X1/m1_994_178# d0.t29 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X185 X2/X1/X1/X1/X1/X2/X1/m1_994_178# d0.t133 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X186 X1/X2/X1/X2/X2/sw_0/m1_994_178# d2.t23 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X187 X1/X1/X2/X2/X2/X2/X1/m1_994_178# d0.t61 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X188 X1/X1/X1/X1/X2/X1/X2/m1_994_178# d0.t11 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X189 X2/X1/X2/X2/X2/X2/X2/m1_994_178# d0.t191 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X190 X1/X2/X1/X1/X2/sw_0/m1_994_178# d2.t19 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X191 X2/X2/X2/X1/X2/X1/X1/m1_994_178# d0.t233 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X192 X2/X2/X1/X1/X2/X1/X1/m1_994_178# d0.t201 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X193 X1/X2/X2/X1/X2/X2/X1/m1_994_178# d0.t109 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X194 X1/X2/X2/X2/X2/X2/X3/m1_994_178# d1.t63 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X195 X2/X1/X2/X1/X2/sw_0/m1_994_178# d2.t43 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X196 X1/X1/X1/X2/X2/sw_0/m1_994_178# d2.t7 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X197 X1/X1/X2/X1/X3/m1_994_178# d3.t5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X198 X1/X1/X2/X1/X2/X1/X3/m1_994_178# d1.t21 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X199 X2/X1/X1/X1/X2/sw_0/m1_994_178# d2.t35 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X200 X1/X1/X1/X1/X3/m1_994_178# d3.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X201 X2/X1/X2/X2/X2/X1/X1/m1_994_178# d0.t185 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X202 X1/X3/m1_994_178# d6.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X203 X1/X2/X1/X2/X1/X1/X1/m1_994_178# d0.t81 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X204 X2/X2/X1/X1/X2/X2/X2/m1_994_178# d0.t207 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X205 X1/X1/X1/X1/X1/sw_0/m1_994_178# d2.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X206 X2/X2/X2/X2/X1/X1/X3/m1_994_178# d1.t121 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X207 X1/X2/X1/X1/X1/X2/X1/m1_994_178# d0.t69 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X208 X2/X2/X2/X2/X1/X2/X1/m1_994_178# d0.t245 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X209 X1/X1/X2/X2/X1/X2/X2/m1_994_178# d0.t55 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X210 X2/X1/X1/X1/X1/X1/X2/m1_994_178# d0.t131 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X211 X2/X2/X1/X2/X1/X2/X3/m1_994_178# d1.t107 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X212 X1/X2/X2/X1/X1/sw_0/m1_994_178# d2.t25 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X213 X1/X1/X2/X2/X2/sw_0/m1_994_178# d2.t15 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X214 X1/X1/X2/X1/X1/X2/X2/m1_994_178# d0.t39 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X215 X2/X1/X1/X2/X1/X1/X3/m1_994_178# d1.t73 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X216 X2/X2/X2/X1/X1/X2/X1/m1_994_178# d0.t229 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X217 X2/X2/X2/X1/X2/X2/X2/m1_994_178# d0.t239 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X218 X1/X1/X1/X2/X1/sw_0/m1_994_178# d2.t5 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X219 X1/X1/X2/X1/X1/X1/X1/m1_994_178# d0.t33 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X220 X1/X2/X3/m1_994_178# d5.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X221 X1/X1/X1/X1/X1/X2/X2/m1_994_178# d0.t7 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X222 X2/X1/X2/X1/X1/sw_0/m1_994_178# d2.t41 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X223 X2/X2/X2/X2/X1/sw_0/m1_994_178# d2.t61 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X224 X1/X1/X2/X2/X1/X2/X3/m1_994_178# d1.t27 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X225 X2/X2/X1/X1/X2/X2/X1/m1_994_178# d0.t205 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X226 X2/X1/X2/X2/X1/X1/X3/m1_994_178# d1.t89 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X227 X1/X2/X2/X1/X2/X1/X1/m1_994_178# d0.t105 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X228 X2/X1/X2/X1/X1/X2/X1/m1_994_178# d0.t165 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X229 X2/X2/X1/X1/X2/X1/X3/m1_994_178# d1.t101 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X230 X2/X2/X2/X2/X3/m1_994_178# d3.t31 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X231 X1/X2/X1/X1/X1/X1/X2/m1_994_178# d0.t67 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X232 X1/X2/X1/X2/X2/X1/X2/m1_994_178# d0.t91 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X233 X2/X2/X1/X1/X1/X1/X1/m1_994_178# d0.t193 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X234 X2/X1/X1/X1/X2/X1/X1/m1_994_178# d0.t137 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X235 X1/X2/X2/X1/X2/sw_0/m1_994_178# d2.t27 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X236 X1/X1/X1/X2/X1/X2/X1/m1_994_178# d0.t21 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X237 X2/X2/X1/X2/X1/X1/X2/m1_994_178# d0.t211 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X238 X2/X2/X2/X2/X2/X1/X2/m1_994_178# d0.t251 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X239 X1/X2/X1/X2/X1/X1/X3/m1_994_178# d1.t41 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X240 X1/X1/X1/X1/X1/X1/X3/m1_994_178# d1.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X241 X2/X1/X2/X2/X1/X1/X2/m1_994_178# d0.t179 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X242 X2/X1/X2/X1/X1/X2/X3/m1_994_178# d1.t83 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X243 X1/X2/X2/X2/X1/X1/X3/m1_994_178# d1.t57 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X244 X2/X1/X1/X1/X2/X2/X2/m1_994_178# d0.t143 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X245 X1/X2/X2/X1/X1/X2/X1/m1_994_178# d0.t101 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X246 X2/X2/X2/X2/X1/X1/X1/m1_994_178# d0.t241 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X247 X2/X2/X2/X3/m1_994_178# d4.t15 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X248 X1/X2/X2/X2/X1/X2/X1/m1_994_178# d0.t117 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X249 X2/X1/X2/X2/X1/sw_0/m1_994_178# d2.t45 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X250 X2/X2/X1/X3/m1_994_178# d4.t13 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X251 X2/X2/X1/X2/X3/m1_994_178# d3.t27 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X252 X2/X1/X2/X1/X2/X2/X1/m1_994_178# d0.t173 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X253 X1/X1/X2/X2/X2/X2/X2/m1_994_178# d0.t63 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
X254 X2/X1/X2/X2/X3/m1_994_178# d3.t23 vss vss sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0 l=0
R0 vrefh vrefh 0.0502685
R1 vrefh vrefh 0.0138102
R2 vrefh vrefh 0.00918056
R3 vrefh vrefh 0.00281481
R4 vrefh vrefh 0.00165741
R5 vrefh vrefh 0.0010787
R6 vss.n15545 vss.n378 183359
R7 vss.n14871 vss.n14870 183359
R8 vss.n9441 vss.n9282 94793.4
R9 vss.n4577 vss.n435 94793.4
R10 vss.n2295 vss.n1214 94793.4
R11 vss.n6252 vss.n6251 94793.4
R12 vss.n12236 vss.n12235 75056.3
R13 vss.n12354 vss.n12353 75056.3
R14 vss.n12473 vss.n12472 75056.3
R15 vss.n6333 vss.n6332 75056.3
R16 vss.n5961 vss.n5960 75056.3
R17 vss.n6200 vss.n6199 75056.3
R18 vss.n5294 vss.n3534 75056.3
R19 vss.n5962 vss.n4001 75056.3
R20 vss.n6201 vss.n3993 75056.3
R21 vss.n7488 vss.n7487 75056.3
R22 vss.n7271 vss.n7270 75056.3
R23 vss.n15094 vss.n986 75056.3
R24 vss.n7490 vss.n7489 75056.3
R25 vss.n7224 vss.n3130 75056.3
R26 vss.n13953 vss.n13952 75056.3
R27 vss.n14070 vss.n14069 75056.3
R28 vss.n14399 vss.n1765 75056.3
R29 vss.n13954 vss.n8223 75056.3
R30 vss.n14071 vss.n8095 75056.3
R31 vss.n14398 vss.n14397 75056.3
R32 vss.n15093 vss.n15092 75056.3
R33 vss.n12237 vss.n9803 75056.3
R34 vss.n12355 vss.n9674 75056.3
R35 vss.n12474 vss.n9545 75056.3
R36 vss.n12905 vss.n9282 64989.1
R37 vss.n6271 vss.n6252 64989.1
R38 vss.n15461 vss.n435 64989.1
R39 vss.n14766 vss.n1214 64989.1
R40 vss.n14870 vss.n14849 62700.1
R41 vss.n15545 vss.n15544 62700.1
R42 vss.n14178 vss.n14177 61403.9
R43 vss.n12236 vss.n9851 60091.4
R44 vss.n12354 vss.n9723 60091.4
R45 vss.n12473 vss.n9593 60091.4
R46 vss.n6333 vss.n3535 60091.4
R47 vss.n5961 vss.n5912 60091.4
R48 vss.n6200 vss.n6151 60091.4
R49 vss.n3534 vss.n3488 60091.4
R50 vss.n5962 vss.n4000 60091.4
R51 vss.n6201 vss.n3992 60091.4
R52 vss.n7488 vss.n7439 60091.4
R53 vss.n7270 vss.n7269 60091.4
R54 vss.n15094 vss.n985 60091.4
R55 vss.n7489 vss.n3012 60091.4
R56 vss.n7224 vss.n3129 60091.4
R57 vss.n13953 vss.n13904 60091.4
R58 vss.n14070 vss.n8143 60091.4
R59 vss.n14399 vss.n1764 60091.4
R60 vss.n13954 vss.n8222 60091.4
R61 vss.n14071 vss.n8094 60091.4
R62 vss.n14398 vss.n1813 60091.4
R63 vss.n15093 vss.n1034 60091.4
R64 vss.n12237 vss.n9802 60091.4
R65 vss.n12355 vss.n9673 60091.4
R66 vss.n12474 vss.n9544 60091.4
R67 vss.n11733 vss.n8835 36300
R68 vss.n14177 vss.n14155 35204.9
R69 vss.n14911 vss.n404 31034.7
R70 vss.n14216 vss.n1183 31034.7
R71 vss.n3591 vss.n352 31034.7
R72 vss.n14177 vss.n14176 27452.2
R73 vss.n13250 vss.n13249 24224
R74 vss.n9818 vss.n9807 23948.6
R75 vss.n9689 vss.n9678 23948.6
R76 vss.n9560 vss.n9549 23948.6
R77 vss.n5603 vss.n5602 23948.6
R78 vss.n5879 vss.n5725 23948.6
R79 vss.n6118 vss.n5965 23948.6
R80 vss.n3523 vss.n3490 23948.6
R81 vss.n4073 vss.n4072 23948.6
R82 vss.n4254 vss.n4253 23948.6
R83 vss.n7406 vss.n7395 23948.6
R84 vss.n7236 vss.n7225 23948.6
R85 vss.n2714 vss.n2713 23948.6
R86 vss.n3047 vss.n3014 23948.6
R87 vss.n7059 vss.n7058 23948.6
R88 vss.n13871 vss.n13860 23948.6
R89 vss.n8110 vss.n8099 23948.6
R90 vss.n13547 vss.n13546 23948.6
R91 vss.n13848 vss.n8225 23948.6
R92 vss.n9032 vss.n9031 23948.6
R93 vss.n1780 vss.n1769 23948.6
R94 vss.n1001 vss.n990 23948.6
R95 vss.n11506 vss.n11505 23948.6
R96 vss.n11101 vss.n11100 23948.6
R97 vss.n10204 vss.n10203 23948.6
R98 vss.n6203 vss.n3989 23892
R99 vss.n7222 vss.n7221 23892
R100 vss.n14074 vss.n14073 23892
R101 vss.n10505 vss.n9543 23892
R102 vss.n12236 vss.n9805 22095.7
R103 vss.n12354 vss.n9676 22095.7
R104 vss.n12473 vss.n9547 22095.7
R105 vss.n12474 vss.n9546 22095.7
R106 vss.n12355 vss.n9675 22095.7
R107 vss.n12237 vss.n9804 22095.7
R108 vss.n6333 vss.n3487 22095.7
R109 vss.n5961 vss.n4003 22095.7
R110 vss.n6200 vss.n3995 22095.7
R111 vss.n5962 vss.n4002 22095.7
R112 vss.n6201 vss.n3994 22095.7
R113 vss.n3534 vss.n3533 22095.7
R114 vss.n7488 vss.n7394 22095.7
R115 vss.n7270 vss.n3128 22095.7
R116 vss.n7489 vss.n3057 22095.7
R117 vss.n7224 vss.n3131 22095.7
R118 vss.n15094 vss.n987 22095.7
R119 vss.n13953 vss.n13859 22095.7
R120 vss.n14070 vss.n8097 22095.7
R121 vss.n14071 vss.n8096 22095.7
R122 vss.n13954 vss.n13858 22095.7
R123 vss.n14399 vss.n1766 22095.7
R124 vss.n14398 vss.n1768 22095.7
R125 vss.n15093 vss.n989 22095.7
R126 vss.n14849 vss.n1158 21784
R127 vss.n15544 vss.n379 21784
R128 vss.n12239 vss.n12238 17233.3
R129 vss.n12357 vss.n12356 17233.3
R130 vss.n12476 vss.n12475 17233.3
R131 vss.n5723 vss.n5535 17233.3
R132 vss.n5963 vss.n3998 17233.3
R133 vss.n6202 vss.n3990 17233.3
R134 vss.n6369 vss.n6334 17233.3
R135 vss.n5724 vss.n5534 17233.3
R136 vss.n5964 vss.n3997 17233.3
R137 vss.n7393 vss.n3058 17233.3
R138 vss.n7223 vss.n3132 17233.3
R139 vss.n2674 vss.n988 17233.3
R140 vss.n2924 vss.n984 17233.3
R141 vss.n7985 vss.n2459 17233.3
R142 vss.n13956 vss.n13955 17233.3
R143 vss.n14072 vss.n2225 17233.3
R144 vss.n13591 vss.n1767 17233.3
R145 vss.n13780 vss.n1763 17233.3
R146 vss.n13068 vss.n8098 17233.3
R147 vss.n14447 vss.n14446 17233.3
R148 vss.n15142 vss.n15141 17233.3
R149 vss.n11549 vss.n9806 17233.3
R150 vss.n11238 vss.n9677 17233.3
R151 vss.n10899 vss.n9548 17233.3
R152 vss.n14789 vss.n14788 16848
R153 vss.n15484 vss.n15483 16848
R154 vss.n15657 vss.n351 16848
R155 vss.n12909 vss.n12908 15248
R156 vss.n12912 vss.n12911 15248
R157 vss.n12915 vss.n12914 15248
R158 vss.n13260 vss.n13259 15248
R159 vss.n13257 vss.n13256 15248
R160 vss.n13254 vss.n13253 15248
R161 vss.n13251 vss.n13250 15248
R162 vss.n14106 vss.n14105 15248
R163 vss.n14109 vss.n14108 15248
R164 vss.n14112 vss.n14111 15248
R165 vss.n14115 vss.n14114 15248
R166 vss.n14118 vss.n14117 15248
R167 vss.n14121 vss.n14120 15248
R168 vss.n14124 vss.n14123 15248
R169 vss.n14770 vss.n14769 15248
R170 vss.n14773 vss.n14772 15248
R171 vss.n14776 vss.n14775 15248
R172 vss.n14779 vss.n14778 15248
R173 vss.n14782 vss.n14781 15248
R174 vss.n14785 vss.n14784 15248
R175 vss.n14788 vss.n14787 15248
R176 vss.n7176 vss.n7175 15248
R177 vss.n7173 vss.n7172 15248
R178 vss.n7170 vss.n2470 15248
R179 vss.n7957 vss.n7956 15248
R180 vss.n7954 vss.n7953 15248
R181 vss.n7951 vss.n7950 15248
R182 vss.n7948 vss.n7947 15248
R183 vss.n15465 vss.n15464 15248
R184 vss.n15468 vss.n15467 15248
R185 vss.n15471 vss.n15470 15248
R186 vss.n15474 vss.n15473 15248
R187 vss.n15477 vss.n15476 15248
R188 vss.n15480 vss.n15479 15248
R189 vss.n15483 vss.n15482 15248
R190 vss.n6724 vss.n6723 15248
R191 vss.n6721 vss.n6720 15248
R192 vss.n6718 vss.n6717 15248
R193 vss.n6715 vss.n6714 15248
R194 vss.n6712 vss.n6711 15248
R195 vss.n6709 vss.n6708 15248
R196 vss.n6706 vss.n6705 15248
R197 vss.n6275 vss.n6274 15248
R198 vss.n6278 vss.n6277 15248
R199 vss.n6281 vss.n6280 15248
R200 vss.n6284 vss.n6283 15248
R201 vss.n6287 vss.n6286 15248
R202 vss.n6290 vss.n6289 15248
R203 vss.n6310 vss.n351 15248
R204 vss.n13202 vss.n13201 15248
R205 vss.n13205 vss.n13204 15248
R206 vss.n13208 vss.n13207 15248
R207 vss.n13211 vss.n13210 15248
R208 vss.n13214 vss.n13213 15248
R209 vss.n13217 vss.n13216 15248
R210 vss.n13220 vss.n13219 15248
R211 vss.n12907 vss.n12906 14872
R212 vss.n12910 vss.n12909 14872
R213 vss.n12913 vss.n12912 14872
R214 vss.n12915 vss.n8637 14872
R215 vss.n13259 vss.n13258 14872
R216 vss.n13256 vss.n13255 14872
R217 vss.n13253 vss.n13252 14872
R218 vss.n14108 vss.n14107 14872
R219 vss.n14111 vss.n14110 14872
R220 vss.n14114 vss.n14113 14872
R221 vss.n14117 vss.n14116 14872
R222 vss.n14120 vss.n14119 14872
R223 vss.n14123 vss.n14122 14872
R224 vss.n14768 vss.n14767 14872
R225 vss.n14771 vss.n14770 14872
R226 vss.n14774 vss.n14773 14872
R227 vss.n14777 vss.n14776 14872
R228 vss.n14780 vss.n14779 14872
R229 vss.n14783 vss.n14782 14872
R230 vss.n14786 vss.n14785 14872
R231 vss.n7174 vss.n7173 14872
R232 vss.n7171 vss.n7170 14872
R233 vss.n7958 vss.n7957 14872
R234 vss.n7955 vss.n7954 14872
R235 vss.n7952 vss.n7951 14872
R236 vss.n7949 vss.n7948 14872
R237 vss.n7946 vss.n1158 14872
R238 vss.n15463 vss.n15462 14872
R239 vss.n15466 vss.n15465 14872
R240 vss.n15469 vss.n15468 14872
R241 vss.n15472 vss.n15471 14872
R242 vss.n15475 vss.n15474 14872
R243 vss.n15478 vss.n15477 14872
R244 vss.n15481 vss.n15480 14872
R245 vss.n6722 vss.n6721 14872
R246 vss.n6719 vss.n6718 14872
R247 vss.n6716 vss.n6715 14872
R248 vss.n6713 vss.n6712 14872
R249 vss.n6710 vss.n6709 14872
R250 vss.n6707 vss.n6706 14872
R251 vss.n6704 vss.n379 14872
R252 vss.n6273 vss.n6272 14872
R253 vss.n6276 vss.n6275 14872
R254 vss.n6279 vss.n6278 14872
R255 vss.n6282 vss.n6281 14872
R256 vss.n6285 vss.n6284 14872
R257 vss.n6288 vss.n6287 14872
R258 vss.n6311 vss.n6290 14872
R259 vss.n13204 vss.n13203 14872
R260 vss.n13207 vss.n13206 14872
R261 vss.n13210 vss.n13209 14872
R262 vss.n13213 vss.n13212 14872
R263 vss.n13216 vss.n13215 14872
R264 vss.n13219 vss.n13218 14872
R265 vss.n13258 vss.n8687 14460.6
R266 vss.n12913 vss.n9207 14460.6
R267 vss.n12907 vss.n9280 14460.6
R268 vss.n13252 vss.n8806 14460.6
R269 vss.n6285 vss.n3730 14460.6
R270 vss.n6279 vss.n3849 14460.6
R271 vss.n6273 vss.n3968 14460.6
R272 vss.n6704 vss.n3334 14460.6
R273 vss.n6710 vss.n3326 14460.6
R274 vss.n6716 vss.n3318 14460.6
R275 vss.n6722 vss.n3310 14460.6
R276 vss.n15481 vss.n409 14460.6
R277 vss.n15475 vss.n417 14460.6
R278 vss.n15469 vss.n425 14460.6
R279 vss.n15463 vss.n433 14460.6
R280 vss.n7946 vss.n7925 14460.6
R281 vss.n7952 vss.n2477 14460.6
R282 vss.n7959 vss.n7958 14460.6
R283 vss.n7174 vss.n6824 14460.6
R284 vss.n14786 vss.n1188 14460.6
R285 vss.n14780 vss.n1196 14460.6
R286 vss.n14774 vss.n1204 14460.6
R287 vss.n14768 vss.n1212 14460.6
R288 vss.n13574 vss.n2053 14460.6
R289 vss.n14119 vss.n2107 14460.6
R290 vss.n14113 vss.n2115 14460.6
R291 vss.n14107 vss.n2123 14460.6
R292 vss.n6311 vss.n3611 14460.6
R293 vss.n13221 vss.n8837 14460.6
R294 vss.n13215 vss.n8845 14460.6
R295 vss.n13209 vss.n8853 14460.6
R296 vss.n13203 vss.n8861 14460.6
R297 vss.n13255 vss.n8737 14161.2
R298 vss.n9702 vss.n8637 14161.2
R299 vss.n12910 vss.n9276 14161.2
R300 vss.n6288 vss.n3662 14161.2
R301 vss.n6282 vss.n3781 14161.2
R302 vss.n6276 vss.n3900 14161.2
R303 vss.n6707 vss.n3330 14161.2
R304 vss.n6713 vss.n3322 14161.2
R305 vss.n6719 vss.n3314 14161.2
R306 vss.n15472 vss.n421 14161.2
R307 vss.n15466 vss.n429 14161.2
R308 vss.n7949 vss.n2481 14161.2
R309 vss.n7955 vss.n2473 14161.2
R310 vss.n7171 vss.n7076 14161.2
R311 vss.n14777 vss.n1200 14161.2
R312 vss.n14771 vss.n1208 14161.2
R313 vss.n14122 vss.n2103 14161.2
R314 vss.n14116 vss.n2111 14161.2
R315 vss.n14110 vss.n2119 14161.2
R316 vss.n14783 vss.n1192 14161.2
R317 vss.n15478 vss.n413 14161.2
R318 vss.n13218 vss.n8841 14161.2
R319 vss.n13212 vss.n8849 14161.2
R320 vss.n13206 vss.n8857 14161.2
R321 vss.n6271 vss.n6270 13907.7
R322 vss.n12238 vss.n9801 13814.6
R323 vss.n12356 vss.n9672 13814.6
R324 vss.n12475 vss.n9542 13814.6
R325 vss.n5723 vss.n5722 13814.6
R326 vss.n5963 vss.n3999 13814.6
R327 vss.n6202 vss.n3991 13814.6
R328 vss.n6334 vss.n3486 13814.6
R329 vss.n5724 vss.n4004 13814.6
R330 vss.n5964 vss.n3996 13814.6
R331 vss.n7393 vss.n7392 13814.6
R332 vss.n7223 vss.n3133 13814.6
R333 vss.n7901 vss.n988 13814.6
R334 vss.n7706 vss.n984 13814.6
R335 vss.n7102 vss.n2459 13814.6
R336 vss.n13955 vss.n8221 13814.6
R337 vss.n14072 vss.n8093 13814.6
R338 vss.n13641 vss.n1767 13814.6
R339 vss.n13830 vss.n1763 13814.6
R340 vss.n13118 vss.n8098 13814.6
R341 vss.n14448 vss.n14447 13814.6
R342 vss.n15143 vss.n15142 13814.6
R343 vss.n11599 vss.n9806 13814.6
R344 vss.n11288 vss.n9677 13814.6
R345 vss.n10853 vss.n9548 13814.6
R346 vss.n14178 vss.n2053 13800
R347 vss.n13222 vss.n13221 13800
R348 vss.n6203 vss.n3988 13770.6
R349 vss.n7222 vss.n3134 13770.6
R350 vss.n14073 vss.n2224 13770.6
R351 vss.n10457 vss.n9543 13770.6
R352 vss.n15484 vss.n404 13684
R353 vss.n14789 vss.n1183 13684
R354 vss.n15657 vss.n352 13684
R355 vss.n11793 vss.n8810 13013
R356 vss.n14105 vss.n14104 12952
R357 vss.n7177 vss.n7176 12952
R358 vss.n6725 vss.n6724 12952
R359 vss.n13201 vss.n13200 12952
R360 vss.n12905 vss.n12904 11309.3
R361 vss.n15461 vss.n15460 11309.3
R362 vss.n14766 vss.n14765 11309.3
R363 vss.n12906 vss.n12905 10512
R364 vss.n14767 vss.n14766 10512
R365 vss.n15462 vss.n15461 10512
R366 vss.n6272 vss.n6271 10512
R367 vss.n14870 vss.n14869 10314.6
R368 vss.n15546 vss.n15545 10314.6
R369 vss.n1767 vss.n1183 10235.7
R370 vss.n988 vss.n404 10235.7
R371 vss.n6334 vss.n352 10235.7
R372 vss.n13255 vss.n8736 10178.7
R373 vss.n13258 vss.n8686 10178.7
R374 vss.n9650 vss.n8637 10178.7
R375 vss.n12913 vss.n9206 10178.7
R376 vss.n12910 vss.n9275 10178.7
R377 vss.n12907 vss.n9279 10178.7
R378 vss.n13252 vss.n8805 10178.7
R379 vss.n6288 vss.n3661 10178.7
R380 vss.n6285 vss.n3729 10178.7
R381 vss.n6282 vss.n3780 10178.7
R382 vss.n6279 vss.n3848 10178.7
R383 vss.n6276 vss.n3899 10178.7
R384 vss.n6273 vss.n3967 10178.7
R385 vss.n6704 vss.n6703 10178.7
R386 vss.n6707 vss.n3331 10178.7
R387 vss.n6710 vss.n3327 10178.7
R388 vss.n6713 vss.n3323 10178.7
R389 vss.n6716 vss.n3319 10178.7
R390 vss.n6719 vss.n3315 10178.7
R391 vss.n6722 vss.n3311 10178.7
R392 vss.n15481 vss.n408 10178.7
R393 vss.n15475 vss.n416 10178.7
R394 vss.n15472 vss.n420 10178.7
R395 vss.n15469 vss.n424 10178.7
R396 vss.n15466 vss.n428 10178.7
R397 vss.n15463 vss.n432 10178.7
R398 vss.n7946 vss.n7945 10178.7
R399 vss.n7949 vss.n2482 10178.7
R400 vss.n7952 vss.n2478 10178.7
R401 vss.n7955 vss.n2474 10178.7
R402 vss.n7958 vss.n2469 10178.7
R403 vss.n7171 vss.n7123 10178.7
R404 vss.n7174 vss.n6919 10178.7
R405 vss.n14786 vss.n1187 10178.7
R406 vss.n14780 vss.n1195 10178.7
R407 vss.n14777 vss.n1199 10178.7
R408 vss.n14774 vss.n1203 10178.7
R409 vss.n14771 vss.n1207 10178.7
R410 vss.n14768 vss.n1211 10178.7
R411 vss.n2074 vss.n2053 10178.7
R412 vss.n14122 vss.n2104 10178.7
R413 vss.n14119 vss.n2108 10178.7
R414 vss.n14116 vss.n2112 10178.7
R415 vss.n14113 vss.n2116 10178.7
R416 vss.n14110 vss.n2120 10178.7
R417 vss.n14107 vss.n2124 10178.7
R418 vss.n14783 vss.n1191 10178.7
R419 vss.n15478 vss.n412 10178.7
R420 vss.n6312 vss.n6311 10178.7
R421 vss.n13221 vss.n8838 10178.7
R422 vss.n13218 vss.n8842 10178.7
R423 vss.n13215 vss.n8846 10178.7
R424 vss.n13212 vss.n8850 10178.7
R425 vss.n13209 vss.n8854 10178.7
R426 vss.n13206 vss.n8858 10178.7
R427 vss.n13203 vss.n8862 10178.7
R428 vss.n14175 vss.n2052 9771.87
R429 vss.n12475 vss.n9543 9131.13
R430 vss.n14073 vss.n14072 9131.13
R431 vss.n7223 vss.n7222 9131.13
R432 vss.n6203 vss.n6202 9131.13
R433 vss.n8835 vss.n8810 8418.67
R434 vss.n12356 vss.n9548 8101.44
R435 vss.n12238 vss.n9677 8101.44
R436 vss.n13955 vss.n8098 8101.44
R437 vss.n14447 vss.n1763 8101.44
R438 vss.n7393 vss.n2459 8101.44
R439 vss.n15142 vss.n984 8101.44
R440 vss.n5964 vss.n5963 8101.44
R441 vss.n5724 vss.n5723 8101.44
R442 vss.n13249 vss.n13248 7771.93
R443 vss.n14869 vss.n14868 7343.64
R444 vss.n15547 vss.n15546 7343.64
R445 vss.n12474 vss.n12473 6926.6
R446 vss.n12355 vss.n12354 6926.6
R447 vss.n12237 vss.n12236 6926.6
R448 vss.n14071 vss.n14070 6926.6
R449 vss.n13954 vss.n13953 6926.6
R450 vss.n14399 vss.n14398 6926.6
R451 vss.n7270 vss.n7224 6926.6
R452 vss.n7489 vss.n7488 6926.6
R453 vss.n15094 vss.n15093 6926.6
R454 vss.n6201 vss.n6200 6926.6
R455 vss.n5962 vss.n5961 6926.6
R456 vss.n6333 vss.n3534 6926.6
R457 vss.n15660 vss.n15659 6569.89
R458 vss.n13224 vss.n8834 5870.11
R459 vss.n12181 vss.n8809 5824.14
R460 vss.n15542 vss.n381 5824.14
R461 vss.n14847 vss.n1160 5824.14
R462 vss.n14175 vss.n14174 5175.08
R463 vss.n14849 vss.n14848 5066.66
R464 vss.n15544 vss.n15543 5066.66
R465 vss.n15658 vss.n303 4992.92
R466 vss.n14791 vss.n14790 4992.92
R467 vss.n15486 vss.n15485 4992.92
R468 vss.n11730 vss.n9806 4774.23
R469 vss.n11677 vss.n9932 4548.38
R470 vss.n11677 vss.n9931 4548.38
R471 vss.n11659 vss.n11658 4548.38
R472 vss.n11659 vss.n11655 4548.38
R473 vss.n11440 vss.n11351 4548.38
R474 vss.n11440 vss.n11350 4548.38
R475 vss.n11422 vss.n11421 4548.38
R476 vss.n11422 vss.n11418 4548.38
R477 vss.n11328 vss.n10054 4548.38
R478 vss.n11326 vss.n10054 4548.38
R479 vss.n11347 vss.n9985 4548.38
R480 vss.n11347 vss.n9986 4548.38
R481 vss.n11035 vss.n11031 4548.38
R482 vss.n11035 vss.n11030 4548.38
R483 vss.n11321 vss.n10057 4548.38
R484 vss.n11321 vss.n10058 4548.38
R485 vss.n10761 vss.n10757 4548.38
R486 vss.n10761 vss.n10756 4548.38
R487 vss.n11027 vss.n10145 4548.38
R488 vss.n11027 vss.n10146 4548.38
R489 vss.n10783 vss.n10638 4548.38
R490 vss.n10783 vss.n10637 4548.38
R491 vss.n10765 vss.n10708 4548.38
R492 vss.n10765 vss.n10706 4548.38
R493 vss.n10393 vss.n10389 4548.38
R494 vss.n10393 vss.n10388 4548.38
R495 vss.n10634 vss.n10232 4548.38
R496 vss.n10634 vss.n10233 4548.38
R497 vss.n12094 vss.n12093 4548.38
R498 vss.n12093 vss.n11884 4548.38
R499 vss.n12130 vss.n11841 4548.38
R500 vss.n12130 vss.n11842 4548.38
R501 vss.n8395 vss.n8388 4548.38
R502 vss.n8396 vss.n8395 4548.38
R503 vss.n12072 vss.n12009 4548.38
R504 vss.n12072 vss.n12010 4548.38
R505 vss.n13398 vss.n13397 4548.38
R506 vss.n13397 vss.n13393 4548.38
R507 vss.n13426 vss.n13423 4548.38
R508 vss.n13428 vss.n13423 4548.38
R509 vss.n8592 vss.n8591 4548.38
R510 vss.n8591 vss.n8584 4548.38
R511 vss.n8572 vss.n8569 4548.38
R512 vss.n8572 vss.n8567 4548.38
R513 vss.n12964 vss.n12960 4548.38
R514 vss.n12967 vss.n12964 4548.38
R515 vss.n13307 vss.n8437 4548.38
R516 vss.n13309 vss.n8437 4548.38
R517 vss.n8939 vss.n8932 4548.38
R518 vss.n8940 vss.n8939 4548.38
R519 vss.n9170 vss.n9107 4548.38
R520 vss.n9170 vss.n9108 4548.38
R521 vss.n12702 vss.n12701 4548.38
R522 vss.n12811 vss.n12702 4548.38
R523 vss.n12783 vss.n12779 4548.38
R524 vss.n12781 vss.n12779 4548.38
R525 vss.n9366 vss.n9365 4548.38
R526 vss.n12888 vss.n9366 4548.38
R527 vss.n12830 vss.n9415 4548.38
R528 vss.n12832 vss.n9415 4548.38
R529 vss.n12875 vss.n9382 4548.38
R530 vss.n12877 vss.n9382 4548.38
R531 vss.n12902 vss.n9303 4548.38
R532 vss.n12902 vss.n9304 4548.38
R533 vss.n12798 vss.n12718 4548.38
R534 vss.n12800 vss.n12718 4548.38
R535 vss.n12825 vss.n12640 4548.38
R536 vss.n12825 vss.n12641 4548.38
R537 vss.n13140 vss.n8923 4548.38
R538 vss.n13142 vss.n8923 4548.38
R539 vss.n13160 vss.n8902 4548.38
R540 vss.n13160 vss.n8903 4548.38
R541 vss.n12981 vss.n12953 4548.38
R542 vss.n12983 vss.n12953 4548.38
R543 vss.n13001 vss.n9174 4548.38
R544 vss.n13001 vss.n9175 4548.38
R545 vss.n8607 vss.n8509 4548.38
R546 vss.n8609 vss.n8509 4548.38
R547 vss.n13302 vss.n8488 4548.38
R548 vss.n13302 vss.n8489 4548.38
R549 vss.n13414 vss.n13380 4548.38
R550 vss.n13380 vss.n13378 4548.38
R551 vss.n13713 vss.n8322 4548.38
R552 vss.n13713 vss.n8323 4548.38
R553 vss.n13663 vss.n8379 4548.38
R554 vss.n13665 vss.n8379 4548.38
R555 vss.n13683 vss.n8358 4548.38
R556 vss.n13683 vss.n8359 4548.38
R557 vss.n15662 vss.n301 4548.38
R558 vss.n15664 vss.n301 4548.38
R559 vss.n15685 vss.n281 4548.38
R560 vss.n15685 vss.n282 4548.38
R561 vss.n278 vss.n260 4548.38
R562 vss.n278 vss.n261 4548.38
R563 vss.n15714 vss.n226 4548.38
R564 vss.n15714 vss.n227 4548.38
R565 vss.n15719 vss.n223 4548.38
R566 vss.n15721 vss.n223 4548.38
R567 vss.n15741 vss.n202 4548.38
R568 vss.n15741 vss.n203 4548.38
R569 vss.n199 vss.n181 4548.38
R570 vss.n199 vss.n182 4548.38
R571 vss.n15770 vss.n148 4548.38
R572 vss.n15770 vss.n149 4548.38
R573 vss.n15775 vss.n145 4548.38
R574 vss.n15777 vss.n145 4548.38
R575 vss.n15797 vss.n124 4548.38
R576 vss.n15797 vss.n125 4548.38
R577 vss.n121 vss.n103 4548.38
R578 vss.n121 vss.n104 4548.38
R579 vss.n15826 vss.n69 4548.38
R580 vss.n15826 vss.n70 4548.38
R581 vss.n15831 vss.n66 4548.38
R582 vss.n15833 vss.n66 4548.38
R583 vss.n15853 vss.n45 4548.38
R584 vss.n15853 vss.n46 4548.38
R585 vss.n15879 vss.n26 4548.38
R586 vss.n26 vss.n22 4548.38
R587 vss.n6269 vss.n6254 4548.38
R588 vss.n6269 vss.n6255 4548.38
R589 vss.n4844 vss.n4807 4548.38
R590 vss.n4844 vss.n4808 4548.38
R591 vss.n15458 vss.n438 4548.38
R592 vss.n15458 vss.n439 4548.38
R593 vss.n4897 vss.n4293 4548.38
R594 vss.n4293 vss.n4291 4548.38
R595 vss.n4867 vss.n4365 4548.38
R596 vss.n4865 vss.n4365 4548.38
R597 vss.n15398 vss.n15394 4548.38
R598 vss.n15398 vss.n15395 4548.38
R599 vss.n15426 vss.n539 4548.38
R600 vss.n15426 vss.n540 4548.38
R601 vss.n5160 vss.n5126 4548.38
R602 vss.n5126 vss.n5124 4548.38
R603 vss.n15383 vss.n645 4548.38
R604 vss.n15383 vss.n646 4548.38
R605 vss.n5372 vss.n5338 4548.38
R606 vss.n5338 vss.n5336 4548.38
R607 vss.n15353 vss.n744 4548.38
R608 vss.n15353 vss.n745 4548.38
R609 vss.n15248 vss.n15244 4548.38
R610 vss.n15248 vss.n15245 4548.38
R611 vss.n15276 vss.n797 4548.38
R612 vss.n15276 vss.n798 4548.38
R613 vss.n6444 vss.n6410 4548.38
R614 vss.n6410 vss.n6408 4548.38
R615 vss.n15233 vss.n902 4548.38
R616 vss.n15233 vss.n903 4548.38
R617 vss.n6559 vss.n6525 4548.38
R618 vss.n6525 vss.n6523 4548.38
R619 vss.n15032 vss.n1077 4548.38
R620 vss.n15032 vss.n1078 4548.38
R621 vss.n6544 vss.n6537 4548.38
R622 vss.n6542 vss.n6537 4548.38
R623 vss.n6572 vss.n6568 4548.38
R624 vss.n6574 vss.n6568 4548.38
R625 vss.n6429 vss.n6422 4548.38
R626 vss.n6427 vss.n6422 4548.38
R627 vss.n6456 vss.n6453 4548.38
R628 vss.n6458 vss.n6453 4548.38
R629 vss.n877 vss.n876 4548.38
R630 vss.n876 vss.n870 4548.38
R631 vss.n15239 vss.n889 4548.38
R632 vss.n898 vss.n889 4548.38
R633 vss.n5357 vss.n5350 4548.38
R634 vss.n5355 vss.n5350 4548.38
R635 vss.n5384 vss.n5381 4548.38
R636 vss.n5386 vss.n5381 4548.38
R637 vss.n5145 vss.n5138 4548.38
R638 vss.n5143 vss.n5138 4548.38
R639 vss.n5172 vss.n5169 4548.38
R640 vss.n5174 vss.n5169 4548.38
R641 vss.n620 vss.n619 4548.38
R642 vss.n619 vss.n613 4548.38
R643 vss.n15389 vss.n632 4548.38
R644 vss.n641 vss.n632 4548.38
R645 vss.n4882 vss.n4303 4548.38
R646 vss.n4880 vss.n4303 4548.38
R647 vss.n4909 vss.n4906 4548.38
R648 vss.n4911 vss.n4906 4548.38
R649 vss.n4829 vss.n4821 4548.38
R650 vss.n4821 vss.n4816 4548.38
R651 vss.n4859 vss.n4746 4548.38
R652 vss.n4859 vss.n4747 4548.38
R653 vss.n3266 vss.n3229 4548.38
R654 vss.n3266 vss.n3230 4548.38
R655 vss.n14763 vss.n1217 4548.38
R656 vss.n14763 vss.n1218 4548.38
R657 vss.n8003 vss.n2439 4548.38
R658 vss.n8005 vss.n2439 4548.38
R659 vss.n8030 vss.n2361 4548.38
R660 vss.n8030 vss.n2362 4548.38
R661 vss.n14703 vss.n14699 4548.38
R662 vss.n14703 vss.n14700 4548.38
R663 vss.n14731 vss.n1318 4548.38
R664 vss.n14731 vss.n1319 4548.38
R665 vss.n7568 vss.n7534 4548.38
R666 vss.n7534 vss.n7532 4548.38
R667 vss.n14688 vss.n1424 4548.38
R668 vss.n14688 vss.n1425 4548.38
R669 vss.n2786 vss.n2752 4548.38
R670 vss.n2752 vss.n2750 4548.38
R671 vss.n14658 vss.n1523 4548.38
R672 vss.n14658 vss.n1524 4548.38
R673 vss.n14553 vss.n14549 4548.38
R674 vss.n14553 vss.n14550 4548.38
R675 vss.n14581 vss.n1576 4548.38
R676 vss.n14581 vss.n1577 4548.38
R677 vss.n2552 vss.n2518 4548.38
R678 vss.n2518 vss.n2516 4548.38
R679 vss.n14538 vss.n1681 4548.38
R680 vss.n14538 vss.n1682 4548.38
R681 vss.n1969 vss.n1965 4548.38
R682 vss.n1969 vss.n1966 4548.38
R683 vss.n14337 vss.n1856 4548.38
R684 vss.n14337 vss.n1857 4548.38
R685 vss.n1890 vss.n1887 4548.38
R686 vss.n1887 vss.n1883 4548.38
R687 vss.n1960 vss.n1948 4548.38
R688 vss.n1957 vss.n1948 4548.38
R689 vss.n2539 vss.n2532 4548.38
R690 vss.n2537 vss.n2532 4548.38
R691 vss.n2563 vss.n2560 4548.38
R692 vss.n2565 vss.n2560 4548.38
R693 vss.n1656 vss.n1655 4548.38
R694 vss.n1655 vss.n1649 4548.38
R695 vss.n14544 vss.n1668 4548.38
R696 vss.n1677 vss.n1668 4548.38
R697 vss.n2771 vss.n2764 4548.38
R698 vss.n2769 vss.n2764 4548.38
R699 vss.n2798 vss.n2795 4548.38
R700 vss.n2800 vss.n2795 4548.38
R701 vss.n7553 vss.n7546 4548.38
R702 vss.n7551 vss.n7546 4548.38
R703 vss.n7580 vss.n7577 4548.38
R704 vss.n7582 vss.n7577 4548.38
R705 vss.n1399 vss.n1398 4548.38
R706 vss.n1398 vss.n1392 4548.38
R707 vss.n14694 vss.n1411 4548.38
R708 vss.n1420 vss.n1411 4548.38
R709 vss.n2423 vss.n2422 4548.38
R710 vss.n8016 vss.n2423 4548.38
R711 vss.n6951 vss.n6948 4548.38
R712 vss.n6953 vss.n6948 4548.38
R713 vss.n3252 vss.n3241 4548.38
R714 vss.n3250 vss.n3241 4548.38
R715 vss.n3218 vss.n3215 4548.38
R716 vss.n3220 vss.n3215 4548.38
R717 vss.n12115 vss.n11873 4548.38
R718 vss.n12115 vss.n11874 4548.38
R719 vss.n12080 vss.n11943 4548.38
R720 vss.n12078 vss.n11943 4548.38
R721 vss.n10385 vss.n10274 4548.38
R722 vss.n10385 vss.n10275 4548.38
R723 vss.n10366 vss.n10342 4548.38
R724 vss.n10364 vss.n10342 4548.38
R725 vss.n14178 vss.n2052 4308.9
R726 vss.n15659 vss.n302 4280
R727 vss.n14176 vss.n14175 4223.46
R728 vss.n11797 vss.n8810 4164.16
R729 vss.n13200 vss.n13199 4137.66
R730 vss.n6726 vss.n6725 4137.66
R731 vss.n7177 vss.n3168 4137.66
R732 vss.n14104 vss.n14103 4137.66
R733 vss.n13249 vss.n8809 4000
R734 vss.n9941 vss.n9940 3789.35
R735 vss.n9940 vss.n9936 3789.35
R736 vss.n9944 vss.n9942 3789.35
R737 vss.n9944 vss.n9937 3789.35
R738 vss.n11653 vss.n9947 3789.35
R739 vss.n11653 vss.n11651 3789.35
R740 vss.n11359 vss.n11358 3789.35
R741 vss.n11358 vss.n11354 3789.35
R742 vss.n11362 vss.n11360 3789.35
R743 vss.n11362 vss.n11355 3789.35
R744 vss.n11416 vss.n11365 3789.35
R745 vss.n11416 vss.n11414 3789.35
R746 vss.n10051 vss.n10046 3789.35
R747 vss.n10051 vss.n10050 3789.35
R748 vss.n10048 vss.n10041 3789.35
R749 vss.n10048 vss.n9990 3789.35
R750 vss.n10043 vss.n10042 3789.35
R751 vss.n10042 vss.n9991 3789.35
R752 vss.n10076 vss.n10071 3789.35
R753 vss.n10076 vss.n10075 3789.35
R754 vss.n10073 vss.n10066 3789.35
R755 vss.n10073 vss.n10062 3789.35
R756 vss.n10068 vss.n10067 3789.35
R757 vss.n10067 vss.n10063 3789.35
R758 vss.n10164 vss.n10159 3789.35
R759 vss.n10164 vss.n10163 3789.35
R760 vss.n10161 vss.n10154 3789.35
R761 vss.n10161 vss.n10150 3789.35
R762 vss.n10156 vss.n10155 3789.35
R763 vss.n10155 vss.n10151 3789.35
R764 vss.n10647 vss.n10646 3789.35
R765 vss.n10646 vss.n10642 3789.35
R766 vss.n10650 vss.n10648 3789.35
R767 vss.n10650 vss.n10643 3789.35
R768 vss.n10704 vss.n10653 3789.35
R769 vss.n10704 vss.n10702 3789.35
R770 vss.n10251 vss.n10246 3789.35
R771 vss.n10251 vss.n10250 3789.35
R772 vss.n10248 vss.n10241 3789.35
R773 vss.n10248 vss.n10237 3789.35
R774 vss.n10243 vss.n10242 3789.35
R775 vss.n10242 vss.n10238 3789.35
R776 vss.n12100 vss.n12099 3789.35
R777 vss.n12099 vss.n11885 3789.35
R778 vss.n12118 vss.n11868 3789.35
R779 vss.n12118 vss.n11845 3789.35
R780 vss.n11870 vss.n11869 3789.35
R781 vss.n11869 vss.n11846 3789.35
R782 vss.n8402 vss.n8389 3789.35
R783 vss.n8403 vss.n8402 3789.35
R784 vss.n13660 vss.n8384 3789.35
R785 vss.n13660 vss.n8385 3789.35
R786 vss.n12067 vss.n12013 3789.35
R787 vss.n12067 vss.n12014 3789.35
R788 vss.n13404 vss.n13388 3789.35
R789 vss.n13404 vss.n13389 3789.35
R790 vss.n13417 vss.n13373 3789.35
R791 vss.n13417 vss.n13376 3789.35
R792 vss.n13430 vss.n13374 3789.35
R793 vss.n13430 vss.n13429 3789.35
R794 vss.n8599 vss.n8598 3789.35
R795 vss.n8598 vss.n8585 3789.35
R796 vss.n8604 vss.n8514 3789.35
R797 vss.n8604 vss.n8515 3789.35
R798 vss.n8575 vss.n8517 3789.35
R799 vss.n8575 vss.n8566 3789.35
R800 vss.n12971 vss.n12970 3789.35
R801 vss.n12971 vss.n12957 3789.35
R802 vss.n12978 vss.n8431 3789.35
R803 vss.n12978 vss.n12976 3789.35
R804 vss.n13311 vss.n8432 3789.35
R805 vss.n13311 vss.n13310 3789.35
R806 vss.n8946 vss.n8933 3789.35
R807 vss.n8947 vss.n8946 3789.35
R808 vss.n13137 vss.n8928 3789.35
R809 vss.n13137 vss.n8929 3789.35
R810 vss.n9165 vss.n9111 3789.35
R811 vss.n9165 vss.n9112 3789.35
R812 vss.n12807 vss.n12703 3789.35
R813 vss.n12807 vss.n12708 3789.35
R814 vss.n12795 vss.n12721 3789.35
R815 vss.n12795 vss.n12722 3789.35
R816 vss.n12785 vss.n12777 3789.35
R817 vss.n12785 vss.n12727 3789.35
R818 vss.n12884 vss.n9367 3789.35
R819 vss.n12884 vss.n9372 3789.35
R820 vss.n12872 vss.n9385 3789.35
R821 vss.n12872 vss.n9386 3789.35
R822 vss.n12834 vss.n9412 3789.35
R823 vss.n12834 vss.n12833 3789.35
R824 vss.n12881 vss.n9374 3789.35
R825 vss.n12881 vss.n9375 3789.35
R826 vss.n12891 vss.n9361 3789.35
R827 vss.n12891 vss.n9309 3789.35
R828 vss.n9360 vss.n9359 3789.35
R829 vss.n9359 vss.n9308 3789.35
R830 vss.n12804 vss.n12710 3789.35
R831 vss.n12804 vss.n12711 3789.35
R832 vss.n12814 vss.n12697 3789.35
R833 vss.n12814 vss.n12646 3789.35
R834 vss.n12696 vss.n12695 3789.35
R835 vss.n12695 vss.n12645 3789.35
R836 vss.n8924 vss.n8917 3789.35
R837 vss.n8924 vss.n8920 3789.35
R838 vss.n8936 vss.n8913 3789.35
R839 vss.n8936 vss.n8908 3789.35
R840 vss.n8912 vss.n8911 3789.35
R841 vss.n8911 vss.n8907 3789.35
R842 vss.n12954 vss.n12947 3789.35
R843 vss.n12954 vss.n12950 3789.35
R844 vss.n12961 vss.n12943 3789.35
R845 vss.n12961 vss.n9180 3789.35
R846 vss.n12942 vss.n12941 3789.35
R847 vss.n12941 vss.n9179 3789.35
R848 vss.n8510 vss.n8503 3789.35
R849 vss.n8510 vss.n8506 3789.35
R850 vss.n8588 vss.n8499 3789.35
R851 vss.n8588 vss.n8494 3789.35
R852 vss.n8498 vss.n8497 3789.35
R853 vss.n8497 vss.n8493 3789.35
R854 vss.n13385 vss.n13379 3789.35
R855 vss.n13385 vss.n13383 3789.35
R856 vss.n13394 vss.n8333 3789.35
R857 vss.n13394 vss.n8328 3789.35
R858 vss.n8332 vss.n8331 3789.35
R859 vss.n8331 vss.n8327 3789.35
R860 vss.n8380 vss.n8373 3789.35
R861 vss.n8380 vss.n8376 3789.35
R862 vss.n8392 vss.n8369 3789.35
R863 vss.n8392 vss.n8364 3789.35
R864 vss.n8368 vss.n8367 3789.35
R865 vss.n8367 vss.n8363 3789.35
R866 vss.n15666 vss.n293 3789.35
R867 vss.n15666 vss.n298 3789.35
R868 vss.n296 vss.n290 3789.35
R869 vss.n297 vss.n296 3789.35
R870 vss.n15680 vss.n286 3789.35
R871 vss.n15680 vss.n287 3789.35
R872 vss.n273 vss.n265 3789.35
R873 vss.n273 vss.n266 3789.35
R874 vss.n267 vss.n237 3789.35
R875 vss.n267 vss.n232 3789.35
R876 vss.n236 vss.n235 3789.35
R877 vss.n235 vss.n231 3789.35
R878 vss.n15723 vss.n217 3789.35
R879 vss.n15723 vss.n221 3789.35
R880 vss.n218 vss.n213 3789.35
R881 vss.n218 vss.n208 3789.35
R882 vss.n212 vss.n211 3789.35
R883 vss.n211 vss.n207 3789.35
R884 vss.n194 vss.n186 3789.35
R885 vss.n194 vss.n187 3789.35
R886 vss.n188 vss.n159 3789.35
R887 vss.n188 vss.n154 3789.35
R888 vss.n158 vss.n157 3789.35
R889 vss.n157 vss.n153 3789.35
R890 vss.n15779 vss.n139 3789.35
R891 vss.n15779 vss.n143 3789.35
R892 vss.n140 vss.n135 3789.35
R893 vss.n140 vss.n130 3789.35
R894 vss.n134 vss.n133 3789.35
R895 vss.n133 vss.n129 3789.35
R896 vss.n116 vss.n108 3789.35
R897 vss.n116 vss.n109 3789.35
R898 vss.n110 vss.n80 3789.35
R899 vss.n110 vss.n75 3789.35
R900 vss.n79 vss.n78 3789.35
R901 vss.n78 vss.n74 3789.35
R902 vss.n15835 vss.n60 3789.35
R903 vss.n15835 vss.n64 3789.35
R904 vss.n61 vss.n56 3789.35
R905 vss.n61 vss.n51 3789.35
R906 vss.n55 vss.n54 3789.35
R907 vss.n54 vss.n50 3789.35
R908 vss.n15882 vss.n23 3789.35
R909 vss.n15883 vss.n15882 3789.35
R910 vss.n15888 vss.n17 3789.35
R911 vss.n15888 vss.n18 3789.35
R912 vss.n6264 vss.n6260 3789.35
R913 vss.n6264 vss.n6262 3789.35
R914 vss.n4839 vss.n4812 3789.35
R915 vss.n4839 vss.n4813 3789.35
R916 vss.n4823 vss.n449 3789.35
R917 vss.n4823 vss.n444 3789.35
R918 vss.n448 vss.n447 3789.35
R919 vss.n447 vss.n443 3789.35
R920 vss.n4891 vss.n4292 3789.35
R921 vss.n4891 vss.n4296 3789.35
R922 vss.n4877 vss.n4307 3789.35
R923 vss.n4877 vss.n4309 3789.35
R924 vss.n4362 vss.n4361 3789.35
R925 vss.n4362 vss.n4312 3789.35
R926 vss.n15408 vss.n601 3789.35
R927 vss.n15408 vss.n604 3789.35
R928 vss.n616 vss.n597 3789.35
R929 vss.n616 vss.n545 3789.35
R930 vss.n596 vss.n595 3789.35
R931 vss.n595 vss.n544 3789.35
R932 vss.n5154 vss.n5125 3789.35
R933 vss.n5154 vss.n5129 3789.35
R934 vss.n5140 vss.n656 3789.35
R935 vss.n5140 vss.n651 3789.35
R936 vss.n655 vss.n654 3789.35
R937 vss.n654 vss.n650 3789.35
R938 vss.n5366 vss.n5337 3789.35
R939 vss.n5366 vss.n5341 3789.35
R940 vss.n5352 vss.n755 3789.35
R941 vss.n5352 vss.n750 3789.35
R942 vss.n754 vss.n753 3789.35
R943 vss.n753 vss.n749 3789.35
R944 vss.n15258 vss.n858 3789.35
R945 vss.n15258 vss.n861 3789.35
R946 vss.n873 vss.n854 3789.35
R947 vss.n873 vss.n803 3789.35
R948 vss.n853 vss.n852 3789.35
R949 vss.n852 vss.n802 3789.35
R950 vss.n6438 vss.n6409 3789.35
R951 vss.n6438 vss.n6413 3789.35
R952 vss.n6424 vss.n913 3789.35
R953 vss.n6424 vss.n908 3789.35
R954 vss.n912 vss.n911 3789.35
R955 vss.n911 vss.n907 3789.35
R956 vss.n6553 vss.n6524 3789.35
R957 vss.n6553 vss.n6528 3789.35
R958 vss.n6539 vss.n1088 3789.35
R959 vss.n6539 vss.n1083 3789.35
R960 vss.n1087 vss.n1086 3789.35
R961 vss.n1086 vss.n1082 3789.35
R962 vss.n6550 vss.n6533 3789.35
R963 vss.n6550 vss.n6534 3789.35
R964 vss.n6562 vss.n6518 3789.35
R965 vss.n6562 vss.n6521 3789.35
R966 vss.n6576 vss.n6519 3789.35
R967 vss.n6576 vss.n6575 3789.35
R968 vss.n6435 vss.n6418 3789.35
R969 vss.n6435 vss.n6419 3789.35
R970 vss.n6447 vss.n6403 3789.35
R971 vss.n6447 vss.n6406 3789.35
R972 vss.n6460 vss.n6404 3789.35
R973 vss.n6460 vss.n6459 3789.35
R974 vss.n879 vss.n865 3789.35
R975 vss.n879 vss.n878 3789.35
R976 vss.n15251 vss.n866 3789.35
R977 vss.n15251 vss.n884 3789.35
R978 vss.n15240 vss.n888 3789.35
R979 vss.n891 vss.n888 3789.35
R980 vss.n5363 vss.n5346 3789.35
R981 vss.n5363 vss.n5347 3789.35
R982 vss.n5375 vss.n5331 3789.35
R983 vss.n5375 vss.n5334 3789.35
R984 vss.n5388 vss.n5332 3789.35
R985 vss.n5388 vss.n5387 3789.35
R986 vss.n5151 vss.n5134 3789.35
R987 vss.n5151 vss.n5135 3789.35
R988 vss.n5163 vss.n5119 3789.35
R989 vss.n5163 vss.n5122 3789.35
R990 vss.n5176 vss.n5120 3789.35
R991 vss.n5176 vss.n5175 3789.35
R992 vss.n622 vss.n608 3789.35
R993 vss.n622 vss.n621 3789.35
R994 vss.n15401 vss.n609 3789.35
R995 vss.n15401 vss.n627 3789.35
R996 vss.n15390 vss.n631 3789.35
R997 vss.n634 vss.n631 3789.35
R998 vss.n4888 vss.n4299 3789.35
R999 vss.n4888 vss.n4300 3789.35
R1000 vss.n4900 vss.n4286 3789.35
R1001 vss.n4900 vss.n4289 3789.35
R1002 vss.n4913 vss.n4287 3789.35
R1003 vss.n4913 vss.n4912 3789.35
R1004 vss.n4835 vss.n4834 3789.35
R1005 vss.n4834 vss.n4817 3789.35
R1006 vss.n4847 vss.n4802 3789.35
R1007 vss.n4847 vss.n4751 3789.35
R1008 vss.n4804 vss.n4803 3789.35
R1009 vss.n4803 vss.n4752 3789.35
R1010 vss.n3261 vss.n3234 3789.35
R1011 vss.n3261 vss.n3235 3789.35
R1012 vss.n3245 vss.n1228 3789.35
R1013 vss.n3245 vss.n1223 3789.35
R1014 vss.n1227 vss.n1226 3789.35
R1015 vss.n1226 vss.n1222 3789.35
R1016 vss.n8009 vss.n2431 3789.35
R1017 vss.n8009 vss.n2432 3789.35
R1018 vss.n8019 vss.n2418 3789.35
R1019 vss.n8019 vss.n2367 3789.35
R1020 vss.n2417 vss.n2416 3789.35
R1021 vss.n2416 vss.n2366 3789.35
R1022 vss.n14713 vss.n1380 3789.35
R1023 vss.n14713 vss.n1383 3789.35
R1024 vss.n1395 vss.n1376 3789.35
R1025 vss.n1395 vss.n1324 3789.35
R1026 vss.n1375 vss.n1374 3789.35
R1027 vss.n1374 vss.n1323 3789.35
R1028 vss.n7562 vss.n7533 3789.35
R1029 vss.n7562 vss.n7537 3789.35
R1030 vss.n7548 vss.n1435 3789.35
R1031 vss.n7548 vss.n1430 3789.35
R1032 vss.n1434 vss.n1433 3789.35
R1033 vss.n1433 vss.n1429 3789.35
R1034 vss.n2780 vss.n2751 3789.35
R1035 vss.n2780 vss.n2755 3789.35
R1036 vss.n2766 vss.n1534 3789.35
R1037 vss.n2766 vss.n1529 3789.35
R1038 vss.n1533 vss.n1532 3789.35
R1039 vss.n1532 vss.n1528 3789.35
R1040 vss.n14563 vss.n1637 3789.35
R1041 vss.n14563 vss.n1640 3789.35
R1042 vss.n1652 vss.n1633 3789.35
R1043 vss.n1652 vss.n1582 3789.35
R1044 vss.n1632 vss.n1631 3789.35
R1045 vss.n1631 vss.n1581 3789.35
R1046 vss.n2546 vss.n2517 3789.35
R1047 vss.n2546 vss.n2521 3789.35
R1048 vss.n2534 vss.n1692 3789.35
R1049 vss.n2534 vss.n1687 3789.35
R1050 vss.n1691 vss.n1690 3789.35
R1051 vss.n1690 vss.n1686 3789.35
R1052 vss.n1979 vss.n1871 3789.35
R1053 vss.n1979 vss.n1874 3789.35
R1054 vss.n1884 vss.n1867 3789.35
R1055 vss.n1884 vss.n1862 3789.35
R1056 vss.n1866 vss.n1865 3789.35
R1057 vss.n1865 vss.n1861 3789.35
R1058 vss.n1892 vss.n1878 3789.35
R1059 vss.n1892 vss.n1891 3789.35
R1060 vss.n1972 vss.n1879 3789.35
R1061 vss.n1972 vss.n1896 3789.35
R1062 vss.n1961 vss.n1947 3789.35
R1063 vss.n1950 vss.n1947 3789.35
R1064 vss.n2543 vss.n2525 3789.35
R1065 vss.n2543 vss.n2527 3789.35
R1066 vss.n2555 vss.n2509 3789.35
R1067 vss.n2555 vss.n2514 3789.35
R1068 vss.n2567 vss.n2510 3789.35
R1069 vss.n2567 vss.n2566 3789.35
R1070 vss.n1658 vss.n1644 3789.35
R1071 vss.n1658 vss.n1657 3789.35
R1072 vss.n14556 vss.n1645 3789.35
R1073 vss.n14556 vss.n1663 3789.35
R1074 vss.n14545 vss.n1667 3789.35
R1075 vss.n1670 vss.n1667 3789.35
R1076 vss.n2777 vss.n2760 3789.35
R1077 vss.n2777 vss.n2761 3789.35
R1078 vss.n2789 vss.n2745 3789.35
R1079 vss.n2789 vss.n2748 3789.35
R1080 vss.n2802 vss.n2746 3789.35
R1081 vss.n2802 vss.n2801 3789.35
R1082 vss.n7559 vss.n7542 3789.35
R1083 vss.n7559 vss.n7543 3789.35
R1084 vss.n7571 vss.n7527 3789.35
R1085 vss.n7571 vss.n7530 3789.35
R1086 vss.n7584 vss.n7528 3789.35
R1087 vss.n7584 vss.n7583 3789.35
R1088 vss.n1401 vss.n1387 3789.35
R1089 vss.n1401 vss.n1400 3789.35
R1090 vss.n14706 vss.n1388 3789.35
R1091 vss.n14706 vss.n1406 3789.35
R1092 vss.n14695 vss.n1410 3789.35
R1093 vss.n1413 vss.n1410 3789.35
R1094 vss.n8012 vss.n2424 3789.35
R1095 vss.n8012 vss.n2429 3789.35
R1096 vss.n8000 vss.n2442 3789.35
R1097 vss.n8000 vss.n2443 3789.35
R1098 vss.n6955 vss.n6945 3789.35
R1099 vss.n6955 vss.n6954 3789.35
R1100 vss.n3254 vss.n3238 3789.35
R1101 vss.n3254 vss.n3253 3789.35
R1102 vss.n3269 vss.n3188 3789.35
R1103 vss.n3269 vss.n3189 3789.35
R1104 vss.n3222 vss.n3212 3789.35
R1105 vss.n3222 vss.n3221 3789.35
R1106 vss.n12105 vss.n12104 3789.35
R1107 vss.n12104 vss.n11879 3789.35
R1108 vss.n12090 vss.n11882 3789.35
R1109 vss.n12090 vss.n11878 3789.35
R1110 vss.n11940 vss.n11937 3789.35
R1111 vss.n11940 vss.n11939 3789.35
R1112 vss.n10331 vss.n10330 3789.35
R1113 vss.n10330 vss.n10280 3789.35
R1114 vss.n10336 vss.n10329 3789.35
R1115 vss.n10336 vss.n10279 3789.35
R1116 vss.n10339 vss.n10334 3789.35
R1117 vss.n10339 vss.n10338 3789.35
R1118 vss.n9780 vss.n8736 3549.33
R1119 vss.n12334 vss.n8686 3549.33
R1120 vss.n9651 vss.n9650 3549.33
R1121 vss.n12453 vss.n9206 3549.33
R1122 vss.n9521 vss.n9275 3549.33
R1123 vss.n9459 vss.n9279 3549.33
R1124 vss.n12216 vss.n8805 3549.33
R1125 vss.n5703 vss.n3661 3549.33
R1126 vss.n5941 vss.n3729 3549.33
R1127 vss.n5811 vss.n3780 3549.33
R1128 vss.n6180 vss.n3848 3549.33
R1129 vss.n6051 vss.n3899 3549.33
R1130 vss.n6232 vss.n3967 3549.33
R1131 vss.n6703 vss.n6702 3549.33
R1132 vss.n3463 vss.n3331 3549.33
R1133 vss.n5280 vss.n3327 3549.33
R1134 vss.n5495 vss.n3323 3549.33
R1135 vss.n5069 vss.n3319 3549.33
R1136 vss.n5021 vss.n3315 3549.33
R1137 vss.n4516 vss.n3311 3549.33
R1138 vss.n15073 vss.n408 3549.33
R1139 vss.n7468 vss.n416 3549.33
R1140 vss.n7371 vss.n420 3549.33
R1141 vss.n7286 vss.n424 3549.33
R1142 vss.n4642 vss.n428 3549.33
R1143 vss.n4595 vss.n432 3549.33
R1144 vss.n7945 vss.n7944 3549.33
R1145 vss.n7887 vss.n2482 3549.33
R1146 vss.n7741 vss.n2478 3549.33
R1147 vss.n7692 vss.n2474 3549.33
R1148 vss.n2998 vss.n2469 3549.33
R1149 vss.n7123 vss.n7122 3549.33
R1150 vss.n6919 vss.n6918 3549.33
R1151 vss.n14378 vss.n1187 3549.33
R1152 vss.n13933 vss.n1195 3549.33
R1153 vss.n8200 vss.n1199 3549.33
R1154 vss.n14050 vss.n1203 3549.33
R1155 vss.n8072 vss.n1207 3549.33
R1156 vss.n2313 vss.n1211 3549.33
R1157 vss.n2077 vss.n2074 3549.33
R1158 vss.n13627 vss.n2104 3549.33
R1159 vss.n8277 vss.n2108 3549.33
R1160 vss.n13816 vss.n2112 3549.33
R1161 vss.n9063 vss.n2116 3549.33
R1162 vss.n13104 vss.n2120 3549.33
R1163 vss.n12601 vss.n2124 3549.33
R1164 vss.n14466 vss.n1191 3549.33
R1165 vss.n15161 vss.n412 3549.33
R1166 vss.n6313 vss.n6312 3549.33
R1167 vss.n9901 vss.n8838 3549.33
R1168 vss.n11585 vss.n8842 3549.33
R1169 vss.n11132 vss.n8846 3549.33
R1170 vss.n11274 vss.n8850 3549.33
R1171 vss.n10935 vss.n8854 3549.33
R1172 vss.n10839 vss.n8858 3549.33
R1173 vss.n10541 vss.n8862 3549.33
R1174 vss.n11726 vss.n8835 3445.36
R1175 vss.n10362 vss.n10361 3444.61
R1176 vss.n15855 vss.n15854 3272.21
R1177 vss.n15828 vss.n15827 3272.21
R1178 vss.n15799 vss.n15798 3272.21
R1179 vss.n15772 vss.n15771 3272.21
R1180 vss.n15743 vss.n15742 3272.21
R1181 vss.n15716 vss.n15715 3272.21
R1182 vss.n15687 vss.n15686 3272.21
R1183 vss.n10395 vss.n10386 3272.21
R1184 vss.n10785 vss.n10635 3272.21
R1185 vss.n10764 vss.n10763 3272.21
R1186 vss.n11037 vss.n11028 3272.21
R1187 vss.n11323 vss.n11322 3272.21
R1188 vss.n11442 vss.n11348 3272.21
R1189 vss.n11679 vss.n9929 3272.21
R1190 vss.n13249 vss.n8810 3245.44
R1191 vss.n14789 vss.n1184 3154.67
R1192 vss.n15484 vss.n405 3154.67
R1193 vss.n15657 vss.n15656 3154.67
R1194 vss.n14790 vss.n14789 2943.95
R1195 vss.n15485 vss.n15484 2943.95
R1196 vss.n15658 vss.n15657 2943.95
R1197 vss.n9781 vss.n9780 2918.71
R1198 vss.n12334 vss.n12333 2918.71
R1199 vss.n9652 vss.n9651 2918.71
R1200 vss.n12453 vss.n12452 2918.71
R1201 vss.n9522 vss.n9521 2918.71
R1202 vss.n9460 vss.n9459 2918.71
R1203 vss.n12216 vss.n12215 2918.71
R1204 vss.n5703 vss.n5702 2918.71
R1205 vss.n5941 vss.n5940 2918.71
R1206 vss.n5812 vss.n5811 2918.71
R1207 vss.n6180 vss.n6179 2918.71
R1208 vss.n6052 vss.n6051 2918.71
R1209 vss.n6232 vss.n6231 2918.71
R1210 vss.n6702 vss.n3336 2918.71
R1211 vss.n3464 vss.n3463 2918.71
R1212 vss.n5280 vss.n5279 2918.71
R1213 vss.n5495 vss.n5494 2918.71
R1214 vss.n5069 vss.n5068 2918.71
R1215 vss.n5021 vss.n5020 2918.71
R1216 vss.n4516 vss.n4515 2918.71
R1217 vss.n15073 vss.n15072 2918.71
R1218 vss.n7468 vss.n7467 2918.71
R1219 vss.n7372 vss.n7371 2918.71
R1220 vss.n7290 vss.n7286 2918.71
R1221 vss.n4643 vss.n4642 2918.71
R1222 vss.n4596 vss.n4595 2918.71
R1223 vss.n7944 vss.n7927 2918.71
R1224 vss.n7887 vss.n7886 2918.71
R1225 vss.n7741 vss.n7740 2918.71
R1226 vss.n7692 vss.n7691 2918.71
R1227 vss.n2998 vss.n2997 2918.71
R1228 vss.n7122 vss.n7078 2918.71
R1229 vss.n6918 vss.n6826 2918.71
R1230 vss.n14378 vss.n14377 2918.71
R1231 vss.n13933 vss.n13932 2918.71
R1232 vss.n8201 vss.n8200 2918.71
R1233 vss.n14050 vss.n14049 2918.71
R1234 vss.n8073 vss.n8072 2918.71
R1235 vss.n2314 vss.n2313 2918.71
R1236 vss.n2078 vss.n2077 2918.71
R1237 vss.n13627 vss.n13626 2918.71
R1238 vss.n8277 vss.n8276 2918.71
R1239 vss.n13816 vss.n13815 2918.71
R1240 vss.n9063 vss.n9062 2918.71
R1241 vss.n13104 vss.n13103 2918.71
R1242 vss.n12601 vss.n12600 2918.71
R1243 vss.n14467 vss.n14466 2918.71
R1244 vss.n15162 vss.n15161 2918.71
R1245 vss.n6313 vss.n3563 2918.71
R1246 vss.n9902 vss.n9901 2918.71
R1247 vss.n11585 vss.n11584 2918.71
R1248 vss.n11132 vss.n11131 2918.71
R1249 vss.n11274 vss.n11273 2918.71
R1250 vss.n10935 vss.n10934 2918.71
R1251 vss.n10839 vss.n10838 2918.71
R1252 vss.n10541 vss.n10540 2918.71
R1253 vss.n14869 vss.n404 2869.13
R1254 vss.n15546 vss.n352 2869.13
R1255 vss.n14790 vss.n1160 2862.9
R1256 vss.n15485 vss.n381 2862.9
R1257 vss.n15659 vss.n15658 2862.9
R1258 vss.n13225 vss.n13224 2820.86
R1259 vss.n15855 vss.n25 2813.68
R1260 vss.n15829 vss.n15828 2813.68
R1261 vss.n15799 vss.n122 2813.68
R1262 vss.n15773 vss.n15772 2813.68
R1263 vss.n15743 vss.n200 2813.68
R1264 vss.n15717 vss.n15716 2813.68
R1265 vss.n15687 vss.n279 2813.68
R1266 vss.n10395 vss.n10394 2813.68
R1267 vss.n10785 vss.n10784 2813.68
R1268 vss.n10763 vss.n10762 2813.68
R1269 vss.n11037 vss.n11036 2813.68
R1270 vss.n11324 vss.n11323 2813.68
R1271 vss.n11442 vss.n11441 2813.68
R1272 vss.n11679 vss.n11678 2813.68
R1273 vss.n13223 vss.n13222 2602
R1274 vss.n12183 vss.n8809 2458.67
R1275 vss.n1160 vss.n1159 2458.67
R1276 vss.n381 vss.n380 2458.67
R1277 vss.n9754 vss.n9753 2376.04
R1278 vss.n9624 vss.n9623 2376.04
R1279 vss.n9495 vss.n9494 2376.04
R1280 vss.n5557 vss.n5556 2376.04
R1281 vss.n5745 vss.n5744 2376.04
R1282 vss.n5985 vss.n5984 2376.04
R1283 vss.n6368 vss.n6367 2376.04
R1284 vss.n5528 vss.n4005 2376.04
R1285 vss.n4212 vss.n4211 2376.04
R1286 vss.n4483 vss.n4479 2376.04
R1287 vss.n14910 vss.n14909 2376.04
R1288 vss.n3080 vss.n3079 2376.04
R1289 vss.n4671 vss.n4670 2376.04
R1290 vss.n2673 vss.n2672 2376.04
R1291 vss.n2923 vss.n2922 2376.04
R1292 vss.n7984 vss.n7983 2376.04
R1293 vss.n7215 vss.n3135 2376.04
R1294 vss.n14215 vss.n14214 2376.04
R1295 vss.n8174 vss.n8173 2376.04
R1296 vss.n2247 vss.n2246 2376.04
R1297 vss.n13594 vss.n13589 2376.04
R1298 vss.n13783 vss.n13778 2376.04
R1299 vss.n13071 vss.n13066 2376.04
R1300 vss.n14077 vss.n2178 2376.04
R1301 vss.n14412 vss.n14400 2376.04
R1302 vss.n15107 vss.n15095 2376.04
R1303 vss.n3590 vss.n3589 2376.04
R1304 vss.n11552 vss.n11547 2376.04
R1305 vss.n11241 vss.n11236 2376.04
R1306 vss.n10902 vss.n10897 2376.04
R1307 vss.n10508 vss.n10503 2376.04
R1308 vss.n11732 vss.n11731 2376
R1309 vss.n12182 vss.n2052 2320.72
R1310 vss.n11793 vss.n11792 2189.03
R1311 vss.n13198 vss.n8867 2172.79
R1312 vss.n13198 vss.n8868 2172.79
R1313 vss.n10360 vss.n10345 2172.79
R1314 vss.n10360 vss.n10344 2172.79
R1315 vss.n10311 vss.n10299 2172.79
R1316 vss.n10309 vss.n10299 2172.79
R1317 vss.n10325 vss.n10283 2172.79
R1318 vss.n10325 vss.n10282 2172.79
R1319 vss.n11633 vss.n11621 2172.79
R1320 vss.n11631 vss.n11621 2172.79
R1321 vss.n11647 vss.n9950 2172.79
R1322 vss.n11647 vss.n9949 2172.79
R1323 vss.n11685 vss.n9925 2172.79
R1324 vss.n11683 vss.n9925 2172.79
R1325 vss.n11697 vss.n11695 2172.79
R1326 vss.n11699 vss.n11695 2172.79
R1327 vss.n11448 vss.n9980 2172.79
R1328 vss.n11446 vss.n9980 2172.79
R1329 vss.n11460 vss.n11458 2172.79
R1330 vss.n11462 vss.n11458 2172.79
R1331 vss.n11410 vss.n11367 2172.79
R1332 vss.n11410 vss.n11368 2172.79
R1333 vss.n11391 vss.n11389 2172.79
R1334 vss.n11393 vss.n11389 2172.79
R1335 vss.n11179 vss.n11171 2172.79
R1336 vss.n11177 vss.n11171 2172.79
R1337 vss.n11191 vss.n11189 2172.79
R1338 vss.n11193 vss.n11189 2172.79
R1339 vss.n11043 vss.n10140 2172.79
R1340 vss.n11041 vss.n10140 2172.79
R1341 vss.n11055 vss.n11053 2172.79
R1342 vss.n11057 vss.n11053 2172.79
R1343 vss.n10103 vss.n10094 2172.79
R1344 vss.n10101 vss.n10094 2172.79
R1345 vss.n10115 vss.n10113 2172.79
R1346 vss.n10117 vss.n10113 2172.79
R1347 vss.n10753 vss.n10711 2172.79
R1348 vss.n10753 vss.n10712 2172.79
R1349 vss.n10734 vss.n10731 2172.79
R1350 vss.n10736 vss.n10731 2172.79
R1351 vss.n10791 vss.n10227 2172.79
R1352 vss.n10789 vss.n10227 2172.79
R1353 vss.n10803 vss.n10801 2172.79
R1354 vss.n10805 vss.n10801 2172.79
R1355 vss.n10698 vss.n10655 2172.79
R1356 vss.n10698 vss.n10656 2172.79
R1357 vss.n10679 vss.n10677 2172.79
R1358 vss.n10681 vss.n10677 2172.79
R1359 vss.n10401 vss.n10269 2172.79
R1360 vss.n10399 vss.n10269 2172.79
R1361 vss.n10413 vss.n10411 2172.79
R1362 vss.n10415 vss.n10411 2172.79
R1363 vss.n10507 vss.n10506 2172.79
R1364 vss.n10491 vss.n10485 2172.79
R1365 vss.n10493 vss.n10485 2172.79
R1366 vss.n10554 vss.n10552 2172.79
R1367 vss.n10556 vss.n10552 2172.79
R1368 vss.n10542 vss.n10533 2172.79
R1369 vss.n10852 vss.n10850 2172.79
R1370 vss.n10855 vss.n10850 2172.79
R1371 vss.n10840 vss.n10831 2172.79
R1372 vss.n10901 vss.n10900 2172.79
R1373 vss.n10885 vss.n10879 2172.79
R1374 vss.n10887 vss.n10879 2172.79
R1375 vss.n10948 vss.n10946 2172.79
R1376 vss.n10950 vss.n10946 2172.79
R1377 vss.n10936 vss.n10927 2172.79
R1378 vss.n11287 vss.n11285 2172.79
R1379 vss.n11290 vss.n11285 2172.79
R1380 vss.n11275 vss.n11266 2172.79
R1381 vss.n11240 vss.n11239 2172.79
R1382 vss.n11224 vss.n11218 2172.79
R1383 vss.n11226 vss.n11218 2172.79
R1384 vss.n11145 vss.n11143 2172.79
R1385 vss.n11147 vss.n11143 2172.79
R1386 vss.n11133 vss.n11124 2172.79
R1387 vss.n11598 vss.n11596 2172.79
R1388 vss.n11601 vss.n11596 2172.79
R1389 vss.n11586 vss.n11577 2172.79
R1390 vss.n11551 vss.n11550 2172.79
R1391 vss.n11535 vss.n11529 2172.79
R1392 vss.n11537 vss.n11529 2172.79
R1393 vss.n11724 vss.n9880 2172.79
R1394 vss.n11724 vss.n9881 2172.79
R1395 vss.n9900 vss.n9898 2172.79
R1396 vss.n13227 vss.n8833 2172.79
R1397 vss.n13229 vss.n8833 2172.79
R1398 vss.n13247 vss.n8812 2172.79
R1399 vss.n13247 vss.n8813 2172.79
R1400 vss.n11794 vss.n11766 2172.79
R1401 vss.n11785 vss.n11777 2172.79
R1402 vss.n11777 vss.n11764 2172.79
R1403 vss.n11816 vss.n11811 2172.79
R1404 vss.n11839 vss.n11811 2172.79
R1405 vss.n11831 vss.n11822 2172.79
R1406 vss.n11822 vss.n11810 2172.79
R1407 vss.n11913 vss.n11911 2172.79
R1408 vss.n11915 vss.n11911 2172.79
R1409 vss.n11933 vss.n11890 2172.79
R1410 vss.n11933 vss.n11891 2172.79
R1411 vss.n11729 vss.n9875 2172.79
R1412 vss.n11734 vss.n9875 2172.79
R1413 vss.n11748 vss.n11744 2172.79
R1414 vss.n11746 vss.n11744 2172.79
R1415 vss.n9444 vss.n9437 2172.79
R1416 vss.n9446 vss.n9437 2172.79
R1417 vss.n9458 vss.n9456 2172.79
R1418 vss.n12477 vss.n9487 2172.79
R1419 vss.n12491 vss.n12487 2172.79
R1420 vss.n12489 vss.n12487 2172.79
R1421 vss.n9541 vss.n9497 2172.79
R1422 vss.n9541 vss.n9498 2172.79
R1423 vss.n9523 vss.n9518 2172.79
R1424 vss.n9560 vss.n9547 2172.79
R1425 vss.n9574 vss.n9572 2172.79
R1426 vss.n9576 vss.n9572 2172.79
R1427 vss.n9592 vss.n9547 2172.79
R1428 vss.n9258 vss.n9256 2172.79
R1429 vss.n13168 vss.n8898 2172.79
R1430 vss.n13166 vss.n8898 2172.79
R1431 vss.n9272 vss.n9256 2172.79
R1432 vss.n12402 vss.n12396 2172.79
R1433 vss.n12419 vss.n12414 2172.79
R1434 vss.n12417 vss.n12414 2172.79
R1435 vss.n12404 vss.n12396 2172.79
R1436 vss.n12358 vss.n9616 2172.79
R1437 vss.n12372 vss.n12368 2172.79
R1438 vss.n12370 vss.n12368 2172.79
R1439 vss.n9671 vss.n9626 2172.79
R1440 vss.n9671 vss.n9627 2172.79
R1441 vss.n9653 vss.n9647 2172.79
R1442 vss.n9689 vss.n9676 2172.79
R1443 vss.n9704 vss.n9701 2172.79
R1444 vss.n9706 vss.n9701 2172.79
R1445 vss.n9722 vss.n9676 2172.79
R1446 vss.n13264 vss.n8633 2172.79
R1447 vss.n13280 vss.n13276 2172.79
R1448 vss.n13278 vss.n13276 2172.79
R1449 vss.n13266 vss.n8633 2172.79
R1450 vss.n12284 vss.n12278 2172.79
R1451 vss.n12301 vss.n12296 2172.79
R1452 vss.n12299 vss.n12296 2172.79
R1453 vss.n12286 vss.n12278 2172.79
R1454 vss.n12240 vss.n9746 2172.79
R1455 vss.n12254 vss.n12250 2172.79
R1456 vss.n12252 vss.n12250 2172.79
R1457 vss.n9800 vss.n9756 2172.79
R1458 vss.n9800 vss.n9757 2172.79
R1459 vss.n9782 vss.n9777 2172.79
R1460 vss.n9818 vss.n9805 2172.79
R1461 vss.n9832 vss.n9830 2172.79
R1462 vss.n9834 vss.n9830 2172.79
R1463 vss.n9850 vss.n9805 2172.79
R1464 vss.n8740 vss.n8738 2172.79
R1465 vss.n13691 vss.n8354 2172.79
R1466 vss.n13689 vss.n8354 2172.79
R1467 vss.n8754 vss.n8738 2172.79
R1468 vss.n11986 vss.n11984 2172.79
R1469 vss.n12006 vss.n11964 2172.79
R1470 vss.n12006 vss.n11965 2172.79
R1471 vss.n11988 vss.n11984 2172.79
R1472 vss.n9854 vss.n9852 2172.79
R1473 vss.n12217 vss.n12212 2172.79
R1474 vss.n12233 vss.n9852 2172.79
R1475 vss.n8759 vss.n8757 2172.79
R1476 vss.n8784 vss.n8781 2172.79
R1477 vss.n8786 vss.n8781 2172.79
R1478 vss.n8802 vss.n8757 2172.79
R1479 vss.n8691 vss.n8689 2172.79
R1480 vss.n8715 vss.n8712 2172.79
R1481 vss.n8717 vss.n8712 2172.79
R1482 vss.n8733 vss.n8689 2172.79
R1483 vss.n9726 vss.n9724 2172.79
R1484 vss.n12335 vss.n12330 2172.79
R1485 vss.n12351 vss.n9724 2172.79
R1486 vss.n8640 vss.n8638 2172.79
R1487 vss.n8665 vss.n8662 2172.79
R1488 vss.n8667 vss.n8662 2172.79
R1489 vss.n8683 vss.n8638 2172.79
R1490 vss.n12918 vss.n9204 2172.79
R1491 vss.n12938 vss.n9183 2172.79
R1492 vss.n12938 vss.n9184 2172.79
R1493 vss.n12920 vss.n9204 2172.79
R1494 vss.n9596 vss.n9594 2172.79
R1495 vss.n12454 vss.n12449 2172.79
R1496 vss.n12470 vss.n9594 2172.79
R1497 vss.n9210 vss.n9208 2172.79
R1498 vss.n9235 vss.n9232 2172.79
R1499 vss.n9237 vss.n9232 2172.79
R1500 vss.n9253 vss.n9208 2172.79
R1501 vss.n9336 vss.n9334 2172.79
R1502 vss.n9356 vss.n9312 2172.79
R1503 vss.n9356 vss.n9313 2172.79
R1504 vss.n9338 vss.n9334 2172.79
R1505 vss.n12522 vss.n12520 2172.79
R1506 vss.n12542 vss.n9419 2172.79
R1507 vss.n12542 vss.n9420 2172.79
R1508 vss.n12524 vss.n12520 2172.79
R1509 vss.n12672 vss.n12670 2172.79
R1510 vss.n12692 vss.n12649 2172.79
R1511 vss.n12692 vss.n12650 2172.79
R1512 vss.n12674 vss.n12670 2172.79
R1513 vss.n10191 vss.n10183 2172.79
R1514 vss.n10189 vss.n10183 2172.79
R1515 vss.n10200 vss.n9546 2172.79
R1516 vss.n10204 vss.n9546 2172.79
R1517 vss.n11088 vss.n11080 2172.79
R1518 vss.n11086 vss.n11080 2172.79
R1519 vss.n11097 vss.n9675 2172.79
R1520 vss.n11101 vss.n9675 2172.79
R1521 vss.n11493 vss.n11485 2172.79
R1522 vss.n11491 vss.n11485 2172.79
R1523 vss.n11502 vss.n9804 2172.79
R1524 vss.n11506 vss.n9804 2172.79
R1525 vss.n12179 vss.n12134 2172.79
R1526 vss.n12179 vss.n12135 2172.79
R1527 vss.n12160 vss.n12158 2172.79
R1528 vss.n12162 vss.n12158 2172.79
R1529 vss.n15639 vss.n15627 2172.79
R1530 vss.n15639 vss.n356 2172.79
R1531 vss.n15650 vss.n15649 2172.79
R1532 vss.n15650 vss.n355 2172.79
R1533 vss.n3592 vss.n3586 2172.79
R1534 vss.n3610 vss.n3565 2172.79
R1535 vss.n3610 vss.n3566 2172.79
R1536 vss.n3986 vss.n3970 2172.79
R1537 vss.n3986 vss.n3971 2172.79
R1538 vss.n15895 vss.n14 2172.79
R1539 vss.n15893 vss.n14 2172.79
R1540 vss.n6308 vss.n6292 2172.79
R1541 vss.n6308 vss.n6293 2172.79
R1542 vss.n15692 vss.n258 2172.79
R1543 vss.n15690 vss.n258 2172.79
R1544 vss.n5652 vss.n5646 2172.79
R1545 vss.n5668 vss.n5664 2172.79
R1546 vss.n5666 vss.n5664 2172.79
R1547 vss.n5654 vss.n5646 2172.79
R1548 vss.n3712 vss.n3710 2172.79
R1549 vss.n15748 vss.n179 2172.79
R1550 vss.n15746 vss.n179 2172.79
R1551 vss.n3726 vss.n3710 2172.79
R1552 vss.n3665 vss.n3663 2172.79
R1553 vss.n3689 vss.n3686 2172.79
R1554 vss.n3691 vss.n3686 2172.79
R1555 vss.n3707 vss.n3663 2172.79
R1556 vss.n5844 vss.n5838 2172.79
R1557 vss.n5860 vss.n5856 2172.79
R1558 vss.n5858 vss.n5856 2172.79
R1559 vss.n5846 vss.n5838 2172.79
R1560 vss.n3831 vss.n3829 2172.79
R1561 vss.n15804 vss.n101 2172.79
R1562 vss.n15802 vss.n101 2172.79
R1563 vss.n3845 vss.n3829 2172.79
R1564 vss.n3784 vss.n3782 2172.79
R1565 vss.n3808 vss.n3805 2172.79
R1566 vss.n3810 vss.n3805 2172.79
R1567 vss.n3826 vss.n3782 2172.79
R1568 vss.n3903 vss.n3901 2172.79
R1569 vss.n3927 vss.n3924 2172.79
R1570 vss.n3929 vss.n3924 2172.79
R1571 vss.n3945 vss.n3901 2172.79
R1572 vss.n6084 vss.n6078 2172.79
R1573 vss.n6100 vss.n6096 2172.79
R1574 vss.n6098 vss.n6096 2172.79
R1575 vss.n6086 vss.n6078 2172.79
R1576 vss.n6036 vss.n6030 2172.79
R1577 vss.n6038 vss.n6030 2172.79
R1578 vss.n6050 vss.n6048 2172.79
R1579 vss.n6198 vss.n6153 2172.79
R1580 vss.n6198 vss.n6154 2172.79
R1581 vss.n6181 vss.n6176 2172.79
R1582 vss.n5752 vss.n5743 2172.79
R1583 vss.n5766 vss.n5762 2172.79
R1584 vss.n5764 vss.n5762 2172.79
R1585 vss.n5796 vss.n5790 2172.79
R1586 vss.n5798 vss.n5790 2172.79
R1587 vss.n5810 vss.n5808 2172.79
R1588 vss.n5959 vss.n5914 2172.79
R1589 vss.n5959 vss.n5915 2172.79
R1590 vss.n5942 vss.n5937 2172.79
R1591 vss.n5564 vss.n5555 2172.79
R1592 vss.n5578 vss.n5574 2172.79
R1593 vss.n5576 vss.n5574 2172.79
R1594 vss.n5721 vss.n5537 2172.79
R1595 vss.n5721 vss.n5538 2172.79
R1596 vss.n5704 vss.n5699 2172.79
R1597 vss.n6331 vss.n3537 2172.79
R1598 vss.n6331 vss.n3538 2172.79
R1599 vss.n6314 vss.n3560 2172.79
R1600 vss.n5603 vss.n3487 2172.79
R1601 vss.n5623 vss.n5619 2172.79
R1602 vss.n5621 vss.n5619 2172.79
R1603 vss.n5609 vss.n3487 2172.79
R1604 vss.n5879 vss.n4003 2172.79
R1605 vss.n5893 vss.n5891 2172.79
R1606 vss.n5895 vss.n5891 2172.79
R1607 vss.n5911 vss.n4003 2172.79
R1608 vss.n6118 vss.n3995 2172.79
R1609 vss.n6132 vss.n6130 2172.79
R1610 vss.n6134 vss.n6130 2172.79
R1611 vss.n6150 vss.n3995 2172.79
R1612 vss.n5992 vss.n5983 2172.79
R1613 vss.n6006 vss.n6002 2172.79
R1614 vss.n6004 vss.n6002 2172.79
R1615 vss.n3296 vss.n3288 2172.79
R1616 vss.n3294 vss.n3288 2172.79
R1617 vss.n6728 vss.n3306 2172.79
R1618 vss.n6730 vss.n3306 2172.79
R1619 vss.n4552 vss.n4367 2172.79
R1620 vss.n4552 vss.n4368 2172.79
R1621 vss.n4391 vss.n4389 2172.79
R1622 vss.n4393 vss.n4389 2172.79
R1623 vss.n4482 vss.n4481 2172.79
R1624 vss.n4467 vss.n4461 2172.79
R1625 vss.n4469 vss.n4461 2172.79
R1626 vss.n4529 vss.n4527 2172.79
R1627 vss.n4531 vss.n4527 2172.79
R1628 vss.n4517 vss.n4508 2172.79
R1629 vss.n5034 vss.n5032 2172.79
R1630 vss.n5036 vss.n5032 2172.79
R1631 vss.n5022 vss.n5013 2172.79
R1632 vss.n4214 vss.n4213 2172.79
R1633 vss.n4192 vss.n4186 2172.79
R1634 vss.n4194 vss.n4186 2172.79
R1635 vss.n5082 vss.n5080 2172.79
R1636 vss.n5084 vss.n5080 2172.79
R1637 vss.n5070 vss.n5061 2172.79
R1638 vss.n5508 vss.n5506 2172.79
R1639 vss.n5510 vss.n5506 2172.79
R1640 vss.n5496 vss.n5487 2172.79
R1641 vss.n5533 vss.n4007 2172.79
R1642 vss.n4029 vss.n4025 2172.79
R1643 vss.n4027 vss.n4025 2172.79
R1644 vss.n5293 vss.n5291 2172.79
R1645 vss.n5296 vss.n5291 2172.79
R1646 vss.n5281 vss.n5272 2172.79
R1647 vss.n3485 vss.n3442 2172.79
R1648 vss.n3485 vss.n3443 2172.79
R1649 vss.n3462 vss.n3459 2172.79
R1650 vss.n6370 vss.n3440 2172.79
R1651 vss.n6353 vss.n6342 2172.79
R1652 vss.n6355 vss.n6342 2172.79
R1653 vss.n6684 vss.n6683 2172.79
R1654 vss.n6683 vss.n6682 2172.79
R1655 vss.n6701 vss.n3337 2172.79
R1656 vss.n6637 vss.n6629 2172.79
R1657 vss.n6635 vss.n6629 2172.79
R1658 vss.n6649 vss.n6647 2172.79
R1659 vss.n6651 vss.n6647 2172.79
R1660 vss.n6588 vss.n6511 2172.79
R1661 vss.n6586 vss.n6511 2172.79
R1662 vss.n6601 vss.n6598 2172.79
R1663 vss.n6603 vss.n6598 2172.79
R1664 vss.n5235 vss.n5227 2172.79
R1665 vss.n5233 vss.n5227 2172.79
R1666 vss.n5247 vss.n5245 2172.79
R1667 vss.n5249 vss.n5245 2172.79
R1668 vss.n4060 vss.n4052 2172.79
R1669 vss.n4058 vss.n4052 2172.79
R1670 vss.n4069 vss.n4002 2172.79
R1671 vss.n4073 vss.n4002 2172.79
R1672 vss.n5447 vss.n5439 2172.79
R1673 vss.n5445 vss.n5439 2172.79
R1674 vss.n5459 vss.n5457 2172.79
R1675 vss.n5461 vss.n5457 2172.79
R1676 vss.n5400 vss.n5324 2172.79
R1677 vss.n5398 vss.n5324 2172.79
R1678 vss.n5412 vss.n5410 2172.79
R1679 vss.n5414 vss.n5410 2172.79
R1680 vss.n4150 vss.n4142 2172.79
R1681 vss.n4148 vss.n4142 2172.79
R1682 vss.n4162 vss.n4160 2172.79
R1683 vss.n4164 vss.n4160 2172.79
R1684 vss.n4241 vss.n4233 2172.79
R1685 vss.n4239 vss.n4233 2172.79
R1686 vss.n4250 vss.n3994 2172.79
R1687 vss.n4254 vss.n3994 2172.79
R1688 vss.n4973 vss.n4965 2172.79
R1689 vss.n4971 vss.n4965 2172.79
R1690 vss.n4985 vss.n4983 2172.79
R1691 vss.n4987 vss.n4983 2172.79
R1692 vss.n4104 vss.n4096 2172.79
R1693 vss.n4102 vss.n4096 2172.79
R1694 vss.n4116 vss.n4114 2172.79
R1695 vss.n4118 vss.n4114 2172.79
R1696 vss.n4925 vss.n4279 2172.79
R1697 vss.n4923 vss.n4279 2172.79
R1698 vss.n4937 vss.n4935 2172.79
R1699 vss.n4939 vss.n4935 2172.79
R1700 vss.n5188 vss.n5112 2172.79
R1701 vss.n5186 vss.n5112 2172.79
R1702 vss.n5200 vss.n5198 2172.79
R1703 vss.n5202 vss.n5198 2172.79
R1704 vss.n3363 vss.n3355 2172.79
R1705 vss.n3361 vss.n3355 2172.79
R1706 vss.n3375 vss.n3373 2172.79
R1707 vss.n3377 vss.n3373 2172.79
R1708 vss.n3410 vss.n3402 2172.79
R1709 vss.n3408 vss.n3402 2172.79
R1710 vss.n3422 vss.n3420 2172.79
R1711 vss.n3424 vss.n3420 2172.79
R1712 vss.n3509 vss.n3507 2172.79
R1713 vss.n3511 vss.n3507 2172.79
R1714 vss.n3533 vss.n3489 2172.79
R1715 vss.n3533 vss.n3490 2172.79
R1716 vss.n6472 vss.n6396 2172.79
R1717 vss.n6470 vss.n6396 2172.79
R1718 vss.n6484 vss.n6482 2172.79
R1719 vss.n6486 vss.n6482 2172.79
R1720 vss.n4423 vss.n4415 2172.79
R1721 vss.n4421 vss.n4415 2172.79
R1722 vss.n4435 vss.n4433 2172.79
R1723 vss.n4437 vss.n4433 2172.79
R1724 vss.n4798 vss.n4754 2172.79
R1725 vss.n4798 vss.n4755 2172.79
R1726 vss.n4778 vss.n4776 2172.79
R1727 vss.n4780 vss.n4776 2172.79
R1728 vss.n14991 vss.n14986 2172.79
R1729 vss.n15014 vss.n14986 2172.79
R1730 vss.n15006 vss.n14997 2172.79
R1731 vss.n14997 vss.n14985 2172.79
R1732 vss.n15520 vss.n15518 2172.79
R1733 vss.n15522 vss.n15518 2172.79
R1734 vss.n15540 vss.n384 2172.79
R1735 vss.n15540 vss.n385 2172.79
R1736 vss.n14867 vss.n14851 2172.79
R1737 vss.n14867 vss.n14852 2172.79
R1738 vss.n15490 vss.n403 2172.79
R1739 vss.n15488 vss.n403 2172.79
R1740 vss.n14958 vss.n14946 2172.79
R1741 vss.n14958 vss.n14957 2172.79
R1742 vss.n14967 vss.n14941 2172.79
R1743 vss.n14971 vss.n14941 2172.79
R1744 vss.n1061 vss.n1055 2172.79
R1745 vss.n15040 vss.n1073 2172.79
R1746 vss.n15038 vss.n1073 2172.79
R1747 vss.n1063 vss.n1055 2172.79
R1748 vss.n15146 vss.n980 2172.79
R1749 vss.n15148 vss.n980 2172.79
R1750 vss.n15160 vss.n15158 2172.79
R1751 vss.n14912 vss.n14902 2172.79
R1752 vss.n14926 vss.n14922 2172.79
R1753 vss.n14924 vss.n14922 2172.79
R1754 vss.n4580 vss.n4573 2172.79
R1755 vss.n4582 vss.n4573 2172.79
R1756 vss.n4594 vss.n4592 2172.79
R1757 vss.n4678 vss.n4669 2172.79
R1758 vss.n4692 vss.n4688 2172.79
R1759 vss.n4690 vss.n4688 2172.79
R1760 vss.n4627 vss.n4621 2172.79
R1761 vss.n4629 vss.n4621 2172.79
R1762 vss.n4641 vss.n4639 2172.79
R1763 vss.n7236 vss.n3128 2172.79
R1764 vss.n7250 vss.n7248 2172.79
R1765 vss.n7252 vss.n7248 2172.79
R1766 vss.n7268 vss.n3128 2172.79
R1767 vss.n523 vss.n517 2172.79
R1768 vss.n15434 vss.n535 2172.79
R1769 vss.n15432 vss.n535 2172.79
R1770 vss.n525 vss.n517 2172.79
R1771 vss.n7321 vss.n7315 2172.79
R1772 vss.n7337 vss.n7333 2172.79
R1773 vss.n7335 vss.n7333 2172.79
R1774 vss.n7323 vss.n7315 2172.79
R1775 vss.n3087 vss.n3078 2172.79
R1776 vss.n3101 vss.n3097 2172.79
R1777 vss.n3099 vss.n3097 2172.79
R1778 vss.n7391 vss.n3060 2172.79
R1779 vss.n7391 vss.n3061 2172.79
R1780 vss.n7373 vss.n7368 2172.79
R1781 vss.n7406 vss.n7394 2172.79
R1782 vss.n7420 vss.n7418 2172.79
R1783 vss.n7422 vss.n7418 2172.79
R1784 vss.n7438 vss.n7394 2172.79
R1785 vss.n728 vss.n722 2172.79
R1786 vss.n15361 vss.n740 2172.79
R1787 vss.n15359 vss.n740 2172.79
R1788 vss.n730 vss.n722 2172.79
R1789 vss.n781 vss.n775 2172.79
R1790 vss.n15284 vss.n793 2172.79
R1791 vss.n15282 vss.n793 2172.79
R1792 vss.n783 vss.n775 2172.79
R1793 vss.n15140 vss.n15096 2172.79
R1794 vss.n15122 vss.n15120 2172.79
R1795 vss.n15124 vss.n15120 2172.79
R1796 vss.n15195 vss.n15189 2172.79
R1797 vss.n15211 vss.n15207 2172.79
R1798 vss.n15209 vss.n15207 2172.79
R1799 vss.n15197 vss.n15189 2172.79
R1800 vss.n938 vss.n932 2172.79
R1801 vss.n955 vss.n950 2172.79
R1802 vss.n953 vss.n950 2172.79
R1803 vss.n940 vss.n932 2172.79
R1804 vss.n829 vss.n827 2172.79
R1805 vss.n849 vss.n806 2172.79
R1806 vss.n849 vss.n807 2172.79
R1807 vss.n831 vss.n827 2172.79
R1808 vss.n7442 vss.n7440 2172.79
R1809 vss.n7469 vss.n7464 2172.79
R1810 vss.n7485 vss.n7440 2172.79
R1811 vss.n15315 vss.n15309 2172.79
R1812 vss.n15332 vss.n15327 2172.79
R1813 vss.n15330 vss.n15327 2172.79
R1814 vss.n15317 vss.n15309 2172.79
R1815 vss.n681 vss.n675 2172.79
R1816 vss.n698 vss.n693 2172.79
R1817 vss.n696 vss.n693 2172.79
R1818 vss.n683 vss.n675 2172.79
R1819 vss.n7274 vss.n3124 2172.79
R1820 vss.n7289 vss.n7288 2172.79
R1821 vss.n7276 vss.n3124 2172.79
R1822 vss.n572 vss.n570 2172.79
R1823 vss.n592 vss.n548 2172.79
R1824 vss.n592 vss.n549 2172.79
R1825 vss.n574 vss.n570 2172.79
R1826 vss.n473 vss.n467 2172.79
R1827 vss.n490 vss.n485 2172.79
R1828 vss.n488 vss.n485 2172.79
R1829 vss.n475 vss.n467 2172.79
R1830 vss.n4723 vss.n4721 2172.79
R1831 vss.n4743 vss.n4555 2172.79
R1832 vss.n4743 vss.n4556 2172.79
R1833 vss.n4725 vss.n4721 2172.79
R1834 vss.n4338 vss.n4336 2172.79
R1835 vss.n4358 vss.n4315 2172.79
R1836 vss.n4358 vss.n4316 2172.79
R1837 vss.n4340 vss.n4336 2172.79
R1838 vss.n6779 vss.n6777 2172.79
R1839 vss.n6781 vss.n6777 2172.79
R1840 vss.n6765 vss.n6759 2172.79
R1841 vss.n6767 vss.n6759 2172.79
R1842 vss.n6853 vss.n6845 2172.79
R1843 vss.n6851 vss.n6845 2172.79
R1844 vss.n6865 vss.n6863 2172.79
R1845 vss.n6867 vss.n6863 2172.79
R1846 vss.n7220 vss.n3137 2172.79
R1847 vss.n6823 vss.n6807 2172.79
R1848 vss.n6823 vss.n6806 2172.79
R1849 vss.n6900 vss.n6899 2172.79
R1850 vss.n6899 vss.n6898 2172.79
R1851 vss.n6917 vss.n6827 2172.79
R1852 vss.n7103 vss.n7099 2172.79
R1853 vss.n7103 vss.n7101 2172.79
R1854 vss.n7121 vss.n7079 2172.79
R1855 vss.n7986 vss.n2458 2172.79
R1856 vss.n7969 vss.n2467 2172.79
R1857 vss.n7971 vss.n2467 2172.79
R1858 vss.n3011 vss.n3009 2172.79
R1859 vss.n7492 vss.n3009 2172.79
R1860 vss.n2999 vss.n2990 2172.79
R1861 vss.n7705 vss.n7703 2172.79
R1862 vss.n7708 vss.n7703 2172.79
R1863 vss.n7693 vss.n7684 2172.79
R1864 vss.n2925 vss.n2889 2172.79
R1865 vss.n2908 vss.n2897 2172.79
R1866 vss.n2910 vss.n2897 2172.79
R1867 vss.n7754 vss.n7752 2172.79
R1868 vss.n7756 vss.n7752 2172.79
R1869 vss.n7742 vss.n7733 2172.79
R1870 vss.n7900 vss.n7898 2172.79
R1871 vss.n7903 vss.n7898 2172.79
R1872 vss.n7888 vss.n7879 2172.79
R1873 vss.n2675 vss.n2663 2172.79
R1874 vss.n7924 vss.n2645 2172.79
R1875 vss.n7924 vss.n2644 2172.79
R1876 vss.n1157 vss.n1155 2172.79
R1877 vss.n14873 vss.n1155 2172.79
R1878 vss.n7943 vss.n7928 2172.79
R1879 vss.n2620 vss.n2617 2172.79
R1880 vss.n2622 vss.n2617 2172.79
R1881 vss.n2641 vss.n2599 2172.79
R1882 vss.n2641 vss.n2600 2172.79
R1883 vss.n1943 vss.n1898 2172.79
R1884 vss.n1943 vss.n1899 2172.79
R1885 vss.n1923 vss.n1920 2172.79
R1886 vss.n1925 vss.n1920 2172.79
R1887 vss.n2860 vss.n2852 2172.79
R1888 vss.n2858 vss.n2852 2172.79
R1889 vss.n2872 vss.n2870 2172.79
R1890 vss.n2874 vss.n2870 2172.79
R1891 vss.n3033 vss.n3031 2172.79
R1892 vss.n3035 vss.n3031 2172.79
R1893 vss.n3057 vss.n3013 2172.79
R1894 vss.n3057 vss.n3014 2172.79
R1895 vss.n7644 vss.n7636 2172.79
R1896 vss.n7642 vss.n7636 2172.79
R1897 vss.n7656 vss.n7654 2172.79
R1898 vss.n7658 vss.n7654 2172.79
R1899 vss.n2814 vss.n2738 2172.79
R1900 vss.n2812 vss.n2738 2172.79
R1901 vss.n2826 vss.n2824 2172.79
R1902 vss.n2828 vss.n2824 2172.79
R1903 vss.n2952 vss.n2944 2172.79
R1904 vss.n2950 vss.n2944 2172.79
R1905 vss.n2965 vss.n2962 2172.79
R1906 vss.n2967 vss.n2962 2172.79
R1907 vss.n7075 vss.n7033 2172.79
R1908 vss.n7075 vss.n7034 2172.79
R1909 vss.n7049 vss.n3131 2172.79
R1910 vss.n7058 vss.n3131 2172.79
R1911 vss.n7009 vss.n7006 2172.79
R1912 vss.n7011 vss.n7006 2172.79
R1913 vss.n7030 vss.n6988 2172.79
R1914 vss.n7030 vss.n6989 2172.79
R1915 vss.n7148 vss.n7146 2172.79
R1916 vss.n7150 vss.n7146 2172.79
R1917 vss.n7168 vss.n7125 2172.79
R1918 vss.n7168 vss.n7126 2172.79
R1919 vss.n6964 vss.n6942 2172.79
R1920 vss.n6966 vss.n6942 2172.79
R1921 vss.n6985 vss.n6921 2172.79
R1922 vss.n6985 vss.n6922 2172.79
R1923 vss.n7596 vss.n7520 2172.79
R1924 vss.n7594 vss.n7520 2172.79
R1925 vss.n7608 vss.n7606 2172.79
R1926 vss.n7610 vss.n7606 2172.79
R1927 vss.n7791 vss.n7783 2172.79
R1928 vss.n7789 vss.n7783 2172.79
R1929 vss.n7803 vss.n7801 2172.79
R1930 vss.n7805 vss.n7801 2172.79
R1931 vss.n7839 vss.n7831 2172.79
R1932 vss.n7837 vss.n7831 2172.79
R1933 vss.n7851 vss.n7849 2172.79
R1934 vss.n7853 vss.n7849 2172.79
R1935 vss.n2701 vss.n2693 2172.79
R1936 vss.n2699 vss.n2693 2172.79
R1937 vss.n2710 vss.n987 2172.79
R1938 vss.n2714 vss.n987 2172.79
R1939 vss.n2576 vss.n2505 2172.79
R1940 vss.n2578 vss.n2505 2172.79
R1941 vss.n2596 vss.n2484 2172.79
R1942 vss.n2596 vss.n2485 2172.79
R1943 vss.n7183 vss.n3164 2172.79
R1944 vss.n7181 vss.n3164 2172.79
R1945 vss.n7195 vss.n7193 2172.79
R1946 vss.n7197 vss.n7193 2172.79
R1947 vss.n3208 vss.n3192 2172.79
R1948 vss.n3208 vss.n3193 2172.79
R1949 vss.n6802 vss.n3170 2172.79
R1950 vss.n6802 vss.n3171 2172.79
R1951 vss.n14296 vss.n14291 2172.79
R1952 vss.n14319 vss.n14291 2172.79
R1953 vss.n14311 vss.n14302 2172.79
R1954 vss.n14302 vss.n14290 2172.79
R1955 vss.n14825 vss.n14823 2172.79
R1956 vss.n14827 vss.n14823 2172.79
R1957 vss.n14845 vss.n1163 2172.79
R1958 vss.n14845 vss.n1164 2172.79
R1959 vss.n14173 vss.n14157 2172.79
R1960 vss.n14173 vss.n14158 2172.79
R1961 vss.n14795 vss.n1182 2172.79
R1962 vss.n14793 vss.n1182 2172.79
R1963 vss.n14263 vss.n14251 2172.79
R1964 vss.n14263 vss.n14262 2172.79
R1965 vss.n14272 vss.n14246 2172.79
R1966 vss.n14276 vss.n14246 2172.79
R1967 vss.n1840 vss.n1834 2172.79
R1968 vss.n14345 vss.n1852 2172.79
R1969 vss.n14343 vss.n1852 2172.79
R1970 vss.n1842 vss.n1834 2172.79
R1971 vss.n14451 vss.n1759 2172.79
R1972 vss.n14453 vss.n1759 2172.79
R1973 vss.n14465 vss.n14463 2172.79
R1974 vss.n14217 vss.n14207 2172.79
R1975 vss.n14231 vss.n14227 2172.79
R1976 vss.n14229 vss.n14227 2172.79
R1977 vss.n2298 vss.n2291 2172.79
R1978 vss.n2300 vss.n2291 2172.79
R1979 vss.n2312 vss.n2310 2172.79
R1980 vss.n2254 vss.n2245 2172.79
R1981 vss.n2268 vss.n2264 2172.79
R1982 vss.n2266 vss.n2264 2172.79
R1983 vss.n8092 vss.n2227 2172.79
R1984 vss.n8092 vss.n2228 2172.79
R1985 vss.n8074 vss.n8069 2172.79
R1986 vss.n8110 vss.n8097 2172.79
R1987 vss.n8124 vss.n8122 2172.79
R1988 vss.n8126 vss.n8122 2172.79
R1989 vss.n8142 vss.n8097 2172.79
R1990 vss.n1302 vss.n1296 2172.79
R1991 vss.n14739 vss.n1314 2172.79
R1992 vss.n14737 vss.n1314 2172.79
R1993 vss.n1304 vss.n1296 2172.79
R1994 vss.n14001 vss.n13995 2172.79
R1995 vss.n14017 vss.n14013 2172.79
R1996 vss.n14015 vss.n14013 2172.79
R1997 vss.n14003 vss.n13995 2172.79
R1998 vss.n13957 vss.n8166 2172.79
R1999 vss.n13971 vss.n13967 2172.79
R2000 vss.n13969 vss.n13967 2172.79
R2001 vss.n8220 vss.n8176 2172.79
R2002 vss.n8220 vss.n8177 2172.79
R2003 vss.n8202 vss.n8197 2172.79
R2004 vss.n13871 vss.n13859 2172.79
R2005 vss.n13885 vss.n13883 2172.79
R2006 vss.n13887 vss.n13883 2172.79
R2007 vss.n13903 vss.n13859 2172.79
R2008 vss.n1507 vss.n1501 2172.79
R2009 vss.n14666 vss.n1519 2172.79
R2010 vss.n14664 vss.n1519 2172.79
R2011 vss.n1509 vss.n1501 2172.79
R2012 vss.n1560 vss.n1554 2172.79
R2013 vss.n14589 vss.n1572 2172.79
R2014 vss.n14587 vss.n1572 2172.79
R2015 vss.n1562 vss.n1554 2172.79
R2016 vss.n14445 vss.n14401 2172.79
R2017 vss.n14427 vss.n14425 2172.79
R2018 vss.n14429 vss.n14425 2172.79
R2019 vss.n14500 vss.n14494 2172.79
R2020 vss.n14516 vss.n14512 2172.79
R2021 vss.n14514 vss.n14512 2172.79
R2022 vss.n14502 vss.n14494 2172.79
R2023 vss.n1717 vss.n1711 2172.79
R2024 vss.n1734 vss.n1729 2172.79
R2025 vss.n1732 vss.n1729 2172.79
R2026 vss.n1719 vss.n1711 2172.79
R2027 vss.n1608 vss.n1606 2172.79
R2028 vss.n1628 vss.n1585 2172.79
R2029 vss.n1628 vss.n1586 2172.79
R2030 vss.n1610 vss.n1606 2172.79
R2031 vss.n13907 vss.n13905 2172.79
R2032 vss.n13934 vss.n13929 2172.79
R2033 vss.n13950 vss.n13905 2172.79
R2034 vss.n14620 vss.n14614 2172.79
R2035 vss.n14637 vss.n14632 2172.79
R2036 vss.n14635 vss.n14632 2172.79
R2037 vss.n14622 vss.n14614 2172.79
R2038 vss.n1460 vss.n1454 2172.79
R2039 vss.n1477 vss.n1472 2172.79
R2040 vss.n1475 vss.n1472 2172.79
R2041 vss.n1462 vss.n1454 2172.79
R2042 vss.n8146 vss.n8144 2172.79
R2043 vss.n14051 vss.n14046 2172.79
R2044 vss.n14067 vss.n8144 2172.79
R2045 vss.n1351 vss.n1349 2172.79
R2046 vss.n1371 vss.n1327 2172.79
R2047 vss.n1371 vss.n1328 2172.79
R2048 vss.n1353 vss.n1349 2172.79
R2049 vss.n1252 vss.n1246 2172.79
R2050 vss.n1269 vss.n1264 2172.79
R2051 vss.n1267 vss.n1264 2172.79
R2052 vss.n1254 vss.n1246 2172.79
R2053 vss.n2345 vss.n2339 2172.79
R2054 vss.n8038 vss.n2357 2172.79
R2055 vss.n8036 vss.n2357 2172.79
R2056 vss.n2347 vss.n2339 2172.79
R2057 vss.n2393 vss.n2391 2172.79
R2058 vss.n2413 vss.n2370 2172.79
R2059 vss.n2413 vss.n2371 2172.79
R2060 vss.n2395 vss.n2391 2172.79
R2061 vss.n2051 vss.n2049 2172.79
R2062 vss.n14181 vss.n2049 2172.79
R2063 vss.n11864 vss.n11849 2172.79
R2064 vss.n11864 vss.n11848 2172.79
R2065 vss.n11961 vss.n11945 2172.79
R2066 vss.n11961 vss.n11946 2172.79
R2067 vss.n14127 vss.n2101 2172.79
R2068 vss.n14129 vss.n2101 2172.79
R2069 vss.n13489 vss.n13481 2172.79
R2070 vss.n13487 vss.n13481 2172.79
R2071 vss.n13501 vss.n13499 2172.79
R2072 vss.n13503 vss.n13499 2172.79
R2073 vss.n12059 vss.n12016 2172.79
R2074 vss.n12059 vss.n12017 2172.79
R2075 vss.n12040 vss.n12038 2172.79
R2076 vss.n12042 vss.n12038 2172.79
R2077 vss.n13721 vss.n8316 2172.79
R2078 vss.n13719 vss.n8316 2172.79
R2079 vss.n13733 vss.n13731 2172.79
R2080 vss.n13735 vss.n13731 2172.79
R2081 vss.n8485 vss.n8442 2172.79
R2082 vss.n8485 vss.n8443 2172.79
R2083 vss.n8466 vss.n8464 2172.79
R2084 vss.n8468 vss.n8464 2172.79
R2085 vss.n8562 vss.n8519 2172.79
R2086 vss.n8562 vss.n8520 2172.79
R2087 vss.n8543 vss.n8541 2172.79
R2088 vss.n8545 vss.n8541 2172.79
R2089 vss.n13009 vss.n9102 2172.79
R2090 vss.n13007 vss.n9102 2172.79
R2091 vss.n13021 vss.n13019 2172.79
R2092 vss.n13023 vss.n13019 2172.79
R2093 vss.n8974 vss.n8966 2172.79
R2094 vss.n8972 vss.n8966 2172.79
R2095 vss.n8986 vss.n8984 2172.79
R2096 vss.n8988 vss.n8984 2172.79
R2097 vss.n9157 vss.n9114 2172.79
R2098 vss.n9157 vss.n9115 2172.79
R2099 vss.n9138 vss.n9136 2172.79
R2100 vss.n9140 vss.n9136 2172.79
R2101 vss.n12637 vss.n12545 2172.79
R2102 vss.n12637 vss.n12546 2172.79
R2103 vss.n12569 vss.n12567 2172.79
R2104 vss.n12571 vss.n12567 2172.79
R2105 vss.n14076 vss.n14075 2172.79
R2106 vss.n2166 vss.n2160 2172.79
R2107 vss.n2168 vss.n2160 2172.79
R2108 vss.n12614 vss.n12612 2172.79
R2109 vss.n12616 vss.n12612 2172.79
R2110 vss.n12602 vss.n12593 2172.79
R2111 vss.n9019 vss.n9011 2172.79
R2112 vss.n9017 vss.n9011 2172.79
R2113 vss.n9028 vss.n8096 2172.79
R2114 vss.n9032 vss.n8096 2172.79
R2115 vss.n13117 vss.n13115 2172.79
R2116 vss.n13120 vss.n13115 2172.79
R2117 vss.n13105 vss.n13096 2172.79
R2118 vss.n13070 vss.n13069 2172.79
R2119 vss.n13054 vss.n13048 2172.79
R2120 vss.n13056 vss.n13048 2172.79
R2121 vss.n9076 vss.n9074 2172.79
R2122 vss.n9078 vss.n9074 2172.79
R2123 vss.n9064 vss.n9055 2172.79
R2124 vss.n8244 vss.n8242 2172.79
R2125 vss.n8246 vss.n8242 2172.79
R2126 vss.n13858 vss.n8224 2172.79
R2127 vss.n13858 vss.n8225 2172.79
R2128 vss.n13829 vss.n13827 2172.79
R2129 vss.n13832 vss.n13827 2172.79
R2130 vss.n13817 vss.n13808 2172.79
R2131 vss.n13782 vss.n13781 2172.79
R2132 vss.n13766 vss.n13760 2172.79
R2133 vss.n13768 vss.n13760 2172.79
R2134 vss.n8290 vss.n8288 2172.79
R2135 vss.n8292 vss.n8288 2172.79
R2136 vss.n8278 vss.n8269 2172.79
R2137 vss.n13534 vss.n13526 2172.79
R2138 vss.n13532 vss.n13526 2172.79
R2139 vss.n13543 vss.n1766 2172.79
R2140 vss.n13547 vss.n1766 2172.79
R2141 vss.n13640 vss.n13638 2172.79
R2142 vss.n13643 vss.n13638 2172.79
R2143 vss.n13628 vss.n13619 2172.79
R2144 vss.n13593 vss.n13592 2172.79
R2145 vss.n13577 vss.n13570 2172.79
R2146 vss.n13579 vss.n13570 2172.79
R2147 vss.n14154 vss.n2055 2172.79
R2148 vss.n14154 vss.n2056 2172.79
R2149 vss.n2076 vss.n2073 2172.79
R2150 vss.n2202 vss.n2199 2172.79
R2151 vss.n2204 vss.n2199 2172.79
R2152 vss.n2223 vss.n2181 2172.79
R2153 vss.n2223 vss.n2182 2172.79
R2154 vss.n9300 vss.n9284 2172.79
R2155 vss.n9300 vss.n9285 2172.79
R2156 vss.n14102 vss.n2129 2172.79
R2157 vss.n14102 vss.n2130 2172.79
R2158 vss.n12846 vss.n9406 2172.79
R2159 vss.n12844 vss.n9406 2172.79
R2160 vss.n12858 vss.n12856 2172.79
R2161 vss.n12860 vss.n12856 2172.79
R2162 vss.n12773 vss.n12729 2172.79
R2163 vss.n12773 vss.n12730 2172.79
R2164 vss.n12753 vss.n12751 2172.79
R2165 vss.n12755 vss.n12751 2172.79
R2166 vss.n13323 vss.n8424 2172.79
R2167 vss.n13321 vss.n8424 2172.79
R2168 vss.n13335 vss.n13333 2172.79
R2169 vss.n13337 vss.n13333 2172.79
R2170 vss.n13442 vss.n13366 2172.79
R2171 vss.n13440 vss.n13366 2172.79
R2172 vss.n13454 vss.n13452 2172.79
R2173 vss.n13456 vss.n13452 2172.79
R2174 vss.n1780 vss.n1768 2172.79
R2175 vss.n1812 vss.n1768 2172.79
R2176 vss.n1794 vss.n1792 2172.79
R2177 vss.n1796 vss.n1792 2172.79
R2178 vss.n1816 vss.n1814 2172.79
R2179 vss.n14379 vss.n14374 2172.79
R2180 vss.n14395 vss.n1814 2172.79
R2181 vss.n2007 vss.n2001 2172.79
R2182 vss.n2024 vss.n2019 2172.79
R2183 vss.n2022 vss.n2019 2172.79
R2184 vss.n2009 vss.n2001 2172.79
R2185 vss.n1001 vss.n989 2172.79
R2186 vss.n1033 vss.n989 2172.79
R2187 vss.n1015 vss.n1013 2172.79
R2188 vss.n1017 vss.n1013 2172.79
R2189 vss.n1037 vss.n1035 2172.79
R2190 vss.n15074 vss.n15069 2172.79
R2191 vss.n15090 vss.n1035 2172.79
R2192 vss.n1112 vss.n1106 2172.79
R2193 vss.n1129 vss.n1124 2172.79
R2194 vss.n1127 vss.n1124 2172.79
R2195 vss.n1114 vss.n1106 2172.79
R2196 vss.n6206 vss.n6204 2172.79
R2197 vss.n6233 vss.n6228 2172.79
R2198 vss.n6249 vss.n6204 2172.79
R2199 vss.n3950 vss.n3948 2172.79
R2200 vss.n15860 vss.n43 2172.79
R2201 vss.n15858 vss.n43 2172.79
R2202 vss.n3964 vss.n3948 2172.79
R2203 vss.n3852 vss.n3850 2172.79
R2204 vss.n3877 vss.n3874 2172.79
R2205 vss.n3879 vss.n3874 2172.79
R2206 vss.n3895 vss.n3850 2172.79
R2207 vss.n3733 vss.n3731 2172.79
R2208 vss.n3758 vss.n3755 2172.79
R2209 vss.n3760 vss.n3755 2172.79
R2210 vss.n3776 vss.n3731 2172.79
R2211 vss.n3614 vss.n3612 2172.79
R2212 vss.n3639 vss.n3636 2172.79
R2213 vss.n3641 vss.n3636 2172.79
R2214 vss.n3657 vss.n3612 2172.79
R2215 vss.n15601 vss.n15589 2172.79
R2216 vss.n15601 vss.n15600 2172.79
R2217 vss.n15610 vss.n15584 2172.79
R2218 vss.n15614 vss.n15584 2172.79
R2219 vss.n306 vss.n304 2172.79
R2220 vss.n330 vss.n327 2172.79
R2221 vss.n332 vss.n327 2172.79
R2222 vss.n348 vss.n304 2172.79
R2223 vss.n15550 vss.n374 2172.79
R2224 vss.n15566 vss.n15562 2172.79
R2225 vss.n15564 vss.n15562 2172.79
R2226 vss.n15552 vss.n374 2172.79
R2227 vss.n10446 vss.n10438 2172.79
R2228 vss.n10444 vss.n10438 2172.79
R2229 vss.n10459 vss.n10456 2172.79
R2230 vss.n10461 vss.n10456 2172.79
R2231 vss.n10592 vss.n10583 2172.79
R2232 vss.n10590 vss.n10583 2172.79
R2233 vss.n10604 vss.n10602 2172.79
R2234 vss.n10606 vss.n10602 2172.79
R2235 vss.n10986 vss.n10977 2172.79
R2236 vss.n10984 vss.n10977 2172.79
R2237 vss.n10998 vss.n10996 2172.79
R2238 vss.n11000 vss.n10996 2172.79
R2239 vss.n10037 vss.n9993 2172.79
R2240 vss.n10037 vss.n9994 2172.79
R2241 vss.n10017 vss.n10015 2172.79
R2242 vss.n10019 vss.n10015 2172.79
R2243 vss.n11730 vss.n11726 1997.67
R2244 vss.n14847 vss.n1161 1987.64
R2245 vss.n13223 vss.n8835 1911.25
R2246 vss.n12184 vss.n12183 1821.33
R2247 vss.n14320 vss.n1159 1821.33
R2248 vss.n15015 vss.n380 1821.33
R2249 vss.n11730 vss.n11729 1554.74
R2250 vss.n15542 vss.n382 1414.97
R2251 vss.n12181 vss.n12180 1414.97
R2252 vss.n1958 vss.n1159 1409
R2253 vss.n6571 vss.n380 1409
R2254 vss.n12183 vss.n12131 1409
R2255 vss.n11731 vss.n11730 1364
R2256 vss.n10540 vss.n10539 1245.55
R2257 vss.n10838 vss.n10837 1245.55
R2258 vss.n10934 vss.n10933 1245.55
R2259 vss.n11273 vss.n11272 1245.55
R2260 vss.n11131 vss.n11130 1245.55
R2261 vss.n11584 vss.n11583 1245.55
R2262 vss.n9903 vss.n9902 1245.55
R2263 vss.n9461 vss.n9460 1245.55
R2264 vss.n9494 vss.n9493 1245.55
R2265 vss.n9522 vss.n9520 1245.55
R2266 vss.n9623 vss.n9622 1245.55
R2267 vss.n9652 vss.n9649 1245.55
R2268 vss.n9753 vss.n9752 1245.55
R2269 vss.n9781 vss.n9779 1245.55
R2270 vss.n12215 vss.n12214 1245.55
R2271 vss.n12333 vss.n12332 1245.55
R2272 vss.n12452 vss.n12451 1245.55
R2273 vss.n3589 vss.n3588 1245.55
R2274 vss.n6053 vss.n6052 1245.55
R2275 vss.n6179 vss.n6178 1245.55
R2276 vss.n5746 vss.n5745 1245.55
R2277 vss.n5813 vss.n5812 1245.55
R2278 vss.n5940 vss.n5939 1245.55
R2279 vss.n5558 vss.n5557 1245.55
R2280 vss.n5702 vss.n5701 1245.55
R2281 vss.n3563 vss.n3562 1245.55
R2282 vss.n5986 vss.n5985 1245.55
R2283 vss.n6231 vss.n6230 1245.55
R2284 vss.n4515 vss.n4514 1245.55
R2285 vss.n5020 vss.n5019 1245.55
R2286 vss.n5068 vss.n5067 1245.55
R2287 vss.n5494 vss.n5493 1245.55
R2288 vss.n5279 vss.n5278 1245.55
R2289 vss.n3465 vss.n3464 1245.55
R2290 vss.n6669 vss.n3336 1245.55
R2291 vss.n6367 vss.n6366 1245.55
R2292 vss.n5529 vss.n5528 1245.55
R2293 vss.n4212 vss.n4179 1245.55
R2294 vss.n4484 vss.n4483 1245.55
R2295 vss.n15163 vss.n15162 1245.55
R2296 vss.n14909 vss.n14908 1245.55
R2297 vss.n15072 vss.n15071 1245.55
R2298 vss.n4597 vss.n4596 1245.55
R2299 vss.n4672 vss.n4671 1245.55
R2300 vss.n4644 vss.n4643 1245.55
R2301 vss.n3081 vss.n3080 1245.55
R2302 vss.n7372 vss.n7370 1245.55
R2303 vss.n15108 vss.n15107 1245.55
R2304 vss.n7467 vss.n7466 1245.55
R2305 vss.n7291 vss.n7290 1245.55
R2306 vss.n6885 vss.n6826 1245.55
R2307 vss.n7088 vss.n7078 1245.55
R2308 vss.n2997 vss.n2996 1245.55
R2309 vss.n7691 vss.n7690 1245.55
R2310 vss.n7740 vss.n7739 1245.55
R2311 vss.n7886 vss.n7885 1245.55
R2312 vss.n7933 vss.n7927 1245.55
R2313 vss.n2672 vss.n2671 1245.55
R2314 vss.n2922 vss.n2921 1245.55
R2315 vss.n7983 vss.n7982 1245.55
R2316 vss.n7216 vss.n7215 1245.55
R2317 vss.n14468 vss.n14467 1245.55
R2318 vss.n14214 vss.n14213 1245.55
R2319 vss.n14377 vss.n14376 1245.55
R2320 vss.n2315 vss.n2314 1245.55
R2321 vss.n2248 vss.n2247 1245.55
R2322 vss.n8073 vss.n8071 1245.55
R2323 vss.n8173 vss.n8172 1245.55
R2324 vss.n8201 vss.n8199 1245.55
R2325 vss.n14413 vss.n14412 1245.55
R2326 vss.n13932 vss.n13931 1245.55
R2327 vss.n14049 vss.n14048 1245.55
R2328 vss.n12600 vss.n12599 1245.55
R2329 vss.n13103 vss.n13102 1245.55
R2330 vss.n9062 vss.n9061 1245.55
R2331 vss.n13815 vss.n13814 1245.55
R2332 vss.n8276 vss.n8275 1245.55
R2333 vss.n13626 vss.n13625 1245.55
R2334 vss.n2079 vss.n2078 1245.55
R2335 vss.n13595 vss.n13594 1245.55
R2336 vss.n13784 vss.n13783 1245.55
R2337 vss.n13072 vss.n13071 1245.55
R2338 vss.n14078 vss.n14077 1245.55
R2339 vss.n11553 vss.n11552 1245.55
R2340 vss.n11242 vss.n11241 1245.55
R2341 vss.n10903 vss.n10902 1245.55
R2342 vss.n10509 vss.n10508 1245.55
R2343 vss.n12475 vss.n12474 1131.75
R2344 vss.n12473 vss.n9548 1131.75
R2345 vss.n12356 vss.n12355 1131.75
R2346 vss.n12354 vss.n9677 1131.75
R2347 vss.n12238 vss.n12237 1131.75
R2348 vss.n12236 vss.n9806 1131.75
R2349 vss.n14072 vss.n14071 1131.75
R2350 vss.n14070 vss.n8098 1131.75
R2351 vss.n13955 vss.n13954 1131.75
R2352 vss.n13953 vss.n1763 1131.75
R2353 vss.n14447 vss.n14399 1131.75
R2354 vss.n14398 vss.n1767 1131.75
R2355 vss.n7224 vss.n7223 1131.75
R2356 vss.n7270 vss.n2459 1131.75
R2357 vss.n7489 vss.n7393 1131.75
R2358 vss.n7488 vss.n984 1131.75
R2359 vss.n15142 vss.n15094 1131.75
R2360 vss.n15093 vss.n988 1131.75
R2361 vss.n6202 vss.n6201 1131.75
R2362 vss.n6200 vss.n5964 1131.75
R2363 vss.n5963 vss.n5962 1131.75
R2364 vss.n5961 vss.n5724 1131.75
R2365 vss.n5723 vss.n3534 1131.75
R2366 vss.n6334 vss.n6333 1131.75
R2367 vss.n10349 vss.n10345 1118.26
R2368 vss.n10355 vss.n10349 1118.26
R2369 vss.n10355 vss.n8872 1118.26
R2370 vss.n13193 vss.n8872 1118.26
R2371 vss.n13193 vss.n8873 1118.26
R2372 vss.n8873 vss.n8868 1118.26
R2373 vss.n10352 vss.n10344 1118.26
R2374 vss.n10353 vss.n10352 1118.26
R2375 vss.n10353 vss.n8875 1118.26
R2376 vss.n13188 vss.n8875 1118.26
R2377 vss.n13189 vss.n13188 1118.26
R2378 vss.n13189 vss.n8867 1118.26
R2379 vss.n10287 vss.n10283 1118.26
R2380 vss.n10320 vss.n10287 1118.26
R2381 vss.n10320 vss.n10288 1118.26
R2382 vss.n10304 vss.n10288 1118.26
R2383 vss.n10304 vss.n10302 1118.26
R2384 vss.n10309 vss.n10302 1118.26
R2385 vss.n10291 vss.n10282 1118.26
R2386 vss.n10292 vss.n10291 1118.26
R2387 vss.n10294 vss.n10292 1118.26
R2388 vss.n10313 vss.n10294 1118.26
R2389 vss.n10313 vss.n10312 1118.26
R2390 vss.n10312 vss.n10311 1118.26
R2391 vss.n9954 vss.n9950 1118.26
R2392 vss.n11642 vss.n9954 1118.26
R2393 vss.n11642 vss.n9955 1118.26
R2394 vss.n11626 vss.n9955 1118.26
R2395 vss.n11626 vss.n11624 1118.26
R2396 vss.n11631 vss.n11624 1118.26
R2397 vss.n9958 vss.n9949 1118.26
R2398 vss.n9959 vss.n9958 1118.26
R2399 vss.n9961 vss.n9959 1118.26
R2400 vss.n11635 vss.n9961 1118.26
R2401 vss.n11635 vss.n11634 1118.26
R2402 vss.n11634 vss.n11633 1118.26
R2403 vss.n11686 vss.n11685 1118.26
R2404 vss.n11687 vss.n11686 1118.26
R2405 vss.n11687 vss.n9914 1118.26
R2406 vss.n11705 vss.n9914 1118.26
R2407 vss.n11705 vss.n9915 1118.26
R2408 vss.n11697 vss.n9915 1118.26
R2409 vss.n11683 vss.n9922 1118.26
R2410 vss.n11689 vss.n9922 1118.26
R2411 vss.n11689 vss.n9919 1118.26
R2412 vss.n11703 vss.n9919 1118.26
R2413 vss.n11703 vss.n9920 1118.26
R2414 vss.n11699 vss.n9920 1118.26
R2415 vss.n11449 vss.n11448 1118.26
R2416 vss.n11450 vss.n11449 1118.26
R2417 vss.n11450 vss.n9969 1118.26
R2418 vss.n11468 vss.n9969 1118.26
R2419 vss.n11468 vss.n9970 1118.26
R2420 vss.n11460 vss.n9970 1118.26
R2421 vss.n11446 vss.n9977 1118.26
R2422 vss.n11452 vss.n9977 1118.26
R2423 vss.n11452 vss.n9974 1118.26
R2424 vss.n11466 vss.n9974 1118.26
R2425 vss.n11466 vss.n9975 1118.26
R2426 vss.n11462 vss.n9975 1118.26
R2427 vss.n11377 vss.n11367 1118.26
R2428 vss.n11403 vss.n11377 1118.26
R2429 vss.n11403 vss.n11378 1118.26
R2430 vss.n11399 vss.n11378 1118.26
R2431 vss.n11399 vss.n11383 1118.26
R2432 vss.n11391 vss.n11383 1118.26
R2433 vss.n11372 vss.n11368 1118.26
R2434 vss.n11405 vss.n11372 1118.26
R2435 vss.n11405 vss.n11373 1118.26
R2436 vss.n11397 vss.n11373 1118.26
R2437 vss.n11397 vss.n11385 1118.26
R2438 vss.n11393 vss.n11385 1118.26
R2439 vss.n11180 vss.n11179 1118.26
R2440 vss.n11181 vss.n11180 1118.26
R2441 vss.n11181 vss.n11160 1118.26
R2442 vss.n11199 vss.n11160 1118.26
R2443 vss.n11199 vss.n11161 1118.26
R2444 vss.n11191 vss.n11161 1118.26
R2445 vss.n11177 vss.n11168 1118.26
R2446 vss.n11183 vss.n11168 1118.26
R2447 vss.n11183 vss.n11165 1118.26
R2448 vss.n11197 vss.n11165 1118.26
R2449 vss.n11197 vss.n11166 1118.26
R2450 vss.n11193 vss.n11166 1118.26
R2451 vss.n11044 vss.n11043 1118.26
R2452 vss.n11045 vss.n11044 1118.26
R2453 vss.n11045 vss.n10129 1118.26
R2454 vss.n11063 vss.n10129 1118.26
R2455 vss.n11063 vss.n10130 1118.26
R2456 vss.n11055 vss.n10130 1118.26
R2457 vss.n11041 vss.n10137 1118.26
R2458 vss.n11047 vss.n10137 1118.26
R2459 vss.n11047 vss.n10134 1118.26
R2460 vss.n11061 vss.n10134 1118.26
R2461 vss.n11061 vss.n10135 1118.26
R2462 vss.n11057 vss.n10135 1118.26
R2463 vss.n10104 vss.n10103 1118.26
R2464 vss.n10105 vss.n10104 1118.26
R2465 vss.n10105 vss.n10083 1118.26
R2466 vss.n10123 vss.n10083 1118.26
R2467 vss.n10123 vss.n10084 1118.26
R2468 vss.n10115 vss.n10084 1118.26
R2469 vss.n10101 vss.n10091 1118.26
R2470 vss.n10107 vss.n10091 1118.26
R2471 vss.n10107 vss.n10088 1118.26
R2472 vss.n10121 vss.n10088 1118.26
R2473 vss.n10121 vss.n10089 1118.26
R2474 vss.n10117 vss.n10089 1118.26
R2475 vss.n10721 vss.n10711 1118.26
R2476 vss.n10746 vss.n10721 1118.26
R2477 vss.n10746 vss.n10743 1118.26
R2478 vss.n10743 vss.n10742 1118.26
R2479 vss.n10742 vss.n10724 1118.26
R2480 vss.n10734 vss.n10724 1118.26
R2481 vss.n10716 vss.n10712 1118.26
R2482 vss.n10748 vss.n10716 1118.26
R2483 vss.n10748 vss.n10717 1118.26
R2484 vss.n10740 vss.n10717 1118.26
R2485 vss.n10740 vss.n10727 1118.26
R2486 vss.n10736 vss.n10727 1118.26
R2487 vss.n10792 vss.n10791 1118.26
R2488 vss.n10793 vss.n10792 1118.26
R2489 vss.n10793 vss.n10216 1118.26
R2490 vss.n10811 vss.n10216 1118.26
R2491 vss.n10811 vss.n10217 1118.26
R2492 vss.n10803 vss.n10217 1118.26
R2493 vss.n10789 vss.n10224 1118.26
R2494 vss.n10795 vss.n10224 1118.26
R2495 vss.n10795 vss.n10221 1118.26
R2496 vss.n10809 vss.n10221 1118.26
R2497 vss.n10809 vss.n10222 1118.26
R2498 vss.n10805 vss.n10222 1118.26
R2499 vss.n10665 vss.n10655 1118.26
R2500 vss.n10691 vss.n10665 1118.26
R2501 vss.n10691 vss.n10666 1118.26
R2502 vss.n10687 vss.n10666 1118.26
R2503 vss.n10687 vss.n10671 1118.26
R2504 vss.n10679 vss.n10671 1118.26
R2505 vss.n10660 vss.n10656 1118.26
R2506 vss.n10693 vss.n10660 1118.26
R2507 vss.n10693 vss.n10661 1118.26
R2508 vss.n10685 vss.n10661 1118.26
R2509 vss.n10685 vss.n10673 1118.26
R2510 vss.n10681 vss.n10673 1118.26
R2511 vss.n10402 vss.n10401 1118.26
R2512 vss.n10403 vss.n10402 1118.26
R2513 vss.n10403 vss.n10258 1118.26
R2514 vss.n10421 vss.n10258 1118.26
R2515 vss.n10421 vss.n10259 1118.26
R2516 vss.n10413 vss.n10259 1118.26
R2517 vss.n10399 vss.n10266 1118.26
R2518 vss.n10405 vss.n10266 1118.26
R2519 vss.n10405 vss.n10263 1118.26
R2520 vss.n10419 vss.n10263 1118.26
R2521 vss.n10419 vss.n10264 1118.26
R2522 vss.n10415 vss.n10264 1118.26
R2523 vss.n10491 vss.n10482 1118.26
R2524 vss.n10497 vss.n10482 1118.26
R2525 vss.n10497 vss.n10479 1118.26
R2526 vss.n10513 vss.n10479 1118.26
R2527 vss.n10513 vss.n10480 1118.26
R2528 vss.n10509 vss.n10480 1118.26
R2529 vss.n10494 vss.n10493 1118.26
R2530 vss.n10495 vss.n10494 1118.26
R2531 vss.n10495 vss.n10474 1118.26
R2532 vss.n10515 vss.n10474 1118.26
R2533 vss.n10515 vss.n10475 1118.26
R2534 vss.n10506 vss.n10475 1118.26
R2535 vss.n10539 vss.n10530 1118.26
R2536 vss.n10546 vss.n10530 1118.26
R2537 vss.n10546 vss.n10527 1118.26
R2538 vss.n10560 vss.n10527 1118.26
R2539 vss.n10560 vss.n10528 1118.26
R2540 vss.n10556 vss.n10528 1118.26
R2541 vss.n10543 vss.n10542 1118.26
R2542 vss.n10544 vss.n10543 1118.26
R2543 vss.n10544 vss.n10522 1118.26
R2544 vss.n10562 vss.n10522 1118.26
R2545 vss.n10562 vss.n10523 1118.26
R2546 vss.n10554 vss.n10523 1118.26
R2547 vss.n10837 vss.n10828 1118.26
R2548 vss.n10844 vss.n10828 1118.26
R2549 vss.n10844 vss.n10825 1118.26
R2550 vss.n10859 vss.n10825 1118.26
R2551 vss.n10859 vss.n10826 1118.26
R2552 vss.n10855 vss.n10826 1118.26
R2553 vss.n10841 vss.n10840 1118.26
R2554 vss.n10842 vss.n10841 1118.26
R2555 vss.n10842 vss.n10820 1118.26
R2556 vss.n10861 vss.n10820 1118.26
R2557 vss.n10861 vss.n10821 1118.26
R2558 vss.n10852 vss.n10821 1118.26
R2559 vss.n10885 vss.n10876 1118.26
R2560 vss.n10891 vss.n10876 1118.26
R2561 vss.n10891 vss.n10873 1118.26
R2562 vss.n10907 vss.n10873 1118.26
R2563 vss.n10907 vss.n10874 1118.26
R2564 vss.n10903 vss.n10874 1118.26
R2565 vss.n10888 vss.n10887 1118.26
R2566 vss.n10889 vss.n10888 1118.26
R2567 vss.n10889 vss.n10868 1118.26
R2568 vss.n10909 vss.n10868 1118.26
R2569 vss.n10909 vss.n10869 1118.26
R2570 vss.n10900 vss.n10869 1118.26
R2571 vss.n10933 vss.n10924 1118.26
R2572 vss.n10940 vss.n10924 1118.26
R2573 vss.n10940 vss.n10921 1118.26
R2574 vss.n10954 vss.n10921 1118.26
R2575 vss.n10954 vss.n10922 1118.26
R2576 vss.n10950 vss.n10922 1118.26
R2577 vss.n10937 vss.n10936 1118.26
R2578 vss.n10938 vss.n10937 1118.26
R2579 vss.n10938 vss.n10916 1118.26
R2580 vss.n10956 vss.n10916 1118.26
R2581 vss.n10956 vss.n10917 1118.26
R2582 vss.n10948 vss.n10917 1118.26
R2583 vss.n11272 vss.n11263 1118.26
R2584 vss.n11279 vss.n11263 1118.26
R2585 vss.n11279 vss.n11260 1118.26
R2586 vss.n11294 vss.n11260 1118.26
R2587 vss.n11294 vss.n11261 1118.26
R2588 vss.n11290 vss.n11261 1118.26
R2589 vss.n11276 vss.n11275 1118.26
R2590 vss.n11277 vss.n11276 1118.26
R2591 vss.n11277 vss.n11255 1118.26
R2592 vss.n11296 vss.n11255 1118.26
R2593 vss.n11296 vss.n11256 1118.26
R2594 vss.n11287 vss.n11256 1118.26
R2595 vss.n11224 vss.n11215 1118.26
R2596 vss.n11230 vss.n11215 1118.26
R2597 vss.n11230 vss.n11212 1118.26
R2598 vss.n11246 vss.n11212 1118.26
R2599 vss.n11246 vss.n11213 1118.26
R2600 vss.n11242 vss.n11213 1118.26
R2601 vss.n11227 vss.n11226 1118.26
R2602 vss.n11228 vss.n11227 1118.26
R2603 vss.n11228 vss.n11207 1118.26
R2604 vss.n11248 vss.n11207 1118.26
R2605 vss.n11248 vss.n11208 1118.26
R2606 vss.n11239 vss.n11208 1118.26
R2607 vss.n11130 vss.n11121 1118.26
R2608 vss.n11137 vss.n11121 1118.26
R2609 vss.n11137 vss.n11118 1118.26
R2610 vss.n11151 vss.n11118 1118.26
R2611 vss.n11151 vss.n11119 1118.26
R2612 vss.n11147 vss.n11119 1118.26
R2613 vss.n11134 vss.n11133 1118.26
R2614 vss.n11135 vss.n11134 1118.26
R2615 vss.n11135 vss.n11113 1118.26
R2616 vss.n11153 vss.n11113 1118.26
R2617 vss.n11153 vss.n11114 1118.26
R2618 vss.n11145 vss.n11114 1118.26
R2619 vss.n11583 vss.n11574 1118.26
R2620 vss.n11590 vss.n11574 1118.26
R2621 vss.n11590 vss.n11571 1118.26
R2622 vss.n11605 vss.n11571 1118.26
R2623 vss.n11605 vss.n11572 1118.26
R2624 vss.n11601 vss.n11572 1118.26
R2625 vss.n11587 vss.n11586 1118.26
R2626 vss.n11588 vss.n11587 1118.26
R2627 vss.n11588 vss.n11566 1118.26
R2628 vss.n11607 vss.n11566 1118.26
R2629 vss.n11607 vss.n11567 1118.26
R2630 vss.n11598 vss.n11567 1118.26
R2631 vss.n11535 vss.n11526 1118.26
R2632 vss.n11541 vss.n11526 1118.26
R2633 vss.n11541 vss.n11523 1118.26
R2634 vss.n11557 vss.n11523 1118.26
R2635 vss.n11557 vss.n11524 1118.26
R2636 vss.n11553 vss.n11524 1118.26
R2637 vss.n11538 vss.n11537 1118.26
R2638 vss.n11539 vss.n11538 1118.26
R2639 vss.n11539 vss.n11518 1118.26
R2640 vss.n11559 vss.n11518 1118.26
R2641 vss.n11559 vss.n11519 1118.26
R2642 vss.n11550 vss.n11519 1118.26
R2643 vss.n9903 vss.n9894 1118.26
R2644 vss.n9907 vss.n9894 1118.26
R2645 vss.n9907 vss.n9885 1118.26
R2646 vss.n11719 vss.n9885 1118.26
R2647 vss.n11719 vss.n9886 1118.26
R2648 vss.n9886 vss.n9881 1118.26
R2649 vss.n9900 vss.n9892 1118.26
R2650 vss.n9909 vss.n9892 1118.26
R2651 vss.n9909 vss.n9888 1118.26
R2652 vss.n11714 vss.n9888 1118.26
R2653 vss.n11715 vss.n11714 1118.26
R2654 vss.n11715 vss.n9880 1118.26
R2655 vss.n13227 vss.n8827 1118.26
R2656 vss.n13235 vss.n8827 1118.26
R2657 vss.n13235 vss.n8821 1118.26
R2658 vss.n13240 vss.n8821 1118.26
R2659 vss.n13240 vss.n8823 1118.26
R2660 vss.n8823 vss.n8812 1118.26
R2661 vss.n13229 vss.n8829 1118.26
R2662 vss.n13233 vss.n8829 1118.26
R2663 vss.n13233 vss.n8817 1118.26
R2664 vss.n13242 vss.n8817 1118.26
R2665 vss.n13242 vss.n8818 1118.26
R2666 vss.n8818 vss.n8813 1118.26
R2667 vss.n11791 vss.n11768 1118.26
R2668 vss.n11787 vss.n11768 1118.26
R2669 vss.n11787 vss.n11774 1118.26
R2670 vss.n11775 vss.n11774 1118.26
R2671 vss.n11776 vss.n11775 1118.26
R2672 vss.n11785 vss.n11776 1118.26
R2673 vss.n11795 vss.n11794 1118.26
R2674 vss.n11796 vss.n11795 1118.26
R2675 vss.n11796 vss.n11761 1118.26
R2676 vss.n11798 vss.n11761 1118.26
R2677 vss.n11798 vss.n11762 1118.26
R2678 vss.n11764 vss.n11762 1118.26
R2679 vss.n11834 vss.n11816 1118.26
R2680 vss.n11834 vss.n11833 1118.26
R2681 vss.n11833 vss.n11818 1118.26
R2682 vss.n11820 vss.n11818 1118.26
R2683 vss.n11821 vss.n11820 1118.26
R2684 vss.n11831 vss.n11821 1118.26
R2685 vss.n11839 vss.n11812 1118.26
R2686 vss.n11812 vss.n11809 1118.26
R2687 vss.n11809 vss.n11806 1118.26
R2688 vss.n12185 vss.n11806 1118.26
R2689 vss.n12185 vss.n11807 1118.26
R2690 vss.n11810 vss.n11807 1118.26
R2691 vss.n11913 vss.n11905 1118.26
R2692 vss.n11921 vss.n11905 1118.26
R2693 vss.n11921 vss.n11899 1118.26
R2694 vss.n11926 vss.n11899 1118.26
R2695 vss.n11926 vss.n11901 1118.26
R2696 vss.n11901 vss.n11890 1118.26
R2697 vss.n11915 vss.n11907 1118.26
R2698 vss.n11919 vss.n11907 1118.26
R2699 vss.n11919 vss.n11895 1118.26
R2700 vss.n11928 vss.n11895 1118.26
R2701 vss.n11928 vss.n11896 1118.26
R2702 vss.n11896 vss.n11891 1118.26
R2703 vss.n11729 vss.n9872 1118.26
R2704 vss.n11738 vss.n9872 1118.26
R2705 vss.n11738 vss.n9869 1118.26
R2706 vss.n11752 vss.n9869 1118.26
R2707 vss.n11752 vss.n9870 1118.26
R2708 vss.n11748 vss.n9870 1118.26
R2709 vss.n11735 vss.n11734 1118.26
R2710 vss.n11736 vss.n11735 1118.26
R2711 vss.n11736 vss.n9864 1118.26
R2712 vss.n11754 vss.n9864 1118.26
R2713 vss.n11754 vss.n9865 1118.26
R2714 vss.n11746 vss.n9865 1118.26
R2715 vss.n9444 vss.n9434 1118.26
R2716 vss.n9450 vss.n9434 1118.26
R2717 vss.n9450 vss.n9431 1118.26
R2718 vss.n9465 vss.n9431 1118.26
R2719 vss.n9465 vss.n9432 1118.26
R2720 vss.n9461 vss.n9432 1118.26
R2721 vss.n9447 vss.n9446 1118.26
R2722 vss.n9448 vss.n9447 1118.26
R2723 vss.n9448 vss.n9426 1118.26
R2724 vss.n9467 vss.n9426 1118.26
R2725 vss.n9467 vss.n9427 1118.26
R2726 vss.n9458 vss.n9427 1118.26
R2727 vss.n9493 vss.n9484 1118.26
R2728 vss.n12481 vss.n9484 1118.26
R2729 vss.n12481 vss.n9481 1118.26
R2730 vss.n12495 vss.n9481 1118.26
R2731 vss.n12495 vss.n9482 1118.26
R2732 vss.n12491 vss.n9482 1118.26
R2733 vss.n12478 vss.n12477 1118.26
R2734 vss.n12479 vss.n12478 1118.26
R2735 vss.n12479 vss.n9476 1118.26
R2736 vss.n12497 vss.n9476 1118.26
R2737 vss.n12497 vss.n9477 1118.26
R2738 vss.n12489 vss.n9477 1118.26
R2739 vss.n9507 vss.n9497 1118.26
R2740 vss.n9534 vss.n9507 1118.26
R2741 vss.n9534 vss.n9508 1118.26
R2742 vss.n9530 vss.n9508 1118.26
R2743 vss.n9530 vss.n9513 1118.26
R2744 vss.n9520 vss.n9513 1118.26
R2745 vss.n9502 vss.n9498 1118.26
R2746 vss.n9536 vss.n9502 1118.26
R2747 vss.n9536 vss.n9503 1118.26
R2748 vss.n9528 vss.n9503 1118.26
R2749 vss.n9528 vss.n9515 1118.26
R2750 vss.n9518 vss.n9515 1118.26
R2751 vss.n9560 vss.n9558 1118.26
R2752 vss.n9586 vss.n9558 1118.26
R2753 vss.n9586 vss.n9559 1118.26
R2754 vss.n9582 vss.n9559 1118.26
R2755 vss.n9582 vss.n9566 1118.26
R2756 vss.n9574 vss.n9566 1118.26
R2757 vss.n9592 vss.n9550 1118.26
R2758 vss.n9588 vss.n9550 1118.26
R2759 vss.n9588 vss.n9554 1118.26
R2760 vss.n9580 vss.n9554 1118.26
R2761 vss.n9580 vss.n9568 1118.26
R2762 vss.n9576 vss.n9568 1118.26
R2763 vss.n9267 vss.n9258 1118.26
R2764 vss.n9267 vss.n9266 1118.26
R2765 vss.n9266 vss.n8892 1118.26
R2766 vss.n13172 vss.n8892 1118.26
R2767 vss.n13172 vss.n8893 1118.26
R2768 vss.n13168 vss.n8893 1118.26
R2769 vss.n9272 vss.n9259 1118.26
R2770 vss.n9264 vss.n9259 1118.26
R2771 vss.n9264 vss.n8887 1118.26
R2772 vss.n13174 vss.n8887 1118.26
R2773 vss.n13174 vss.n8888 1118.26
R2774 vss.n13166 vss.n8888 1118.26
R2775 vss.n12402 vss.n12393 1118.26
R2776 vss.n12408 vss.n12393 1118.26
R2777 vss.n12408 vss.n12390 1118.26
R2778 vss.n12423 vss.n12390 1118.26
R2779 vss.n12423 vss.n12391 1118.26
R2780 vss.n12419 vss.n12391 1118.26
R2781 vss.n12405 vss.n12404 1118.26
R2782 vss.n12406 vss.n12405 1118.26
R2783 vss.n12406 vss.n12385 1118.26
R2784 vss.n12425 vss.n12385 1118.26
R2785 vss.n12425 vss.n12386 1118.26
R2786 vss.n12417 vss.n12386 1118.26
R2787 vss.n9622 vss.n9613 1118.26
R2788 vss.n12362 vss.n9613 1118.26
R2789 vss.n12362 vss.n9610 1118.26
R2790 vss.n12376 vss.n9610 1118.26
R2791 vss.n12376 vss.n9611 1118.26
R2792 vss.n12372 vss.n9611 1118.26
R2793 vss.n12359 vss.n12358 1118.26
R2794 vss.n12360 vss.n12359 1118.26
R2795 vss.n12360 vss.n9605 1118.26
R2796 vss.n12378 vss.n9605 1118.26
R2797 vss.n12378 vss.n9606 1118.26
R2798 vss.n12370 vss.n9606 1118.26
R2799 vss.n9636 vss.n9626 1118.26
R2800 vss.n9664 vss.n9636 1118.26
R2801 vss.n9664 vss.n9637 1118.26
R2802 vss.n9660 vss.n9637 1118.26
R2803 vss.n9660 vss.n9642 1118.26
R2804 vss.n9649 vss.n9642 1118.26
R2805 vss.n9631 vss.n9627 1118.26
R2806 vss.n9666 vss.n9631 1118.26
R2807 vss.n9666 vss.n9632 1118.26
R2808 vss.n9658 vss.n9632 1118.26
R2809 vss.n9658 vss.n9644 1118.26
R2810 vss.n9647 vss.n9644 1118.26
R2811 vss.n9689 vss.n9687 1118.26
R2812 vss.n9716 vss.n9687 1118.26
R2813 vss.n9716 vss.n9688 1118.26
R2814 vss.n9712 vss.n9688 1118.26
R2815 vss.n9712 vss.n9695 1118.26
R2816 vss.n9704 vss.n9695 1118.26
R2817 vss.n9722 vss.n9679 1118.26
R2818 vss.n9718 vss.n9679 1118.26
R2819 vss.n9718 vss.n9683 1118.26
R2820 vss.n9710 vss.n9683 1118.26
R2821 vss.n9710 vss.n9697 1118.26
R2822 vss.n9706 vss.n9697 1118.26
R2823 vss.n13264 vss.n8630 1118.26
R2824 vss.n13270 vss.n8630 1118.26
R2825 vss.n13270 vss.n8627 1118.26
R2826 vss.n13284 vss.n8627 1118.26
R2827 vss.n13284 vss.n8628 1118.26
R2828 vss.n13280 vss.n8628 1118.26
R2829 vss.n13267 vss.n13266 1118.26
R2830 vss.n13268 vss.n13267 1118.26
R2831 vss.n13268 vss.n8622 1118.26
R2832 vss.n13286 vss.n8622 1118.26
R2833 vss.n13286 vss.n8623 1118.26
R2834 vss.n13278 vss.n8623 1118.26
R2835 vss.n12284 vss.n12275 1118.26
R2836 vss.n12290 vss.n12275 1118.26
R2837 vss.n12290 vss.n12272 1118.26
R2838 vss.n12305 vss.n12272 1118.26
R2839 vss.n12305 vss.n12273 1118.26
R2840 vss.n12301 vss.n12273 1118.26
R2841 vss.n12287 vss.n12286 1118.26
R2842 vss.n12288 vss.n12287 1118.26
R2843 vss.n12288 vss.n12267 1118.26
R2844 vss.n12307 vss.n12267 1118.26
R2845 vss.n12307 vss.n12268 1118.26
R2846 vss.n12299 vss.n12268 1118.26
R2847 vss.n9752 vss.n9743 1118.26
R2848 vss.n12244 vss.n9743 1118.26
R2849 vss.n12244 vss.n9740 1118.26
R2850 vss.n12258 vss.n9740 1118.26
R2851 vss.n12258 vss.n9741 1118.26
R2852 vss.n12254 vss.n9741 1118.26
R2853 vss.n12241 vss.n12240 1118.26
R2854 vss.n12242 vss.n12241 1118.26
R2855 vss.n12242 vss.n9735 1118.26
R2856 vss.n12260 vss.n9735 1118.26
R2857 vss.n12260 vss.n9736 1118.26
R2858 vss.n12252 vss.n9736 1118.26
R2859 vss.n9766 vss.n9756 1118.26
R2860 vss.n9793 vss.n9766 1118.26
R2861 vss.n9793 vss.n9767 1118.26
R2862 vss.n9789 vss.n9767 1118.26
R2863 vss.n9789 vss.n9772 1118.26
R2864 vss.n9779 vss.n9772 1118.26
R2865 vss.n9761 vss.n9757 1118.26
R2866 vss.n9795 vss.n9761 1118.26
R2867 vss.n9795 vss.n9762 1118.26
R2868 vss.n9787 vss.n9762 1118.26
R2869 vss.n9787 vss.n9774 1118.26
R2870 vss.n9777 vss.n9774 1118.26
R2871 vss.n9818 vss.n9816 1118.26
R2872 vss.n9844 vss.n9816 1118.26
R2873 vss.n9844 vss.n9817 1118.26
R2874 vss.n9840 vss.n9817 1118.26
R2875 vss.n9840 vss.n9824 1118.26
R2876 vss.n9832 vss.n9824 1118.26
R2877 vss.n9850 vss.n9808 1118.26
R2878 vss.n9846 vss.n9808 1118.26
R2879 vss.n9846 vss.n9812 1118.26
R2880 vss.n9838 vss.n9812 1118.26
R2881 vss.n9838 vss.n9826 1118.26
R2882 vss.n9834 vss.n9826 1118.26
R2883 vss.n8749 vss.n8740 1118.26
R2884 vss.n8749 vss.n8748 1118.26
R2885 vss.n8748 vss.n8348 1118.26
R2886 vss.n13695 vss.n8348 1118.26
R2887 vss.n13695 vss.n8349 1118.26
R2888 vss.n13691 vss.n8349 1118.26
R2889 vss.n8754 vss.n8741 1118.26
R2890 vss.n8746 vss.n8741 1118.26
R2891 vss.n8746 vss.n8343 1118.26
R2892 vss.n13697 vss.n8343 1118.26
R2893 vss.n13697 vss.n8344 1118.26
R2894 vss.n13689 vss.n8344 1118.26
R2895 vss.n11986 vss.n11978 1118.26
R2896 vss.n11994 vss.n11978 1118.26
R2897 vss.n11994 vss.n11972 1118.26
R2898 vss.n11999 vss.n11972 1118.26
R2899 vss.n11999 vss.n11974 1118.26
R2900 vss.n11974 vss.n11964 1118.26
R2901 vss.n11988 vss.n11980 1118.26
R2902 vss.n11992 vss.n11980 1118.26
R2903 vss.n11992 vss.n11968 1118.26
R2904 vss.n12001 vss.n11968 1118.26
R2905 vss.n12001 vss.n11969 1118.26
R2906 vss.n11969 vss.n11965 1118.26
R2907 vss.n12199 vss.n9854 1118.26
R2908 vss.n12227 vss.n12199 1118.26
R2909 vss.n12227 vss.n12200 1118.26
R2910 vss.n12223 vss.n12200 1118.26
R2911 vss.n12223 vss.n12206 1118.26
R2912 vss.n12214 vss.n12206 1118.26
R2913 vss.n12233 vss.n9855 1118.26
R2914 vss.n12229 vss.n9855 1118.26
R2915 vss.n12229 vss.n12196 1118.26
R2916 vss.n12221 vss.n12196 1118.26
R2917 vss.n12221 vss.n12208 1118.26
R2918 vss.n12217 vss.n12208 1118.26
R2919 vss.n8768 vss.n8759 1118.26
R2920 vss.n8796 vss.n8768 1118.26
R2921 vss.n8796 vss.n8769 1118.26
R2922 vss.n8792 vss.n8769 1118.26
R2923 vss.n8792 vss.n8775 1118.26
R2924 vss.n8784 vss.n8775 1118.26
R2925 vss.n8802 vss.n8760 1118.26
R2926 vss.n8798 vss.n8760 1118.26
R2927 vss.n8798 vss.n8765 1118.26
R2928 vss.n8790 vss.n8765 1118.26
R2929 vss.n8790 vss.n8777 1118.26
R2930 vss.n8786 vss.n8777 1118.26
R2931 vss.n8699 vss.n8691 1118.26
R2932 vss.n8727 vss.n8699 1118.26
R2933 vss.n8727 vss.n8700 1118.26
R2934 vss.n8723 vss.n8700 1118.26
R2935 vss.n8723 vss.n8706 1118.26
R2936 vss.n8715 vss.n8706 1118.26
R2937 vss.n8733 vss.n8692 1118.26
R2938 vss.n8729 vss.n8692 1118.26
R2939 vss.n8729 vss.n8696 1118.26
R2940 vss.n8721 vss.n8696 1118.26
R2941 vss.n8721 vss.n8708 1118.26
R2942 vss.n8717 vss.n8708 1118.26
R2943 vss.n12317 vss.n9726 1118.26
R2944 vss.n12345 vss.n12317 1118.26
R2945 vss.n12345 vss.n12318 1118.26
R2946 vss.n12341 vss.n12318 1118.26
R2947 vss.n12341 vss.n12324 1118.26
R2948 vss.n12332 vss.n12324 1118.26
R2949 vss.n12351 vss.n9727 1118.26
R2950 vss.n12347 vss.n9727 1118.26
R2951 vss.n12347 vss.n12314 1118.26
R2952 vss.n12339 vss.n12314 1118.26
R2953 vss.n12339 vss.n12326 1118.26
R2954 vss.n12335 vss.n12326 1118.26
R2955 vss.n8649 vss.n8640 1118.26
R2956 vss.n8677 vss.n8649 1118.26
R2957 vss.n8677 vss.n8650 1118.26
R2958 vss.n8673 vss.n8650 1118.26
R2959 vss.n8673 vss.n8656 1118.26
R2960 vss.n8665 vss.n8656 1118.26
R2961 vss.n8683 vss.n8641 1118.26
R2962 vss.n8679 vss.n8641 1118.26
R2963 vss.n8679 vss.n8646 1118.26
R2964 vss.n8671 vss.n8646 1118.26
R2965 vss.n8671 vss.n8658 1118.26
R2966 vss.n8667 vss.n8658 1118.26
R2967 vss.n12918 vss.n9198 1118.26
R2968 vss.n12926 vss.n9198 1118.26
R2969 vss.n12926 vss.n9192 1118.26
R2970 vss.n12931 vss.n9192 1118.26
R2971 vss.n12931 vss.n9194 1118.26
R2972 vss.n9194 vss.n9183 1118.26
R2973 vss.n12920 vss.n9200 1118.26
R2974 vss.n12924 vss.n9200 1118.26
R2975 vss.n12924 vss.n9188 1118.26
R2976 vss.n12933 vss.n9188 1118.26
R2977 vss.n12933 vss.n9189 1118.26
R2978 vss.n9189 vss.n9184 1118.26
R2979 vss.n12436 vss.n9596 1118.26
R2980 vss.n12464 vss.n12436 1118.26
R2981 vss.n12464 vss.n12437 1118.26
R2982 vss.n12460 vss.n12437 1118.26
R2983 vss.n12460 vss.n12443 1118.26
R2984 vss.n12451 vss.n12443 1118.26
R2985 vss.n12470 vss.n9597 1118.26
R2986 vss.n12466 vss.n9597 1118.26
R2987 vss.n12466 vss.n12433 1118.26
R2988 vss.n12458 vss.n12433 1118.26
R2989 vss.n12458 vss.n12445 1118.26
R2990 vss.n12454 vss.n12445 1118.26
R2991 vss.n9219 vss.n9210 1118.26
R2992 vss.n9247 vss.n9219 1118.26
R2993 vss.n9247 vss.n9220 1118.26
R2994 vss.n9243 vss.n9220 1118.26
R2995 vss.n9243 vss.n9226 1118.26
R2996 vss.n9235 vss.n9226 1118.26
R2997 vss.n9253 vss.n9211 1118.26
R2998 vss.n9249 vss.n9211 1118.26
R2999 vss.n9249 vss.n9216 1118.26
R3000 vss.n9241 vss.n9216 1118.26
R3001 vss.n9241 vss.n9228 1118.26
R3002 vss.n9237 vss.n9228 1118.26
R3003 vss.n9336 vss.n9328 1118.26
R3004 vss.n9344 vss.n9328 1118.26
R3005 vss.n9344 vss.n9322 1118.26
R3006 vss.n9349 vss.n9322 1118.26
R3007 vss.n9349 vss.n9324 1118.26
R3008 vss.n9324 vss.n9312 1118.26
R3009 vss.n9338 vss.n9330 1118.26
R3010 vss.n9342 vss.n9330 1118.26
R3011 vss.n9342 vss.n9318 1118.26
R3012 vss.n9351 vss.n9318 1118.26
R3013 vss.n9351 vss.n9319 1118.26
R3014 vss.n9319 vss.n9313 1118.26
R3015 vss.n12522 vss.n12514 1118.26
R3016 vss.n12530 vss.n12514 1118.26
R3017 vss.n12530 vss.n12508 1118.26
R3018 vss.n12535 vss.n12508 1118.26
R3019 vss.n12535 vss.n12510 1118.26
R3020 vss.n12510 vss.n9419 1118.26
R3021 vss.n12524 vss.n12516 1118.26
R3022 vss.n12528 vss.n12516 1118.26
R3023 vss.n12528 vss.n12504 1118.26
R3024 vss.n12537 vss.n12504 1118.26
R3025 vss.n12537 vss.n12505 1118.26
R3026 vss.n12505 vss.n9420 1118.26
R3027 vss.n12672 vss.n12664 1118.26
R3028 vss.n12680 vss.n12664 1118.26
R3029 vss.n12680 vss.n12658 1118.26
R3030 vss.n12685 vss.n12658 1118.26
R3031 vss.n12685 vss.n12660 1118.26
R3032 vss.n12660 vss.n12649 1118.26
R3033 vss.n12674 vss.n12666 1118.26
R3034 vss.n12678 vss.n12666 1118.26
R3035 vss.n12678 vss.n12654 1118.26
R3036 vss.n12687 vss.n12654 1118.26
R3037 vss.n12687 vss.n12655 1118.26
R3038 vss.n12655 vss.n12650 1118.26
R3039 vss.n10192 vss.n10191 1118.26
R3040 vss.n10193 vss.n10192 1118.26
R3041 vss.n10193 vss.n10172 1118.26
R3042 vss.n10210 vss.n10172 1118.26
R3043 vss.n10210 vss.n10173 1118.26
R3044 vss.n10200 vss.n10173 1118.26
R3045 vss.n10189 vss.n10180 1118.26
R3046 vss.n10195 vss.n10180 1118.26
R3047 vss.n10195 vss.n10177 1118.26
R3048 vss.n10208 vss.n10177 1118.26
R3049 vss.n10208 vss.n10178 1118.26
R3050 vss.n10204 vss.n10178 1118.26
R3051 vss.n11089 vss.n11088 1118.26
R3052 vss.n11090 vss.n11089 1118.26
R3053 vss.n11090 vss.n11069 1118.26
R3054 vss.n11107 vss.n11069 1118.26
R3055 vss.n11107 vss.n11070 1118.26
R3056 vss.n11097 vss.n11070 1118.26
R3057 vss.n11086 vss.n11077 1118.26
R3058 vss.n11092 vss.n11077 1118.26
R3059 vss.n11092 vss.n11074 1118.26
R3060 vss.n11105 vss.n11074 1118.26
R3061 vss.n11105 vss.n11075 1118.26
R3062 vss.n11101 vss.n11075 1118.26
R3063 vss.n11494 vss.n11493 1118.26
R3064 vss.n11495 vss.n11494 1118.26
R3065 vss.n11495 vss.n11474 1118.26
R3066 vss.n11512 vss.n11474 1118.26
R3067 vss.n11512 vss.n11475 1118.26
R3068 vss.n11502 vss.n11475 1118.26
R3069 vss.n11491 vss.n11482 1118.26
R3070 vss.n11497 vss.n11482 1118.26
R3071 vss.n11497 vss.n11479 1118.26
R3072 vss.n11510 vss.n11479 1118.26
R3073 vss.n11510 vss.n11480 1118.26
R3074 vss.n11506 vss.n11480 1118.26
R3075 vss.n12146 vss.n12134 1118.26
R3076 vss.n12172 vss.n12146 1118.26
R3077 vss.n12172 vss.n12147 1118.26
R3078 vss.n12168 vss.n12147 1118.26
R3079 vss.n12168 vss.n12152 1118.26
R3080 vss.n12160 vss.n12152 1118.26
R3081 vss.n12141 vss.n12135 1118.26
R3082 vss.n12174 vss.n12141 1118.26
R3083 vss.n12174 vss.n12142 1118.26
R3084 vss.n12166 vss.n12142 1118.26
R3085 vss.n12166 vss.n12154 1118.26
R3086 vss.n12162 vss.n12154 1118.26
R3087 vss.n15632 vss.n15627 1118.26
R3088 vss.n15632 vss.n15628 1118.26
R3089 vss.n15629 vss.n15628 1118.26
R3090 vss.n15647 vss.n15629 1118.26
R3091 vss.n15647 vss.n15626 1118.26
R3092 vss.n15649 vss.n15626 1118.26
R3093 vss.n15633 vss.n356 1118.26
R3094 vss.n15633 vss.n354 1118.26
R3095 vss.n357 vss.n354 1118.26
R3096 vss.n15655 vss.n357 1118.26
R3097 vss.n15655 vss.n358 1118.26
R3098 vss.n358 vss.n355 1118.26
R3099 vss.n3588 vss.n3580 1118.26
R3100 vss.n3598 vss.n3580 1118.26
R3101 vss.n3598 vss.n3574 1118.26
R3102 vss.n3603 vss.n3574 1118.26
R3103 vss.n3603 vss.n3576 1118.26
R3104 vss.n3576 vss.n3565 1118.26
R3105 vss.n3592 vss.n3582 1118.26
R3106 vss.n3596 vss.n3582 1118.26
R3107 vss.n3596 vss.n3570 1118.26
R3108 vss.n3605 vss.n3570 1118.26
R3109 vss.n3605 vss.n3571 1118.26
R3110 vss.n3571 vss.n3566 1118.26
R3111 vss.n3974 vss.n3970 1118.26
R3112 vss.n3978 vss.n3974 1118.26
R3113 vss.n3978 vss.n8 1118.26
R3114 vss.n15899 vss.n8 1118.26
R3115 vss.n15899 vss.n9 1118.26
R3116 vss.n15895 vss.n9 1118.26
R3117 vss.n3975 vss.n3971 1118.26
R3118 vss.n3976 vss.n3975 1118.26
R3119 vss.n3976 vss.n3 1118.26
R3120 vss.n15901 vss.n3 1118.26
R3121 vss.n15901 vss.n4 1118.26
R3122 vss.n15893 vss.n4 1118.26
R3123 vss.n6296 vss.n6292 1118.26
R3124 vss.n6300 vss.n6296 1118.26
R3125 vss.n6300 vss.n252 1118.26
R3126 vss.n15696 vss.n252 1118.26
R3127 vss.n15696 vss.n253 1118.26
R3128 vss.n15692 vss.n253 1118.26
R3129 vss.n6297 vss.n6293 1118.26
R3130 vss.n6298 vss.n6297 1118.26
R3131 vss.n6298 vss.n247 1118.26
R3132 vss.n15698 vss.n247 1118.26
R3133 vss.n15698 vss.n248 1118.26
R3134 vss.n15690 vss.n248 1118.26
R3135 vss.n5652 vss.n5643 1118.26
R3136 vss.n5658 vss.n5643 1118.26
R3137 vss.n5658 vss.n5640 1118.26
R3138 vss.n5672 vss.n5640 1118.26
R3139 vss.n5672 vss.n5641 1118.26
R3140 vss.n5668 vss.n5641 1118.26
R3141 vss.n5655 vss.n5654 1118.26
R3142 vss.n5656 vss.n5655 1118.26
R3143 vss.n5656 vss.n5635 1118.26
R3144 vss.n5674 vss.n5635 1118.26
R3145 vss.n5674 vss.n5636 1118.26
R3146 vss.n5666 vss.n5636 1118.26
R3147 vss.n3721 vss.n3712 1118.26
R3148 vss.n3721 vss.n3720 1118.26
R3149 vss.n3720 vss.n173 1118.26
R3150 vss.n15752 vss.n173 1118.26
R3151 vss.n15752 vss.n174 1118.26
R3152 vss.n15748 vss.n174 1118.26
R3153 vss.n3726 vss.n3713 1118.26
R3154 vss.n3718 vss.n3713 1118.26
R3155 vss.n3718 vss.n168 1118.26
R3156 vss.n15754 vss.n168 1118.26
R3157 vss.n15754 vss.n169 1118.26
R3158 vss.n15746 vss.n169 1118.26
R3159 vss.n3673 vss.n3665 1118.26
R3160 vss.n3701 vss.n3673 1118.26
R3161 vss.n3701 vss.n3674 1118.26
R3162 vss.n3697 vss.n3674 1118.26
R3163 vss.n3697 vss.n3680 1118.26
R3164 vss.n3689 vss.n3680 1118.26
R3165 vss.n3707 vss.n3666 1118.26
R3166 vss.n3703 vss.n3666 1118.26
R3167 vss.n3703 vss.n3670 1118.26
R3168 vss.n3695 vss.n3670 1118.26
R3169 vss.n3695 vss.n3682 1118.26
R3170 vss.n3691 vss.n3682 1118.26
R3171 vss.n5844 vss.n5835 1118.26
R3172 vss.n5850 vss.n5835 1118.26
R3173 vss.n5850 vss.n5832 1118.26
R3174 vss.n5864 vss.n5832 1118.26
R3175 vss.n5864 vss.n5833 1118.26
R3176 vss.n5860 vss.n5833 1118.26
R3177 vss.n5847 vss.n5846 1118.26
R3178 vss.n5848 vss.n5847 1118.26
R3179 vss.n5848 vss.n5827 1118.26
R3180 vss.n5866 vss.n5827 1118.26
R3181 vss.n5866 vss.n5828 1118.26
R3182 vss.n5858 vss.n5828 1118.26
R3183 vss.n3840 vss.n3831 1118.26
R3184 vss.n3840 vss.n3839 1118.26
R3185 vss.n3839 vss.n95 1118.26
R3186 vss.n15808 vss.n95 1118.26
R3187 vss.n15808 vss.n96 1118.26
R3188 vss.n15804 vss.n96 1118.26
R3189 vss.n3845 vss.n3832 1118.26
R3190 vss.n3837 vss.n3832 1118.26
R3191 vss.n3837 vss.n90 1118.26
R3192 vss.n15810 vss.n90 1118.26
R3193 vss.n15810 vss.n91 1118.26
R3194 vss.n15802 vss.n91 1118.26
R3195 vss.n3792 vss.n3784 1118.26
R3196 vss.n3820 vss.n3792 1118.26
R3197 vss.n3820 vss.n3793 1118.26
R3198 vss.n3816 vss.n3793 1118.26
R3199 vss.n3816 vss.n3799 1118.26
R3200 vss.n3808 vss.n3799 1118.26
R3201 vss.n3826 vss.n3785 1118.26
R3202 vss.n3822 vss.n3785 1118.26
R3203 vss.n3822 vss.n3789 1118.26
R3204 vss.n3814 vss.n3789 1118.26
R3205 vss.n3814 vss.n3801 1118.26
R3206 vss.n3810 vss.n3801 1118.26
R3207 vss.n3911 vss.n3903 1118.26
R3208 vss.n3939 vss.n3911 1118.26
R3209 vss.n3939 vss.n3912 1118.26
R3210 vss.n3935 vss.n3912 1118.26
R3211 vss.n3935 vss.n3918 1118.26
R3212 vss.n3927 vss.n3918 1118.26
R3213 vss.n3945 vss.n3904 1118.26
R3214 vss.n3941 vss.n3904 1118.26
R3215 vss.n3941 vss.n3908 1118.26
R3216 vss.n3933 vss.n3908 1118.26
R3217 vss.n3933 vss.n3920 1118.26
R3218 vss.n3929 vss.n3920 1118.26
R3219 vss.n6084 vss.n6075 1118.26
R3220 vss.n6090 vss.n6075 1118.26
R3221 vss.n6090 vss.n6072 1118.26
R3222 vss.n6104 vss.n6072 1118.26
R3223 vss.n6104 vss.n6073 1118.26
R3224 vss.n6100 vss.n6073 1118.26
R3225 vss.n6087 vss.n6086 1118.26
R3226 vss.n6088 vss.n6087 1118.26
R3227 vss.n6088 vss.n6067 1118.26
R3228 vss.n6106 vss.n6067 1118.26
R3229 vss.n6106 vss.n6068 1118.26
R3230 vss.n6098 vss.n6068 1118.26
R3231 vss.n6036 vss.n6027 1118.26
R3232 vss.n6042 vss.n6027 1118.26
R3233 vss.n6042 vss.n6024 1118.26
R3234 vss.n6057 vss.n6024 1118.26
R3235 vss.n6057 vss.n6025 1118.26
R3236 vss.n6053 vss.n6025 1118.26
R3237 vss.n6039 vss.n6038 1118.26
R3238 vss.n6040 vss.n6039 1118.26
R3239 vss.n6040 vss.n6019 1118.26
R3240 vss.n6059 vss.n6019 1118.26
R3241 vss.n6059 vss.n6020 1118.26
R3242 vss.n6050 vss.n6020 1118.26
R3243 vss.n6164 vss.n6153 1118.26
R3244 vss.n6191 vss.n6164 1118.26
R3245 vss.n6191 vss.n6165 1118.26
R3246 vss.n6187 vss.n6165 1118.26
R3247 vss.n6187 vss.n6170 1118.26
R3248 vss.n6178 vss.n6170 1118.26
R3249 vss.n6159 vss.n6154 1118.26
R3250 vss.n6193 vss.n6159 1118.26
R3251 vss.n6193 vss.n6160 1118.26
R3252 vss.n6185 vss.n6160 1118.26
R3253 vss.n6185 vss.n6172 1118.26
R3254 vss.n6181 vss.n6172 1118.26
R3255 vss.n5746 vss.n5740 1118.26
R3256 vss.n5756 vss.n5740 1118.26
R3257 vss.n5756 vss.n5737 1118.26
R3258 vss.n5770 vss.n5737 1118.26
R3259 vss.n5770 vss.n5738 1118.26
R3260 vss.n5766 vss.n5738 1118.26
R3261 vss.n5753 vss.n5752 1118.26
R3262 vss.n5754 vss.n5753 1118.26
R3263 vss.n5754 vss.n5732 1118.26
R3264 vss.n5772 vss.n5732 1118.26
R3265 vss.n5772 vss.n5733 1118.26
R3266 vss.n5764 vss.n5733 1118.26
R3267 vss.n5796 vss.n5787 1118.26
R3268 vss.n5802 vss.n5787 1118.26
R3269 vss.n5802 vss.n5784 1118.26
R3270 vss.n5817 vss.n5784 1118.26
R3271 vss.n5817 vss.n5785 1118.26
R3272 vss.n5813 vss.n5785 1118.26
R3273 vss.n5799 vss.n5798 1118.26
R3274 vss.n5800 vss.n5799 1118.26
R3275 vss.n5800 vss.n5779 1118.26
R3276 vss.n5819 vss.n5779 1118.26
R3277 vss.n5819 vss.n5780 1118.26
R3278 vss.n5810 vss.n5780 1118.26
R3279 vss.n5925 vss.n5914 1118.26
R3280 vss.n5952 vss.n5925 1118.26
R3281 vss.n5952 vss.n5926 1118.26
R3282 vss.n5948 vss.n5926 1118.26
R3283 vss.n5948 vss.n5931 1118.26
R3284 vss.n5939 vss.n5931 1118.26
R3285 vss.n5920 vss.n5915 1118.26
R3286 vss.n5954 vss.n5920 1118.26
R3287 vss.n5954 vss.n5921 1118.26
R3288 vss.n5946 vss.n5921 1118.26
R3289 vss.n5946 vss.n5933 1118.26
R3290 vss.n5942 vss.n5933 1118.26
R3291 vss.n5558 vss.n5552 1118.26
R3292 vss.n5568 vss.n5552 1118.26
R3293 vss.n5568 vss.n5549 1118.26
R3294 vss.n5582 vss.n5549 1118.26
R3295 vss.n5582 vss.n5550 1118.26
R3296 vss.n5578 vss.n5550 1118.26
R3297 vss.n5565 vss.n5564 1118.26
R3298 vss.n5566 vss.n5565 1118.26
R3299 vss.n5566 vss.n5544 1118.26
R3300 vss.n5584 vss.n5544 1118.26
R3301 vss.n5584 vss.n5545 1118.26
R3302 vss.n5576 vss.n5545 1118.26
R3303 vss.n5687 vss.n5537 1118.26
R3304 vss.n5714 vss.n5687 1118.26
R3305 vss.n5714 vss.n5688 1118.26
R3306 vss.n5710 vss.n5688 1118.26
R3307 vss.n5710 vss.n5693 1118.26
R3308 vss.n5701 vss.n5693 1118.26
R3309 vss.n5682 vss.n5538 1118.26
R3310 vss.n5716 vss.n5682 1118.26
R3311 vss.n5716 vss.n5683 1118.26
R3312 vss.n5708 vss.n5683 1118.26
R3313 vss.n5708 vss.n5695 1118.26
R3314 vss.n5704 vss.n5695 1118.26
R3315 vss.n3548 vss.n3537 1118.26
R3316 vss.n6324 vss.n3548 1118.26
R3317 vss.n6324 vss.n3549 1118.26
R3318 vss.n6320 vss.n3549 1118.26
R3319 vss.n6320 vss.n3554 1118.26
R3320 vss.n3562 vss.n3554 1118.26
R3321 vss.n3543 vss.n3538 1118.26
R3322 vss.n6326 vss.n3543 1118.26
R3323 vss.n6326 vss.n3544 1118.26
R3324 vss.n6318 vss.n3544 1118.26
R3325 vss.n6318 vss.n3556 1118.26
R3326 vss.n6314 vss.n3556 1118.26
R3327 vss.n5603 vss.n5599 1118.26
R3328 vss.n5613 vss.n5599 1118.26
R3329 vss.n5613 vss.n5596 1118.26
R3330 vss.n5627 vss.n5596 1118.26
R3331 vss.n5627 vss.n5597 1118.26
R3332 vss.n5623 vss.n5597 1118.26
R3333 vss.n5610 vss.n5609 1118.26
R3334 vss.n5611 vss.n5610 1118.26
R3335 vss.n5611 vss.n5591 1118.26
R3336 vss.n5629 vss.n5591 1118.26
R3337 vss.n5629 vss.n5592 1118.26
R3338 vss.n5621 vss.n5592 1118.26
R3339 vss.n5879 vss.n5877 1118.26
R3340 vss.n5905 vss.n5877 1118.26
R3341 vss.n5905 vss.n5878 1118.26
R3342 vss.n5901 vss.n5878 1118.26
R3343 vss.n5901 vss.n5885 1118.26
R3344 vss.n5893 vss.n5885 1118.26
R3345 vss.n5911 vss.n5726 1118.26
R3346 vss.n5907 vss.n5726 1118.26
R3347 vss.n5907 vss.n5873 1118.26
R3348 vss.n5899 vss.n5873 1118.26
R3349 vss.n5899 vss.n5887 1118.26
R3350 vss.n5895 vss.n5887 1118.26
R3351 vss.n6118 vss.n6116 1118.26
R3352 vss.n6144 vss.n6116 1118.26
R3353 vss.n6144 vss.n6117 1118.26
R3354 vss.n6140 vss.n6117 1118.26
R3355 vss.n6140 vss.n6124 1118.26
R3356 vss.n6132 vss.n6124 1118.26
R3357 vss.n6150 vss.n5966 1118.26
R3358 vss.n6146 vss.n5966 1118.26
R3359 vss.n6146 vss.n6112 1118.26
R3360 vss.n6138 vss.n6112 1118.26
R3361 vss.n6138 vss.n6126 1118.26
R3362 vss.n6134 vss.n6126 1118.26
R3363 vss.n5986 vss.n5980 1118.26
R3364 vss.n5996 vss.n5980 1118.26
R3365 vss.n5996 vss.n5977 1118.26
R3366 vss.n6010 vss.n5977 1118.26
R3367 vss.n6010 vss.n5978 1118.26
R3368 vss.n6006 vss.n5978 1118.26
R3369 vss.n5993 vss.n5992 1118.26
R3370 vss.n5994 vss.n5993 1118.26
R3371 vss.n5994 vss.n5972 1118.26
R3372 vss.n6012 vss.n5972 1118.26
R3373 vss.n6012 vss.n5973 1118.26
R3374 vss.n6004 vss.n5973 1118.26
R3375 vss.n3297 vss.n3296 1118.26
R3376 vss.n3298 vss.n3297 1118.26
R3377 vss.n3298 vss.n3277 1118.26
R3378 vss.n6736 vss.n3277 1118.26
R3379 vss.n6736 vss.n3278 1118.26
R3380 vss.n6728 vss.n3278 1118.26
R3381 vss.n3294 vss.n3285 1118.26
R3382 vss.n3300 vss.n3285 1118.26
R3383 vss.n3300 vss.n3282 1118.26
R3384 vss.n6734 vss.n3282 1118.26
R3385 vss.n6734 vss.n3283 1118.26
R3386 vss.n6730 vss.n3283 1118.26
R3387 vss.n4377 vss.n4367 1118.26
R3388 vss.n4545 vss.n4377 1118.26
R3389 vss.n4545 vss.n4378 1118.26
R3390 vss.n4399 vss.n4378 1118.26
R3391 vss.n4399 vss.n4383 1118.26
R3392 vss.n4391 vss.n4383 1118.26
R3393 vss.n4372 vss.n4368 1118.26
R3394 vss.n4547 vss.n4372 1118.26
R3395 vss.n4547 vss.n4373 1118.26
R3396 vss.n4397 vss.n4373 1118.26
R3397 vss.n4397 vss.n4385 1118.26
R3398 vss.n4393 vss.n4385 1118.26
R3399 vss.n4467 vss.n4458 1118.26
R3400 vss.n4473 vss.n4458 1118.26
R3401 vss.n4473 vss.n4455 1118.26
R3402 vss.n4488 vss.n4455 1118.26
R3403 vss.n4488 vss.n4456 1118.26
R3404 vss.n4484 vss.n4456 1118.26
R3405 vss.n4470 vss.n4469 1118.26
R3406 vss.n4471 vss.n4470 1118.26
R3407 vss.n4471 vss.n4450 1118.26
R3408 vss.n4490 vss.n4450 1118.26
R3409 vss.n4490 vss.n4451 1118.26
R3410 vss.n4481 vss.n4451 1118.26
R3411 vss.n4514 vss.n4505 1118.26
R3412 vss.n4521 vss.n4505 1118.26
R3413 vss.n4521 vss.n4502 1118.26
R3414 vss.n4535 vss.n4502 1118.26
R3415 vss.n4535 vss.n4503 1118.26
R3416 vss.n4531 vss.n4503 1118.26
R3417 vss.n4518 vss.n4517 1118.26
R3418 vss.n4519 vss.n4518 1118.26
R3419 vss.n4519 vss.n4497 1118.26
R3420 vss.n4537 vss.n4497 1118.26
R3421 vss.n4537 vss.n4498 1118.26
R3422 vss.n4529 vss.n4498 1118.26
R3423 vss.n5019 vss.n5010 1118.26
R3424 vss.n5026 vss.n5010 1118.26
R3425 vss.n5026 vss.n5007 1118.26
R3426 vss.n5040 vss.n5007 1118.26
R3427 vss.n5040 vss.n5008 1118.26
R3428 vss.n5036 vss.n5008 1118.26
R3429 vss.n5023 vss.n5022 1118.26
R3430 vss.n5024 vss.n5023 1118.26
R3431 vss.n5024 vss.n5002 1118.26
R3432 vss.n5042 vss.n5002 1118.26
R3433 vss.n5042 vss.n5003 1118.26
R3434 vss.n5034 vss.n5003 1118.26
R3435 vss.n4192 vss.n4183 1118.26
R3436 vss.n4201 vss.n4183 1118.26
R3437 vss.n4201 vss.n4181 1118.26
R3438 vss.n4207 vss.n4181 1118.26
R3439 vss.n4208 vss.n4207 1118.26
R3440 vss.n4208 vss.n4179 1118.26
R3441 vss.n4195 vss.n4194 1118.26
R3442 vss.n4196 vss.n4195 1118.26
R3443 vss.n4197 vss.n4196 1118.26
R3444 vss.n4197 vss.n4175 1118.26
R3445 vss.n4178 vss.n4175 1118.26
R3446 vss.n4214 vss.n4178 1118.26
R3447 vss.n5067 vss.n5058 1118.26
R3448 vss.n5074 vss.n5058 1118.26
R3449 vss.n5074 vss.n5055 1118.26
R3450 vss.n5088 vss.n5055 1118.26
R3451 vss.n5088 vss.n5056 1118.26
R3452 vss.n5084 vss.n5056 1118.26
R3453 vss.n5071 vss.n5070 1118.26
R3454 vss.n5072 vss.n5071 1118.26
R3455 vss.n5072 vss.n5050 1118.26
R3456 vss.n5090 vss.n5050 1118.26
R3457 vss.n5090 vss.n5051 1118.26
R3458 vss.n5082 vss.n5051 1118.26
R3459 vss.n5493 vss.n5484 1118.26
R3460 vss.n5500 vss.n5484 1118.26
R3461 vss.n5500 vss.n5481 1118.26
R3462 vss.n5514 vss.n5481 1118.26
R3463 vss.n5514 vss.n5482 1118.26
R3464 vss.n5510 vss.n5482 1118.26
R3465 vss.n5497 vss.n5496 1118.26
R3466 vss.n5498 vss.n5497 1118.26
R3467 vss.n5498 vss.n5476 1118.26
R3468 vss.n5516 vss.n5476 1118.26
R3469 vss.n5516 vss.n5477 1118.26
R3470 vss.n5508 vss.n5477 1118.26
R3471 vss.n4029 vss.n4021 1118.26
R3472 vss.n4034 vss.n4021 1118.26
R3473 vss.n4034 vss.n4012 1118.26
R3474 vss.n5526 vss.n4012 1118.26
R3475 vss.n5527 vss.n5526 1118.26
R3476 vss.n5529 vss.n5527 1118.26
R3477 vss.n4027 vss.n4019 1118.26
R3478 vss.n4036 vss.n4019 1118.26
R3479 vss.n4036 vss.n4015 1118.26
R3480 vss.n5523 vss.n4015 1118.26
R3481 vss.n5523 vss.n4006 1118.26
R3482 vss.n5533 vss.n4006 1118.26
R3483 vss.n5278 vss.n5269 1118.26
R3484 vss.n5285 vss.n5269 1118.26
R3485 vss.n5285 vss.n5266 1118.26
R3486 vss.n5300 vss.n5266 1118.26
R3487 vss.n5300 vss.n5267 1118.26
R3488 vss.n5296 vss.n5267 1118.26
R3489 vss.n5282 vss.n5281 1118.26
R3490 vss.n5283 vss.n5282 1118.26
R3491 vss.n5283 vss.n5261 1118.26
R3492 vss.n5302 vss.n5261 1118.26
R3493 vss.n5302 vss.n5262 1118.26
R3494 vss.n5293 vss.n5262 1118.26
R3495 vss.n3465 vss.n3455 1118.26
R3496 vss.n3469 vss.n3455 1118.26
R3497 vss.n3469 vss.n3447 1118.26
R3498 vss.n3480 vss.n3447 1118.26
R3499 vss.n3480 vss.n3448 1118.26
R3500 vss.n3448 vss.n3443 1118.26
R3501 vss.n3462 vss.n3452 1118.26
R3502 vss.n3471 vss.n3452 1118.26
R3503 vss.n3472 vss.n3471 1118.26
R3504 vss.n3475 vss.n3472 1118.26
R3505 vss.n3476 vss.n3475 1118.26
R3506 vss.n3476 vss.n3442 1118.26
R3507 vss.n6353 vss.n6345 1118.26
R3508 vss.n6349 vss.n6345 1118.26
R3509 vss.n6349 vss.n6339 1118.26
R3510 vss.n6362 vss.n6339 1118.26
R3511 vss.n6362 vss.n6337 1118.26
R3512 vss.n6366 vss.n6337 1118.26
R3513 vss.n6356 vss.n6355 1118.26
R3514 vss.n6357 vss.n6356 1118.26
R3515 vss.n6358 vss.n6357 1118.26
R3516 vss.n6358 vss.n3436 1118.26
R3517 vss.n3439 vss.n3436 1118.26
R3518 vss.n6370 vss.n3439 1118.26
R3519 vss.n6669 vss.n6667 1118.26
R3520 vss.n6695 vss.n6667 1118.26
R3521 vss.n6695 vss.n6668 1118.26
R3522 vss.n6691 vss.n6668 1118.26
R3523 vss.n6691 vss.n6675 1118.26
R3524 vss.n6682 vss.n6675 1118.26
R3525 vss.n6701 vss.n3338 1118.26
R3526 vss.n6697 vss.n3338 1118.26
R3527 vss.n6697 vss.n6664 1118.26
R3528 vss.n6676 vss.n6664 1118.26
R3529 vss.n6678 vss.n6676 1118.26
R3530 vss.n6684 vss.n6678 1118.26
R3531 vss.n6638 vss.n6637 1118.26
R3532 vss.n6639 vss.n6638 1118.26
R3533 vss.n6639 vss.n6618 1118.26
R3534 vss.n6657 vss.n6618 1118.26
R3535 vss.n6657 vss.n6619 1118.26
R3536 vss.n6649 vss.n6619 1118.26
R3537 vss.n6635 vss.n6626 1118.26
R3538 vss.n6641 vss.n6626 1118.26
R3539 vss.n6641 vss.n6623 1118.26
R3540 vss.n6655 vss.n6623 1118.26
R3541 vss.n6655 vss.n6624 1118.26
R3542 vss.n6651 vss.n6624 1118.26
R3543 vss.n6589 vss.n6588 1118.26
R3544 vss.n6590 vss.n6589 1118.26
R3545 vss.n6590 vss.n6500 1118.26
R3546 vss.n6609 vss.n6500 1118.26
R3547 vss.n6609 vss.n6501 1118.26
R3548 vss.n6601 vss.n6501 1118.26
R3549 vss.n6586 vss.n6508 1118.26
R3550 vss.n6592 vss.n6508 1118.26
R3551 vss.n6592 vss.n6505 1118.26
R3552 vss.n6607 vss.n6505 1118.26
R3553 vss.n6607 vss.n6506 1118.26
R3554 vss.n6603 vss.n6506 1118.26
R3555 vss.n5236 vss.n5235 1118.26
R3556 vss.n5237 vss.n5236 1118.26
R3557 vss.n5237 vss.n5216 1118.26
R3558 vss.n5255 vss.n5216 1118.26
R3559 vss.n5255 vss.n5217 1118.26
R3560 vss.n5247 vss.n5217 1118.26
R3561 vss.n5233 vss.n5224 1118.26
R3562 vss.n5239 vss.n5224 1118.26
R3563 vss.n5239 vss.n5221 1118.26
R3564 vss.n5253 vss.n5221 1118.26
R3565 vss.n5253 vss.n5222 1118.26
R3566 vss.n5249 vss.n5222 1118.26
R3567 vss.n4061 vss.n4060 1118.26
R3568 vss.n4062 vss.n4061 1118.26
R3569 vss.n4062 vss.n4041 1118.26
R3570 vss.n4079 vss.n4041 1118.26
R3571 vss.n4079 vss.n4042 1118.26
R3572 vss.n4069 vss.n4042 1118.26
R3573 vss.n4058 vss.n4049 1118.26
R3574 vss.n4064 vss.n4049 1118.26
R3575 vss.n4064 vss.n4046 1118.26
R3576 vss.n4077 vss.n4046 1118.26
R3577 vss.n4077 vss.n4047 1118.26
R3578 vss.n4073 vss.n4047 1118.26
R3579 vss.n5448 vss.n5447 1118.26
R3580 vss.n5449 vss.n5448 1118.26
R3581 vss.n5449 vss.n5428 1118.26
R3582 vss.n5467 vss.n5428 1118.26
R3583 vss.n5467 vss.n5429 1118.26
R3584 vss.n5459 vss.n5429 1118.26
R3585 vss.n5445 vss.n5436 1118.26
R3586 vss.n5451 vss.n5436 1118.26
R3587 vss.n5451 vss.n5433 1118.26
R3588 vss.n5465 vss.n5433 1118.26
R3589 vss.n5465 vss.n5434 1118.26
R3590 vss.n5461 vss.n5434 1118.26
R3591 vss.n5401 vss.n5400 1118.26
R3592 vss.n5402 vss.n5401 1118.26
R3593 vss.n5402 vss.n5313 1118.26
R3594 vss.n5420 vss.n5313 1118.26
R3595 vss.n5420 vss.n5314 1118.26
R3596 vss.n5412 vss.n5314 1118.26
R3597 vss.n5398 vss.n5321 1118.26
R3598 vss.n5404 vss.n5321 1118.26
R3599 vss.n5404 vss.n5318 1118.26
R3600 vss.n5418 vss.n5318 1118.26
R3601 vss.n5418 vss.n5319 1118.26
R3602 vss.n5414 vss.n5319 1118.26
R3603 vss.n4151 vss.n4150 1118.26
R3604 vss.n4152 vss.n4151 1118.26
R3605 vss.n4152 vss.n4131 1118.26
R3606 vss.n4170 vss.n4131 1118.26
R3607 vss.n4170 vss.n4132 1118.26
R3608 vss.n4162 vss.n4132 1118.26
R3609 vss.n4148 vss.n4139 1118.26
R3610 vss.n4154 vss.n4139 1118.26
R3611 vss.n4154 vss.n4136 1118.26
R3612 vss.n4168 vss.n4136 1118.26
R3613 vss.n4168 vss.n4137 1118.26
R3614 vss.n4164 vss.n4137 1118.26
R3615 vss.n4242 vss.n4241 1118.26
R3616 vss.n4243 vss.n4242 1118.26
R3617 vss.n4243 vss.n4222 1118.26
R3618 vss.n4260 vss.n4222 1118.26
R3619 vss.n4260 vss.n4223 1118.26
R3620 vss.n4250 vss.n4223 1118.26
R3621 vss.n4239 vss.n4230 1118.26
R3622 vss.n4245 vss.n4230 1118.26
R3623 vss.n4245 vss.n4227 1118.26
R3624 vss.n4258 vss.n4227 1118.26
R3625 vss.n4258 vss.n4228 1118.26
R3626 vss.n4254 vss.n4228 1118.26
R3627 vss.n4974 vss.n4973 1118.26
R3628 vss.n4975 vss.n4974 1118.26
R3629 vss.n4975 vss.n4954 1118.26
R3630 vss.n4993 vss.n4954 1118.26
R3631 vss.n4993 vss.n4955 1118.26
R3632 vss.n4985 vss.n4955 1118.26
R3633 vss.n4971 vss.n4962 1118.26
R3634 vss.n4977 vss.n4962 1118.26
R3635 vss.n4977 vss.n4959 1118.26
R3636 vss.n4991 vss.n4959 1118.26
R3637 vss.n4991 vss.n4960 1118.26
R3638 vss.n4987 vss.n4960 1118.26
R3639 vss.n4105 vss.n4104 1118.26
R3640 vss.n4106 vss.n4105 1118.26
R3641 vss.n4106 vss.n4085 1118.26
R3642 vss.n4124 vss.n4085 1118.26
R3643 vss.n4124 vss.n4086 1118.26
R3644 vss.n4116 vss.n4086 1118.26
R3645 vss.n4102 vss.n4093 1118.26
R3646 vss.n4108 vss.n4093 1118.26
R3647 vss.n4108 vss.n4090 1118.26
R3648 vss.n4122 vss.n4090 1118.26
R3649 vss.n4122 vss.n4091 1118.26
R3650 vss.n4118 vss.n4091 1118.26
R3651 vss.n4926 vss.n4925 1118.26
R3652 vss.n4927 vss.n4926 1118.26
R3653 vss.n4927 vss.n4268 1118.26
R3654 vss.n4945 vss.n4268 1118.26
R3655 vss.n4945 vss.n4269 1118.26
R3656 vss.n4937 vss.n4269 1118.26
R3657 vss.n4923 vss.n4276 1118.26
R3658 vss.n4929 vss.n4276 1118.26
R3659 vss.n4929 vss.n4273 1118.26
R3660 vss.n4943 vss.n4273 1118.26
R3661 vss.n4943 vss.n4274 1118.26
R3662 vss.n4939 vss.n4274 1118.26
R3663 vss.n5189 vss.n5188 1118.26
R3664 vss.n5190 vss.n5189 1118.26
R3665 vss.n5190 vss.n5101 1118.26
R3666 vss.n5208 vss.n5101 1118.26
R3667 vss.n5208 vss.n5102 1118.26
R3668 vss.n5200 vss.n5102 1118.26
R3669 vss.n5186 vss.n5109 1118.26
R3670 vss.n5192 vss.n5109 1118.26
R3671 vss.n5192 vss.n5106 1118.26
R3672 vss.n5206 vss.n5106 1118.26
R3673 vss.n5206 vss.n5107 1118.26
R3674 vss.n5202 vss.n5107 1118.26
R3675 vss.n3364 vss.n3363 1118.26
R3676 vss.n3365 vss.n3364 1118.26
R3677 vss.n3365 vss.n3344 1118.26
R3678 vss.n3383 vss.n3344 1118.26
R3679 vss.n3383 vss.n3345 1118.26
R3680 vss.n3375 vss.n3345 1118.26
R3681 vss.n3361 vss.n3352 1118.26
R3682 vss.n3367 vss.n3352 1118.26
R3683 vss.n3367 vss.n3349 1118.26
R3684 vss.n3381 vss.n3349 1118.26
R3685 vss.n3381 vss.n3350 1118.26
R3686 vss.n3377 vss.n3350 1118.26
R3687 vss.n3411 vss.n3410 1118.26
R3688 vss.n3412 vss.n3411 1118.26
R3689 vss.n3412 vss.n3391 1118.26
R3690 vss.n3430 vss.n3391 1118.26
R3691 vss.n3430 vss.n3392 1118.26
R3692 vss.n3422 vss.n3392 1118.26
R3693 vss.n3408 vss.n3399 1118.26
R3694 vss.n3414 vss.n3399 1118.26
R3695 vss.n3414 vss.n3396 1118.26
R3696 vss.n3428 vss.n3396 1118.26
R3697 vss.n3428 vss.n3397 1118.26
R3698 vss.n3424 vss.n3397 1118.26
R3699 vss.n3509 vss.n3501 1118.26
R3700 vss.n3517 vss.n3501 1118.26
R3701 vss.n3517 vss.n3497 1118.26
R3702 vss.n3522 vss.n3497 1118.26
R3703 vss.n3524 vss.n3522 1118.26
R3704 vss.n3524 vss.n3489 1118.26
R3705 vss.n3511 vss.n3503 1118.26
R3706 vss.n3515 vss.n3503 1118.26
R3707 vss.n3515 vss.n3494 1118.26
R3708 vss.n3528 vss.n3494 1118.26
R3709 vss.n3528 vss.n3495 1118.26
R3710 vss.n3495 vss.n3490 1118.26
R3711 vss.n6473 vss.n6472 1118.26
R3712 vss.n6474 vss.n6473 1118.26
R3713 vss.n6474 vss.n6385 1118.26
R3714 vss.n6492 vss.n6385 1118.26
R3715 vss.n6492 vss.n6386 1118.26
R3716 vss.n6484 vss.n6386 1118.26
R3717 vss.n6470 vss.n6393 1118.26
R3718 vss.n6476 vss.n6393 1118.26
R3719 vss.n6476 vss.n6390 1118.26
R3720 vss.n6490 vss.n6390 1118.26
R3721 vss.n6490 vss.n6391 1118.26
R3722 vss.n6486 vss.n6391 1118.26
R3723 vss.n4424 vss.n4423 1118.26
R3724 vss.n4425 vss.n4424 1118.26
R3725 vss.n4425 vss.n4404 1118.26
R3726 vss.n4443 vss.n4404 1118.26
R3727 vss.n4443 vss.n4405 1118.26
R3728 vss.n4435 vss.n4405 1118.26
R3729 vss.n4421 vss.n4412 1118.26
R3730 vss.n4427 vss.n4412 1118.26
R3731 vss.n4427 vss.n4409 1118.26
R3732 vss.n4441 vss.n4409 1118.26
R3733 vss.n4441 vss.n4410 1118.26
R3734 vss.n4437 vss.n4410 1118.26
R3735 vss.n4764 vss.n4754 1118.26
R3736 vss.n4791 vss.n4764 1118.26
R3737 vss.n4791 vss.n4765 1118.26
R3738 vss.n4786 vss.n4765 1118.26
R3739 vss.n4786 vss.n4770 1118.26
R3740 vss.n4778 vss.n4770 1118.26
R3741 vss.n4759 vss.n4755 1118.26
R3742 vss.n4793 vss.n4759 1118.26
R3743 vss.n4793 vss.n4760 1118.26
R3744 vss.n4784 vss.n4760 1118.26
R3745 vss.n4784 vss.n4772 1118.26
R3746 vss.n4780 vss.n4772 1118.26
R3747 vss.n15009 vss.n14991 1118.26
R3748 vss.n15009 vss.n15008 1118.26
R3749 vss.n15008 vss.n14993 1118.26
R3750 vss.n14995 vss.n14993 1118.26
R3751 vss.n14996 vss.n14995 1118.26
R3752 vss.n15006 vss.n14996 1118.26
R3753 vss.n15014 vss.n14987 1118.26
R3754 vss.n14987 vss.n14984 1118.26
R3755 vss.n14984 vss.n14981 1118.26
R3756 vss.n15016 vss.n14981 1118.26
R3757 vss.n15016 vss.n14982 1118.26
R3758 vss.n14985 vss.n14982 1118.26
R3759 vss.n15520 vss.n15512 1118.26
R3760 vss.n15528 vss.n15512 1118.26
R3761 vss.n15528 vss.n15506 1118.26
R3762 vss.n15533 vss.n15506 1118.26
R3763 vss.n15533 vss.n15508 1118.26
R3764 vss.n15508 vss.n384 1118.26
R3765 vss.n15522 vss.n15514 1118.26
R3766 vss.n15526 vss.n15514 1118.26
R3767 vss.n15526 vss.n15502 1118.26
R3768 vss.n15535 vss.n15502 1118.26
R3769 vss.n15535 vss.n15503 1118.26
R3770 vss.n15503 vss.n385 1118.26
R3771 vss.n14855 vss.n14851 1118.26
R3772 vss.n14859 vss.n14855 1118.26
R3773 vss.n14859 vss.n397 1118.26
R3774 vss.n15494 vss.n397 1118.26
R3775 vss.n15494 vss.n398 1118.26
R3776 vss.n15490 vss.n398 1118.26
R3777 vss.n14856 vss.n14852 1118.26
R3778 vss.n14857 vss.n14856 1118.26
R3779 vss.n14857 vss.n392 1118.26
R3780 vss.n15496 vss.n392 1118.26
R3781 vss.n15496 vss.n393 1118.26
R3782 vss.n15488 vss.n393 1118.26
R3783 vss.n14953 vss.n14946 1118.26
R3784 vss.n14953 vss.n14947 1118.26
R3785 vss.n14949 vss.n14947 1118.26
R3786 vss.n14965 vss.n14949 1118.26
R3787 vss.n14965 vss.n14944 1118.26
R3788 vss.n14967 vss.n14944 1118.26
R3789 vss.n14957 vss.n14956 1118.26
R3790 vss.n14956 vss.n14955 1118.26
R3791 vss.n14955 vss.n14939 1118.26
R3792 vss.n14973 vss.n14939 1118.26
R3793 vss.n14973 vss.n14972 1118.26
R3794 vss.n14972 vss.n14971 1118.26
R3795 vss.n1061 vss.n1052 1118.26
R3796 vss.n1067 vss.n1052 1118.26
R3797 vss.n1067 vss.n1049 1118.26
R3798 vss.n15044 vss.n1049 1118.26
R3799 vss.n15044 vss.n1050 1118.26
R3800 vss.n15040 vss.n1050 1118.26
R3801 vss.n1064 vss.n1063 1118.26
R3802 vss.n1065 vss.n1064 1118.26
R3803 vss.n1065 vss.n1044 1118.26
R3804 vss.n15046 vss.n1044 1118.26
R3805 vss.n15046 vss.n1045 1118.26
R3806 vss.n15038 vss.n1045 1118.26
R3807 vss.n15146 vss.n977 1118.26
R3808 vss.n15152 vss.n977 1118.26
R3809 vss.n15152 vss.n974 1118.26
R3810 vss.n15167 vss.n974 1118.26
R3811 vss.n15167 vss.n975 1118.26
R3812 vss.n15163 vss.n975 1118.26
R3813 vss.n15149 vss.n15148 1118.26
R3814 vss.n15150 vss.n15149 1118.26
R3815 vss.n15150 vss.n969 1118.26
R3816 vss.n15169 vss.n969 1118.26
R3817 vss.n15169 vss.n970 1118.26
R3818 vss.n15160 vss.n970 1118.26
R3819 vss.n14908 vss.n14899 1118.26
R3820 vss.n14916 vss.n14899 1118.26
R3821 vss.n14916 vss.n14896 1118.26
R3822 vss.n14930 vss.n14896 1118.26
R3823 vss.n14930 vss.n14897 1118.26
R3824 vss.n14926 vss.n14897 1118.26
R3825 vss.n14913 vss.n14912 1118.26
R3826 vss.n14914 vss.n14913 1118.26
R3827 vss.n14914 vss.n14891 1118.26
R3828 vss.n14932 vss.n14891 1118.26
R3829 vss.n14932 vss.n14892 1118.26
R3830 vss.n14924 vss.n14892 1118.26
R3831 vss.n4580 vss.n4570 1118.26
R3832 vss.n4586 vss.n4570 1118.26
R3833 vss.n4586 vss.n4567 1118.26
R3834 vss.n4601 vss.n4567 1118.26
R3835 vss.n4601 vss.n4568 1118.26
R3836 vss.n4597 vss.n4568 1118.26
R3837 vss.n4583 vss.n4582 1118.26
R3838 vss.n4584 vss.n4583 1118.26
R3839 vss.n4584 vss.n4562 1118.26
R3840 vss.n4603 vss.n4562 1118.26
R3841 vss.n4603 vss.n4563 1118.26
R3842 vss.n4594 vss.n4563 1118.26
R3843 vss.n4672 vss.n4666 1118.26
R3844 vss.n4682 vss.n4666 1118.26
R3845 vss.n4682 vss.n4663 1118.26
R3846 vss.n4696 vss.n4663 1118.26
R3847 vss.n4696 vss.n4664 1118.26
R3848 vss.n4692 vss.n4664 1118.26
R3849 vss.n4679 vss.n4678 1118.26
R3850 vss.n4680 vss.n4679 1118.26
R3851 vss.n4680 vss.n4658 1118.26
R3852 vss.n4698 vss.n4658 1118.26
R3853 vss.n4698 vss.n4659 1118.26
R3854 vss.n4690 vss.n4659 1118.26
R3855 vss.n4627 vss.n4618 1118.26
R3856 vss.n4633 vss.n4618 1118.26
R3857 vss.n4633 vss.n4615 1118.26
R3858 vss.n4648 vss.n4615 1118.26
R3859 vss.n4648 vss.n4616 1118.26
R3860 vss.n4644 vss.n4616 1118.26
R3861 vss.n4630 vss.n4629 1118.26
R3862 vss.n4631 vss.n4630 1118.26
R3863 vss.n4631 vss.n4610 1118.26
R3864 vss.n4650 vss.n4610 1118.26
R3865 vss.n4650 vss.n4611 1118.26
R3866 vss.n4641 vss.n4611 1118.26
R3867 vss.n7236 vss.n7234 1118.26
R3868 vss.n7262 vss.n7234 1118.26
R3869 vss.n7262 vss.n7235 1118.26
R3870 vss.n7258 vss.n7235 1118.26
R3871 vss.n7258 vss.n7242 1118.26
R3872 vss.n7250 vss.n7242 1118.26
R3873 vss.n7268 vss.n7226 1118.26
R3874 vss.n7264 vss.n7226 1118.26
R3875 vss.n7264 vss.n7230 1118.26
R3876 vss.n7256 vss.n7230 1118.26
R3877 vss.n7256 vss.n7244 1118.26
R3878 vss.n7252 vss.n7244 1118.26
R3879 vss.n523 vss.n514 1118.26
R3880 vss.n529 vss.n514 1118.26
R3881 vss.n529 vss.n511 1118.26
R3882 vss.n15438 vss.n511 1118.26
R3883 vss.n15438 vss.n512 1118.26
R3884 vss.n15434 vss.n512 1118.26
R3885 vss.n526 vss.n525 1118.26
R3886 vss.n527 vss.n526 1118.26
R3887 vss.n527 vss.n506 1118.26
R3888 vss.n15440 vss.n506 1118.26
R3889 vss.n15440 vss.n507 1118.26
R3890 vss.n15432 vss.n507 1118.26
R3891 vss.n7321 vss.n7312 1118.26
R3892 vss.n7327 vss.n7312 1118.26
R3893 vss.n7327 vss.n7309 1118.26
R3894 vss.n7341 vss.n7309 1118.26
R3895 vss.n7341 vss.n7310 1118.26
R3896 vss.n7337 vss.n7310 1118.26
R3897 vss.n7324 vss.n7323 1118.26
R3898 vss.n7325 vss.n7324 1118.26
R3899 vss.n7325 vss.n7304 1118.26
R3900 vss.n7343 vss.n7304 1118.26
R3901 vss.n7343 vss.n7305 1118.26
R3902 vss.n7335 vss.n7305 1118.26
R3903 vss.n3081 vss.n3075 1118.26
R3904 vss.n3091 vss.n3075 1118.26
R3905 vss.n3091 vss.n3072 1118.26
R3906 vss.n3105 vss.n3072 1118.26
R3907 vss.n3105 vss.n3073 1118.26
R3908 vss.n3101 vss.n3073 1118.26
R3909 vss.n3088 vss.n3087 1118.26
R3910 vss.n3089 vss.n3088 1118.26
R3911 vss.n3089 vss.n3067 1118.26
R3912 vss.n3107 vss.n3067 1118.26
R3913 vss.n3107 vss.n3068 1118.26
R3914 vss.n3099 vss.n3068 1118.26
R3915 vss.n7357 vss.n3060 1118.26
R3916 vss.n7384 vss.n7357 1118.26
R3917 vss.n7384 vss.n7358 1118.26
R3918 vss.n7380 vss.n7358 1118.26
R3919 vss.n7380 vss.n7363 1118.26
R3920 vss.n7370 vss.n7363 1118.26
R3921 vss.n7352 vss.n3061 1118.26
R3922 vss.n7386 vss.n7352 1118.26
R3923 vss.n7386 vss.n7353 1118.26
R3924 vss.n7378 vss.n7353 1118.26
R3925 vss.n7378 vss.n7365 1118.26
R3926 vss.n7368 vss.n7365 1118.26
R3927 vss.n7406 vss.n7404 1118.26
R3928 vss.n7432 vss.n7404 1118.26
R3929 vss.n7432 vss.n7405 1118.26
R3930 vss.n7428 vss.n7405 1118.26
R3931 vss.n7428 vss.n7412 1118.26
R3932 vss.n7420 vss.n7412 1118.26
R3933 vss.n7438 vss.n7396 1118.26
R3934 vss.n7434 vss.n7396 1118.26
R3935 vss.n7434 vss.n7400 1118.26
R3936 vss.n7426 vss.n7400 1118.26
R3937 vss.n7426 vss.n7414 1118.26
R3938 vss.n7422 vss.n7414 1118.26
R3939 vss.n728 vss.n719 1118.26
R3940 vss.n734 vss.n719 1118.26
R3941 vss.n734 vss.n716 1118.26
R3942 vss.n15365 vss.n716 1118.26
R3943 vss.n15365 vss.n717 1118.26
R3944 vss.n15361 vss.n717 1118.26
R3945 vss.n731 vss.n730 1118.26
R3946 vss.n732 vss.n731 1118.26
R3947 vss.n732 vss.n711 1118.26
R3948 vss.n15367 vss.n711 1118.26
R3949 vss.n15367 vss.n712 1118.26
R3950 vss.n15359 vss.n712 1118.26
R3951 vss.n781 vss.n772 1118.26
R3952 vss.n787 vss.n772 1118.26
R3953 vss.n787 vss.n769 1118.26
R3954 vss.n15288 vss.n769 1118.26
R3955 vss.n15288 vss.n770 1118.26
R3956 vss.n15284 vss.n770 1118.26
R3957 vss.n784 vss.n783 1118.26
R3958 vss.n785 vss.n784 1118.26
R3959 vss.n785 vss.n764 1118.26
R3960 vss.n15290 vss.n764 1118.26
R3961 vss.n15290 vss.n765 1118.26
R3962 vss.n15282 vss.n765 1118.26
R3963 vss.n15108 vss.n15105 1118.26
R3964 vss.n15134 vss.n15105 1118.26
R3965 vss.n15134 vss.n15106 1118.26
R3966 vss.n15130 vss.n15106 1118.26
R3967 vss.n15130 vss.n15114 1118.26
R3968 vss.n15122 vss.n15114 1118.26
R3969 vss.n15140 vss.n15097 1118.26
R3970 vss.n15136 vss.n15097 1118.26
R3971 vss.n15136 vss.n15101 1118.26
R3972 vss.n15128 vss.n15101 1118.26
R3973 vss.n15128 vss.n15116 1118.26
R3974 vss.n15124 vss.n15116 1118.26
R3975 vss.n15195 vss.n15186 1118.26
R3976 vss.n15201 vss.n15186 1118.26
R3977 vss.n15201 vss.n15183 1118.26
R3978 vss.n15215 vss.n15183 1118.26
R3979 vss.n15215 vss.n15184 1118.26
R3980 vss.n15211 vss.n15184 1118.26
R3981 vss.n15198 vss.n15197 1118.26
R3982 vss.n15199 vss.n15198 1118.26
R3983 vss.n15199 vss.n15178 1118.26
R3984 vss.n15217 vss.n15178 1118.26
R3985 vss.n15217 vss.n15179 1118.26
R3986 vss.n15209 vss.n15179 1118.26
R3987 vss.n938 vss.n929 1118.26
R3988 vss.n944 vss.n929 1118.26
R3989 vss.n944 vss.n926 1118.26
R3990 vss.n959 vss.n926 1118.26
R3991 vss.n959 vss.n927 1118.26
R3992 vss.n955 vss.n927 1118.26
R3993 vss.n941 vss.n940 1118.26
R3994 vss.n942 vss.n941 1118.26
R3995 vss.n942 vss.n921 1118.26
R3996 vss.n961 vss.n921 1118.26
R3997 vss.n961 vss.n922 1118.26
R3998 vss.n953 vss.n922 1118.26
R3999 vss.n829 vss.n821 1118.26
R4000 vss.n837 vss.n821 1118.26
R4001 vss.n837 vss.n815 1118.26
R4002 vss.n842 vss.n815 1118.26
R4003 vss.n842 vss.n817 1118.26
R4004 vss.n817 vss.n806 1118.26
R4005 vss.n831 vss.n823 1118.26
R4006 vss.n835 vss.n823 1118.26
R4007 vss.n835 vss.n811 1118.26
R4008 vss.n844 vss.n811 1118.26
R4009 vss.n844 vss.n812 1118.26
R4010 vss.n812 vss.n807 1118.26
R4011 vss.n7451 vss.n7442 1118.26
R4012 vss.n7479 vss.n7451 1118.26
R4013 vss.n7479 vss.n7452 1118.26
R4014 vss.n7475 vss.n7452 1118.26
R4015 vss.n7475 vss.n7458 1118.26
R4016 vss.n7466 vss.n7458 1118.26
R4017 vss.n7485 vss.n7443 1118.26
R4018 vss.n7481 vss.n7443 1118.26
R4019 vss.n7481 vss.n7448 1118.26
R4020 vss.n7473 vss.n7448 1118.26
R4021 vss.n7473 vss.n7460 1118.26
R4022 vss.n7469 vss.n7460 1118.26
R4023 vss.n15315 vss.n15306 1118.26
R4024 vss.n15321 vss.n15306 1118.26
R4025 vss.n15321 vss.n15303 1118.26
R4026 vss.n15336 vss.n15303 1118.26
R4027 vss.n15336 vss.n15304 1118.26
R4028 vss.n15332 vss.n15304 1118.26
R4029 vss.n15318 vss.n15317 1118.26
R4030 vss.n15319 vss.n15318 1118.26
R4031 vss.n15319 vss.n15298 1118.26
R4032 vss.n15338 vss.n15298 1118.26
R4033 vss.n15338 vss.n15299 1118.26
R4034 vss.n15330 vss.n15299 1118.26
R4035 vss.n681 vss.n672 1118.26
R4036 vss.n687 vss.n672 1118.26
R4037 vss.n687 vss.n669 1118.26
R4038 vss.n702 vss.n669 1118.26
R4039 vss.n702 vss.n670 1118.26
R4040 vss.n698 vss.n670 1118.26
R4041 vss.n684 vss.n683 1118.26
R4042 vss.n685 vss.n684 1118.26
R4043 vss.n685 vss.n664 1118.26
R4044 vss.n704 vss.n664 1118.26
R4045 vss.n704 vss.n665 1118.26
R4046 vss.n696 vss.n665 1118.26
R4047 vss.n7274 vss.n3121 1118.26
R4048 vss.n7280 vss.n3121 1118.26
R4049 vss.n7280 vss.n3118 1118.26
R4050 vss.n7295 vss.n3118 1118.26
R4051 vss.n7295 vss.n3119 1118.26
R4052 vss.n7291 vss.n3119 1118.26
R4053 vss.n7277 vss.n7276 1118.26
R4054 vss.n7278 vss.n7277 1118.26
R4055 vss.n7278 vss.n3113 1118.26
R4056 vss.n7297 vss.n3113 1118.26
R4057 vss.n7297 vss.n3114 1118.26
R4058 vss.n7288 vss.n3114 1118.26
R4059 vss.n572 vss.n564 1118.26
R4060 vss.n580 vss.n564 1118.26
R4061 vss.n580 vss.n558 1118.26
R4062 vss.n585 vss.n558 1118.26
R4063 vss.n585 vss.n560 1118.26
R4064 vss.n560 vss.n548 1118.26
R4065 vss.n574 vss.n566 1118.26
R4066 vss.n578 vss.n566 1118.26
R4067 vss.n578 vss.n554 1118.26
R4068 vss.n587 vss.n554 1118.26
R4069 vss.n587 vss.n555 1118.26
R4070 vss.n555 vss.n549 1118.26
R4071 vss.n473 vss.n464 1118.26
R4072 vss.n479 vss.n464 1118.26
R4073 vss.n479 vss.n461 1118.26
R4074 vss.n494 vss.n461 1118.26
R4075 vss.n494 vss.n462 1118.26
R4076 vss.n490 vss.n462 1118.26
R4077 vss.n476 vss.n475 1118.26
R4078 vss.n477 vss.n476 1118.26
R4079 vss.n477 vss.n456 1118.26
R4080 vss.n496 vss.n456 1118.26
R4081 vss.n496 vss.n457 1118.26
R4082 vss.n488 vss.n457 1118.26
R4083 vss.n4723 vss.n4715 1118.26
R4084 vss.n4731 vss.n4715 1118.26
R4085 vss.n4731 vss.n4709 1118.26
R4086 vss.n4736 vss.n4709 1118.26
R4087 vss.n4736 vss.n4711 1118.26
R4088 vss.n4711 vss.n4555 1118.26
R4089 vss.n4725 vss.n4717 1118.26
R4090 vss.n4729 vss.n4717 1118.26
R4091 vss.n4729 vss.n4705 1118.26
R4092 vss.n4738 vss.n4705 1118.26
R4093 vss.n4738 vss.n4706 1118.26
R4094 vss.n4706 vss.n4556 1118.26
R4095 vss.n4338 vss.n4330 1118.26
R4096 vss.n4346 vss.n4330 1118.26
R4097 vss.n4346 vss.n4324 1118.26
R4098 vss.n4351 vss.n4324 1118.26
R4099 vss.n4351 vss.n4326 1118.26
R4100 vss.n4326 vss.n4315 1118.26
R4101 vss.n4340 vss.n4332 1118.26
R4102 vss.n4344 vss.n4332 1118.26
R4103 vss.n4344 vss.n4320 1118.26
R4104 vss.n4353 vss.n4320 1118.26
R4105 vss.n4353 vss.n4321 1118.26
R4106 vss.n4321 vss.n4316 1118.26
R4107 vss.n6765 vss.n6756 1118.26
R4108 vss.n6771 vss.n6756 1118.26
R4109 vss.n6771 vss.n6753 1118.26
R4110 vss.n6785 vss.n6753 1118.26
R4111 vss.n6785 vss.n6754 1118.26
R4112 vss.n6781 vss.n6754 1118.26
R4113 vss.n6768 vss.n6767 1118.26
R4114 vss.n6769 vss.n6768 1118.26
R4115 vss.n6769 vss.n6748 1118.26
R4116 vss.n6787 vss.n6748 1118.26
R4117 vss.n6787 vss.n6749 1118.26
R4118 vss.n6779 vss.n6749 1118.26
R4119 vss.n6854 vss.n6853 1118.26
R4120 vss.n6855 vss.n6854 1118.26
R4121 vss.n6855 vss.n6834 1118.26
R4122 vss.n6873 vss.n6834 1118.26
R4123 vss.n6873 vss.n6835 1118.26
R4124 vss.n6865 vss.n6835 1118.26
R4125 vss.n6851 vss.n6842 1118.26
R4126 vss.n6857 vss.n6842 1118.26
R4127 vss.n6857 vss.n6839 1118.26
R4128 vss.n6871 vss.n6839 1118.26
R4129 vss.n6871 vss.n6840 1118.26
R4130 vss.n6867 vss.n6840 1118.26
R4131 vss.n6812 vss.n6807 1118.26
R4132 vss.n6818 vss.n6812 1118.26
R4133 vss.n6818 vss.n3142 1118.26
R4134 vss.n7213 vss.n3142 1118.26
R4135 vss.n7214 vss.n7213 1118.26
R4136 vss.n7216 vss.n7214 1118.26
R4137 vss.n6815 vss.n6806 1118.26
R4138 vss.n6816 vss.n6815 1118.26
R4139 vss.n6816 vss.n3145 1118.26
R4140 vss.n7210 vss.n3145 1118.26
R4141 vss.n7210 vss.n3136 1118.26
R4142 vss.n7220 vss.n3136 1118.26
R4143 vss.n6885 vss.n6883 1118.26
R4144 vss.n6911 vss.n6883 1118.26
R4145 vss.n6911 vss.n6884 1118.26
R4146 vss.n6907 vss.n6884 1118.26
R4147 vss.n6907 vss.n6891 1118.26
R4148 vss.n6898 vss.n6891 1118.26
R4149 vss.n6917 vss.n6828 1118.26
R4150 vss.n6913 vss.n6828 1118.26
R4151 vss.n6913 vss.n6880 1118.26
R4152 vss.n6892 vss.n6880 1118.26
R4153 vss.n6894 vss.n6892 1118.26
R4154 vss.n6900 vss.n6894 1118.26
R4155 vss.n7088 vss.n7086 1118.26
R4156 vss.n7115 vss.n7086 1118.26
R4157 vss.n7115 vss.n7087 1118.26
R4158 vss.n7111 vss.n7087 1118.26
R4159 vss.n7111 vss.n7094 1118.26
R4160 vss.n7101 vss.n7094 1118.26
R4161 vss.n7121 vss.n7080 1118.26
R4162 vss.n7117 vss.n7080 1118.26
R4163 vss.n7117 vss.n7083 1118.26
R4164 vss.n7095 vss.n7083 1118.26
R4165 vss.n7097 vss.n7095 1118.26
R4166 vss.n7099 vss.n7097 1118.26
R4167 vss.n7969 vss.n7961 1118.26
R4168 vss.n7965 vss.n7961 1118.26
R4169 vss.n7965 vss.n2464 1118.26
R4170 vss.n7978 vss.n2464 1118.26
R4171 vss.n7978 vss.n2462 1118.26
R4172 vss.n7982 vss.n2462 1118.26
R4173 vss.n7972 vss.n7971 1118.26
R4174 vss.n7973 vss.n7972 1118.26
R4175 vss.n7974 vss.n7973 1118.26
R4176 vss.n7974 vss.n2454 1118.26
R4177 vss.n2457 vss.n2454 1118.26
R4178 vss.n7986 vss.n2457 1118.26
R4179 vss.n2996 vss.n2987 1118.26
R4180 vss.n3003 vss.n2987 1118.26
R4181 vss.n3003 vss.n2984 1118.26
R4182 vss.n7496 vss.n2984 1118.26
R4183 vss.n7496 vss.n2985 1118.26
R4184 vss.n7492 vss.n2985 1118.26
R4185 vss.n3000 vss.n2999 1118.26
R4186 vss.n3001 vss.n3000 1118.26
R4187 vss.n3001 vss.n2979 1118.26
R4188 vss.n7498 vss.n2979 1118.26
R4189 vss.n7498 vss.n2980 1118.26
R4190 vss.n3011 vss.n2980 1118.26
R4191 vss.n7690 vss.n7681 1118.26
R4192 vss.n7697 vss.n7681 1118.26
R4193 vss.n7697 vss.n7678 1118.26
R4194 vss.n7712 vss.n7678 1118.26
R4195 vss.n7712 vss.n7679 1118.26
R4196 vss.n7708 vss.n7679 1118.26
R4197 vss.n7694 vss.n7693 1118.26
R4198 vss.n7695 vss.n7694 1118.26
R4199 vss.n7695 vss.n7673 1118.26
R4200 vss.n7714 vss.n7673 1118.26
R4201 vss.n7714 vss.n7674 1118.26
R4202 vss.n7705 vss.n7674 1118.26
R4203 vss.n2908 vss.n2900 1118.26
R4204 vss.n2904 vss.n2900 1118.26
R4205 vss.n2904 vss.n2894 1118.26
R4206 vss.n2917 vss.n2894 1118.26
R4207 vss.n2917 vss.n2892 1118.26
R4208 vss.n2921 vss.n2892 1118.26
R4209 vss.n2911 vss.n2910 1118.26
R4210 vss.n2912 vss.n2911 1118.26
R4211 vss.n2913 vss.n2912 1118.26
R4212 vss.n2913 vss.n2885 1118.26
R4213 vss.n2888 vss.n2885 1118.26
R4214 vss.n2925 vss.n2888 1118.26
R4215 vss.n7739 vss.n7730 1118.26
R4216 vss.n7746 vss.n7730 1118.26
R4217 vss.n7746 vss.n7727 1118.26
R4218 vss.n7760 vss.n7727 1118.26
R4219 vss.n7760 vss.n7728 1118.26
R4220 vss.n7756 vss.n7728 1118.26
R4221 vss.n7743 vss.n7742 1118.26
R4222 vss.n7744 vss.n7743 1118.26
R4223 vss.n7744 vss.n7722 1118.26
R4224 vss.n7762 vss.n7722 1118.26
R4225 vss.n7762 vss.n7723 1118.26
R4226 vss.n7754 vss.n7723 1118.26
R4227 vss.n7885 vss.n7876 1118.26
R4228 vss.n7892 vss.n7876 1118.26
R4229 vss.n7892 vss.n7873 1118.26
R4230 vss.n7907 vss.n7873 1118.26
R4231 vss.n7907 vss.n7874 1118.26
R4232 vss.n7903 vss.n7874 1118.26
R4233 vss.n7889 vss.n7888 1118.26
R4234 vss.n7890 vss.n7889 1118.26
R4235 vss.n7890 vss.n7868 1118.26
R4236 vss.n7909 vss.n7868 1118.26
R4237 vss.n7909 vss.n7869 1118.26
R4238 vss.n7900 vss.n7869 1118.26
R4239 vss.n2649 vss.n2645 1118.26
R4240 vss.n7919 vss.n2649 1118.26
R4241 vss.n7919 vss.n2650 1118.26
R4242 vss.n2667 vss.n2650 1118.26
R4243 vss.n2667 vss.n2666 1118.26
R4244 vss.n2671 vss.n2666 1118.26
R4245 vss.n2653 vss.n2644 1118.26
R4246 vss.n2654 vss.n2653 1118.26
R4247 vss.n2656 vss.n2654 1118.26
R4248 vss.n2659 vss.n2656 1118.26
R4249 vss.n2662 vss.n2659 1118.26
R4250 vss.n2675 vss.n2662 1118.26
R4251 vss.n7938 vss.n7933 1118.26
R4252 vss.n7938 vss.n7937 1118.26
R4253 vss.n7937 vss.n1149 1118.26
R4254 vss.n14877 vss.n1149 1118.26
R4255 vss.n14877 vss.n1150 1118.26
R4256 vss.n14873 vss.n1150 1118.26
R4257 vss.n7943 vss.n7929 1118.26
R4258 vss.n7935 vss.n7929 1118.26
R4259 vss.n7935 vss.n1144 1118.26
R4260 vss.n14879 vss.n1144 1118.26
R4261 vss.n14879 vss.n1145 1118.26
R4262 vss.n1157 vss.n1145 1118.26
R4263 vss.n2620 vss.n2610 1118.26
R4264 vss.n2628 vss.n2610 1118.26
R4265 vss.n2629 vss.n2628 1118.26
R4266 vss.n2634 vss.n2629 1118.26
R4267 vss.n2634 vss.n2631 1118.26
R4268 vss.n2631 vss.n2599 1118.26
R4269 vss.n2622 vss.n2613 1118.26
R4270 vss.n2626 vss.n2613 1118.26
R4271 vss.n2626 vss.n2604 1118.26
R4272 vss.n2636 vss.n2604 1118.26
R4273 vss.n2636 vss.n2605 1118.26
R4274 vss.n2605 vss.n2600 1118.26
R4275 vss.n1908 vss.n1898 1118.26
R4276 vss.n1936 vss.n1908 1118.26
R4277 vss.n1936 vss.n1909 1118.26
R4278 vss.n1931 vss.n1909 1118.26
R4279 vss.n1931 vss.n1914 1118.26
R4280 vss.n1923 vss.n1914 1118.26
R4281 vss.n1903 vss.n1899 1118.26
R4282 vss.n1938 vss.n1903 1118.26
R4283 vss.n1938 vss.n1904 1118.26
R4284 vss.n1929 vss.n1904 1118.26
R4285 vss.n1929 vss.n1916 1118.26
R4286 vss.n1925 vss.n1916 1118.26
R4287 vss.n2861 vss.n2860 1118.26
R4288 vss.n2862 vss.n2861 1118.26
R4289 vss.n2862 vss.n2841 1118.26
R4290 vss.n2880 vss.n2841 1118.26
R4291 vss.n2880 vss.n2842 1118.26
R4292 vss.n2872 vss.n2842 1118.26
R4293 vss.n2858 vss.n2849 1118.26
R4294 vss.n2864 vss.n2849 1118.26
R4295 vss.n2864 vss.n2846 1118.26
R4296 vss.n2878 vss.n2846 1118.26
R4297 vss.n2878 vss.n2847 1118.26
R4298 vss.n2874 vss.n2847 1118.26
R4299 vss.n3033 vss.n3025 1118.26
R4300 vss.n3041 vss.n3025 1118.26
R4301 vss.n3041 vss.n3021 1118.26
R4302 vss.n3046 vss.n3021 1118.26
R4303 vss.n3048 vss.n3046 1118.26
R4304 vss.n3048 vss.n3013 1118.26
R4305 vss.n3035 vss.n3027 1118.26
R4306 vss.n3039 vss.n3027 1118.26
R4307 vss.n3039 vss.n3018 1118.26
R4308 vss.n3052 vss.n3018 1118.26
R4309 vss.n3052 vss.n3019 1118.26
R4310 vss.n3019 vss.n3014 1118.26
R4311 vss.n7645 vss.n7644 1118.26
R4312 vss.n7646 vss.n7645 1118.26
R4313 vss.n7646 vss.n7625 1118.26
R4314 vss.n7664 vss.n7625 1118.26
R4315 vss.n7664 vss.n7626 1118.26
R4316 vss.n7656 vss.n7626 1118.26
R4317 vss.n7642 vss.n7633 1118.26
R4318 vss.n7648 vss.n7633 1118.26
R4319 vss.n7648 vss.n7630 1118.26
R4320 vss.n7662 vss.n7630 1118.26
R4321 vss.n7662 vss.n7631 1118.26
R4322 vss.n7658 vss.n7631 1118.26
R4323 vss.n2815 vss.n2814 1118.26
R4324 vss.n2816 vss.n2815 1118.26
R4325 vss.n2816 vss.n2727 1118.26
R4326 vss.n2834 vss.n2727 1118.26
R4327 vss.n2834 vss.n2728 1118.26
R4328 vss.n2826 vss.n2728 1118.26
R4329 vss.n2812 vss.n2735 1118.26
R4330 vss.n2818 vss.n2735 1118.26
R4331 vss.n2818 vss.n2732 1118.26
R4332 vss.n2832 vss.n2732 1118.26
R4333 vss.n2832 vss.n2733 1118.26
R4334 vss.n2828 vss.n2733 1118.26
R4335 vss.n2953 vss.n2952 1118.26
R4336 vss.n2954 vss.n2953 1118.26
R4337 vss.n2954 vss.n2933 1118.26
R4338 vss.n2973 vss.n2933 1118.26
R4339 vss.n2973 vss.n2934 1118.26
R4340 vss.n2965 vss.n2934 1118.26
R4341 vss.n2950 vss.n2941 1118.26
R4342 vss.n2956 vss.n2941 1118.26
R4343 vss.n2956 vss.n2938 1118.26
R4344 vss.n2971 vss.n2938 1118.26
R4345 vss.n2971 vss.n2939 1118.26
R4346 vss.n2967 vss.n2939 1118.26
R4347 vss.n7042 vss.n7033 1118.26
R4348 vss.n7043 vss.n7042 1118.26
R4349 vss.n7045 vss.n7043 1118.26
R4350 vss.n7063 vss.n7045 1118.26
R4351 vss.n7063 vss.n7062 1118.26
R4352 vss.n7062 vss.n7049 1118.26
R4353 vss.n7038 vss.n7034 1118.26
R4354 vss.n7070 vss.n7038 1118.26
R4355 vss.n7070 vss.n7039 1118.26
R4356 vss.n7052 vss.n7039 1118.26
R4357 vss.n7052 vss.n7050 1118.26
R4358 vss.n7058 vss.n7050 1118.26
R4359 vss.n7009 vss.n6999 1118.26
R4360 vss.n7017 vss.n6999 1118.26
R4361 vss.n7018 vss.n7017 1118.26
R4362 vss.n7023 vss.n7018 1118.26
R4363 vss.n7023 vss.n7020 1118.26
R4364 vss.n7020 vss.n6988 1118.26
R4365 vss.n7011 vss.n7002 1118.26
R4366 vss.n7015 vss.n7002 1118.26
R4367 vss.n7015 vss.n6993 1118.26
R4368 vss.n7025 vss.n6993 1118.26
R4369 vss.n7025 vss.n6994 1118.26
R4370 vss.n6994 vss.n6989 1118.26
R4371 vss.n7148 vss.n7140 1118.26
R4372 vss.n7156 vss.n7140 1118.26
R4373 vss.n7156 vss.n7134 1118.26
R4374 vss.n7161 vss.n7134 1118.26
R4375 vss.n7161 vss.n7136 1118.26
R4376 vss.n7136 vss.n7125 1118.26
R4377 vss.n7150 vss.n7142 1118.26
R4378 vss.n7154 vss.n7142 1118.26
R4379 vss.n7154 vss.n7130 1118.26
R4380 vss.n7163 vss.n7130 1118.26
R4381 vss.n7163 vss.n7131 1118.26
R4382 vss.n7131 vss.n7126 1118.26
R4383 vss.n6964 vss.n6936 1118.26
R4384 vss.n6972 vss.n6936 1118.26
R4385 vss.n6972 vss.n6930 1118.26
R4386 vss.n6978 vss.n6930 1118.26
R4387 vss.n6978 vss.n6932 1118.26
R4388 vss.n6932 vss.n6921 1118.26
R4389 vss.n6966 vss.n6938 1118.26
R4390 vss.n6970 vss.n6938 1118.26
R4391 vss.n6970 vss.n6926 1118.26
R4392 vss.n6980 vss.n6926 1118.26
R4393 vss.n6980 vss.n6927 1118.26
R4394 vss.n6927 vss.n6922 1118.26
R4395 vss.n7597 vss.n7596 1118.26
R4396 vss.n7598 vss.n7597 1118.26
R4397 vss.n7598 vss.n7509 1118.26
R4398 vss.n7616 vss.n7509 1118.26
R4399 vss.n7616 vss.n7510 1118.26
R4400 vss.n7608 vss.n7510 1118.26
R4401 vss.n7594 vss.n7517 1118.26
R4402 vss.n7600 vss.n7517 1118.26
R4403 vss.n7600 vss.n7514 1118.26
R4404 vss.n7614 vss.n7514 1118.26
R4405 vss.n7614 vss.n7515 1118.26
R4406 vss.n7610 vss.n7515 1118.26
R4407 vss.n7792 vss.n7791 1118.26
R4408 vss.n7793 vss.n7792 1118.26
R4409 vss.n7793 vss.n7772 1118.26
R4410 vss.n7811 vss.n7772 1118.26
R4411 vss.n7811 vss.n7773 1118.26
R4412 vss.n7803 vss.n7773 1118.26
R4413 vss.n7789 vss.n7780 1118.26
R4414 vss.n7795 vss.n7780 1118.26
R4415 vss.n7795 vss.n7777 1118.26
R4416 vss.n7809 vss.n7777 1118.26
R4417 vss.n7809 vss.n7778 1118.26
R4418 vss.n7805 vss.n7778 1118.26
R4419 vss.n7840 vss.n7839 1118.26
R4420 vss.n7841 vss.n7840 1118.26
R4421 vss.n7841 vss.n7820 1118.26
R4422 vss.n7859 vss.n7820 1118.26
R4423 vss.n7859 vss.n7821 1118.26
R4424 vss.n7851 vss.n7821 1118.26
R4425 vss.n7837 vss.n7828 1118.26
R4426 vss.n7843 vss.n7828 1118.26
R4427 vss.n7843 vss.n7825 1118.26
R4428 vss.n7857 vss.n7825 1118.26
R4429 vss.n7857 vss.n7826 1118.26
R4430 vss.n7853 vss.n7826 1118.26
R4431 vss.n2702 vss.n2701 1118.26
R4432 vss.n2703 vss.n2702 1118.26
R4433 vss.n2703 vss.n2682 1118.26
R4434 vss.n2720 vss.n2682 1118.26
R4435 vss.n2720 vss.n2683 1118.26
R4436 vss.n2710 vss.n2683 1118.26
R4437 vss.n2699 vss.n2690 1118.26
R4438 vss.n2705 vss.n2690 1118.26
R4439 vss.n2705 vss.n2687 1118.26
R4440 vss.n2718 vss.n2687 1118.26
R4441 vss.n2718 vss.n2688 1118.26
R4442 vss.n2714 vss.n2688 1118.26
R4443 vss.n2576 vss.n2499 1118.26
R4444 vss.n2584 vss.n2499 1118.26
R4445 vss.n2584 vss.n2493 1118.26
R4446 vss.n2589 vss.n2493 1118.26
R4447 vss.n2589 vss.n2495 1118.26
R4448 vss.n2495 vss.n2484 1118.26
R4449 vss.n2578 vss.n2501 1118.26
R4450 vss.n2582 vss.n2501 1118.26
R4451 vss.n2582 vss.n2489 1118.26
R4452 vss.n2591 vss.n2489 1118.26
R4453 vss.n2591 vss.n2490 1118.26
R4454 vss.n2490 vss.n2485 1118.26
R4455 vss.n7184 vss.n7183 1118.26
R4456 vss.n7185 vss.n7184 1118.26
R4457 vss.n7185 vss.n3153 1118.26
R4458 vss.n7203 vss.n3153 1118.26
R4459 vss.n7203 vss.n3154 1118.26
R4460 vss.n7195 vss.n3154 1118.26
R4461 vss.n7181 vss.n3161 1118.26
R4462 vss.n7187 vss.n3161 1118.26
R4463 vss.n7187 vss.n3158 1118.26
R4464 vss.n7201 vss.n3158 1118.26
R4465 vss.n7201 vss.n3159 1118.26
R4466 vss.n7197 vss.n3159 1118.26
R4467 vss.n3200 vss.n3192 1118.26
R4468 vss.n3201 vss.n3200 1118.26
R4469 vss.n3201 vss.n3179 1118.26
R4470 vss.n6795 vss.n3179 1118.26
R4471 vss.n6795 vss.n3181 1118.26
R4472 vss.n3181 vss.n3170 1118.26
R4473 vss.n3197 vss.n3193 1118.26
R4474 vss.n3203 vss.n3197 1118.26
R4475 vss.n3203 vss.n3175 1118.26
R4476 vss.n6797 vss.n3175 1118.26
R4477 vss.n6797 vss.n3176 1118.26
R4478 vss.n3176 vss.n3171 1118.26
R4479 vss.n14314 vss.n14296 1118.26
R4480 vss.n14314 vss.n14313 1118.26
R4481 vss.n14313 vss.n14298 1118.26
R4482 vss.n14300 vss.n14298 1118.26
R4483 vss.n14301 vss.n14300 1118.26
R4484 vss.n14311 vss.n14301 1118.26
R4485 vss.n14319 vss.n14292 1118.26
R4486 vss.n14292 vss.n14289 1118.26
R4487 vss.n14289 vss.n14286 1118.26
R4488 vss.n14321 vss.n14286 1118.26
R4489 vss.n14321 vss.n14287 1118.26
R4490 vss.n14290 vss.n14287 1118.26
R4491 vss.n14825 vss.n14817 1118.26
R4492 vss.n14833 vss.n14817 1118.26
R4493 vss.n14833 vss.n14811 1118.26
R4494 vss.n14838 vss.n14811 1118.26
R4495 vss.n14838 vss.n14813 1118.26
R4496 vss.n14813 vss.n1163 1118.26
R4497 vss.n14827 vss.n14819 1118.26
R4498 vss.n14831 vss.n14819 1118.26
R4499 vss.n14831 vss.n14807 1118.26
R4500 vss.n14840 vss.n14807 1118.26
R4501 vss.n14840 vss.n14808 1118.26
R4502 vss.n14808 vss.n1164 1118.26
R4503 vss.n14161 vss.n14157 1118.26
R4504 vss.n14165 vss.n14161 1118.26
R4505 vss.n14165 vss.n1176 1118.26
R4506 vss.n14799 vss.n1176 1118.26
R4507 vss.n14799 vss.n1177 1118.26
R4508 vss.n14795 vss.n1177 1118.26
R4509 vss.n14162 vss.n14158 1118.26
R4510 vss.n14163 vss.n14162 1118.26
R4511 vss.n14163 vss.n1171 1118.26
R4512 vss.n14801 vss.n1171 1118.26
R4513 vss.n14801 vss.n1172 1118.26
R4514 vss.n14793 vss.n1172 1118.26
R4515 vss.n14258 vss.n14251 1118.26
R4516 vss.n14258 vss.n14252 1118.26
R4517 vss.n14254 vss.n14252 1118.26
R4518 vss.n14270 vss.n14254 1118.26
R4519 vss.n14270 vss.n14249 1118.26
R4520 vss.n14272 vss.n14249 1118.26
R4521 vss.n14262 vss.n14261 1118.26
R4522 vss.n14261 vss.n14260 1118.26
R4523 vss.n14260 vss.n14244 1118.26
R4524 vss.n14278 vss.n14244 1118.26
R4525 vss.n14278 vss.n14277 1118.26
R4526 vss.n14277 vss.n14276 1118.26
R4527 vss.n1840 vss.n1831 1118.26
R4528 vss.n1846 vss.n1831 1118.26
R4529 vss.n1846 vss.n1828 1118.26
R4530 vss.n14349 vss.n1828 1118.26
R4531 vss.n14349 vss.n1829 1118.26
R4532 vss.n14345 vss.n1829 1118.26
R4533 vss.n1843 vss.n1842 1118.26
R4534 vss.n1844 vss.n1843 1118.26
R4535 vss.n1844 vss.n1823 1118.26
R4536 vss.n14351 vss.n1823 1118.26
R4537 vss.n14351 vss.n1824 1118.26
R4538 vss.n14343 vss.n1824 1118.26
R4539 vss.n14451 vss.n1756 1118.26
R4540 vss.n14457 vss.n1756 1118.26
R4541 vss.n14457 vss.n1753 1118.26
R4542 vss.n14472 vss.n1753 1118.26
R4543 vss.n14472 vss.n1754 1118.26
R4544 vss.n14468 vss.n1754 1118.26
R4545 vss.n14454 vss.n14453 1118.26
R4546 vss.n14455 vss.n14454 1118.26
R4547 vss.n14455 vss.n1748 1118.26
R4548 vss.n14474 vss.n1748 1118.26
R4549 vss.n14474 vss.n1749 1118.26
R4550 vss.n14465 vss.n1749 1118.26
R4551 vss.n14213 vss.n14204 1118.26
R4552 vss.n14221 vss.n14204 1118.26
R4553 vss.n14221 vss.n14201 1118.26
R4554 vss.n14235 vss.n14201 1118.26
R4555 vss.n14235 vss.n14202 1118.26
R4556 vss.n14231 vss.n14202 1118.26
R4557 vss.n14218 vss.n14217 1118.26
R4558 vss.n14219 vss.n14218 1118.26
R4559 vss.n14219 vss.n14196 1118.26
R4560 vss.n14237 vss.n14196 1118.26
R4561 vss.n14237 vss.n14197 1118.26
R4562 vss.n14229 vss.n14197 1118.26
R4563 vss.n2298 vss.n2288 1118.26
R4564 vss.n2304 vss.n2288 1118.26
R4565 vss.n2304 vss.n2285 1118.26
R4566 vss.n2319 vss.n2285 1118.26
R4567 vss.n2319 vss.n2286 1118.26
R4568 vss.n2315 vss.n2286 1118.26
R4569 vss.n2301 vss.n2300 1118.26
R4570 vss.n2302 vss.n2301 1118.26
R4571 vss.n2302 vss.n2280 1118.26
R4572 vss.n2321 vss.n2280 1118.26
R4573 vss.n2321 vss.n2281 1118.26
R4574 vss.n2312 vss.n2281 1118.26
R4575 vss.n2248 vss.n2242 1118.26
R4576 vss.n2258 vss.n2242 1118.26
R4577 vss.n2258 vss.n2239 1118.26
R4578 vss.n2272 vss.n2239 1118.26
R4579 vss.n2272 vss.n2240 1118.26
R4580 vss.n2268 vss.n2240 1118.26
R4581 vss.n2255 vss.n2254 1118.26
R4582 vss.n2256 vss.n2255 1118.26
R4583 vss.n2256 vss.n2234 1118.26
R4584 vss.n2274 vss.n2234 1118.26
R4585 vss.n2274 vss.n2235 1118.26
R4586 vss.n2266 vss.n2235 1118.26
R4587 vss.n8058 vss.n2227 1118.26
R4588 vss.n8085 vss.n8058 1118.26
R4589 vss.n8085 vss.n8059 1118.26
R4590 vss.n8081 vss.n8059 1118.26
R4591 vss.n8081 vss.n8064 1118.26
R4592 vss.n8071 vss.n8064 1118.26
R4593 vss.n8053 vss.n2228 1118.26
R4594 vss.n8087 vss.n8053 1118.26
R4595 vss.n8087 vss.n8054 1118.26
R4596 vss.n8079 vss.n8054 1118.26
R4597 vss.n8079 vss.n8066 1118.26
R4598 vss.n8069 vss.n8066 1118.26
R4599 vss.n8110 vss.n8108 1118.26
R4600 vss.n8136 vss.n8108 1118.26
R4601 vss.n8136 vss.n8109 1118.26
R4602 vss.n8132 vss.n8109 1118.26
R4603 vss.n8132 vss.n8116 1118.26
R4604 vss.n8124 vss.n8116 1118.26
R4605 vss.n8142 vss.n8100 1118.26
R4606 vss.n8138 vss.n8100 1118.26
R4607 vss.n8138 vss.n8104 1118.26
R4608 vss.n8130 vss.n8104 1118.26
R4609 vss.n8130 vss.n8118 1118.26
R4610 vss.n8126 vss.n8118 1118.26
R4611 vss.n1302 vss.n1293 1118.26
R4612 vss.n1308 vss.n1293 1118.26
R4613 vss.n1308 vss.n1290 1118.26
R4614 vss.n14743 vss.n1290 1118.26
R4615 vss.n14743 vss.n1291 1118.26
R4616 vss.n14739 vss.n1291 1118.26
R4617 vss.n1305 vss.n1304 1118.26
R4618 vss.n1306 vss.n1305 1118.26
R4619 vss.n1306 vss.n1285 1118.26
R4620 vss.n14745 vss.n1285 1118.26
R4621 vss.n14745 vss.n1286 1118.26
R4622 vss.n14737 vss.n1286 1118.26
R4623 vss.n14001 vss.n13992 1118.26
R4624 vss.n14007 vss.n13992 1118.26
R4625 vss.n14007 vss.n13989 1118.26
R4626 vss.n14021 vss.n13989 1118.26
R4627 vss.n14021 vss.n13990 1118.26
R4628 vss.n14017 vss.n13990 1118.26
R4629 vss.n14004 vss.n14003 1118.26
R4630 vss.n14005 vss.n14004 1118.26
R4631 vss.n14005 vss.n13984 1118.26
R4632 vss.n14023 vss.n13984 1118.26
R4633 vss.n14023 vss.n13985 1118.26
R4634 vss.n14015 vss.n13985 1118.26
R4635 vss.n8172 vss.n8163 1118.26
R4636 vss.n13961 vss.n8163 1118.26
R4637 vss.n13961 vss.n8160 1118.26
R4638 vss.n13975 vss.n8160 1118.26
R4639 vss.n13975 vss.n8161 1118.26
R4640 vss.n13971 vss.n8161 1118.26
R4641 vss.n13958 vss.n13957 1118.26
R4642 vss.n13959 vss.n13958 1118.26
R4643 vss.n13959 vss.n8155 1118.26
R4644 vss.n13977 vss.n8155 1118.26
R4645 vss.n13977 vss.n8156 1118.26
R4646 vss.n13969 vss.n8156 1118.26
R4647 vss.n8186 vss.n8176 1118.26
R4648 vss.n8213 vss.n8186 1118.26
R4649 vss.n8213 vss.n8187 1118.26
R4650 vss.n8209 vss.n8187 1118.26
R4651 vss.n8209 vss.n8192 1118.26
R4652 vss.n8199 vss.n8192 1118.26
R4653 vss.n8181 vss.n8177 1118.26
R4654 vss.n8215 vss.n8181 1118.26
R4655 vss.n8215 vss.n8182 1118.26
R4656 vss.n8207 vss.n8182 1118.26
R4657 vss.n8207 vss.n8194 1118.26
R4658 vss.n8197 vss.n8194 1118.26
R4659 vss.n13871 vss.n13869 1118.26
R4660 vss.n13897 vss.n13869 1118.26
R4661 vss.n13897 vss.n13870 1118.26
R4662 vss.n13893 vss.n13870 1118.26
R4663 vss.n13893 vss.n13877 1118.26
R4664 vss.n13885 vss.n13877 1118.26
R4665 vss.n13903 vss.n13861 1118.26
R4666 vss.n13899 vss.n13861 1118.26
R4667 vss.n13899 vss.n13865 1118.26
R4668 vss.n13891 vss.n13865 1118.26
R4669 vss.n13891 vss.n13879 1118.26
R4670 vss.n13887 vss.n13879 1118.26
R4671 vss.n1507 vss.n1498 1118.26
R4672 vss.n1513 vss.n1498 1118.26
R4673 vss.n1513 vss.n1495 1118.26
R4674 vss.n14670 vss.n1495 1118.26
R4675 vss.n14670 vss.n1496 1118.26
R4676 vss.n14666 vss.n1496 1118.26
R4677 vss.n1510 vss.n1509 1118.26
R4678 vss.n1511 vss.n1510 1118.26
R4679 vss.n1511 vss.n1490 1118.26
R4680 vss.n14672 vss.n1490 1118.26
R4681 vss.n14672 vss.n1491 1118.26
R4682 vss.n14664 vss.n1491 1118.26
R4683 vss.n1560 vss.n1551 1118.26
R4684 vss.n1566 vss.n1551 1118.26
R4685 vss.n1566 vss.n1548 1118.26
R4686 vss.n14593 vss.n1548 1118.26
R4687 vss.n14593 vss.n1549 1118.26
R4688 vss.n14589 vss.n1549 1118.26
R4689 vss.n1563 vss.n1562 1118.26
R4690 vss.n1564 vss.n1563 1118.26
R4691 vss.n1564 vss.n1543 1118.26
R4692 vss.n14595 vss.n1543 1118.26
R4693 vss.n14595 vss.n1544 1118.26
R4694 vss.n14587 vss.n1544 1118.26
R4695 vss.n14413 vss.n14410 1118.26
R4696 vss.n14439 vss.n14410 1118.26
R4697 vss.n14439 vss.n14411 1118.26
R4698 vss.n14435 vss.n14411 1118.26
R4699 vss.n14435 vss.n14419 1118.26
R4700 vss.n14427 vss.n14419 1118.26
R4701 vss.n14445 vss.n14402 1118.26
R4702 vss.n14441 vss.n14402 1118.26
R4703 vss.n14441 vss.n14406 1118.26
R4704 vss.n14433 vss.n14406 1118.26
R4705 vss.n14433 vss.n14421 1118.26
R4706 vss.n14429 vss.n14421 1118.26
R4707 vss.n14500 vss.n14491 1118.26
R4708 vss.n14506 vss.n14491 1118.26
R4709 vss.n14506 vss.n14488 1118.26
R4710 vss.n14520 vss.n14488 1118.26
R4711 vss.n14520 vss.n14489 1118.26
R4712 vss.n14516 vss.n14489 1118.26
R4713 vss.n14503 vss.n14502 1118.26
R4714 vss.n14504 vss.n14503 1118.26
R4715 vss.n14504 vss.n14483 1118.26
R4716 vss.n14522 vss.n14483 1118.26
R4717 vss.n14522 vss.n14484 1118.26
R4718 vss.n14514 vss.n14484 1118.26
R4719 vss.n1717 vss.n1708 1118.26
R4720 vss.n1723 vss.n1708 1118.26
R4721 vss.n1723 vss.n1705 1118.26
R4722 vss.n1738 vss.n1705 1118.26
R4723 vss.n1738 vss.n1706 1118.26
R4724 vss.n1734 vss.n1706 1118.26
R4725 vss.n1720 vss.n1719 1118.26
R4726 vss.n1721 vss.n1720 1118.26
R4727 vss.n1721 vss.n1700 1118.26
R4728 vss.n1740 vss.n1700 1118.26
R4729 vss.n1740 vss.n1701 1118.26
R4730 vss.n1732 vss.n1701 1118.26
R4731 vss.n1608 vss.n1600 1118.26
R4732 vss.n1616 vss.n1600 1118.26
R4733 vss.n1616 vss.n1594 1118.26
R4734 vss.n1621 vss.n1594 1118.26
R4735 vss.n1621 vss.n1596 1118.26
R4736 vss.n1596 vss.n1585 1118.26
R4737 vss.n1610 vss.n1602 1118.26
R4738 vss.n1614 vss.n1602 1118.26
R4739 vss.n1614 vss.n1590 1118.26
R4740 vss.n1623 vss.n1590 1118.26
R4741 vss.n1623 vss.n1591 1118.26
R4742 vss.n1591 vss.n1586 1118.26
R4743 vss.n13916 vss.n13907 1118.26
R4744 vss.n13944 vss.n13916 1118.26
R4745 vss.n13944 vss.n13917 1118.26
R4746 vss.n13940 vss.n13917 1118.26
R4747 vss.n13940 vss.n13923 1118.26
R4748 vss.n13931 vss.n13923 1118.26
R4749 vss.n13950 vss.n13908 1118.26
R4750 vss.n13946 vss.n13908 1118.26
R4751 vss.n13946 vss.n13913 1118.26
R4752 vss.n13938 vss.n13913 1118.26
R4753 vss.n13938 vss.n13925 1118.26
R4754 vss.n13934 vss.n13925 1118.26
R4755 vss.n14620 vss.n14611 1118.26
R4756 vss.n14626 vss.n14611 1118.26
R4757 vss.n14626 vss.n14608 1118.26
R4758 vss.n14641 vss.n14608 1118.26
R4759 vss.n14641 vss.n14609 1118.26
R4760 vss.n14637 vss.n14609 1118.26
R4761 vss.n14623 vss.n14622 1118.26
R4762 vss.n14624 vss.n14623 1118.26
R4763 vss.n14624 vss.n14603 1118.26
R4764 vss.n14643 vss.n14603 1118.26
R4765 vss.n14643 vss.n14604 1118.26
R4766 vss.n14635 vss.n14604 1118.26
R4767 vss.n1460 vss.n1451 1118.26
R4768 vss.n1466 vss.n1451 1118.26
R4769 vss.n1466 vss.n1448 1118.26
R4770 vss.n1481 vss.n1448 1118.26
R4771 vss.n1481 vss.n1449 1118.26
R4772 vss.n1477 vss.n1449 1118.26
R4773 vss.n1463 vss.n1462 1118.26
R4774 vss.n1464 vss.n1463 1118.26
R4775 vss.n1464 vss.n1443 1118.26
R4776 vss.n1483 vss.n1443 1118.26
R4777 vss.n1483 vss.n1444 1118.26
R4778 vss.n1475 vss.n1444 1118.26
R4779 vss.n14033 vss.n8146 1118.26
R4780 vss.n14061 vss.n14033 1118.26
R4781 vss.n14061 vss.n14034 1118.26
R4782 vss.n14057 vss.n14034 1118.26
R4783 vss.n14057 vss.n14040 1118.26
R4784 vss.n14048 vss.n14040 1118.26
R4785 vss.n14067 vss.n8147 1118.26
R4786 vss.n14063 vss.n8147 1118.26
R4787 vss.n14063 vss.n14030 1118.26
R4788 vss.n14055 vss.n14030 1118.26
R4789 vss.n14055 vss.n14042 1118.26
R4790 vss.n14051 vss.n14042 1118.26
R4791 vss.n1351 vss.n1343 1118.26
R4792 vss.n1359 vss.n1343 1118.26
R4793 vss.n1359 vss.n1337 1118.26
R4794 vss.n1364 vss.n1337 1118.26
R4795 vss.n1364 vss.n1339 1118.26
R4796 vss.n1339 vss.n1327 1118.26
R4797 vss.n1353 vss.n1345 1118.26
R4798 vss.n1357 vss.n1345 1118.26
R4799 vss.n1357 vss.n1333 1118.26
R4800 vss.n1366 vss.n1333 1118.26
R4801 vss.n1366 vss.n1334 1118.26
R4802 vss.n1334 vss.n1328 1118.26
R4803 vss.n1252 vss.n1243 1118.26
R4804 vss.n1258 vss.n1243 1118.26
R4805 vss.n1258 vss.n1240 1118.26
R4806 vss.n1273 vss.n1240 1118.26
R4807 vss.n1273 vss.n1241 1118.26
R4808 vss.n1269 vss.n1241 1118.26
R4809 vss.n1255 vss.n1254 1118.26
R4810 vss.n1256 vss.n1255 1118.26
R4811 vss.n1256 vss.n1235 1118.26
R4812 vss.n1275 vss.n1235 1118.26
R4813 vss.n1275 vss.n1236 1118.26
R4814 vss.n1267 vss.n1236 1118.26
R4815 vss.n2345 vss.n2336 1118.26
R4816 vss.n2351 vss.n2336 1118.26
R4817 vss.n2351 vss.n2333 1118.26
R4818 vss.n8042 vss.n2333 1118.26
R4819 vss.n8042 vss.n2334 1118.26
R4820 vss.n8038 vss.n2334 1118.26
R4821 vss.n2348 vss.n2347 1118.26
R4822 vss.n2349 vss.n2348 1118.26
R4823 vss.n2349 vss.n2328 1118.26
R4824 vss.n8044 vss.n2328 1118.26
R4825 vss.n8044 vss.n2329 1118.26
R4826 vss.n8036 vss.n2329 1118.26
R4827 vss.n2393 vss.n2385 1118.26
R4828 vss.n2401 vss.n2385 1118.26
R4829 vss.n2401 vss.n2379 1118.26
R4830 vss.n2406 vss.n2379 1118.26
R4831 vss.n2406 vss.n2381 1118.26
R4832 vss.n2381 vss.n2370 1118.26
R4833 vss.n2395 vss.n2387 1118.26
R4834 vss.n2399 vss.n2387 1118.26
R4835 vss.n2399 vss.n2375 1118.26
R4836 vss.n2408 vss.n2375 1118.26
R4837 vss.n2408 vss.n2376 1118.26
R4838 vss.n2376 vss.n2371 1118.26
R4839 vss.n11853 vss.n11849 1118.26
R4840 vss.n11859 vss.n11853 1118.26
R4841 vss.n11859 vss.n2043 1118.26
R4842 vss.n14185 vss.n2043 1118.26
R4843 vss.n14185 vss.n2044 1118.26
R4844 vss.n14181 vss.n2044 1118.26
R4845 vss.n11856 vss.n11848 1118.26
R4846 vss.n11857 vss.n11856 1118.26
R4847 vss.n11857 vss.n2038 1118.26
R4848 vss.n14187 vss.n2038 1118.26
R4849 vss.n14187 vss.n2039 1118.26
R4850 vss.n2051 vss.n2039 1118.26
R4851 vss.n11953 vss.n11945 1118.26
R4852 vss.n11954 vss.n11953 1118.26
R4853 vss.n11954 vss.n2090 1118.26
R4854 vss.n14135 vss.n2090 1118.26
R4855 vss.n14135 vss.n2091 1118.26
R4856 vss.n14127 vss.n2091 1118.26
R4857 vss.n11950 vss.n11946 1118.26
R4858 vss.n11956 vss.n11950 1118.26
R4859 vss.n11956 vss.n2095 1118.26
R4860 vss.n14133 vss.n2095 1118.26
R4861 vss.n14133 vss.n2096 1118.26
R4862 vss.n14129 vss.n2096 1118.26
R4863 vss.n13490 vss.n13489 1118.26
R4864 vss.n13491 vss.n13490 1118.26
R4865 vss.n13491 vss.n13470 1118.26
R4866 vss.n13509 vss.n13470 1118.26
R4867 vss.n13509 vss.n13471 1118.26
R4868 vss.n13501 vss.n13471 1118.26
R4869 vss.n13487 vss.n13478 1118.26
R4870 vss.n13493 vss.n13478 1118.26
R4871 vss.n13493 vss.n13475 1118.26
R4872 vss.n13507 vss.n13475 1118.26
R4873 vss.n13507 vss.n13476 1118.26
R4874 vss.n13503 vss.n13476 1118.26
R4875 vss.n12026 vss.n12016 1118.26
R4876 vss.n12052 vss.n12026 1118.26
R4877 vss.n12052 vss.n12027 1118.26
R4878 vss.n12048 vss.n12027 1118.26
R4879 vss.n12048 vss.n12032 1118.26
R4880 vss.n12040 vss.n12032 1118.26
R4881 vss.n12021 vss.n12017 1118.26
R4882 vss.n12054 vss.n12021 1118.26
R4883 vss.n12054 vss.n12022 1118.26
R4884 vss.n12046 vss.n12022 1118.26
R4885 vss.n12046 vss.n12034 1118.26
R4886 vss.n12042 vss.n12034 1118.26
R4887 vss.n13722 vss.n13721 1118.26
R4888 vss.n13723 vss.n13722 1118.26
R4889 vss.n13723 vss.n8305 1118.26
R4890 vss.n13741 vss.n8305 1118.26
R4891 vss.n13741 vss.n8306 1118.26
R4892 vss.n13733 vss.n8306 1118.26
R4893 vss.n13719 vss.n8313 1118.26
R4894 vss.n13725 vss.n8313 1118.26
R4895 vss.n13725 vss.n8310 1118.26
R4896 vss.n13739 vss.n8310 1118.26
R4897 vss.n13739 vss.n8311 1118.26
R4898 vss.n13735 vss.n8311 1118.26
R4899 vss.n8452 vss.n8442 1118.26
R4900 vss.n8478 vss.n8452 1118.26
R4901 vss.n8478 vss.n8453 1118.26
R4902 vss.n8474 vss.n8453 1118.26
R4903 vss.n8474 vss.n8458 1118.26
R4904 vss.n8466 vss.n8458 1118.26
R4905 vss.n8447 vss.n8443 1118.26
R4906 vss.n8480 vss.n8447 1118.26
R4907 vss.n8480 vss.n8448 1118.26
R4908 vss.n8472 vss.n8448 1118.26
R4909 vss.n8472 vss.n8460 1118.26
R4910 vss.n8468 vss.n8460 1118.26
R4911 vss.n8529 vss.n8519 1118.26
R4912 vss.n8555 vss.n8529 1118.26
R4913 vss.n8555 vss.n8530 1118.26
R4914 vss.n8551 vss.n8530 1118.26
R4915 vss.n8551 vss.n8535 1118.26
R4916 vss.n8543 vss.n8535 1118.26
R4917 vss.n8524 vss.n8520 1118.26
R4918 vss.n8557 vss.n8524 1118.26
R4919 vss.n8557 vss.n8525 1118.26
R4920 vss.n8549 vss.n8525 1118.26
R4921 vss.n8549 vss.n8537 1118.26
R4922 vss.n8545 vss.n8537 1118.26
R4923 vss.n13010 vss.n13009 1118.26
R4924 vss.n13011 vss.n13010 1118.26
R4925 vss.n13011 vss.n9091 1118.26
R4926 vss.n13029 vss.n9091 1118.26
R4927 vss.n13029 vss.n9092 1118.26
R4928 vss.n13021 vss.n9092 1118.26
R4929 vss.n13007 vss.n9099 1118.26
R4930 vss.n13013 vss.n9099 1118.26
R4931 vss.n13013 vss.n9096 1118.26
R4932 vss.n13027 vss.n9096 1118.26
R4933 vss.n13027 vss.n9097 1118.26
R4934 vss.n13023 vss.n9097 1118.26
R4935 vss.n8975 vss.n8974 1118.26
R4936 vss.n8976 vss.n8975 1118.26
R4937 vss.n8976 vss.n8955 1118.26
R4938 vss.n8994 vss.n8955 1118.26
R4939 vss.n8994 vss.n8956 1118.26
R4940 vss.n8986 vss.n8956 1118.26
R4941 vss.n8972 vss.n8963 1118.26
R4942 vss.n8978 vss.n8963 1118.26
R4943 vss.n8978 vss.n8960 1118.26
R4944 vss.n8992 vss.n8960 1118.26
R4945 vss.n8992 vss.n8961 1118.26
R4946 vss.n8988 vss.n8961 1118.26
R4947 vss.n9124 vss.n9114 1118.26
R4948 vss.n9150 vss.n9124 1118.26
R4949 vss.n9150 vss.n9125 1118.26
R4950 vss.n9146 vss.n9125 1118.26
R4951 vss.n9146 vss.n9130 1118.26
R4952 vss.n9138 vss.n9130 1118.26
R4953 vss.n9119 vss.n9115 1118.26
R4954 vss.n9152 vss.n9119 1118.26
R4955 vss.n9152 vss.n9120 1118.26
R4956 vss.n9144 vss.n9120 1118.26
R4957 vss.n9144 vss.n9132 1118.26
R4958 vss.n9140 vss.n9132 1118.26
R4959 vss.n12555 vss.n12545 1118.26
R4960 vss.n12630 vss.n12555 1118.26
R4961 vss.n12630 vss.n12556 1118.26
R4962 vss.n12577 vss.n12556 1118.26
R4963 vss.n12577 vss.n12561 1118.26
R4964 vss.n12569 vss.n12561 1118.26
R4965 vss.n12550 vss.n12546 1118.26
R4966 vss.n12632 vss.n12550 1118.26
R4967 vss.n12632 vss.n12551 1118.26
R4968 vss.n12575 vss.n12551 1118.26
R4969 vss.n12575 vss.n12563 1118.26
R4970 vss.n12571 vss.n12563 1118.26
R4971 vss.n2166 vss.n2157 1118.26
R4972 vss.n2172 vss.n2157 1118.26
R4973 vss.n2172 vss.n2154 1118.26
R4974 vss.n14082 vss.n2154 1118.26
R4975 vss.n14082 vss.n2155 1118.26
R4976 vss.n14078 vss.n2155 1118.26
R4977 vss.n2169 vss.n2168 1118.26
R4978 vss.n2170 vss.n2169 1118.26
R4979 vss.n2170 vss.n2149 1118.26
R4980 vss.n14084 vss.n2149 1118.26
R4981 vss.n14084 vss.n2150 1118.26
R4982 vss.n14075 vss.n2150 1118.26
R4983 vss.n12599 vss.n12590 1118.26
R4984 vss.n12606 vss.n12590 1118.26
R4985 vss.n12606 vss.n12587 1118.26
R4986 vss.n12620 vss.n12587 1118.26
R4987 vss.n12620 vss.n12588 1118.26
R4988 vss.n12616 vss.n12588 1118.26
R4989 vss.n12603 vss.n12602 1118.26
R4990 vss.n12604 vss.n12603 1118.26
R4991 vss.n12604 vss.n12582 1118.26
R4992 vss.n12622 vss.n12582 1118.26
R4993 vss.n12622 vss.n12583 1118.26
R4994 vss.n12614 vss.n12583 1118.26
R4995 vss.n9020 vss.n9019 1118.26
R4996 vss.n9021 vss.n9020 1118.26
R4997 vss.n9021 vss.n9000 1118.26
R4998 vss.n9038 vss.n9000 1118.26
R4999 vss.n9038 vss.n9001 1118.26
R5000 vss.n9028 vss.n9001 1118.26
R5001 vss.n9017 vss.n9008 1118.26
R5002 vss.n9023 vss.n9008 1118.26
R5003 vss.n9023 vss.n9005 1118.26
R5004 vss.n9036 vss.n9005 1118.26
R5005 vss.n9036 vss.n9006 1118.26
R5006 vss.n9032 vss.n9006 1118.26
R5007 vss.n13102 vss.n13093 1118.26
R5008 vss.n13109 vss.n13093 1118.26
R5009 vss.n13109 vss.n13090 1118.26
R5010 vss.n13124 vss.n13090 1118.26
R5011 vss.n13124 vss.n13091 1118.26
R5012 vss.n13120 vss.n13091 1118.26
R5013 vss.n13106 vss.n13105 1118.26
R5014 vss.n13107 vss.n13106 1118.26
R5015 vss.n13107 vss.n13085 1118.26
R5016 vss.n13126 vss.n13085 1118.26
R5017 vss.n13126 vss.n13086 1118.26
R5018 vss.n13117 vss.n13086 1118.26
R5019 vss.n13054 vss.n13045 1118.26
R5020 vss.n13060 vss.n13045 1118.26
R5021 vss.n13060 vss.n13042 1118.26
R5022 vss.n13076 vss.n13042 1118.26
R5023 vss.n13076 vss.n13043 1118.26
R5024 vss.n13072 vss.n13043 1118.26
R5025 vss.n13057 vss.n13056 1118.26
R5026 vss.n13058 vss.n13057 1118.26
R5027 vss.n13058 vss.n13037 1118.26
R5028 vss.n13078 vss.n13037 1118.26
R5029 vss.n13078 vss.n13038 1118.26
R5030 vss.n13069 vss.n13038 1118.26
R5031 vss.n9061 vss.n9052 1118.26
R5032 vss.n9068 vss.n9052 1118.26
R5033 vss.n9068 vss.n9049 1118.26
R5034 vss.n9082 vss.n9049 1118.26
R5035 vss.n9082 vss.n9050 1118.26
R5036 vss.n9078 vss.n9050 1118.26
R5037 vss.n9065 vss.n9064 1118.26
R5038 vss.n9066 vss.n9065 1118.26
R5039 vss.n9066 vss.n9044 1118.26
R5040 vss.n9084 vss.n9044 1118.26
R5041 vss.n9084 vss.n9045 1118.26
R5042 vss.n9076 vss.n9045 1118.26
R5043 vss.n8244 vss.n8236 1118.26
R5044 vss.n8252 vss.n8236 1118.26
R5045 vss.n8252 vss.n8232 1118.26
R5046 vss.n13847 vss.n8232 1118.26
R5047 vss.n13849 vss.n13847 1118.26
R5048 vss.n13849 vss.n8224 1118.26
R5049 vss.n8246 vss.n8238 1118.26
R5050 vss.n8250 vss.n8238 1118.26
R5051 vss.n8250 vss.n8229 1118.26
R5052 vss.n13853 vss.n8229 1118.26
R5053 vss.n13853 vss.n8230 1118.26
R5054 vss.n8230 vss.n8225 1118.26
R5055 vss.n13814 vss.n13805 1118.26
R5056 vss.n13821 vss.n13805 1118.26
R5057 vss.n13821 vss.n13802 1118.26
R5058 vss.n13836 vss.n13802 1118.26
R5059 vss.n13836 vss.n13803 1118.26
R5060 vss.n13832 vss.n13803 1118.26
R5061 vss.n13818 vss.n13817 1118.26
R5062 vss.n13819 vss.n13818 1118.26
R5063 vss.n13819 vss.n13797 1118.26
R5064 vss.n13838 vss.n13797 1118.26
R5065 vss.n13838 vss.n13798 1118.26
R5066 vss.n13829 vss.n13798 1118.26
R5067 vss.n13766 vss.n13757 1118.26
R5068 vss.n13772 vss.n13757 1118.26
R5069 vss.n13772 vss.n13754 1118.26
R5070 vss.n13788 vss.n13754 1118.26
R5071 vss.n13788 vss.n13755 1118.26
R5072 vss.n13784 vss.n13755 1118.26
R5073 vss.n13769 vss.n13768 1118.26
R5074 vss.n13770 vss.n13769 1118.26
R5075 vss.n13770 vss.n13749 1118.26
R5076 vss.n13790 vss.n13749 1118.26
R5077 vss.n13790 vss.n13750 1118.26
R5078 vss.n13781 vss.n13750 1118.26
R5079 vss.n8275 vss.n8266 1118.26
R5080 vss.n8282 vss.n8266 1118.26
R5081 vss.n8282 vss.n8263 1118.26
R5082 vss.n8296 vss.n8263 1118.26
R5083 vss.n8296 vss.n8264 1118.26
R5084 vss.n8292 vss.n8264 1118.26
R5085 vss.n8279 vss.n8278 1118.26
R5086 vss.n8280 vss.n8279 1118.26
R5087 vss.n8280 vss.n8258 1118.26
R5088 vss.n8298 vss.n8258 1118.26
R5089 vss.n8298 vss.n8259 1118.26
R5090 vss.n8290 vss.n8259 1118.26
R5091 vss.n13535 vss.n13534 1118.26
R5092 vss.n13536 vss.n13535 1118.26
R5093 vss.n13536 vss.n13515 1118.26
R5094 vss.n13553 vss.n13515 1118.26
R5095 vss.n13553 vss.n13516 1118.26
R5096 vss.n13543 vss.n13516 1118.26
R5097 vss.n13532 vss.n13523 1118.26
R5098 vss.n13538 vss.n13523 1118.26
R5099 vss.n13538 vss.n13520 1118.26
R5100 vss.n13551 vss.n13520 1118.26
R5101 vss.n13551 vss.n13521 1118.26
R5102 vss.n13547 vss.n13521 1118.26
R5103 vss.n13625 vss.n13616 1118.26
R5104 vss.n13632 vss.n13616 1118.26
R5105 vss.n13632 vss.n13613 1118.26
R5106 vss.n13647 vss.n13613 1118.26
R5107 vss.n13647 vss.n13614 1118.26
R5108 vss.n13643 vss.n13614 1118.26
R5109 vss.n13629 vss.n13628 1118.26
R5110 vss.n13630 vss.n13629 1118.26
R5111 vss.n13630 vss.n13608 1118.26
R5112 vss.n13649 vss.n13608 1118.26
R5113 vss.n13649 vss.n13609 1118.26
R5114 vss.n13640 vss.n13609 1118.26
R5115 vss.n13577 vss.n13567 1118.26
R5116 vss.n13583 vss.n13567 1118.26
R5117 vss.n13583 vss.n13564 1118.26
R5118 vss.n13599 vss.n13564 1118.26
R5119 vss.n13599 vss.n13565 1118.26
R5120 vss.n13595 vss.n13565 1118.26
R5121 vss.n13580 vss.n13579 1118.26
R5122 vss.n13581 vss.n13580 1118.26
R5123 vss.n13581 vss.n13559 1118.26
R5124 vss.n13601 vss.n13559 1118.26
R5125 vss.n13601 vss.n13560 1118.26
R5126 vss.n13592 vss.n13560 1118.26
R5127 vss.n2079 vss.n2069 1118.26
R5128 vss.n2083 vss.n2069 1118.26
R5129 vss.n2083 vss.n2060 1118.26
R5130 vss.n14149 vss.n2060 1118.26
R5131 vss.n14149 vss.n2061 1118.26
R5132 vss.n2061 vss.n2056 1118.26
R5133 vss.n2076 vss.n2067 1118.26
R5134 vss.n2085 vss.n2067 1118.26
R5135 vss.n2085 vss.n2063 1118.26
R5136 vss.n14144 vss.n2063 1118.26
R5137 vss.n14145 vss.n14144 1118.26
R5138 vss.n14145 vss.n2055 1118.26
R5139 vss.n2202 vss.n2192 1118.26
R5140 vss.n2210 vss.n2192 1118.26
R5141 vss.n2211 vss.n2210 1118.26
R5142 vss.n2216 vss.n2211 1118.26
R5143 vss.n2216 vss.n2213 1118.26
R5144 vss.n2213 vss.n2181 1118.26
R5145 vss.n2204 vss.n2195 1118.26
R5146 vss.n2208 vss.n2195 1118.26
R5147 vss.n2208 vss.n2186 1118.26
R5148 vss.n2218 vss.n2186 1118.26
R5149 vss.n2218 vss.n2187 1118.26
R5150 vss.n2187 vss.n2182 1118.26
R5151 vss.n9292 vss.n9284 1118.26
R5152 vss.n9293 vss.n9292 1118.26
R5153 vss.n9293 vss.n2138 1118.26
R5154 vss.n14095 vss.n2138 1118.26
R5155 vss.n14095 vss.n2140 1118.26
R5156 vss.n2140 vss.n2129 1118.26
R5157 vss.n9289 vss.n9285 1118.26
R5158 vss.n9295 vss.n9289 1118.26
R5159 vss.n9295 vss.n2134 1118.26
R5160 vss.n14097 vss.n2134 1118.26
R5161 vss.n14097 vss.n2135 1118.26
R5162 vss.n2135 vss.n2130 1118.26
R5163 vss.n12847 vss.n12846 1118.26
R5164 vss.n12848 vss.n12847 1118.26
R5165 vss.n12848 vss.n9395 1118.26
R5166 vss.n12866 vss.n9395 1118.26
R5167 vss.n12866 vss.n9396 1118.26
R5168 vss.n12858 vss.n9396 1118.26
R5169 vss.n12844 vss.n9403 1118.26
R5170 vss.n12850 vss.n9403 1118.26
R5171 vss.n12850 vss.n9400 1118.26
R5172 vss.n12864 vss.n9400 1118.26
R5173 vss.n12864 vss.n9401 1118.26
R5174 vss.n12860 vss.n9401 1118.26
R5175 vss.n12739 vss.n12729 1118.26
R5176 vss.n12766 vss.n12739 1118.26
R5177 vss.n12766 vss.n12740 1118.26
R5178 vss.n12761 vss.n12740 1118.26
R5179 vss.n12761 vss.n12745 1118.26
R5180 vss.n12753 vss.n12745 1118.26
R5181 vss.n12734 vss.n12730 1118.26
R5182 vss.n12768 vss.n12734 1118.26
R5183 vss.n12768 vss.n12735 1118.26
R5184 vss.n12759 vss.n12735 1118.26
R5185 vss.n12759 vss.n12747 1118.26
R5186 vss.n12755 vss.n12747 1118.26
R5187 vss.n13324 vss.n13323 1118.26
R5188 vss.n13325 vss.n13324 1118.26
R5189 vss.n13325 vss.n8413 1118.26
R5190 vss.n13343 vss.n8413 1118.26
R5191 vss.n13343 vss.n8414 1118.26
R5192 vss.n13335 vss.n8414 1118.26
R5193 vss.n13321 vss.n8421 1118.26
R5194 vss.n13327 vss.n8421 1118.26
R5195 vss.n13327 vss.n8418 1118.26
R5196 vss.n13341 vss.n8418 1118.26
R5197 vss.n13341 vss.n8419 1118.26
R5198 vss.n13337 vss.n8419 1118.26
R5199 vss.n13443 vss.n13442 1118.26
R5200 vss.n13444 vss.n13443 1118.26
R5201 vss.n13444 vss.n13355 1118.26
R5202 vss.n13462 vss.n13355 1118.26
R5203 vss.n13462 vss.n13356 1118.26
R5204 vss.n13454 vss.n13356 1118.26
R5205 vss.n13440 vss.n13363 1118.26
R5206 vss.n13446 vss.n13363 1118.26
R5207 vss.n13446 vss.n13360 1118.26
R5208 vss.n13460 vss.n13360 1118.26
R5209 vss.n13460 vss.n13361 1118.26
R5210 vss.n13456 vss.n13361 1118.26
R5211 vss.n1780 vss.n1778 1118.26
R5212 vss.n1806 vss.n1778 1118.26
R5213 vss.n1806 vss.n1779 1118.26
R5214 vss.n1802 vss.n1779 1118.26
R5215 vss.n1802 vss.n1786 1118.26
R5216 vss.n1794 vss.n1786 1118.26
R5217 vss.n1812 vss.n1770 1118.26
R5218 vss.n1808 vss.n1770 1118.26
R5219 vss.n1808 vss.n1774 1118.26
R5220 vss.n1800 vss.n1774 1118.26
R5221 vss.n1800 vss.n1788 1118.26
R5222 vss.n1796 vss.n1788 1118.26
R5223 vss.n14361 vss.n1816 1118.26
R5224 vss.n14389 vss.n14361 1118.26
R5225 vss.n14389 vss.n14362 1118.26
R5226 vss.n14385 vss.n14362 1118.26
R5227 vss.n14385 vss.n14368 1118.26
R5228 vss.n14376 vss.n14368 1118.26
R5229 vss.n14395 vss.n1817 1118.26
R5230 vss.n14391 vss.n1817 1118.26
R5231 vss.n14391 vss.n14358 1118.26
R5232 vss.n14383 vss.n14358 1118.26
R5233 vss.n14383 vss.n14370 1118.26
R5234 vss.n14379 vss.n14370 1118.26
R5235 vss.n2007 vss.n1998 1118.26
R5236 vss.n2013 vss.n1998 1118.26
R5237 vss.n2013 vss.n1995 1118.26
R5238 vss.n2028 vss.n1995 1118.26
R5239 vss.n2028 vss.n1996 1118.26
R5240 vss.n2024 vss.n1996 1118.26
R5241 vss.n2010 vss.n2009 1118.26
R5242 vss.n2011 vss.n2010 1118.26
R5243 vss.n2011 vss.n1990 1118.26
R5244 vss.n2030 vss.n1990 1118.26
R5245 vss.n2030 vss.n1991 1118.26
R5246 vss.n2022 vss.n1991 1118.26
R5247 vss.n1001 vss.n999 1118.26
R5248 vss.n1027 vss.n999 1118.26
R5249 vss.n1027 vss.n1000 1118.26
R5250 vss.n1023 vss.n1000 1118.26
R5251 vss.n1023 vss.n1007 1118.26
R5252 vss.n1015 vss.n1007 1118.26
R5253 vss.n1033 vss.n991 1118.26
R5254 vss.n1029 vss.n991 1118.26
R5255 vss.n1029 vss.n995 1118.26
R5256 vss.n1021 vss.n995 1118.26
R5257 vss.n1021 vss.n1009 1118.26
R5258 vss.n1017 vss.n1009 1118.26
R5259 vss.n15056 vss.n1037 1118.26
R5260 vss.n15084 vss.n15056 1118.26
R5261 vss.n15084 vss.n15057 1118.26
R5262 vss.n15080 vss.n15057 1118.26
R5263 vss.n15080 vss.n15063 1118.26
R5264 vss.n15071 vss.n15063 1118.26
R5265 vss.n15090 vss.n1038 1118.26
R5266 vss.n15086 vss.n1038 1118.26
R5267 vss.n15086 vss.n15053 1118.26
R5268 vss.n15078 vss.n15053 1118.26
R5269 vss.n15078 vss.n15065 1118.26
R5270 vss.n15074 vss.n15065 1118.26
R5271 vss.n1112 vss.n1103 1118.26
R5272 vss.n1118 vss.n1103 1118.26
R5273 vss.n1118 vss.n1100 1118.26
R5274 vss.n1133 vss.n1100 1118.26
R5275 vss.n1133 vss.n1101 1118.26
R5276 vss.n1129 vss.n1101 1118.26
R5277 vss.n1115 vss.n1114 1118.26
R5278 vss.n1116 vss.n1115 1118.26
R5279 vss.n1116 vss.n1095 1118.26
R5280 vss.n1135 vss.n1095 1118.26
R5281 vss.n1135 vss.n1096 1118.26
R5282 vss.n1127 vss.n1096 1118.26
R5283 vss.n6215 vss.n6206 1118.26
R5284 vss.n6243 vss.n6215 1118.26
R5285 vss.n6243 vss.n6216 1118.26
R5286 vss.n6239 vss.n6216 1118.26
R5287 vss.n6239 vss.n6222 1118.26
R5288 vss.n6230 vss.n6222 1118.26
R5289 vss.n6249 vss.n6207 1118.26
R5290 vss.n6245 vss.n6207 1118.26
R5291 vss.n6245 vss.n6212 1118.26
R5292 vss.n6237 vss.n6212 1118.26
R5293 vss.n6237 vss.n6224 1118.26
R5294 vss.n6233 vss.n6224 1118.26
R5295 vss.n3959 vss.n3950 1118.26
R5296 vss.n3959 vss.n3958 1118.26
R5297 vss.n3958 vss.n37 1118.26
R5298 vss.n15864 vss.n37 1118.26
R5299 vss.n15864 vss.n38 1118.26
R5300 vss.n15860 vss.n38 1118.26
R5301 vss.n3964 vss.n3951 1118.26
R5302 vss.n3956 vss.n3951 1118.26
R5303 vss.n3956 vss.n32 1118.26
R5304 vss.n15866 vss.n32 1118.26
R5305 vss.n15866 vss.n33 1118.26
R5306 vss.n15858 vss.n33 1118.26
R5307 vss.n3861 vss.n3852 1118.26
R5308 vss.n3889 vss.n3861 1118.26
R5309 vss.n3889 vss.n3862 1118.26
R5310 vss.n3885 vss.n3862 1118.26
R5311 vss.n3885 vss.n3868 1118.26
R5312 vss.n3877 vss.n3868 1118.26
R5313 vss.n3895 vss.n3853 1118.26
R5314 vss.n3891 vss.n3853 1118.26
R5315 vss.n3891 vss.n3858 1118.26
R5316 vss.n3883 vss.n3858 1118.26
R5317 vss.n3883 vss.n3870 1118.26
R5318 vss.n3879 vss.n3870 1118.26
R5319 vss.n3742 vss.n3733 1118.26
R5320 vss.n3770 vss.n3742 1118.26
R5321 vss.n3770 vss.n3743 1118.26
R5322 vss.n3766 vss.n3743 1118.26
R5323 vss.n3766 vss.n3749 1118.26
R5324 vss.n3758 vss.n3749 1118.26
R5325 vss.n3776 vss.n3734 1118.26
R5326 vss.n3772 vss.n3734 1118.26
R5327 vss.n3772 vss.n3739 1118.26
R5328 vss.n3764 vss.n3739 1118.26
R5329 vss.n3764 vss.n3751 1118.26
R5330 vss.n3760 vss.n3751 1118.26
R5331 vss.n3623 vss.n3614 1118.26
R5332 vss.n3651 vss.n3623 1118.26
R5333 vss.n3651 vss.n3624 1118.26
R5334 vss.n3647 vss.n3624 1118.26
R5335 vss.n3647 vss.n3630 1118.26
R5336 vss.n3639 vss.n3630 1118.26
R5337 vss.n3657 vss.n3615 1118.26
R5338 vss.n3653 vss.n3615 1118.26
R5339 vss.n3653 vss.n3620 1118.26
R5340 vss.n3645 vss.n3620 1118.26
R5341 vss.n3645 vss.n3632 1118.26
R5342 vss.n3641 vss.n3632 1118.26
R5343 vss.n15596 vss.n15589 1118.26
R5344 vss.n15596 vss.n15590 1118.26
R5345 vss.n15592 vss.n15590 1118.26
R5346 vss.n15608 vss.n15592 1118.26
R5347 vss.n15608 vss.n15587 1118.26
R5348 vss.n15610 vss.n15587 1118.26
R5349 vss.n15600 vss.n15599 1118.26
R5350 vss.n15599 vss.n15598 1118.26
R5351 vss.n15598 vss.n15582 1118.26
R5352 vss.n15616 vss.n15582 1118.26
R5353 vss.n15616 vss.n15615 1118.26
R5354 vss.n15615 vss.n15614 1118.26
R5355 vss.n314 vss.n306 1118.26
R5356 vss.n342 vss.n314 1118.26
R5357 vss.n342 vss.n315 1118.26
R5358 vss.n338 vss.n315 1118.26
R5359 vss.n338 vss.n321 1118.26
R5360 vss.n330 vss.n321 1118.26
R5361 vss.n348 vss.n307 1118.26
R5362 vss.n344 vss.n307 1118.26
R5363 vss.n344 vss.n311 1118.26
R5364 vss.n336 vss.n311 1118.26
R5365 vss.n336 vss.n323 1118.26
R5366 vss.n332 vss.n323 1118.26
R5367 vss.n15550 vss.n371 1118.26
R5368 vss.n15556 vss.n371 1118.26
R5369 vss.n15556 vss.n368 1118.26
R5370 vss.n15570 vss.n368 1118.26
R5371 vss.n15570 vss.n369 1118.26
R5372 vss.n15566 vss.n369 1118.26
R5373 vss.n15553 vss.n15552 1118.26
R5374 vss.n15554 vss.n15553 1118.26
R5375 vss.n15554 vss.n363 1118.26
R5376 vss.n15572 vss.n363 1118.26
R5377 vss.n15572 vss.n364 1118.26
R5378 vss.n15564 vss.n364 1118.26
R5379 vss.n10447 vss.n10446 1118.26
R5380 vss.n10448 vss.n10447 1118.26
R5381 vss.n10448 vss.n10427 1118.26
R5382 vss.n10467 vss.n10427 1118.26
R5383 vss.n10467 vss.n10428 1118.26
R5384 vss.n10459 vss.n10428 1118.26
R5385 vss.n10444 vss.n10435 1118.26
R5386 vss.n10450 vss.n10435 1118.26
R5387 vss.n10450 vss.n10432 1118.26
R5388 vss.n10465 vss.n10432 1118.26
R5389 vss.n10465 vss.n10433 1118.26
R5390 vss.n10461 vss.n10433 1118.26
R5391 vss.n10593 vss.n10592 1118.26
R5392 vss.n10594 vss.n10593 1118.26
R5393 vss.n10594 vss.n10572 1118.26
R5394 vss.n10612 vss.n10572 1118.26
R5395 vss.n10612 vss.n10573 1118.26
R5396 vss.n10604 vss.n10573 1118.26
R5397 vss.n10590 vss.n10580 1118.26
R5398 vss.n10596 vss.n10580 1118.26
R5399 vss.n10596 vss.n10577 1118.26
R5400 vss.n10610 vss.n10577 1118.26
R5401 vss.n10610 vss.n10578 1118.26
R5402 vss.n10606 vss.n10578 1118.26
R5403 vss.n10987 vss.n10986 1118.26
R5404 vss.n10988 vss.n10987 1118.26
R5405 vss.n10988 vss.n10966 1118.26
R5406 vss.n11006 vss.n10966 1118.26
R5407 vss.n11006 vss.n10967 1118.26
R5408 vss.n10998 vss.n10967 1118.26
R5409 vss.n10984 vss.n10974 1118.26
R5410 vss.n10990 vss.n10974 1118.26
R5411 vss.n10990 vss.n10971 1118.26
R5412 vss.n11004 vss.n10971 1118.26
R5413 vss.n11004 vss.n10972 1118.26
R5414 vss.n11000 vss.n10972 1118.26
R5415 vss.n10003 vss.n9993 1118.26
R5416 vss.n10030 vss.n10003 1118.26
R5417 vss.n10030 vss.n10004 1118.26
R5418 vss.n10025 vss.n10004 1118.26
R5419 vss.n10025 vss.n10009 1118.26
R5420 vss.n10017 vss.n10009 1118.26
R5421 vss.n9998 vss.n9994 1118.26
R5422 vss.n10032 vss.n9998 1118.26
R5423 vss.n10032 vss.n9999 1118.26
R5424 vss.n10023 vss.n9999 1118.26
R5425 vss.n10023 vss.n10011 1118.26
R5426 vss.n10019 vss.n10011 1118.26
R5427 vss.n11792 vss.n11791 1090.43
R5428 vss.n9543 vss.n9282 1077.63
R5429 vss.n7222 vss.n435 1077.63
R5430 vss.n14073 vss.n1214 1077.63
R5431 vss.n6252 vss.n6203 1077.63
R5432 vss.n9851 vss.n9807 1068.57
R5433 vss.n9723 vss.n9678 1068.57
R5434 vss.n9593 vss.n9549 1068.57
R5435 vss.n5602 vss.n3535 1068.57
R5436 vss.n5912 vss.n5725 1068.57
R5437 vss.n6151 vss.n5965 1068.57
R5438 vss.n3523 vss.n3488 1068.57
R5439 vss.n4072 vss.n4000 1068.57
R5440 vss.n4253 vss.n3992 1068.57
R5441 vss.n7439 vss.n7395 1068.57
R5442 vss.n7269 vss.n7225 1068.57
R5443 vss.n2713 vss.n985 1068.57
R5444 vss.n3047 vss.n3012 1068.57
R5445 vss.n7059 vss.n3129 1068.57
R5446 vss.n13904 vss.n13860 1068.57
R5447 vss.n8143 vss.n8099 1068.57
R5448 vss.n13546 vss.n1764 1068.57
R5449 vss.n13848 vss.n8222 1068.57
R5450 vss.n9031 vss.n8094 1068.57
R5451 vss.n1813 vss.n1769 1068.57
R5452 vss.n1034 vss.n990 1068.57
R5453 vss.n11505 vss.n9802 1068.57
R5454 vss.n11100 vss.n9673 1068.57
R5455 vss.n10203 vss.n9544 1068.57
R5456 vss.n10352 vss.n10351 1054.53
R5457 vss.n10351 vss.n10349 1054.53
R5458 vss.n8876 vss.n8875 1054.53
R5459 vss.n8876 vss.n8872 1054.53
R5460 vss.n13190 vss.n13189 1054.53
R5461 vss.n13190 vss.n8873 1054.53
R5462 vss.n10291 vss.n10290 1054.53
R5463 vss.n10290 vss.n10287 1054.53
R5464 vss.n10317 vss.n10294 1054.53
R5465 vss.n10317 vss.n10288 1054.53
R5466 vss.n10312 vss.n10298 1054.53
R5467 vss.n10302 vss.n10298 1054.53
R5468 vss.n9958 vss.n9957 1054.53
R5469 vss.n9957 vss.n9954 1054.53
R5470 vss.n11639 vss.n9961 1054.53
R5471 vss.n11639 vss.n9955 1054.53
R5472 vss.n11634 vss.n11620 1054.53
R5473 vss.n11624 vss.n11620 1054.53
R5474 vss.n9918 vss.n9914 1054.53
R5475 vss.n9919 vss.n9918 1054.53
R5476 vss.n11686 vss.n9924 1054.53
R5477 vss.n9924 vss.n9922 1054.53
R5478 vss.n11692 vss.n9915 1054.53
R5479 vss.n11692 vss.n9920 1054.53
R5480 vss.n9973 vss.n9969 1054.53
R5481 vss.n9974 vss.n9973 1054.53
R5482 vss.n11449 vss.n9979 1054.53
R5483 vss.n9979 vss.n9977 1054.53
R5484 vss.n11455 vss.n9970 1054.53
R5485 vss.n11455 vss.n9975 1054.53
R5486 vss.n11380 vss.n11378 1054.53
R5487 vss.n11380 vss.n11373 1054.53
R5488 vss.n11377 vss.n11376 1054.53
R5489 vss.n11376 vss.n11372 1054.53
R5490 vss.n11386 vss.n11383 1054.53
R5491 vss.n11386 vss.n11385 1054.53
R5492 vss.n11164 vss.n11160 1054.53
R5493 vss.n11165 vss.n11164 1054.53
R5494 vss.n11180 vss.n11170 1054.53
R5495 vss.n11170 vss.n11168 1054.53
R5496 vss.n11186 vss.n11161 1054.53
R5497 vss.n11186 vss.n11166 1054.53
R5498 vss.n10133 vss.n10129 1054.53
R5499 vss.n10134 vss.n10133 1054.53
R5500 vss.n11044 vss.n10139 1054.53
R5501 vss.n10139 vss.n10137 1054.53
R5502 vss.n11050 vss.n10130 1054.53
R5503 vss.n11050 vss.n10135 1054.53
R5504 vss.n10087 vss.n10083 1054.53
R5505 vss.n10088 vss.n10087 1054.53
R5506 vss.n10104 vss.n10093 1054.53
R5507 vss.n10093 vss.n10091 1054.53
R5508 vss.n10110 vss.n10084 1054.53
R5509 vss.n10110 vss.n10089 1054.53
R5510 vss.n10743 vss.n10723 1054.53
R5511 vss.n10723 vss.n10717 1054.53
R5512 vss.n10721 vss.n10720 1054.53
R5513 vss.n10720 vss.n10716 1054.53
R5514 vss.n10728 vss.n10724 1054.53
R5515 vss.n10728 vss.n10727 1054.53
R5516 vss.n10220 vss.n10216 1054.53
R5517 vss.n10221 vss.n10220 1054.53
R5518 vss.n10792 vss.n10226 1054.53
R5519 vss.n10226 vss.n10224 1054.53
R5520 vss.n10798 vss.n10217 1054.53
R5521 vss.n10798 vss.n10222 1054.53
R5522 vss.n10668 vss.n10666 1054.53
R5523 vss.n10668 vss.n10661 1054.53
R5524 vss.n10665 vss.n10664 1054.53
R5525 vss.n10664 vss.n10660 1054.53
R5526 vss.n10674 vss.n10671 1054.53
R5527 vss.n10674 vss.n10673 1054.53
R5528 vss.n10262 vss.n10258 1054.53
R5529 vss.n10263 vss.n10262 1054.53
R5530 vss.n10402 vss.n10268 1054.53
R5531 vss.n10268 vss.n10266 1054.53
R5532 vss.n10408 vss.n10259 1054.53
R5533 vss.n10408 vss.n10264 1054.53
R5534 vss.n10431 vss.n10427 1054.53
R5535 vss.n10432 vss.n10431 1054.53
R5536 vss.n10494 vss.n10484 1054.53
R5537 vss.n10484 vss.n10482 1054.53
R5538 vss.n10478 vss.n10474 1054.53
R5539 vss.n10479 vss.n10478 1054.53
R5540 vss.n10500 vss.n10475 1054.53
R5541 vss.n10500 vss.n10480 1054.53
R5542 vss.n10543 vss.n10532 1054.53
R5543 vss.n10532 vss.n10530 1054.53
R5544 vss.n10526 vss.n10522 1054.53
R5545 vss.n10527 vss.n10526 1054.53
R5546 vss.n10549 vss.n10523 1054.53
R5547 vss.n10549 vss.n10528 1054.53
R5548 vss.n10841 vss.n10830 1054.53
R5549 vss.n10830 vss.n10828 1054.53
R5550 vss.n10824 vss.n10820 1054.53
R5551 vss.n10825 vss.n10824 1054.53
R5552 vss.n10847 vss.n10821 1054.53
R5553 vss.n10847 vss.n10826 1054.53
R5554 vss.n10888 vss.n10878 1054.53
R5555 vss.n10878 vss.n10876 1054.53
R5556 vss.n10872 vss.n10868 1054.53
R5557 vss.n10873 vss.n10872 1054.53
R5558 vss.n10894 vss.n10869 1054.53
R5559 vss.n10894 vss.n10874 1054.53
R5560 vss.n10937 vss.n10926 1054.53
R5561 vss.n10926 vss.n10924 1054.53
R5562 vss.n10920 vss.n10916 1054.53
R5563 vss.n10921 vss.n10920 1054.53
R5564 vss.n10943 vss.n10917 1054.53
R5565 vss.n10943 vss.n10922 1054.53
R5566 vss.n11276 vss.n11265 1054.53
R5567 vss.n11265 vss.n11263 1054.53
R5568 vss.n11259 vss.n11255 1054.53
R5569 vss.n11260 vss.n11259 1054.53
R5570 vss.n11282 vss.n11256 1054.53
R5571 vss.n11282 vss.n11261 1054.53
R5572 vss.n11227 vss.n11217 1054.53
R5573 vss.n11217 vss.n11215 1054.53
R5574 vss.n11211 vss.n11207 1054.53
R5575 vss.n11212 vss.n11211 1054.53
R5576 vss.n11233 vss.n11208 1054.53
R5577 vss.n11233 vss.n11213 1054.53
R5578 vss.n11134 vss.n11123 1054.53
R5579 vss.n11123 vss.n11121 1054.53
R5580 vss.n11117 vss.n11113 1054.53
R5581 vss.n11118 vss.n11117 1054.53
R5582 vss.n11140 vss.n11114 1054.53
R5583 vss.n11140 vss.n11119 1054.53
R5584 vss.n11587 vss.n11576 1054.53
R5585 vss.n11576 vss.n11574 1054.53
R5586 vss.n11570 vss.n11566 1054.53
R5587 vss.n11571 vss.n11570 1054.53
R5588 vss.n11593 vss.n11567 1054.53
R5589 vss.n11593 vss.n11572 1054.53
R5590 vss.n11538 vss.n11528 1054.53
R5591 vss.n11528 vss.n11526 1054.53
R5592 vss.n11522 vss.n11518 1054.53
R5593 vss.n11523 vss.n11522 1054.53
R5594 vss.n11544 vss.n11519 1054.53
R5595 vss.n11544 vss.n11524 1054.53
R5596 vss.n9895 vss.n9892 1054.53
R5597 vss.n9895 vss.n9894 1054.53
R5598 vss.n9889 vss.n9888 1054.53
R5599 vss.n9889 vss.n9885 1054.53
R5600 vss.n11716 vss.n11715 1054.53
R5601 vss.n11716 vss.n9886 1054.53
R5602 vss.n8823 vss.n8822 1054.53
R5603 vss.n8822 vss.n8818 1054.53
R5604 vss.n8824 vss.n8821 1054.53
R5605 vss.n8824 vss.n8817 1054.53
R5606 vss.n8830 vss.n8827 1054.53
R5607 vss.n8830 vss.n8829 1054.53
R5608 vss.n11778 vss.n11776 1054.53
R5609 vss.n11778 vss.n11762 1054.53
R5610 vss.n11774 vss.n11773 1054.53
R5611 vss.n11773 vss.n11761 1054.53
R5612 vss.n11768 vss.n11765 1054.53
R5613 vss.n11795 vss.n11765 1054.53
R5614 vss.n11823 vss.n11821 1054.53
R5615 vss.n11823 vss.n11807 1054.53
R5616 vss.n11818 vss.n11817 1054.53
R5617 vss.n11817 vss.n11806 1054.53
R5618 vss.n11835 vss.n11834 1054.53
R5619 vss.n11835 vss.n11812 1054.53
R5620 vss.n11901 vss.n11900 1054.53
R5621 vss.n11900 vss.n11896 1054.53
R5622 vss.n11902 vss.n11899 1054.53
R5623 vss.n11902 vss.n11895 1054.53
R5624 vss.n11908 vss.n11905 1054.53
R5625 vss.n11908 vss.n11907 1054.53
R5626 vss.n11741 vss.n9870 1054.53
R5627 vss.n11741 vss.n9865 1054.53
R5628 vss.n9869 vss.n9868 1054.53
R5629 vss.n9868 vss.n9864 1054.53
R5630 vss.n9874 vss.n9872 1054.53
R5631 vss.n11735 vss.n9874 1054.53
R5632 vss.n9453 vss.n9432 1054.53
R5633 vss.n9453 vss.n9427 1054.53
R5634 vss.n9431 vss.n9430 1054.53
R5635 vss.n9430 vss.n9426 1054.53
R5636 vss.n9436 vss.n9434 1054.53
R5637 vss.n9447 vss.n9436 1054.53
R5638 vss.n12484 vss.n9482 1054.53
R5639 vss.n12484 vss.n9477 1054.53
R5640 vss.n9481 vss.n9480 1054.53
R5641 vss.n9480 vss.n9476 1054.53
R5642 vss.n9486 vss.n9484 1054.53
R5643 vss.n12478 vss.n9486 1054.53
R5644 vss.n9516 vss.n9513 1054.53
R5645 vss.n9516 vss.n9515 1054.53
R5646 vss.n9510 vss.n9508 1054.53
R5647 vss.n9510 vss.n9503 1054.53
R5648 vss.n9507 vss.n9506 1054.53
R5649 vss.n9506 vss.n9502 1054.53
R5650 vss.n9569 vss.n9566 1054.53
R5651 vss.n9569 vss.n9568 1054.53
R5652 vss.n9563 vss.n9559 1054.53
R5653 vss.n9563 vss.n9554 1054.53
R5654 vss.n9558 vss.n9557 1054.53
R5655 vss.n9557 vss.n9550 1054.53
R5656 vss.n8895 vss.n8893 1054.53
R5657 vss.n8895 vss.n8888 1054.53
R5658 vss.n8892 vss.n8891 1054.53
R5659 vss.n8891 vss.n8887 1054.53
R5660 vss.n9268 vss.n9267 1054.53
R5661 vss.n9268 vss.n9259 1054.53
R5662 vss.n12411 vss.n12391 1054.53
R5663 vss.n12411 vss.n12386 1054.53
R5664 vss.n12390 vss.n12389 1054.53
R5665 vss.n12389 vss.n12385 1054.53
R5666 vss.n12395 vss.n12393 1054.53
R5667 vss.n12405 vss.n12395 1054.53
R5668 vss.n12446 vss.n12443 1054.53
R5669 vss.n12446 vss.n12445 1054.53
R5670 vss.n12440 vss.n12437 1054.53
R5671 vss.n12440 vss.n12433 1054.53
R5672 vss.n12365 vss.n9611 1054.53
R5673 vss.n12365 vss.n9606 1054.53
R5674 vss.n9610 vss.n9609 1054.53
R5675 vss.n9609 vss.n9605 1054.53
R5676 vss.n9615 vss.n9613 1054.53
R5677 vss.n12359 vss.n9615 1054.53
R5678 vss.n9645 vss.n9642 1054.53
R5679 vss.n9645 vss.n9644 1054.53
R5680 vss.n9639 vss.n9637 1054.53
R5681 vss.n9639 vss.n9632 1054.53
R5682 vss.n9636 vss.n9635 1054.53
R5683 vss.n9635 vss.n9631 1054.53
R5684 vss.n9698 vss.n9695 1054.53
R5685 vss.n9698 vss.n9697 1054.53
R5686 vss.n9692 vss.n9688 1054.53
R5687 vss.n9692 vss.n9683 1054.53
R5688 vss.n9687 vss.n9686 1054.53
R5689 vss.n9686 vss.n9679 1054.53
R5690 vss.n13273 vss.n8628 1054.53
R5691 vss.n13273 vss.n8623 1054.53
R5692 vss.n8627 vss.n8626 1054.53
R5693 vss.n8626 vss.n8622 1054.53
R5694 vss.n8632 vss.n8630 1054.53
R5695 vss.n13267 vss.n8632 1054.53
R5696 vss.n12293 vss.n12273 1054.53
R5697 vss.n12293 vss.n12268 1054.53
R5698 vss.n12272 vss.n12271 1054.53
R5699 vss.n12271 vss.n12267 1054.53
R5700 vss.n12277 vss.n12275 1054.53
R5701 vss.n12287 vss.n12277 1054.53
R5702 vss.n12327 vss.n12324 1054.53
R5703 vss.n12327 vss.n12326 1054.53
R5704 vss.n12321 vss.n12318 1054.53
R5705 vss.n12321 vss.n12314 1054.53
R5706 vss.n12247 vss.n9741 1054.53
R5707 vss.n12247 vss.n9736 1054.53
R5708 vss.n9740 vss.n9739 1054.53
R5709 vss.n9739 vss.n9735 1054.53
R5710 vss.n9745 vss.n9743 1054.53
R5711 vss.n12241 vss.n9745 1054.53
R5712 vss.n9775 vss.n9772 1054.53
R5713 vss.n9775 vss.n9774 1054.53
R5714 vss.n9769 vss.n9767 1054.53
R5715 vss.n9769 vss.n9762 1054.53
R5716 vss.n9766 vss.n9765 1054.53
R5717 vss.n9765 vss.n9761 1054.53
R5718 vss.n9827 vss.n9824 1054.53
R5719 vss.n9827 vss.n9826 1054.53
R5720 vss.n9821 vss.n9817 1054.53
R5721 vss.n9821 vss.n9812 1054.53
R5722 vss.n9816 vss.n9815 1054.53
R5723 vss.n9815 vss.n9808 1054.53
R5724 vss.n8351 vss.n8349 1054.53
R5725 vss.n8351 vss.n8344 1054.53
R5726 vss.n8348 vss.n8347 1054.53
R5727 vss.n8347 vss.n8343 1054.53
R5728 vss.n8750 vss.n8749 1054.53
R5729 vss.n8750 vss.n8741 1054.53
R5730 vss.n11974 vss.n11973 1054.53
R5731 vss.n11973 vss.n11969 1054.53
R5732 vss.n11975 vss.n11972 1054.53
R5733 vss.n11975 vss.n11968 1054.53
R5734 vss.n11981 vss.n11978 1054.53
R5735 vss.n11981 vss.n11980 1054.53
R5736 vss.n12209 vss.n12206 1054.53
R5737 vss.n12209 vss.n12208 1054.53
R5738 vss.n12203 vss.n12200 1054.53
R5739 vss.n12203 vss.n12196 1054.53
R5740 vss.n12199 vss.n12198 1054.53
R5741 vss.n12198 vss.n9855 1054.53
R5742 vss.n8778 vss.n8775 1054.53
R5743 vss.n8778 vss.n8777 1054.53
R5744 vss.n8772 vss.n8769 1054.53
R5745 vss.n8772 vss.n8765 1054.53
R5746 vss.n8768 vss.n8767 1054.53
R5747 vss.n8767 vss.n8760 1054.53
R5748 vss.n8709 vss.n8706 1054.53
R5749 vss.n8709 vss.n8708 1054.53
R5750 vss.n8703 vss.n8700 1054.53
R5751 vss.n8703 vss.n8696 1054.53
R5752 vss.n8699 vss.n8698 1054.53
R5753 vss.n8698 vss.n8692 1054.53
R5754 vss.n12317 vss.n12316 1054.53
R5755 vss.n12316 vss.n9727 1054.53
R5756 vss.n8659 vss.n8656 1054.53
R5757 vss.n8659 vss.n8658 1054.53
R5758 vss.n8653 vss.n8650 1054.53
R5759 vss.n8653 vss.n8646 1054.53
R5760 vss.n8649 vss.n8648 1054.53
R5761 vss.n8648 vss.n8641 1054.53
R5762 vss.n9194 vss.n9193 1054.53
R5763 vss.n9193 vss.n9189 1054.53
R5764 vss.n9195 vss.n9192 1054.53
R5765 vss.n9195 vss.n9188 1054.53
R5766 vss.n9201 vss.n9198 1054.53
R5767 vss.n9201 vss.n9200 1054.53
R5768 vss.n12436 vss.n12435 1054.53
R5769 vss.n12435 vss.n9597 1054.53
R5770 vss.n9229 vss.n9226 1054.53
R5771 vss.n9229 vss.n9228 1054.53
R5772 vss.n9223 vss.n9220 1054.53
R5773 vss.n9223 vss.n9216 1054.53
R5774 vss.n9219 vss.n9218 1054.53
R5775 vss.n9218 vss.n9211 1054.53
R5776 vss.n9324 vss.n9323 1054.53
R5777 vss.n9323 vss.n9319 1054.53
R5778 vss.n9325 vss.n9322 1054.53
R5779 vss.n9325 vss.n9318 1054.53
R5780 vss.n9331 vss.n9328 1054.53
R5781 vss.n9331 vss.n9330 1054.53
R5782 vss.n12510 vss.n12509 1054.53
R5783 vss.n12509 vss.n12505 1054.53
R5784 vss.n12511 vss.n12508 1054.53
R5785 vss.n12511 vss.n12504 1054.53
R5786 vss.n12517 vss.n12514 1054.53
R5787 vss.n12517 vss.n12516 1054.53
R5788 vss.n12660 vss.n12659 1054.53
R5789 vss.n12659 vss.n12655 1054.53
R5790 vss.n12661 vss.n12658 1054.53
R5791 vss.n12661 vss.n12654 1054.53
R5792 vss.n12667 vss.n12664 1054.53
R5793 vss.n12667 vss.n12666 1054.53
R5794 vss.n10176 vss.n10172 1054.53
R5795 vss.n10177 vss.n10176 1054.53
R5796 vss.n10192 vss.n10182 1054.53
R5797 vss.n10182 vss.n10180 1054.53
R5798 vss.n10198 vss.n10173 1054.53
R5799 vss.n10198 vss.n10178 1054.53
R5800 vss.n11073 vss.n11069 1054.53
R5801 vss.n11074 vss.n11073 1054.53
R5802 vss.n11089 vss.n11079 1054.53
R5803 vss.n11079 vss.n11077 1054.53
R5804 vss.n11095 vss.n11070 1054.53
R5805 vss.n11095 vss.n11075 1054.53
R5806 vss.n11478 vss.n11474 1054.53
R5807 vss.n11479 vss.n11478 1054.53
R5808 vss.n11494 vss.n11484 1054.53
R5809 vss.n11484 vss.n11482 1054.53
R5810 vss.n11500 vss.n11475 1054.53
R5811 vss.n11500 vss.n11480 1054.53
R5812 vss.n12155 vss.n12152 1054.53
R5813 vss.n12155 vss.n12154 1054.53
R5814 vss.n12149 vss.n12147 1054.53
R5815 vss.n12149 vss.n12142 1054.53
R5816 vss.n12146 vss.n12145 1054.53
R5817 vss.n12145 vss.n12141 1054.53
R5818 vss.n15559 vss.n369 1054.53
R5819 vss.n15559 vss.n364 1054.53
R5820 vss.n368 vss.n367 1054.53
R5821 vss.n367 vss.n363 1054.53
R5822 vss.n15626 vss.n15625 1054.53
R5823 vss.n15625 vss.n358 1054.53
R5824 vss.n15630 vss.n15629 1054.53
R5825 vss.n15630 vss.n357 1054.53
R5826 vss.n15634 vss.n15632 1054.53
R5827 vss.n15634 vss.n15633 1054.53
R5828 vss.n3576 vss.n3575 1054.53
R5829 vss.n3575 vss.n3571 1054.53
R5830 vss.n3577 vss.n3574 1054.53
R5831 vss.n3577 vss.n3570 1054.53
R5832 vss.n3583 vss.n3580 1054.53
R5833 vss.n3583 vss.n3582 1054.53
R5834 vss.n324 vss.n321 1054.53
R5835 vss.n324 vss.n323 1054.53
R5836 vss.n318 vss.n315 1054.53
R5837 vss.n318 vss.n311 1054.53
R5838 vss.n11 vss.n9 1054.53
R5839 vss.n11 vss.n4 1054.53
R5840 vss.n8 vss.n7 1054.53
R5841 vss.n7 vss.n3 1054.53
R5842 vss.n3981 vss.n3974 1054.53
R5843 vss.n3981 vss.n3975 1054.53
R5844 vss.n255 vss.n253 1054.53
R5845 vss.n255 vss.n248 1054.53
R5846 vss.n252 vss.n251 1054.53
R5847 vss.n251 vss.n247 1054.53
R5848 vss.n6303 vss.n6296 1054.53
R5849 vss.n6303 vss.n6297 1054.53
R5850 vss.n5661 vss.n5641 1054.53
R5851 vss.n5661 vss.n5636 1054.53
R5852 vss.n5640 vss.n5639 1054.53
R5853 vss.n5639 vss.n5635 1054.53
R5854 vss.n5645 vss.n5643 1054.53
R5855 vss.n5655 vss.n5645 1054.53
R5856 vss.n176 vss.n174 1054.53
R5857 vss.n176 vss.n169 1054.53
R5858 vss.n173 vss.n172 1054.53
R5859 vss.n172 vss.n168 1054.53
R5860 vss.n3722 vss.n3721 1054.53
R5861 vss.n3722 vss.n3713 1054.53
R5862 vss.n3683 vss.n3680 1054.53
R5863 vss.n3683 vss.n3682 1054.53
R5864 vss.n3677 vss.n3674 1054.53
R5865 vss.n3677 vss.n3670 1054.53
R5866 vss.n3673 vss.n3672 1054.53
R5867 vss.n3672 vss.n3666 1054.53
R5868 vss.n5853 vss.n5833 1054.53
R5869 vss.n5853 vss.n5828 1054.53
R5870 vss.n5832 vss.n5831 1054.53
R5871 vss.n5831 vss.n5827 1054.53
R5872 vss.n5837 vss.n5835 1054.53
R5873 vss.n5847 vss.n5837 1054.53
R5874 vss.n98 vss.n96 1054.53
R5875 vss.n98 vss.n91 1054.53
R5876 vss.n95 vss.n94 1054.53
R5877 vss.n94 vss.n90 1054.53
R5878 vss.n3841 vss.n3840 1054.53
R5879 vss.n3841 vss.n3832 1054.53
R5880 vss.n3802 vss.n3799 1054.53
R5881 vss.n3802 vss.n3801 1054.53
R5882 vss.n3796 vss.n3793 1054.53
R5883 vss.n3796 vss.n3789 1054.53
R5884 vss.n3792 vss.n3791 1054.53
R5885 vss.n3791 vss.n3785 1054.53
R5886 vss.n3921 vss.n3918 1054.53
R5887 vss.n3921 vss.n3920 1054.53
R5888 vss.n3915 vss.n3912 1054.53
R5889 vss.n3915 vss.n3908 1054.53
R5890 vss.n3911 vss.n3910 1054.53
R5891 vss.n3910 vss.n3904 1054.53
R5892 vss.n6093 vss.n6073 1054.53
R5893 vss.n6093 vss.n6068 1054.53
R5894 vss.n6072 vss.n6071 1054.53
R5895 vss.n6071 vss.n6067 1054.53
R5896 vss.n6077 vss.n6075 1054.53
R5897 vss.n6087 vss.n6077 1054.53
R5898 vss.n6225 vss.n6222 1054.53
R5899 vss.n6225 vss.n6224 1054.53
R5900 vss.n6219 vss.n6216 1054.53
R5901 vss.n6219 vss.n6212 1054.53
R5902 vss.n6045 vss.n6025 1054.53
R5903 vss.n6045 vss.n6020 1054.53
R5904 vss.n6024 vss.n6023 1054.53
R5905 vss.n6023 vss.n6019 1054.53
R5906 vss.n6029 vss.n6027 1054.53
R5907 vss.n6039 vss.n6029 1054.53
R5908 vss.n6173 vss.n6170 1054.53
R5909 vss.n6173 vss.n6172 1054.53
R5910 vss.n6167 vss.n6165 1054.53
R5911 vss.n6167 vss.n6160 1054.53
R5912 vss.n6164 vss.n6163 1054.53
R5913 vss.n6163 vss.n6159 1054.53
R5914 vss.n5759 vss.n5738 1054.53
R5915 vss.n5759 vss.n5733 1054.53
R5916 vss.n5737 vss.n5736 1054.53
R5917 vss.n5736 vss.n5732 1054.53
R5918 vss.n5742 vss.n5740 1054.53
R5919 vss.n5753 vss.n5742 1054.53
R5920 vss.n5805 vss.n5785 1054.53
R5921 vss.n5805 vss.n5780 1054.53
R5922 vss.n5784 vss.n5783 1054.53
R5923 vss.n5783 vss.n5779 1054.53
R5924 vss.n5789 vss.n5787 1054.53
R5925 vss.n5799 vss.n5789 1054.53
R5926 vss.n5934 vss.n5931 1054.53
R5927 vss.n5934 vss.n5933 1054.53
R5928 vss.n5928 vss.n5926 1054.53
R5929 vss.n5928 vss.n5921 1054.53
R5930 vss.n5925 vss.n5924 1054.53
R5931 vss.n5924 vss.n5920 1054.53
R5932 vss.n5571 vss.n5550 1054.53
R5933 vss.n5571 vss.n5545 1054.53
R5934 vss.n5549 vss.n5548 1054.53
R5935 vss.n5548 vss.n5544 1054.53
R5936 vss.n5554 vss.n5552 1054.53
R5937 vss.n5565 vss.n5554 1054.53
R5938 vss.n5696 vss.n5693 1054.53
R5939 vss.n5696 vss.n5695 1054.53
R5940 vss.n5690 vss.n5688 1054.53
R5941 vss.n5690 vss.n5683 1054.53
R5942 vss.n5687 vss.n5686 1054.53
R5943 vss.n5686 vss.n5682 1054.53
R5944 vss.n3557 vss.n3554 1054.53
R5945 vss.n3557 vss.n3556 1054.53
R5946 vss.n3551 vss.n3549 1054.53
R5947 vss.n3551 vss.n3544 1054.53
R5948 vss.n3548 vss.n3547 1054.53
R5949 vss.n3547 vss.n3543 1054.53
R5950 vss.n5616 vss.n5597 1054.53
R5951 vss.n5616 vss.n5592 1054.53
R5952 vss.n5596 vss.n5595 1054.53
R5953 vss.n5595 vss.n5591 1054.53
R5954 vss.n5601 vss.n5599 1054.53
R5955 vss.n5610 vss.n5601 1054.53
R5956 vss.n5888 vss.n5885 1054.53
R5957 vss.n5888 vss.n5887 1054.53
R5958 vss.n5882 vss.n5878 1054.53
R5959 vss.n5882 vss.n5873 1054.53
R5960 vss.n5877 vss.n5876 1054.53
R5961 vss.n5876 vss.n5726 1054.53
R5962 vss.n6127 vss.n6124 1054.53
R5963 vss.n6127 vss.n6126 1054.53
R5964 vss.n6121 vss.n6117 1054.53
R5965 vss.n6121 vss.n6112 1054.53
R5966 vss.n6116 vss.n6115 1054.53
R5967 vss.n6115 vss.n5966 1054.53
R5968 vss.n5999 vss.n5978 1054.53
R5969 vss.n5999 vss.n5973 1054.53
R5970 vss.n5977 vss.n5976 1054.53
R5971 vss.n5976 vss.n5972 1054.53
R5972 vss.n5982 vss.n5980 1054.53
R5973 vss.n5993 vss.n5982 1054.53
R5974 vss.n3303 vss.n3278 1054.53
R5975 vss.n3303 vss.n3283 1054.53
R5976 vss.n3281 vss.n3277 1054.53
R5977 vss.n3282 vss.n3281 1054.53
R5978 vss.n3297 vss.n3287 1054.53
R5979 vss.n3287 vss.n3285 1054.53
R5980 vss.n4380 vss.n4378 1054.53
R5981 vss.n4380 vss.n4373 1054.53
R5982 vss.n4377 vss.n4376 1054.53
R5983 vss.n4376 vss.n4372 1054.53
R5984 vss.n4386 vss.n4383 1054.53
R5985 vss.n4386 vss.n4385 1054.53
R5986 vss.n4408 vss.n4404 1054.53
R5987 vss.n4409 vss.n4408 1054.53
R5988 vss.n4470 vss.n4460 1054.53
R5989 vss.n4460 vss.n4458 1054.53
R5990 vss.n4454 vss.n4450 1054.53
R5991 vss.n4455 vss.n4454 1054.53
R5992 vss.n4476 vss.n4451 1054.53
R5993 vss.n4476 vss.n4456 1054.53
R5994 vss.n4518 vss.n4507 1054.53
R5995 vss.n4507 vss.n4505 1054.53
R5996 vss.n4501 vss.n4497 1054.53
R5997 vss.n4502 vss.n4501 1054.53
R5998 vss.n4524 vss.n4498 1054.53
R5999 vss.n4524 vss.n4503 1054.53
R6000 vss.n5023 vss.n5012 1054.53
R6001 vss.n5012 vss.n5010 1054.53
R6002 vss.n5006 vss.n5002 1054.53
R6003 vss.n5007 vss.n5006 1054.53
R6004 vss.n5029 vss.n5003 1054.53
R6005 vss.n5029 vss.n5008 1054.53
R6006 vss.n4195 vss.n4185 1054.53
R6007 vss.n4185 vss.n4183 1054.53
R6008 vss.n4198 vss.n4197 1054.53
R6009 vss.n4198 vss.n4181 1054.53
R6010 vss.n4209 vss.n4178 1054.53
R6011 vss.n4209 vss.n4208 1054.53
R6012 vss.n5071 vss.n5060 1054.53
R6013 vss.n5060 vss.n5058 1054.53
R6014 vss.n5054 vss.n5050 1054.53
R6015 vss.n5055 vss.n5054 1054.53
R6016 vss.n5077 vss.n5051 1054.53
R6017 vss.n5077 vss.n5056 1054.53
R6018 vss.n5497 vss.n5486 1054.53
R6019 vss.n5486 vss.n5484 1054.53
R6020 vss.n5480 vss.n5476 1054.53
R6021 vss.n5481 vss.n5480 1054.53
R6022 vss.n5503 vss.n5477 1054.53
R6023 vss.n5503 vss.n5482 1054.53
R6024 vss.n4022 vss.n4019 1054.53
R6025 vss.n4022 vss.n4021 1054.53
R6026 vss.n4016 vss.n4015 1054.53
R6027 vss.n4016 vss.n4012 1054.53
R6028 vss.n4011 vss.n4006 1054.53
R6029 vss.n5527 vss.n4011 1054.53
R6030 vss.n5282 vss.n5271 1054.53
R6031 vss.n5271 vss.n5269 1054.53
R6032 vss.n5265 vss.n5261 1054.53
R6033 vss.n5266 vss.n5265 1054.53
R6034 vss.n5288 vss.n5262 1054.53
R6035 vss.n5288 vss.n5267 1054.53
R6036 vss.n3456 vss.n3452 1054.53
R6037 vss.n3456 vss.n3455 1054.53
R6038 vss.n3472 vss.n3451 1054.53
R6039 vss.n3451 vss.n3447 1054.53
R6040 vss.n3477 vss.n3476 1054.53
R6041 vss.n3477 vss.n3448 1054.53
R6042 vss.n6356 vss.n6341 1054.53
R6043 vss.n6345 vss.n6341 1054.53
R6044 vss.n6359 vss.n6358 1054.53
R6045 vss.n6359 vss.n6339 1054.53
R6046 vss.n6336 vss.n3439 1054.53
R6047 vss.n6337 vss.n6336 1054.53
R6048 vss.n6666 vss.n3338 1054.53
R6049 vss.n6667 vss.n6666 1054.53
R6050 vss.n6672 vss.n6664 1054.53
R6051 vss.n6672 vss.n6668 1054.53
R6052 vss.n6688 vss.n6678 1054.53
R6053 vss.n6688 vss.n6675 1054.53
R6054 vss.n6622 vss.n6618 1054.53
R6055 vss.n6623 vss.n6622 1054.53
R6056 vss.n6638 vss.n6628 1054.53
R6057 vss.n6628 vss.n6626 1054.53
R6058 vss.n6644 vss.n6619 1054.53
R6059 vss.n6644 vss.n6624 1054.53
R6060 vss.n6504 vss.n6500 1054.53
R6061 vss.n6505 vss.n6504 1054.53
R6062 vss.n6589 vss.n6510 1054.53
R6063 vss.n6510 vss.n6508 1054.53
R6064 vss.n6595 vss.n6501 1054.53
R6065 vss.n6595 vss.n6506 1054.53
R6066 vss.n5220 vss.n5216 1054.53
R6067 vss.n5221 vss.n5220 1054.53
R6068 vss.n5236 vss.n5226 1054.53
R6069 vss.n5226 vss.n5224 1054.53
R6070 vss.n5242 vss.n5217 1054.53
R6071 vss.n5242 vss.n5222 1054.53
R6072 vss.n4045 vss.n4041 1054.53
R6073 vss.n4046 vss.n4045 1054.53
R6074 vss.n4061 vss.n4051 1054.53
R6075 vss.n4051 vss.n4049 1054.53
R6076 vss.n4067 vss.n4042 1054.53
R6077 vss.n4067 vss.n4047 1054.53
R6078 vss.n5432 vss.n5428 1054.53
R6079 vss.n5433 vss.n5432 1054.53
R6080 vss.n5448 vss.n5438 1054.53
R6081 vss.n5438 vss.n5436 1054.53
R6082 vss.n5454 vss.n5429 1054.53
R6083 vss.n5454 vss.n5434 1054.53
R6084 vss.n5317 vss.n5313 1054.53
R6085 vss.n5318 vss.n5317 1054.53
R6086 vss.n5401 vss.n5323 1054.53
R6087 vss.n5323 vss.n5321 1054.53
R6088 vss.n5407 vss.n5314 1054.53
R6089 vss.n5407 vss.n5319 1054.53
R6090 vss.n4135 vss.n4131 1054.53
R6091 vss.n4136 vss.n4135 1054.53
R6092 vss.n4151 vss.n4141 1054.53
R6093 vss.n4141 vss.n4139 1054.53
R6094 vss.n4157 vss.n4132 1054.53
R6095 vss.n4157 vss.n4137 1054.53
R6096 vss.n4226 vss.n4222 1054.53
R6097 vss.n4227 vss.n4226 1054.53
R6098 vss.n4242 vss.n4232 1054.53
R6099 vss.n4232 vss.n4230 1054.53
R6100 vss.n4248 vss.n4223 1054.53
R6101 vss.n4248 vss.n4228 1054.53
R6102 vss.n4958 vss.n4954 1054.53
R6103 vss.n4959 vss.n4958 1054.53
R6104 vss.n4974 vss.n4964 1054.53
R6105 vss.n4964 vss.n4962 1054.53
R6106 vss.n4980 vss.n4955 1054.53
R6107 vss.n4980 vss.n4960 1054.53
R6108 vss.n4089 vss.n4085 1054.53
R6109 vss.n4090 vss.n4089 1054.53
R6110 vss.n4105 vss.n4095 1054.53
R6111 vss.n4095 vss.n4093 1054.53
R6112 vss.n4111 vss.n4086 1054.53
R6113 vss.n4111 vss.n4091 1054.53
R6114 vss.n4272 vss.n4268 1054.53
R6115 vss.n4273 vss.n4272 1054.53
R6116 vss.n4926 vss.n4278 1054.53
R6117 vss.n4278 vss.n4276 1054.53
R6118 vss.n4932 vss.n4269 1054.53
R6119 vss.n4932 vss.n4274 1054.53
R6120 vss.n5105 vss.n5101 1054.53
R6121 vss.n5106 vss.n5105 1054.53
R6122 vss.n5189 vss.n5111 1054.53
R6123 vss.n5111 vss.n5109 1054.53
R6124 vss.n5195 vss.n5102 1054.53
R6125 vss.n5195 vss.n5107 1054.53
R6126 vss.n3348 vss.n3344 1054.53
R6127 vss.n3349 vss.n3348 1054.53
R6128 vss.n3364 vss.n3354 1054.53
R6129 vss.n3354 vss.n3352 1054.53
R6130 vss.n3370 vss.n3345 1054.53
R6131 vss.n3370 vss.n3350 1054.53
R6132 vss.n3395 vss.n3391 1054.53
R6133 vss.n3396 vss.n3395 1054.53
R6134 vss.n3411 vss.n3401 1054.53
R6135 vss.n3401 vss.n3399 1054.53
R6136 vss.n3417 vss.n3392 1054.53
R6137 vss.n3417 vss.n3397 1054.53
R6138 vss.n3498 vss.n3497 1054.53
R6139 vss.n3498 vss.n3494 1054.53
R6140 vss.n3504 vss.n3501 1054.53
R6141 vss.n3504 vss.n3503 1054.53
R6142 vss.n3525 vss.n3524 1054.53
R6143 vss.n3525 vss.n3495 1054.53
R6144 vss.n6389 vss.n6385 1054.53
R6145 vss.n6390 vss.n6389 1054.53
R6146 vss.n6473 vss.n6395 1054.53
R6147 vss.n6395 vss.n6393 1054.53
R6148 vss.n6479 vss.n6386 1054.53
R6149 vss.n6479 vss.n6391 1054.53
R6150 vss.n4424 vss.n4414 1054.53
R6151 vss.n4414 vss.n4412 1054.53
R6152 vss.n4430 vss.n4405 1054.53
R6153 vss.n4430 vss.n4410 1054.53
R6154 vss.n4767 vss.n4765 1054.53
R6155 vss.n4767 vss.n4760 1054.53
R6156 vss.n4764 vss.n4763 1054.53
R6157 vss.n4763 vss.n4759 1054.53
R6158 vss.n4773 vss.n4770 1054.53
R6159 vss.n4773 vss.n4772 1054.53
R6160 vss.n14998 vss.n14996 1054.53
R6161 vss.n14998 vss.n14982 1054.53
R6162 vss.n14993 vss.n14992 1054.53
R6163 vss.n14992 vss.n14981 1054.53
R6164 vss.n15010 vss.n15009 1054.53
R6165 vss.n15010 vss.n14987 1054.53
R6166 vss.n15508 vss.n15507 1054.53
R6167 vss.n15507 vss.n15503 1054.53
R6168 vss.n15509 vss.n15506 1054.53
R6169 vss.n15509 vss.n15502 1054.53
R6170 vss.n15515 vss.n15512 1054.53
R6171 vss.n15515 vss.n15514 1054.53
R6172 vss.n400 vss.n398 1054.53
R6173 vss.n400 vss.n393 1054.53
R6174 vss.n397 vss.n396 1054.53
R6175 vss.n396 vss.n392 1054.53
R6176 vss.n14862 vss.n14855 1054.53
R6177 vss.n14862 vss.n14856 1054.53
R6178 vss.n14944 vss.n14940 1054.53
R6179 vss.n14972 vss.n14940 1054.53
R6180 vss.n14949 vss.n14948 1054.53
R6181 vss.n14948 vss.n14939 1054.53
R6182 vss.n14954 vss.n14953 1054.53
R6183 vss.n14956 vss.n14954 1054.53
R6184 vss.n1070 vss.n1050 1054.53
R6185 vss.n1070 vss.n1045 1054.53
R6186 vss.n1049 vss.n1048 1054.53
R6187 vss.n1048 vss.n1044 1054.53
R6188 vss.n1054 vss.n1052 1054.53
R6189 vss.n1064 vss.n1054 1054.53
R6190 vss.n15066 vss.n15063 1054.53
R6191 vss.n15066 vss.n15065 1054.53
R6192 vss.n15060 vss.n15057 1054.53
R6193 vss.n15060 vss.n15053 1054.53
R6194 vss.n1010 vss.n1007 1054.53
R6195 vss.n1010 vss.n1009 1054.53
R6196 vss.n15155 vss.n975 1054.53
R6197 vss.n15155 vss.n970 1054.53
R6198 vss.n974 vss.n973 1054.53
R6199 vss.n973 vss.n969 1054.53
R6200 vss.n979 vss.n977 1054.53
R6201 vss.n15149 vss.n979 1054.53
R6202 vss.n14919 vss.n14897 1054.53
R6203 vss.n14919 vss.n14892 1054.53
R6204 vss.n14896 vss.n14895 1054.53
R6205 vss.n14895 vss.n14891 1054.53
R6206 vss.n14901 vss.n14899 1054.53
R6207 vss.n14913 vss.n14901 1054.53
R6208 vss.n4589 vss.n4568 1054.53
R6209 vss.n4589 vss.n4563 1054.53
R6210 vss.n4567 vss.n4566 1054.53
R6211 vss.n4566 vss.n4562 1054.53
R6212 vss.n4572 vss.n4570 1054.53
R6213 vss.n4583 vss.n4572 1054.53
R6214 vss.n4685 vss.n4664 1054.53
R6215 vss.n4685 vss.n4659 1054.53
R6216 vss.n4663 vss.n4662 1054.53
R6217 vss.n4662 vss.n4658 1054.53
R6218 vss.n4668 vss.n4666 1054.53
R6219 vss.n4679 vss.n4668 1054.53
R6220 vss.n4636 vss.n4616 1054.53
R6221 vss.n4636 vss.n4611 1054.53
R6222 vss.n4615 vss.n4614 1054.53
R6223 vss.n4614 vss.n4610 1054.53
R6224 vss.n4620 vss.n4618 1054.53
R6225 vss.n4630 vss.n4620 1054.53
R6226 vss.n7245 vss.n7242 1054.53
R6227 vss.n7245 vss.n7244 1054.53
R6228 vss.n7239 vss.n7235 1054.53
R6229 vss.n7239 vss.n7230 1054.53
R6230 vss.n7234 vss.n7233 1054.53
R6231 vss.n7233 vss.n7226 1054.53
R6232 vss.n532 vss.n512 1054.53
R6233 vss.n532 vss.n507 1054.53
R6234 vss.n511 vss.n510 1054.53
R6235 vss.n510 vss.n506 1054.53
R6236 vss.n516 vss.n514 1054.53
R6237 vss.n526 vss.n516 1054.53
R6238 vss.n7330 vss.n7310 1054.53
R6239 vss.n7330 vss.n7305 1054.53
R6240 vss.n7309 vss.n7308 1054.53
R6241 vss.n7308 vss.n7304 1054.53
R6242 vss.n7314 vss.n7312 1054.53
R6243 vss.n7324 vss.n7314 1054.53
R6244 vss.n7283 vss.n3119 1054.53
R6245 vss.n7283 vss.n3114 1054.53
R6246 vss.n3118 vss.n3117 1054.53
R6247 vss.n3117 vss.n3113 1054.53
R6248 vss.n3094 vss.n3073 1054.53
R6249 vss.n3094 vss.n3068 1054.53
R6250 vss.n3072 vss.n3071 1054.53
R6251 vss.n3071 vss.n3067 1054.53
R6252 vss.n3077 vss.n3075 1054.53
R6253 vss.n3088 vss.n3077 1054.53
R6254 vss.n7366 vss.n7363 1054.53
R6255 vss.n7366 vss.n7365 1054.53
R6256 vss.n7360 vss.n7358 1054.53
R6257 vss.n7360 vss.n7353 1054.53
R6258 vss.n7357 vss.n7356 1054.53
R6259 vss.n7356 vss.n7352 1054.53
R6260 vss.n7415 vss.n7412 1054.53
R6261 vss.n7415 vss.n7414 1054.53
R6262 vss.n7409 vss.n7405 1054.53
R6263 vss.n7409 vss.n7400 1054.53
R6264 vss.n7404 vss.n7403 1054.53
R6265 vss.n7403 vss.n7396 1054.53
R6266 vss.n737 vss.n717 1054.53
R6267 vss.n737 vss.n712 1054.53
R6268 vss.n716 vss.n715 1054.53
R6269 vss.n715 vss.n711 1054.53
R6270 vss.n721 vss.n719 1054.53
R6271 vss.n731 vss.n721 1054.53
R6272 vss.n790 vss.n770 1054.53
R6273 vss.n790 vss.n765 1054.53
R6274 vss.n769 vss.n768 1054.53
R6275 vss.n768 vss.n764 1054.53
R6276 vss.n774 vss.n772 1054.53
R6277 vss.n784 vss.n774 1054.53
R6278 vss.n7461 vss.n7458 1054.53
R6279 vss.n7461 vss.n7460 1054.53
R6280 vss.n7455 vss.n7452 1054.53
R6281 vss.n7455 vss.n7448 1054.53
R6282 vss.n15117 vss.n15114 1054.53
R6283 vss.n15117 vss.n15116 1054.53
R6284 vss.n15111 vss.n15106 1054.53
R6285 vss.n15111 vss.n15101 1054.53
R6286 vss.n15105 vss.n15104 1054.53
R6287 vss.n15104 vss.n15097 1054.53
R6288 vss.n15204 vss.n15184 1054.53
R6289 vss.n15204 vss.n15179 1054.53
R6290 vss.n15183 vss.n15182 1054.53
R6291 vss.n15182 vss.n15178 1054.53
R6292 vss.n15188 vss.n15186 1054.53
R6293 vss.n15198 vss.n15188 1054.53
R6294 vss.n947 vss.n927 1054.53
R6295 vss.n947 vss.n922 1054.53
R6296 vss.n926 vss.n925 1054.53
R6297 vss.n925 vss.n921 1054.53
R6298 vss.n931 vss.n929 1054.53
R6299 vss.n941 vss.n931 1054.53
R6300 vss.n817 vss.n816 1054.53
R6301 vss.n816 vss.n812 1054.53
R6302 vss.n818 vss.n815 1054.53
R6303 vss.n818 vss.n811 1054.53
R6304 vss.n824 vss.n821 1054.53
R6305 vss.n824 vss.n823 1054.53
R6306 vss.n7451 vss.n7450 1054.53
R6307 vss.n7450 vss.n7443 1054.53
R6308 vss.n15324 vss.n15304 1054.53
R6309 vss.n15324 vss.n15299 1054.53
R6310 vss.n15303 vss.n15302 1054.53
R6311 vss.n15302 vss.n15298 1054.53
R6312 vss.n15308 vss.n15306 1054.53
R6313 vss.n15318 vss.n15308 1054.53
R6314 vss.n690 vss.n670 1054.53
R6315 vss.n690 vss.n665 1054.53
R6316 vss.n669 vss.n668 1054.53
R6317 vss.n668 vss.n664 1054.53
R6318 vss.n674 vss.n672 1054.53
R6319 vss.n684 vss.n674 1054.53
R6320 vss.n3123 vss.n3121 1054.53
R6321 vss.n7277 vss.n3123 1054.53
R6322 vss.n560 vss.n559 1054.53
R6323 vss.n559 vss.n555 1054.53
R6324 vss.n561 vss.n558 1054.53
R6325 vss.n561 vss.n554 1054.53
R6326 vss.n567 vss.n564 1054.53
R6327 vss.n567 vss.n566 1054.53
R6328 vss.n482 vss.n462 1054.53
R6329 vss.n482 vss.n457 1054.53
R6330 vss.n461 vss.n460 1054.53
R6331 vss.n460 vss.n456 1054.53
R6332 vss.n466 vss.n464 1054.53
R6333 vss.n476 vss.n466 1054.53
R6334 vss.n4711 vss.n4710 1054.53
R6335 vss.n4710 vss.n4706 1054.53
R6336 vss.n4712 vss.n4709 1054.53
R6337 vss.n4712 vss.n4705 1054.53
R6338 vss.n4718 vss.n4715 1054.53
R6339 vss.n4718 vss.n4717 1054.53
R6340 vss.n4326 vss.n4325 1054.53
R6341 vss.n4325 vss.n4321 1054.53
R6342 vss.n4327 vss.n4324 1054.53
R6343 vss.n4327 vss.n4320 1054.53
R6344 vss.n4333 vss.n4330 1054.53
R6345 vss.n4333 vss.n4332 1054.53
R6346 vss.n6768 vss.n6758 1054.53
R6347 vss.n6758 vss.n6756 1054.53
R6348 vss.n6752 vss.n6748 1054.53
R6349 vss.n6753 vss.n6752 1054.53
R6350 vss.n6774 vss.n6749 1054.53
R6351 vss.n6774 vss.n6754 1054.53
R6352 vss.n6838 vss.n6834 1054.53
R6353 vss.n6839 vss.n6838 1054.53
R6354 vss.n6854 vss.n6844 1054.53
R6355 vss.n6844 vss.n6842 1054.53
R6356 vss.n6860 vss.n6835 1054.53
R6357 vss.n6860 vss.n6840 1054.53
R6358 vss.n3157 vss.n3153 1054.53
R6359 vss.n3158 vss.n3157 1054.53
R6360 vss.n6815 vss.n6814 1054.53
R6361 vss.n6814 vss.n6812 1054.53
R6362 vss.n3146 vss.n3145 1054.53
R6363 vss.n3146 vss.n3142 1054.53
R6364 vss.n3141 vss.n3136 1054.53
R6365 vss.n7214 vss.n3141 1054.53
R6366 vss.n6882 vss.n6828 1054.53
R6367 vss.n6883 vss.n6882 1054.53
R6368 vss.n6888 vss.n6880 1054.53
R6369 vss.n6888 vss.n6884 1054.53
R6370 vss.n6904 vss.n6894 1054.53
R6371 vss.n6904 vss.n6891 1054.53
R6372 vss.n7085 vss.n7080 1054.53
R6373 vss.n7086 vss.n7085 1054.53
R6374 vss.n7091 vss.n7083 1054.53
R6375 vss.n7091 vss.n7087 1054.53
R6376 vss.n7108 vss.n7097 1054.53
R6377 vss.n7108 vss.n7094 1054.53
R6378 vss.n7972 vss.n2466 1054.53
R6379 vss.n7961 vss.n2466 1054.53
R6380 vss.n7975 vss.n7974 1054.53
R6381 vss.n7975 vss.n2464 1054.53
R6382 vss.n2461 vss.n2457 1054.53
R6383 vss.n2462 vss.n2461 1054.53
R6384 vss.n3000 vss.n2989 1054.53
R6385 vss.n2989 vss.n2987 1054.53
R6386 vss.n2983 vss.n2979 1054.53
R6387 vss.n2984 vss.n2983 1054.53
R6388 vss.n3006 vss.n2980 1054.53
R6389 vss.n3006 vss.n2985 1054.53
R6390 vss.n7694 vss.n7683 1054.53
R6391 vss.n7683 vss.n7681 1054.53
R6392 vss.n7677 vss.n7673 1054.53
R6393 vss.n7678 vss.n7677 1054.53
R6394 vss.n7700 vss.n7674 1054.53
R6395 vss.n7700 vss.n7679 1054.53
R6396 vss.n2911 vss.n2896 1054.53
R6397 vss.n2900 vss.n2896 1054.53
R6398 vss.n2914 vss.n2913 1054.53
R6399 vss.n2914 vss.n2894 1054.53
R6400 vss.n2891 vss.n2888 1054.53
R6401 vss.n2892 vss.n2891 1054.53
R6402 vss.n7743 vss.n7732 1054.53
R6403 vss.n7732 vss.n7730 1054.53
R6404 vss.n7726 vss.n7722 1054.53
R6405 vss.n7727 vss.n7726 1054.53
R6406 vss.n7749 vss.n7723 1054.53
R6407 vss.n7749 vss.n7728 1054.53
R6408 vss.n7889 vss.n7878 1054.53
R6409 vss.n7878 vss.n7876 1054.53
R6410 vss.n7872 vss.n7868 1054.53
R6411 vss.n7873 vss.n7872 1054.53
R6412 vss.n7895 vss.n7869 1054.53
R6413 vss.n7895 vss.n7874 1054.53
R6414 vss.n2653 vss.n2652 1054.53
R6415 vss.n2652 vss.n2649 1054.53
R6416 vss.n7916 vss.n2656 1054.53
R6417 vss.n7916 vss.n2650 1054.53
R6418 vss.n2665 vss.n2662 1054.53
R6419 vss.n2666 vss.n2665 1054.53
R6420 vss.n7939 vss.n7929 1054.53
R6421 vss.n7939 vss.n7938 1054.53
R6422 vss.n1148 vss.n1144 1054.53
R6423 vss.n1149 vss.n1148 1054.53
R6424 vss.n1152 vss.n1145 1054.53
R6425 vss.n1152 vss.n1150 1054.53
R6426 vss.n2629 vss.n2609 1054.53
R6427 vss.n2609 vss.n2604 1054.53
R6428 vss.n2614 vss.n2610 1054.53
R6429 vss.n2614 vss.n2613 1054.53
R6430 vss.n2631 vss.n2630 1054.53
R6431 vss.n2630 vss.n2605 1054.53
R6432 vss.n1911 vss.n1909 1054.53
R6433 vss.n1911 vss.n1904 1054.53
R6434 vss.n1908 vss.n1907 1054.53
R6435 vss.n1907 vss.n1903 1054.53
R6436 vss.n1917 vss.n1914 1054.53
R6437 vss.n1917 vss.n1916 1054.53
R6438 vss.n2845 vss.n2841 1054.53
R6439 vss.n2846 vss.n2845 1054.53
R6440 vss.n2861 vss.n2851 1054.53
R6441 vss.n2851 vss.n2849 1054.53
R6442 vss.n2867 vss.n2842 1054.53
R6443 vss.n2867 vss.n2847 1054.53
R6444 vss.n3022 vss.n3021 1054.53
R6445 vss.n3022 vss.n3018 1054.53
R6446 vss.n3028 vss.n3025 1054.53
R6447 vss.n3028 vss.n3027 1054.53
R6448 vss.n3049 vss.n3048 1054.53
R6449 vss.n3049 vss.n3019 1054.53
R6450 vss.n7629 vss.n7625 1054.53
R6451 vss.n7630 vss.n7629 1054.53
R6452 vss.n7645 vss.n7635 1054.53
R6453 vss.n7635 vss.n7633 1054.53
R6454 vss.n7651 vss.n7626 1054.53
R6455 vss.n7651 vss.n7631 1054.53
R6456 vss.n2731 vss.n2727 1054.53
R6457 vss.n2732 vss.n2731 1054.53
R6458 vss.n2815 vss.n2737 1054.53
R6459 vss.n2737 vss.n2735 1054.53
R6460 vss.n2821 vss.n2728 1054.53
R6461 vss.n2821 vss.n2733 1054.53
R6462 vss.n2937 vss.n2933 1054.53
R6463 vss.n2938 vss.n2937 1054.53
R6464 vss.n2953 vss.n2943 1054.53
R6465 vss.n2943 vss.n2941 1054.53
R6466 vss.n2959 vss.n2934 1054.53
R6467 vss.n2959 vss.n2939 1054.53
R6468 vss.n7067 vss.n7045 1054.53
R6469 vss.n7067 vss.n7039 1054.53
R6470 vss.n7042 vss.n7041 1054.53
R6471 vss.n7041 vss.n7038 1054.53
R6472 vss.n7062 vss.n7061 1054.53
R6473 vss.n7061 vss.n7050 1054.53
R6474 vss.n7018 vss.n6998 1054.53
R6475 vss.n6998 vss.n6993 1054.53
R6476 vss.n7003 vss.n6999 1054.53
R6477 vss.n7003 vss.n7002 1054.53
R6478 vss.n7020 vss.n7019 1054.53
R6479 vss.n7019 vss.n6994 1054.53
R6480 vss.n7137 vss.n7134 1054.53
R6481 vss.n7137 vss.n7130 1054.53
R6482 vss.n7143 vss.n7140 1054.53
R6483 vss.n7143 vss.n7142 1054.53
R6484 vss.n7136 vss.n7135 1054.53
R6485 vss.n7135 vss.n7131 1054.53
R6486 vss.n6933 vss.n6930 1054.53
R6487 vss.n6933 vss.n6926 1054.53
R6488 vss.n6939 vss.n6936 1054.53
R6489 vss.n6939 vss.n6938 1054.53
R6490 vss.n6932 vss.n6931 1054.53
R6491 vss.n6931 vss.n6927 1054.53
R6492 vss.n7513 vss.n7509 1054.53
R6493 vss.n7514 vss.n7513 1054.53
R6494 vss.n7597 vss.n7519 1054.53
R6495 vss.n7519 vss.n7517 1054.53
R6496 vss.n7603 vss.n7510 1054.53
R6497 vss.n7603 vss.n7515 1054.53
R6498 vss.n7776 vss.n7772 1054.53
R6499 vss.n7777 vss.n7776 1054.53
R6500 vss.n7792 vss.n7782 1054.53
R6501 vss.n7782 vss.n7780 1054.53
R6502 vss.n7798 vss.n7773 1054.53
R6503 vss.n7798 vss.n7778 1054.53
R6504 vss.n7824 vss.n7820 1054.53
R6505 vss.n7825 vss.n7824 1054.53
R6506 vss.n7840 vss.n7830 1054.53
R6507 vss.n7830 vss.n7828 1054.53
R6508 vss.n7846 vss.n7821 1054.53
R6509 vss.n7846 vss.n7826 1054.53
R6510 vss.n2686 vss.n2682 1054.53
R6511 vss.n2687 vss.n2686 1054.53
R6512 vss.n2702 vss.n2692 1054.53
R6513 vss.n2692 vss.n2690 1054.53
R6514 vss.n2708 vss.n2683 1054.53
R6515 vss.n2708 vss.n2688 1054.53
R6516 vss.n2496 vss.n2493 1054.53
R6517 vss.n2496 vss.n2489 1054.53
R6518 vss.n2502 vss.n2499 1054.53
R6519 vss.n2502 vss.n2501 1054.53
R6520 vss.n2495 vss.n2494 1054.53
R6521 vss.n2494 vss.n2490 1054.53
R6522 vss.n7184 vss.n3163 1054.53
R6523 vss.n3163 vss.n3161 1054.53
R6524 vss.n7190 vss.n3154 1054.53
R6525 vss.n7190 vss.n3159 1054.53
R6526 vss.n3182 vss.n3179 1054.53
R6527 vss.n3182 vss.n3175 1054.53
R6528 vss.n3200 vss.n3199 1054.53
R6529 vss.n3199 vss.n3197 1054.53
R6530 vss.n3181 vss.n3180 1054.53
R6531 vss.n3180 vss.n3176 1054.53
R6532 vss.n14303 vss.n14301 1054.53
R6533 vss.n14303 vss.n14287 1054.53
R6534 vss.n14298 vss.n14297 1054.53
R6535 vss.n14297 vss.n14286 1054.53
R6536 vss.n14315 vss.n14314 1054.53
R6537 vss.n14315 vss.n14292 1054.53
R6538 vss.n14813 vss.n14812 1054.53
R6539 vss.n14812 vss.n14808 1054.53
R6540 vss.n14814 vss.n14811 1054.53
R6541 vss.n14814 vss.n14807 1054.53
R6542 vss.n14820 vss.n14817 1054.53
R6543 vss.n14820 vss.n14819 1054.53
R6544 vss.n1179 vss.n1177 1054.53
R6545 vss.n1179 vss.n1172 1054.53
R6546 vss.n1176 vss.n1175 1054.53
R6547 vss.n1175 vss.n1171 1054.53
R6548 vss.n14168 vss.n14161 1054.53
R6549 vss.n14168 vss.n14162 1054.53
R6550 vss.n14249 vss.n14245 1054.53
R6551 vss.n14277 vss.n14245 1054.53
R6552 vss.n14254 vss.n14253 1054.53
R6553 vss.n14253 vss.n14244 1054.53
R6554 vss.n14259 vss.n14258 1054.53
R6555 vss.n14261 vss.n14259 1054.53
R6556 vss.n1849 vss.n1829 1054.53
R6557 vss.n1849 vss.n1824 1054.53
R6558 vss.n1828 vss.n1827 1054.53
R6559 vss.n1827 vss.n1823 1054.53
R6560 vss.n1833 vss.n1831 1054.53
R6561 vss.n1843 vss.n1833 1054.53
R6562 vss.n14371 vss.n14368 1054.53
R6563 vss.n14371 vss.n14370 1054.53
R6564 vss.n14365 vss.n14362 1054.53
R6565 vss.n14365 vss.n14358 1054.53
R6566 vss.n1789 vss.n1786 1054.53
R6567 vss.n1789 vss.n1788 1054.53
R6568 vss.n14460 vss.n1754 1054.53
R6569 vss.n14460 vss.n1749 1054.53
R6570 vss.n1753 vss.n1752 1054.53
R6571 vss.n1752 vss.n1748 1054.53
R6572 vss.n1758 vss.n1756 1054.53
R6573 vss.n14454 vss.n1758 1054.53
R6574 vss.n14224 vss.n14202 1054.53
R6575 vss.n14224 vss.n14197 1054.53
R6576 vss.n14201 vss.n14200 1054.53
R6577 vss.n14200 vss.n14196 1054.53
R6578 vss.n14206 vss.n14204 1054.53
R6579 vss.n14218 vss.n14206 1054.53
R6580 vss.n2307 vss.n2286 1054.53
R6581 vss.n2307 vss.n2281 1054.53
R6582 vss.n2285 vss.n2284 1054.53
R6583 vss.n2284 vss.n2280 1054.53
R6584 vss.n2290 vss.n2288 1054.53
R6585 vss.n2301 vss.n2290 1054.53
R6586 vss.n2261 vss.n2240 1054.53
R6587 vss.n2261 vss.n2235 1054.53
R6588 vss.n2239 vss.n2238 1054.53
R6589 vss.n2238 vss.n2234 1054.53
R6590 vss.n2244 vss.n2242 1054.53
R6591 vss.n2255 vss.n2244 1054.53
R6592 vss.n8067 vss.n8064 1054.53
R6593 vss.n8067 vss.n8066 1054.53
R6594 vss.n8061 vss.n8059 1054.53
R6595 vss.n8061 vss.n8054 1054.53
R6596 vss.n8058 vss.n8057 1054.53
R6597 vss.n8057 vss.n8053 1054.53
R6598 vss.n8119 vss.n8116 1054.53
R6599 vss.n8119 vss.n8118 1054.53
R6600 vss.n8113 vss.n8109 1054.53
R6601 vss.n8113 vss.n8104 1054.53
R6602 vss.n8108 vss.n8107 1054.53
R6603 vss.n8107 vss.n8100 1054.53
R6604 vss.n1311 vss.n1291 1054.53
R6605 vss.n1311 vss.n1286 1054.53
R6606 vss.n1290 vss.n1289 1054.53
R6607 vss.n1289 vss.n1285 1054.53
R6608 vss.n1295 vss.n1293 1054.53
R6609 vss.n1305 vss.n1295 1054.53
R6610 vss.n14010 vss.n13990 1054.53
R6611 vss.n14010 vss.n13985 1054.53
R6612 vss.n13989 vss.n13988 1054.53
R6613 vss.n13988 vss.n13984 1054.53
R6614 vss.n13994 vss.n13992 1054.53
R6615 vss.n14004 vss.n13994 1054.53
R6616 vss.n14043 vss.n14040 1054.53
R6617 vss.n14043 vss.n14042 1054.53
R6618 vss.n14037 vss.n14034 1054.53
R6619 vss.n14037 vss.n14030 1054.53
R6620 vss.n13964 vss.n8161 1054.53
R6621 vss.n13964 vss.n8156 1054.53
R6622 vss.n8160 vss.n8159 1054.53
R6623 vss.n8159 vss.n8155 1054.53
R6624 vss.n8165 vss.n8163 1054.53
R6625 vss.n13958 vss.n8165 1054.53
R6626 vss.n8195 vss.n8192 1054.53
R6627 vss.n8195 vss.n8194 1054.53
R6628 vss.n8189 vss.n8187 1054.53
R6629 vss.n8189 vss.n8182 1054.53
R6630 vss.n8186 vss.n8185 1054.53
R6631 vss.n8185 vss.n8181 1054.53
R6632 vss.n13880 vss.n13877 1054.53
R6633 vss.n13880 vss.n13879 1054.53
R6634 vss.n13874 vss.n13870 1054.53
R6635 vss.n13874 vss.n13865 1054.53
R6636 vss.n13869 vss.n13868 1054.53
R6637 vss.n13868 vss.n13861 1054.53
R6638 vss.n1516 vss.n1496 1054.53
R6639 vss.n1516 vss.n1491 1054.53
R6640 vss.n1495 vss.n1494 1054.53
R6641 vss.n1494 vss.n1490 1054.53
R6642 vss.n1500 vss.n1498 1054.53
R6643 vss.n1510 vss.n1500 1054.53
R6644 vss.n1569 vss.n1549 1054.53
R6645 vss.n1569 vss.n1544 1054.53
R6646 vss.n1548 vss.n1547 1054.53
R6647 vss.n1547 vss.n1543 1054.53
R6648 vss.n1553 vss.n1551 1054.53
R6649 vss.n1563 vss.n1553 1054.53
R6650 vss.n13926 vss.n13923 1054.53
R6651 vss.n13926 vss.n13925 1054.53
R6652 vss.n13920 vss.n13917 1054.53
R6653 vss.n13920 vss.n13913 1054.53
R6654 vss.n14422 vss.n14419 1054.53
R6655 vss.n14422 vss.n14421 1054.53
R6656 vss.n14416 vss.n14411 1054.53
R6657 vss.n14416 vss.n14406 1054.53
R6658 vss.n14410 vss.n14409 1054.53
R6659 vss.n14409 vss.n14402 1054.53
R6660 vss.n14509 vss.n14489 1054.53
R6661 vss.n14509 vss.n14484 1054.53
R6662 vss.n14488 vss.n14487 1054.53
R6663 vss.n14487 vss.n14483 1054.53
R6664 vss.n14493 vss.n14491 1054.53
R6665 vss.n14503 vss.n14493 1054.53
R6666 vss.n1726 vss.n1706 1054.53
R6667 vss.n1726 vss.n1701 1054.53
R6668 vss.n1705 vss.n1704 1054.53
R6669 vss.n1704 vss.n1700 1054.53
R6670 vss.n1710 vss.n1708 1054.53
R6671 vss.n1720 vss.n1710 1054.53
R6672 vss.n1596 vss.n1595 1054.53
R6673 vss.n1595 vss.n1591 1054.53
R6674 vss.n1597 vss.n1594 1054.53
R6675 vss.n1597 vss.n1590 1054.53
R6676 vss.n1603 vss.n1600 1054.53
R6677 vss.n1603 vss.n1602 1054.53
R6678 vss.n13916 vss.n13915 1054.53
R6679 vss.n13915 vss.n13908 1054.53
R6680 vss.n14629 vss.n14609 1054.53
R6681 vss.n14629 vss.n14604 1054.53
R6682 vss.n14608 vss.n14607 1054.53
R6683 vss.n14607 vss.n14603 1054.53
R6684 vss.n14613 vss.n14611 1054.53
R6685 vss.n14623 vss.n14613 1054.53
R6686 vss.n1469 vss.n1449 1054.53
R6687 vss.n1469 vss.n1444 1054.53
R6688 vss.n1448 vss.n1447 1054.53
R6689 vss.n1447 vss.n1443 1054.53
R6690 vss.n1453 vss.n1451 1054.53
R6691 vss.n1463 vss.n1453 1054.53
R6692 vss.n14033 vss.n14032 1054.53
R6693 vss.n14032 vss.n8147 1054.53
R6694 vss.n1339 vss.n1338 1054.53
R6695 vss.n1338 vss.n1334 1054.53
R6696 vss.n1340 vss.n1337 1054.53
R6697 vss.n1340 vss.n1333 1054.53
R6698 vss.n1346 vss.n1343 1054.53
R6699 vss.n1346 vss.n1345 1054.53
R6700 vss.n1261 vss.n1241 1054.53
R6701 vss.n1261 vss.n1236 1054.53
R6702 vss.n1240 vss.n1239 1054.53
R6703 vss.n1239 vss.n1235 1054.53
R6704 vss.n1245 vss.n1243 1054.53
R6705 vss.n1255 vss.n1245 1054.53
R6706 vss.n2354 vss.n2334 1054.53
R6707 vss.n2354 vss.n2329 1054.53
R6708 vss.n2333 vss.n2332 1054.53
R6709 vss.n2332 vss.n2328 1054.53
R6710 vss.n2338 vss.n2336 1054.53
R6711 vss.n2348 vss.n2338 1054.53
R6712 vss.n2381 vss.n2380 1054.53
R6713 vss.n2380 vss.n2376 1054.53
R6714 vss.n2382 vss.n2379 1054.53
R6715 vss.n2382 vss.n2375 1054.53
R6716 vss.n2388 vss.n2385 1054.53
R6717 vss.n2388 vss.n2387 1054.53
R6718 vss.n11856 vss.n11855 1054.53
R6719 vss.n11855 vss.n11853 1054.53
R6720 vss.n2042 vss.n2038 1054.53
R6721 vss.n2043 vss.n2042 1054.53
R6722 vss.n2046 vss.n2039 1054.53
R6723 vss.n2046 vss.n2044 1054.53
R6724 vss.n2094 vss.n2090 1054.53
R6725 vss.n2095 vss.n2094 1054.53
R6726 vss.n11953 vss.n11952 1054.53
R6727 vss.n11952 vss.n11950 1054.53
R6728 vss.n2098 vss.n2091 1054.53
R6729 vss.n2098 vss.n2096 1054.53
R6730 vss.n13474 vss.n13470 1054.53
R6731 vss.n13475 vss.n13474 1054.53
R6732 vss.n13490 vss.n13480 1054.53
R6733 vss.n13480 vss.n13478 1054.53
R6734 vss.n13496 vss.n13471 1054.53
R6735 vss.n13496 vss.n13476 1054.53
R6736 vss.n12029 vss.n12027 1054.53
R6737 vss.n12029 vss.n12022 1054.53
R6738 vss.n12026 vss.n12025 1054.53
R6739 vss.n12025 vss.n12021 1054.53
R6740 vss.n12035 vss.n12032 1054.53
R6741 vss.n12035 vss.n12034 1054.53
R6742 vss.n8309 vss.n8305 1054.53
R6743 vss.n8310 vss.n8309 1054.53
R6744 vss.n13722 vss.n8315 1054.53
R6745 vss.n8315 vss.n8313 1054.53
R6746 vss.n13728 vss.n8306 1054.53
R6747 vss.n13728 vss.n8311 1054.53
R6748 vss.n8455 vss.n8453 1054.53
R6749 vss.n8455 vss.n8448 1054.53
R6750 vss.n8452 vss.n8451 1054.53
R6751 vss.n8451 vss.n8447 1054.53
R6752 vss.n8461 vss.n8458 1054.53
R6753 vss.n8461 vss.n8460 1054.53
R6754 vss.n8532 vss.n8530 1054.53
R6755 vss.n8532 vss.n8525 1054.53
R6756 vss.n8529 vss.n8528 1054.53
R6757 vss.n8528 vss.n8524 1054.53
R6758 vss.n8538 vss.n8535 1054.53
R6759 vss.n8538 vss.n8537 1054.53
R6760 vss.n9095 vss.n9091 1054.53
R6761 vss.n9096 vss.n9095 1054.53
R6762 vss.n13010 vss.n9101 1054.53
R6763 vss.n9101 vss.n9099 1054.53
R6764 vss.n13016 vss.n9092 1054.53
R6765 vss.n13016 vss.n9097 1054.53
R6766 vss.n8959 vss.n8955 1054.53
R6767 vss.n8960 vss.n8959 1054.53
R6768 vss.n8975 vss.n8965 1054.53
R6769 vss.n8965 vss.n8963 1054.53
R6770 vss.n8981 vss.n8956 1054.53
R6771 vss.n8981 vss.n8961 1054.53
R6772 vss.n9127 vss.n9125 1054.53
R6773 vss.n9127 vss.n9120 1054.53
R6774 vss.n9124 vss.n9123 1054.53
R6775 vss.n9123 vss.n9119 1054.53
R6776 vss.n9133 vss.n9130 1054.53
R6777 vss.n9133 vss.n9132 1054.53
R6778 vss.n12558 vss.n12556 1054.53
R6779 vss.n12558 vss.n12551 1054.53
R6780 vss.n12555 vss.n12554 1054.53
R6781 vss.n12554 vss.n12550 1054.53
R6782 vss.n12564 vss.n12561 1054.53
R6783 vss.n12564 vss.n12563 1054.53
R6784 vss.n2211 vss.n2191 1054.53
R6785 vss.n2191 vss.n2186 1054.53
R6786 vss.n2169 vss.n2159 1054.53
R6787 vss.n2159 vss.n2157 1054.53
R6788 vss.n2153 vss.n2149 1054.53
R6789 vss.n2154 vss.n2153 1054.53
R6790 vss.n2175 vss.n2150 1054.53
R6791 vss.n2175 vss.n2155 1054.53
R6792 vss.n12603 vss.n12592 1054.53
R6793 vss.n12592 vss.n12590 1054.53
R6794 vss.n12586 vss.n12582 1054.53
R6795 vss.n12587 vss.n12586 1054.53
R6796 vss.n12609 vss.n12583 1054.53
R6797 vss.n12609 vss.n12588 1054.53
R6798 vss.n9004 vss.n9000 1054.53
R6799 vss.n9005 vss.n9004 1054.53
R6800 vss.n9020 vss.n9010 1054.53
R6801 vss.n9010 vss.n9008 1054.53
R6802 vss.n9026 vss.n9001 1054.53
R6803 vss.n9026 vss.n9006 1054.53
R6804 vss.n13106 vss.n13095 1054.53
R6805 vss.n13095 vss.n13093 1054.53
R6806 vss.n13089 vss.n13085 1054.53
R6807 vss.n13090 vss.n13089 1054.53
R6808 vss.n13112 vss.n13086 1054.53
R6809 vss.n13112 vss.n13091 1054.53
R6810 vss.n13057 vss.n13047 1054.53
R6811 vss.n13047 vss.n13045 1054.53
R6812 vss.n13041 vss.n13037 1054.53
R6813 vss.n13042 vss.n13041 1054.53
R6814 vss.n13063 vss.n13038 1054.53
R6815 vss.n13063 vss.n13043 1054.53
R6816 vss.n9065 vss.n9054 1054.53
R6817 vss.n9054 vss.n9052 1054.53
R6818 vss.n9048 vss.n9044 1054.53
R6819 vss.n9049 vss.n9048 1054.53
R6820 vss.n9071 vss.n9045 1054.53
R6821 vss.n9071 vss.n9050 1054.53
R6822 vss.n8233 vss.n8232 1054.53
R6823 vss.n8233 vss.n8229 1054.53
R6824 vss.n8239 vss.n8236 1054.53
R6825 vss.n8239 vss.n8238 1054.53
R6826 vss.n13850 vss.n13849 1054.53
R6827 vss.n13850 vss.n8230 1054.53
R6828 vss.n13818 vss.n13807 1054.53
R6829 vss.n13807 vss.n13805 1054.53
R6830 vss.n13801 vss.n13797 1054.53
R6831 vss.n13802 vss.n13801 1054.53
R6832 vss.n13824 vss.n13798 1054.53
R6833 vss.n13824 vss.n13803 1054.53
R6834 vss.n13769 vss.n13759 1054.53
R6835 vss.n13759 vss.n13757 1054.53
R6836 vss.n13753 vss.n13749 1054.53
R6837 vss.n13754 vss.n13753 1054.53
R6838 vss.n13775 vss.n13750 1054.53
R6839 vss.n13775 vss.n13755 1054.53
R6840 vss.n8279 vss.n8268 1054.53
R6841 vss.n8268 vss.n8266 1054.53
R6842 vss.n8262 vss.n8258 1054.53
R6843 vss.n8263 vss.n8262 1054.53
R6844 vss.n8285 vss.n8259 1054.53
R6845 vss.n8285 vss.n8264 1054.53
R6846 vss.n13519 vss.n13515 1054.53
R6847 vss.n13520 vss.n13519 1054.53
R6848 vss.n13535 vss.n13525 1054.53
R6849 vss.n13525 vss.n13523 1054.53
R6850 vss.n13541 vss.n13516 1054.53
R6851 vss.n13541 vss.n13521 1054.53
R6852 vss.n13629 vss.n13618 1054.53
R6853 vss.n13618 vss.n13616 1054.53
R6854 vss.n13612 vss.n13608 1054.53
R6855 vss.n13613 vss.n13612 1054.53
R6856 vss.n13635 vss.n13609 1054.53
R6857 vss.n13635 vss.n13614 1054.53
R6858 vss.n13580 vss.n13569 1054.53
R6859 vss.n13569 vss.n13567 1054.53
R6860 vss.n13563 vss.n13559 1054.53
R6861 vss.n13564 vss.n13563 1054.53
R6862 vss.n13586 vss.n13560 1054.53
R6863 vss.n13586 vss.n13565 1054.53
R6864 vss.n2070 vss.n2067 1054.53
R6865 vss.n2070 vss.n2069 1054.53
R6866 vss.n2064 vss.n2063 1054.53
R6867 vss.n2064 vss.n2060 1054.53
R6868 vss.n14146 vss.n14145 1054.53
R6869 vss.n14146 vss.n2061 1054.53
R6870 vss.n2196 vss.n2192 1054.53
R6871 vss.n2196 vss.n2195 1054.53
R6872 vss.n2213 vss.n2212 1054.53
R6873 vss.n2212 vss.n2187 1054.53
R6874 vss.n2141 vss.n2138 1054.53
R6875 vss.n2141 vss.n2134 1054.53
R6876 vss.n9292 vss.n9291 1054.53
R6877 vss.n9291 vss.n9289 1054.53
R6878 vss.n2140 vss.n2139 1054.53
R6879 vss.n2139 vss.n2135 1054.53
R6880 vss.n9399 vss.n9395 1054.53
R6881 vss.n9400 vss.n9399 1054.53
R6882 vss.n12847 vss.n9405 1054.53
R6883 vss.n9405 vss.n9403 1054.53
R6884 vss.n12853 vss.n9396 1054.53
R6885 vss.n12853 vss.n9401 1054.53
R6886 vss.n12742 vss.n12740 1054.53
R6887 vss.n12742 vss.n12735 1054.53
R6888 vss.n12739 vss.n12738 1054.53
R6889 vss.n12738 vss.n12734 1054.53
R6890 vss.n12748 vss.n12745 1054.53
R6891 vss.n12748 vss.n12747 1054.53
R6892 vss.n8417 vss.n8413 1054.53
R6893 vss.n8418 vss.n8417 1054.53
R6894 vss.n13324 vss.n8423 1054.53
R6895 vss.n8423 vss.n8421 1054.53
R6896 vss.n13330 vss.n8414 1054.53
R6897 vss.n13330 vss.n8419 1054.53
R6898 vss.n13359 vss.n13355 1054.53
R6899 vss.n13360 vss.n13359 1054.53
R6900 vss.n13443 vss.n13365 1054.53
R6901 vss.n13365 vss.n13363 1054.53
R6902 vss.n13449 vss.n13356 1054.53
R6903 vss.n13449 vss.n13361 1054.53
R6904 vss.n1783 vss.n1779 1054.53
R6905 vss.n1783 vss.n1774 1054.53
R6906 vss.n1778 vss.n1777 1054.53
R6907 vss.n1777 vss.n1770 1054.53
R6908 vss.n14361 vss.n14360 1054.53
R6909 vss.n14360 vss.n1817 1054.53
R6910 vss.n2016 vss.n1996 1054.53
R6911 vss.n2016 vss.n1991 1054.53
R6912 vss.n1995 vss.n1994 1054.53
R6913 vss.n1994 vss.n1990 1054.53
R6914 vss.n2000 vss.n1998 1054.53
R6915 vss.n2010 vss.n2000 1054.53
R6916 vss.n1004 vss.n1000 1054.53
R6917 vss.n1004 vss.n995 1054.53
R6918 vss.n999 vss.n998 1054.53
R6919 vss.n998 vss.n991 1054.53
R6920 vss.n15056 vss.n15055 1054.53
R6921 vss.n15055 vss.n1038 1054.53
R6922 vss.n1121 vss.n1101 1054.53
R6923 vss.n1121 vss.n1096 1054.53
R6924 vss.n1100 vss.n1099 1054.53
R6925 vss.n1099 vss.n1095 1054.53
R6926 vss.n1105 vss.n1103 1054.53
R6927 vss.n1115 vss.n1105 1054.53
R6928 vss.n6215 vss.n6214 1054.53
R6929 vss.n6214 vss.n6207 1054.53
R6930 vss.n40 vss.n38 1054.53
R6931 vss.n40 vss.n33 1054.53
R6932 vss.n37 vss.n36 1054.53
R6933 vss.n36 vss.n32 1054.53
R6934 vss.n3960 vss.n3959 1054.53
R6935 vss.n3960 vss.n3951 1054.53
R6936 vss.n3871 vss.n3868 1054.53
R6937 vss.n3871 vss.n3870 1054.53
R6938 vss.n3865 vss.n3862 1054.53
R6939 vss.n3865 vss.n3858 1054.53
R6940 vss.n3861 vss.n3860 1054.53
R6941 vss.n3860 vss.n3853 1054.53
R6942 vss.n3752 vss.n3749 1054.53
R6943 vss.n3752 vss.n3751 1054.53
R6944 vss.n3746 vss.n3743 1054.53
R6945 vss.n3746 vss.n3739 1054.53
R6946 vss.n3742 vss.n3741 1054.53
R6947 vss.n3741 vss.n3734 1054.53
R6948 vss.n3633 vss.n3630 1054.53
R6949 vss.n3633 vss.n3632 1054.53
R6950 vss.n3627 vss.n3624 1054.53
R6951 vss.n3627 vss.n3620 1054.53
R6952 vss.n3623 vss.n3622 1054.53
R6953 vss.n3622 vss.n3615 1054.53
R6954 vss.n15587 vss.n15583 1054.53
R6955 vss.n15615 vss.n15583 1054.53
R6956 vss.n15592 vss.n15591 1054.53
R6957 vss.n15591 vss.n15582 1054.53
R6958 vss.n15597 vss.n15596 1054.53
R6959 vss.n15599 vss.n15597 1054.53
R6960 vss.n314 vss.n313 1054.53
R6961 vss.n313 vss.n307 1054.53
R6962 vss.n373 vss.n371 1054.53
R6963 vss.n15553 vss.n373 1054.53
R6964 vss.n10447 vss.n10437 1054.53
R6965 vss.n10437 vss.n10435 1054.53
R6966 vss.n10453 vss.n10428 1054.53
R6967 vss.n10453 vss.n10433 1054.53
R6968 vss.n10576 vss.n10572 1054.53
R6969 vss.n10577 vss.n10576 1054.53
R6970 vss.n10593 vss.n10582 1054.53
R6971 vss.n10582 vss.n10580 1054.53
R6972 vss.n10599 vss.n10573 1054.53
R6973 vss.n10599 vss.n10578 1054.53
R6974 vss.n10970 vss.n10966 1054.53
R6975 vss.n10971 vss.n10970 1054.53
R6976 vss.n10987 vss.n10976 1054.53
R6977 vss.n10976 vss.n10974 1054.53
R6978 vss.n10993 vss.n10967 1054.53
R6979 vss.n10993 vss.n10972 1054.53
R6980 vss.n10006 vss.n10004 1054.53
R6981 vss.n10006 vss.n9999 1054.53
R6982 vss.n10003 vss.n10002 1054.53
R6983 vss.n10002 vss.n9998 1054.53
R6984 vss.n10012 vss.n10009 1054.53
R6985 vss.n10012 vss.n10011 1054.53
R6986 vss.n14765 vss.n14764 922
R6987 vss.n15460 vss.n15459 922
R6988 vss.n12904 vss.n12903 922
R6989 vss.n15542 vss.n15541 866.162
R6990 vss.n12181 vss.n12132 866.162
R6991 vss.n13224 vss.n13223 854.47
R6992 vss.n14176 vss.n1183 814.227
R6993 vss.n9936 vss.n9932 759.029
R6994 vss.n9941 vss.n9931 759.029
R6995 vss.n11670 vss.n9941 759.029
R6996 vss.n11670 vss.n9942 759.029
R6997 vss.n11672 vss.n9936 759.029
R6998 vss.n11672 vss.n9937 759.029
R6999 vss.n11664 vss.n9937 759.029
R7000 vss.n11664 vss.n11651 759.029
R7001 vss.n11666 vss.n9942 759.029
R7002 vss.n11666 vss.n9947 759.029
R7003 vss.n11658 vss.n9947 759.029
R7004 vss.n11655 vss.n11651 759.029
R7005 vss.n11354 vss.n11351 759.029
R7006 vss.n11359 vss.n11350 759.029
R7007 vss.n11433 vss.n11359 759.029
R7008 vss.n11433 vss.n11360 759.029
R7009 vss.n11435 vss.n11354 759.029
R7010 vss.n11435 vss.n11355 759.029
R7011 vss.n11427 vss.n11355 759.029
R7012 vss.n11427 vss.n11414 759.029
R7013 vss.n11429 vss.n11360 759.029
R7014 vss.n11429 vss.n11365 759.029
R7015 vss.n11421 vss.n11365 759.029
R7016 vss.n11418 vss.n11414 759.029
R7017 vss.n11328 vss.n10050 759.029
R7018 vss.n11326 vss.n10046 759.029
R7019 vss.n11335 vss.n10046 759.029
R7020 vss.n11335 vss.n10041 759.029
R7021 vss.n11333 vss.n10050 759.029
R7022 vss.n11333 vss.n9990 759.029
R7023 vss.n11342 vss.n9990 759.029
R7024 vss.n11342 vss.n9991 759.029
R7025 vss.n11340 vss.n10041 759.029
R7026 vss.n11340 vss.n10043 759.029
R7027 vss.n10043 vss.n9985 759.029
R7028 vss.n9991 vss.n9986 759.029
R7029 vss.n11031 vss.n10075 759.029
R7030 vss.n11030 vss.n10071 759.029
R7031 vss.n11309 vss.n10071 759.029
R7032 vss.n11309 vss.n10066 759.029
R7033 vss.n11307 vss.n10075 759.029
R7034 vss.n11307 vss.n10062 759.029
R7035 vss.n11316 vss.n10062 759.029
R7036 vss.n11316 vss.n10063 759.029
R7037 vss.n11314 vss.n10066 759.029
R7038 vss.n11314 vss.n10068 759.029
R7039 vss.n10068 vss.n10057 759.029
R7040 vss.n10063 vss.n10058 759.029
R7041 vss.n10757 vss.n10163 759.029
R7042 vss.n10756 vss.n10159 759.029
R7043 vss.n11015 vss.n10159 759.029
R7044 vss.n11015 vss.n10154 759.029
R7045 vss.n11013 vss.n10163 759.029
R7046 vss.n11013 vss.n10150 759.029
R7047 vss.n11022 vss.n10150 759.029
R7048 vss.n11022 vss.n10151 759.029
R7049 vss.n11020 vss.n10154 759.029
R7050 vss.n11020 vss.n10156 759.029
R7051 vss.n10156 vss.n10145 759.029
R7052 vss.n10151 vss.n10146 759.029
R7053 vss.n10642 vss.n10638 759.029
R7054 vss.n10647 vss.n10637 759.029
R7055 vss.n10776 vss.n10647 759.029
R7056 vss.n10776 vss.n10648 759.029
R7057 vss.n10778 vss.n10642 759.029
R7058 vss.n10778 vss.n10643 759.029
R7059 vss.n10770 vss.n10643 759.029
R7060 vss.n10770 vss.n10702 759.029
R7061 vss.n10772 vss.n10648 759.029
R7062 vss.n10772 vss.n10653 759.029
R7063 vss.n10708 vss.n10653 759.029
R7064 vss.n10706 vss.n10702 759.029
R7065 vss.n10389 vss.n10250 759.029
R7066 vss.n10388 vss.n10246 759.029
R7067 vss.n10622 vss.n10246 759.029
R7068 vss.n10622 vss.n10241 759.029
R7069 vss.n10620 vss.n10250 759.029
R7070 vss.n10620 vss.n10237 759.029
R7071 vss.n10629 vss.n10237 759.029
R7072 vss.n10629 vss.n10238 759.029
R7073 vss.n10627 vss.n10241 759.029
R7074 vss.n10627 vss.n10243 759.029
R7075 vss.n10243 vss.n10232 759.029
R7076 vss.n10238 vss.n10233 759.029
R7077 vss.n12094 vss.n11885 759.029
R7078 vss.n12100 vss.n11884 759.029
R7079 vss.n12101 vss.n12100 759.029
R7080 vss.n12101 vss.n11868 759.029
R7081 vss.n11885 vss.n11883 759.029
R7082 vss.n11883 vss.n11845 759.029
R7083 vss.n12125 vss.n11845 759.029
R7084 vss.n12125 vss.n11846 759.029
R7085 vss.n12123 vss.n11868 759.029
R7086 vss.n12123 vss.n11870 759.029
R7087 vss.n11870 vss.n11841 759.029
R7088 vss.n11846 vss.n11842 759.029
R7089 vss.n8403 vss.n8388 759.029
R7090 vss.n8396 vss.n8389 759.029
R7091 vss.n8398 vss.n8389 759.029
R7092 vss.n8398 vss.n8384 759.029
R7093 vss.n8404 vss.n8403 759.029
R7094 vss.n8404 vss.n8385 759.029
R7095 vss.n12062 vss.n8385 759.029
R7096 vss.n12062 vss.n12014 759.029
R7097 vss.n12064 vss.n8384 759.029
R7098 vss.n12064 vss.n12013 759.029
R7099 vss.n12013 vss.n12009 759.029
R7100 vss.n12014 vss.n12010 759.029
R7101 vss.n13398 vss.n13389 759.029
R7102 vss.n13393 vss.n13388 759.029
R7103 vss.n13388 vss.n13387 759.029
R7104 vss.n13387 vss.n13373 759.029
R7105 vss.n13400 vss.n13389 759.029
R7106 vss.n13400 vss.n13376 759.029
R7107 vss.n13376 vss.n13372 759.029
R7108 vss.n13429 vss.n13372 759.029
R7109 vss.n13434 vss.n13373 759.029
R7110 vss.n13434 vss.n13374 759.029
R7111 vss.n13426 vss.n13374 759.029
R7112 vss.n13429 vss.n13428 759.029
R7113 vss.n8592 vss.n8585 759.029
R7114 vss.n8599 vss.n8584 759.029
R7115 vss.n8600 vss.n8599 759.029
R7116 vss.n8600 vss.n8514 759.029
R7117 vss.n8594 vss.n8585 759.029
R7118 vss.n8594 vss.n8515 759.029
R7119 vss.n8579 vss.n8515 759.029
R7120 vss.n8579 vss.n8566 759.029
R7121 vss.n8581 vss.n8514 759.029
R7122 vss.n8581 vss.n8517 759.029
R7123 vss.n8569 vss.n8517 759.029
R7124 vss.n8567 vss.n8566 759.029
R7125 vss.n12960 vss.n12957 759.029
R7126 vss.n12970 vss.n12967 759.029
R7127 vss.n12970 vss.n12969 759.029
R7128 vss.n12969 vss.n8431 759.029
R7129 vss.n12975 vss.n12957 759.029
R7130 vss.n12976 vss.n12975 759.029
R7131 vss.n12976 vss.n8430 759.029
R7132 vss.n13310 vss.n8430 759.029
R7133 vss.n13315 vss.n8431 759.029
R7134 vss.n13315 vss.n8432 759.029
R7135 vss.n13307 vss.n8432 759.029
R7136 vss.n13310 vss.n13309 759.029
R7137 vss.n8947 vss.n8932 759.029
R7138 vss.n8940 vss.n8933 759.029
R7139 vss.n8942 vss.n8933 759.029
R7140 vss.n8942 vss.n8928 759.029
R7141 vss.n8948 vss.n8947 759.029
R7142 vss.n8948 vss.n8929 759.029
R7143 vss.n9160 vss.n8929 759.029
R7144 vss.n9160 vss.n9112 759.029
R7145 vss.n9162 vss.n8928 759.029
R7146 vss.n9162 vss.n9111 759.029
R7147 vss.n9111 vss.n9107 759.029
R7148 vss.n9112 vss.n9108 759.029
R7149 vss.n12708 vss.n12701 759.029
R7150 vss.n12811 vss.n12703 759.029
R7151 vss.n12720 vss.n12703 759.029
R7152 vss.n12721 vss.n12720 759.029
R7153 vss.n12724 vss.n12708 759.029
R7154 vss.n12724 vss.n12722 759.029
R7155 vss.n12791 vss.n12722 759.029
R7156 vss.n12791 vss.n12727 759.029
R7157 vss.n12789 vss.n12721 759.029
R7158 vss.n12789 vss.n12777 759.029
R7159 vss.n12783 vss.n12777 759.029
R7160 vss.n12781 vss.n12727 759.029
R7161 vss.n9372 vss.n9365 759.029
R7162 vss.n12888 vss.n9367 759.029
R7163 vss.n9384 vss.n9367 759.029
R7164 vss.n9385 vss.n9384 759.029
R7165 vss.n9388 vss.n9372 759.029
R7166 vss.n9388 vss.n9386 759.029
R7167 vss.n9411 vss.n9386 759.029
R7168 vss.n12833 vss.n9411 759.029
R7169 vss.n12838 vss.n9385 759.029
R7170 vss.n12838 vss.n9412 759.029
R7171 vss.n12830 vss.n9412 759.029
R7172 vss.n12833 vss.n12832 759.029
R7173 vss.n12875 vss.n9374 759.029
R7174 vss.n9379 vss.n9309 759.029
R7175 vss.n9379 vss.n9375 759.029
R7176 vss.n12877 vss.n9375 759.029
R7177 vss.n12895 vss.n9360 759.029
R7178 vss.n12895 vss.n9361 759.029
R7179 vss.n9376 vss.n9361 759.029
R7180 vss.n9376 vss.n9374 759.029
R7181 vss.n9360 vss.n9303 759.029
R7182 vss.n9308 vss.n9304 759.029
R7183 vss.n12897 vss.n9308 759.029
R7184 vss.n12897 vss.n9309 759.029
R7185 vss.n12798 vss.n12710 759.029
R7186 vss.n12715 vss.n12646 759.029
R7187 vss.n12715 vss.n12711 759.029
R7188 vss.n12800 vss.n12711 759.029
R7189 vss.n12818 vss.n12696 759.029
R7190 vss.n12818 vss.n12697 759.029
R7191 vss.n12712 vss.n12697 759.029
R7192 vss.n12712 vss.n12710 759.029
R7193 vss.n12696 vss.n12640 759.029
R7194 vss.n12645 vss.n12641 759.029
R7195 vss.n12820 vss.n12645 759.029
R7196 vss.n12820 vss.n12646 759.029
R7197 vss.n13140 vss.n8917 759.029
R7198 vss.n13146 vss.n8908 759.029
R7199 vss.n13146 vss.n8920 759.029
R7200 vss.n13142 vss.n8920 759.029
R7201 vss.n13153 vss.n8912 759.029
R7202 vss.n13153 vss.n8913 759.029
R7203 vss.n13148 vss.n8913 759.029
R7204 vss.n13148 vss.n8917 759.029
R7205 vss.n8912 vss.n8902 759.029
R7206 vss.n8907 vss.n8903 759.029
R7207 vss.n13155 vss.n8907 759.029
R7208 vss.n13155 vss.n8908 759.029
R7209 vss.n12981 vss.n12947 759.029
R7210 vss.n12987 vss.n9180 759.029
R7211 vss.n12987 vss.n12950 759.029
R7212 vss.n12983 vss.n12950 759.029
R7213 vss.n12994 vss.n12942 759.029
R7214 vss.n12994 vss.n12943 759.029
R7215 vss.n12989 vss.n12943 759.029
R7216 vss.n12989 vss.n12947 759.029
R7217 vss.n12942 vss.n9174 759.029
R7218 vss.n9179 vss.n9175 759.029
R7219 vss.n12996 vss.n9179 759.029
R7220 vss.n12996 vss.n9180 759.029
R7221 vss.n8607 vss.n8503 759.029
R7222 vss.n8613 vss.n8494 759.029
R7223 vss.n8613 vss.n8506 759.029
R7224 vss.n8609 vss.n8506 759.029
R7225 vss.n13295 vss.n8498 759.029
R7226 vss.n13295 vss.n8499 759.029
R7227 vss.n8615 vss.n8499 759.029
R7228 vss.n8615 vss.n8503 759.029
R7229 vss.n8498 vss.n8488 759.029
R7230 vss.n8493 vss.n8489 759.029
R7231 vss.n13297 vss.n8493 759.029
R7232 vss.n13297 vss.n8494 759.029
R7233 vss.n13414 vss.n13379 759.029
R7234 vss.n13408 vss.n8328 759.029
R7235 vss.n13408 vss.n13383 759.029
R7236 vss.n13383 vss.n13378 759.029
R7237 vss.n13706 vss.n8332 759.029
R7238 vss.n13706 vss.n8333 759.029
R7239 vss.n13406 vss.n8333 759.029
R7240 vss.n13406 vss.n13379 759.029
R7241 vss.n8332 vss.n8322 759.029
R7242 vss.n8327 vss.n8323 759.029
R7243 vss.n13708 vss.n8327 759.029
R7244 vss.n13708 vss.n8328 759.029
R7245 vss.n13663 vss.n8373 759.029
R7246 vss.n13669 vss.n8364 759.029
R7247 vss.n13669 vss.n8376 759.029
R7248 vss.n13665 vss.n8376 759.029
R7249 vss.n13676 vss.n8368 759.029
R7250 vss.n13676 vss.n8369 759.029
R7251 vss.n13671 vss.n8369 759.029
R7252 vss.n13671 vss.n8373 759.029
R7253 vss.n8368 vss.n8358 759.029
R7254 vss.n8363 vss.n8359 759.029
R7255 vss.n13678 vss.n8363 759.029
R7256 vss.n13678 vss.n8364 759.029
R7257 vss.n15662 vss.n293 759.029
R7258 vss.n15670 vss.n297 759.029
R7259 vss.n15670 vss.n298 759.029
R7260 vss.n15664 vss.n298 759.029
R7261 vss.n15677 vss.n286 759.029
R7262 vss.n15677 vss.n290 759.029
R7263 vss.n15672 vss.n290 759.029
R7264 vss.n15672 vss.n293 759.029
R7265 vss.n286 vss.n281 759.029
R7266 vss.n287 vss.n282 759.029
R7267 vss.n289 vss.n287 759.029
R7268 vss.n297 vss.n289 759.029
R7269 vss.n265 vss.n260 759.029
R7270 vss.n269 vss.n232 759.029
R7271 vss.n269 vss.n266 759.029
R7272 vss.n266 vss.n261 759.029
R7273 vss.n15707 vss.n236 759.029
R7274 vss.n15707 vss.n237 759.029
R7275 vss.n270 vss.n237 759.029
R7276 vss.n270 vss.n265 759.029
R7277 vss.n236 vss.n226 759.029
R7278 vss.n231 vss.n227 759.029
R7279 vss.n15709 vss.n231 759.029
R7280 vss.n15709 vss.n232 759.029
R7281 vss.n15719 vss.n217 759.029
R7282 vss.n15727 vss.n208 759.029
R7283 vss.n15727 vss.n221 759.029
R7284 vss.n15721 vss.n221 759.029
R7285 vss.n15734 vss.n212 759.029
R7286 vss.n15734 vss.n213 759.029
R7287 vss.n15729 vss.n213 759.029
R7288 vss.n15729 vss.n217 759.029
R7289 vss.n212 vss.n202 759.029
R7290 vss.n207 vss.n203 759.029
R7291 vss.n15736 vss.n207 759.029
R7292 vss.n15736 vss.n208 759.029
R7293 vss.n186 vss.n181 759.029
R7294 vss.n190 vss.n154 759.029
R7295 vss.n190 vss.n187 759.029
R7296 vss.n187 vss.n182 759.029
R7297 vss.n15763 vss.n158 759.029
R7298 vss.n15763 vss.n159 759.029
R7299 vss.n191 vss.n159 759.029
R7300 vss.n191 vss.n186 759.029
R7301 vss.n158 vss.n148 759.029
R7302 vss.n153 vss.n149 759.029
R7303 vss.n15765 vss.n153 759.029
R7304 vss.n15765 vss.n154 759.029
R7305 vss.n15775 vss.n139 759.029
R7306 vss.n15783 vss.n130 759.029
R7307 vss.n15783 vss.n143 759.029
R7308 vss.n15777 vss.n143 759.029
R7309 vss.n15790 vss.n134 759.029
R7310 vss.n15790 vss.n135 759.029
R7311 vss.n15785 vss.n135 759.029
R7312 vss.n15785 vss.n139 759.029
R7313 vss.n134 vss.n124 759.029
R7314 vss.n129 vss.n125 759.029
R7315 vss.n15792 vss.n129 759.029
R7316 vss.n15792 vss.n130 759.029
R7317 vss.n108 vss.n103 759.029
R7318 vss.n112 vss.n75 759.029
R7319 vss.n112 vss.n109 759.029
R7320 vss.n109 vss.n104 759.029
R7321 vss.n15819 vss.n79 759.029
R7322 vss.n15819 vss.n80 759.029
R7323 vss.n113 vss.n80 759.029
R7324 vss.n113 vss.n108 759.029
R7325 vss.n79 vss.n69 759.029
R7326 vss.n74 vss.n70 759.029
R7327 vss.n15821 vss.n74 759.029
R7328 vss.n15821 vss.n75 759.029
R7329 vss.n15831 vss.n60 759.029
R7330 vss.n15839 vss.n51 759.029
R7331 vss.n15839 vss.n64 759.029
R7332 vss.n15833 vss.n64 759.029
R7333 vss.n15846 vss.n55 759.029
R7334 vss.n15846 vss.n56 759.029
R7335 vss.n15841 vss.n56 759.029
R7336 vss.n15841 vss.n60 759.029
R7337 vss.n55 vss.n45 759.029
R7338 vss.n50 vss.n46 759.029
R7339 vss.n15848 vss.n50 759.029
R7340 vss.n15848 vss.n51 759.029
R7341 vss.n15879 vss.n23 759.029
R7342 vss.n15884 vss.n18 759.029
R7343 vss.n15884 vss.n15883 759.029
R7344 vss.n15883 vss.n22 759.029
R7345 vss.n6260 vss.n6259 759.029
R7346 vss.n6259 vss.n17 759.029
R7347 vss.n15873 vss.n17 759.029
R7348 vss.n15873 vss.n23 759.029
R7349 vss.n6260 vss.n6254 759.029
R7350 vss.n6262 vss.n6255 759.029
R7351 vss.n6262 vss.n6261 759.029
R7352 vss.n6261 vss.n18 759.029
R7353 vss.n4812 vss.n4807 759.029
R7354 vss.n4825 vss.n444 759.029
R7355 vss.n4825 vss.n4813 759.029
R7356 vss.n4813 vss.n4808 759.029
R7357 vss.n15451 vss.n448 759.029
R7358 vss.n15451 vss.n449 759.029
R7359 vss.n4826 vss.n449 759.029
R7360 vss.n4826 vss.n4812 759.029
R7361 vss.n448 vss.n438 759.029
R7362 vss.n443 vss.n439 759.029
R7363 vss.n15453 vss.n443 759.029
R7364 vss.n15453 vss.n444 759.029
R7365 vss.n4897 vss.n4292 759.029
R7366 vss.n4309 vss.n4308 759.029
R7367 vss.n4308 vss.n4296 759.029
R7368 vss.n4296 vss.n4291 759.029
R7369 vss.n4871 vss.n4361 759.029
R7370 vss.n4871 vss.n4307 759.029
R7371 vss.n4307 vss.n4306 759.029
R7372 vss.n4306 vss.n4292 759.029
R7373 vss.n4867 vss.n4361 759.029
R7374 vss.n4865 vss.n4312 759.029
R7375 vss.n4873 vss.n4312 759.029
R7376 vss.n4873 vss.n4309 759.029
R7377 vss.n15394 vss.n601 759.029
R7378 vss.n15412 vss.n545 759.029
R7379 vss.n15412 vss.n604 759.029
R7380 vss.n15395 vss.n604 759.029
R7381 vss.n15419 vss.n596 759.029
R7382 vss.n15419 vss.n597 759.029
R7383 vss.n15414 vss.n597 759.029
R7384 vss.n15414 vss.n601 759.029
R7385 vss.n596 vss.n539 759.029
R7386 vss.n544 vss.n540 759.029
R7387 vss.n15421 vss.n544 759.029
R7388 vss.n15421 vss.n545 759.029
R7389 vss.n5160 vss.n5125 759.029
R7390 vss.n5130 vss.n651 759.029
R7391 vss.n5130 vss.n5129 759.029
R7392 vss.n5129 vss.n5124 759.029
R7393 vss.n15376 vss.n655 759.029
R7394 vss.n15376 vss.n656 759.029
R7395 vss.n5131 vss.n656 759.029
R7396 vss.n5131 vss.n5125 759.029
R7397 vss.n655 vss.n645 759.029
R7398 vss.n650 vss.n646 759.029
R7399 vss.n15378 vss.n650 759.029
R7400 vss.n15378 vss.n651 759.029
R7401 vss.n5372 vss.n5337 759.029
R7402 vss.n5342 vss.n750 759.029
R7403 vss.n5342 vss.n5341 759.029
R7404 vss.n5341 vss.n5336 759.029
R7405 vss.n15346 vss.n754 759.029
R7406 vss.n15346 vss.n755 759.029
R7407 vss.n5343 vss.n755 759.029
R7408 vss.n5343 vss.n5337 759.029
R7409 vss.n754 vss.n744 759.029
R7410 vss.n749 vss.n745 759.029
R7411 vss.n15348 vss.n749 759.029
R7412 vss.n15348 vss.n750 759.029
R7413 vss.n15244 vss.n858 759.029
R7414 vss.n15262 vss.n803 759.029
R7415 vss.n15262 vss.n861 759.029
R7416 vss.n15245 vss.n861 759.029
R7417 vss.n15269 vss.n853 759.029
R7418 vss.n15269 vss.n854 759.029
R7419 vss.n15264 vss.n854 759.029
R7420 vss.n15264 vss.n858 759.029
R7421 vss.n853 vss.n797 759.029
R7422 vss.n802 vss.n798 759.029
R7423 vss.n15271 vss.n802 759.029
R7424 vss.n15271 vss.n803 759.029
R7425 vss.n6444 vss.n6409 759.029
R7426 vss.n6414 vss.n908 759.029
R7427 vss.n6414 vss.n6413 759.029
R7428 vss.n6413 vss.n6408 759.029
R7429 vss.n15226 vss.n912 759.029
R7430 vss.n15226 vss.n913 759.029
R7431 vss.n6415 vss.n913 759.029
R7432 vss.n6415 vss.n6409 759.029
R7433 vss.n912 vss.n902 759.029
R7434 vss.n907 vss.n903 759.029
R7435 vss.n15228 vss.n907 759.029
R7436 vss.n15228 vss.n908 759.029
R7437 vss.n6559 vss.n6524 759.029
R7438 vss.n6529 vss.n1083 759.029
R7439 vss.n6529 vss.n6528 759.029
R7440 vss.n6528 vss.n6523 759.029
R7441 vss.n15025 vss.n1087 759.029
R7442 vss.n15025 vss.n1088 759.029
R7443 vss.n6530 vss.n1088 759.029
R7444 vss.n6530 vss.n6524 759.029
R7445 vss.n1087 vss.n1077 759.029
R7446 vss.n1082 vss.n1078 759.029
R7447 vss.n15027 vss.n1082 759.029
R7448 vss.n15027 vss.n1083 759.029
R7449 vss.n6544 vss.n6534 759.029
R7450 vss.n6542 vss.n6533 759.029
R7451 vss.n6533 vss.n6532 759.029
R7452 vss.n6532 vss.n6518 759.029
R7453 vss.n6546 vss.n6534 759.029
R7454 vss.n6546 vss.n6521 759.029
R7455 vss.n6521 vss.n6517 759.029
R7456 vss.n6575 vss.n6517 759.029
R7457 vss.n6580 vss.n6518 759.029
R7458 vss.n6580 vss.n6519 759.029
R7459 vss.n6572 vss.n6519 759.029
R7460 vss.n6575 vss.n6574 759.029
R7461 vss.n6429 vss.n6419 759.029
R7462 vss.n6427 vss.n6418 759.029
R7463 vss.n6418 vss.n6417 759.029
R7464 vss.n6417 vss.n6403 759.029
R7465 vss.n6431 vss.n6419 759.029
R7466 vss.n6431 vss.n6406 759.029
R7467 vss.n6406 vss.n6402 759.029
R7468 vss.n6459 vss.n6402 759.029
R7469 vss.n6464 vss.n6403 759.029
R7470 vss.n6464 vss.n6404 759.029
R7471 vss.n6456 vss.n6404 759.029
R7472 vss.n6459 vss.n6458 759.029
R7473 vss.n878 vss.n877 759.029
R7474 vss.n870 vss.n865 759.029
R7475 vss.n15255 vss.n865 759.029
R7476 vss.n15255 vss.n866 759.029
R7477 vss.n878 vss.n864 759.029
R7478 vss.n884 vss.n864 759.029
R7479 vss.n887 vss.n884 759.029
R7480 vss.n891 vss.n887 759.029
R7481 vss.n15241 vss.n866 759.029
R7482 vss.n15241 vss.n15240 759.029
R7483 vss.n15240 vss.n15239 759.029
R7484 vss.n898 vss.n891 759.029
R7485 vss.n5357 vss.n5347 759.029
R7486 vss.n5355 vss.n5346 759.029
R7487 vss.n5346 vss.n5345 759.029
R7488 vss.n5345 vss.n5331 759.029
R7489 vss.n5359 vss.n5347 759.029
R7490 vss.n5359 vss.n5334 759.029
R7491 vss.n5334 vss.n5330 759.029
R7492 vss.n5387 vss.n5330 759.029
R7493 vss.n5392 vss.n5331 759.029
R7494 vss.n5392 vss.n5332 759.029
R7495 vss.n5384 vss.n5332 759.029
R7496 vss.n5387 vss.n5386 759.029
R7497 vss.n5145 vss.n5135 759.029
R7498 vss.n5143 vss.n5134 759.029
R7499 vss.n5134 vss.n5133 759.029
R7500 vss.n5133 vss.n5119 759.029
R7501 vss.n5147 vss.n5135 759.029
R7502 vss.n5147 vss.n5122 759.029
R7503 vss.n5122 vss.n5118 759.029
R7504 vss.n5175 vss.n5118 759.029
R7505 vss.n5180 vss.n5119 759.029
R7506 vss.n5180 vss.n5120 759.029
R7507 vss.n5172 vss.n5120 759.029
R7508 vss.n5175 vss.n5174 759.029
R7509 vss.n621 vss.n620 759.029
R7510 vss.n613 vss.n608 759.029
R7511 vss.n15405 vss.n608 759.029
R7512 vss.n15405 vss.n609 759.029
R7513 vss.n621 vss.n607 759.029
R7514 vss.n627 vss.n607 759.029
R7515 vss.n630 vss.n627 759.029
R7516 vss.n634 vss.n630 759.029
R7517 vss.n15391 vss.n609 759.029
R7518 vss.n15391 vss.n15390 759.029
R7519 vss.n15390 vss.n15389 759.029
R7520 vss.n641 vss.n634 759.029
R7521 vss.n4882 vss.n4300 759.029
R7522 vss.n4880 vss.n4299 759.029
R7523 vss.n4299 vss.n4298 759.029
R7524 vss.n4298 vss.n4286 759.029
R7525 vss.n4884 vss.n4300 759.029
R7526 vss.n4884 vss.n4289 759.029
R7527 vss.n4289 vss.n4285 759.029
R7528 vss.n4912 vss.n4285 759.029
R7529 vss.n4917 vss.n4286 759.029
R7530 vss.n4917 vss.n4287 759.029
R7531 vss.n4909 vss.n4287 759.029
R7532 vss.n4912 vss.n4911 759.029
R7533 vss.n4829 vss.n4817 759.029
R7534 vss.n4835 vss.n4816 759.029
R7535 vss.n4836 vss.n4835 759.029
R7536 vss.n4836 vss.n4802 759.029
R7537 vss.n4817 vss.n4815 759.029
R7538 vss.n4815 vss.n4751 759.029
R7539 vss.n4854 vss.n4751 759.029
R7540 vss.n4854 vss.n4752 759.029
R7541 vss.n4852 vss.n4802 759.029
R7542 vss.n4852 vss.n4804 759.029
R7543 vss.n4804 vss.n4746 759.029
R7544 vss.n4752 vss.n4747 759.029
R7545 vss.n3234 vss.n3229 759.029
R7546 vss.n3247 vss.n1223 759.029
R7547 vss.n3247 vss.n3235 759.029
R7548 vss.n3235 vss.n3230 759.029
R7549 vss.n14756 vss.n1227 759.029
R7550 vss.n14756 vss.n1228 759.029
R7551 vss.n3248 vss.n1228 759.029
R7552 vss.n3248 vss.n3234 759.029
R7553 vss.n1227 vss.n1217 759.029
R7554 vss.n1222 vss.n1218 759.029
R7555 vss.n14758 vss.n1222 759.029
R7556 vss.n14758 vss.n1223 759.029
R7557 vss.n8003 vss.n2431 759.029
R7558 vss.n2436 vss.n2367 759.029
R7559 vss.n2436 vss.n2432 759.029
R7560 vss.n8005 vss.n2432 759.029
R7561 vss.n8023 vss.n2417 759.029
R7562 vss.n8023 vss.n2418 759.029
R7563 vss.n2433 vss.n2418 759.029
R7564 vss.n2433 vss.n2431 759.029
R7565 vss.n2417 vss.n2361 759.029
R7566 vss.n2366 vss.n2362 759.029
R7567 vss.n8025 vss.n2366 759.029
R7568 vss.n8025 vss.n2367 759.029
R7569 vss.n14699 vss.n1380 759.029
R7570 vss.n14717 vss.n1324 759.029
R7571 vss.n14717 vss.n1383 759.029
R7572 vss.n14700 vss.n1383 759.029
R7573 vss.n14724 vss.n1375 759.029
R7574 vss.n14724 vss.n1376 759.029
R7575 vss.n14719 vss.n1376 759.029
R7576 vss.n14719 vss.n1380 759.029
R7577 vss.n1375 vss.n1318 759.029
R7578 vss.n1323 vss.n1319 759.029
R7579 vss.n14726 vss.n1323 759.029
R7580 vss.n14726 vss.n1324 759.029
R7581 vss.n7568 vss.n7533 759.029
R7582 vss.n7538 vss.n1430 759.029
R7583 vss.n7538 vss.n7537 759.029
R7584 vss.n7537 vss.n7532 759.029
R7585 vss.n14681 vss.n1434 759.029
R7586 vss.n14681 vss.n1435 759.029
R7587 vss.n7539 vss.n1435 759.029
R7588 vss.n7539 vss.n7533 759.029
R7589 vss.n1434 vss.n1424 759.029
R7590 vss.n1429 vss.n1425 759.029
R7591 vss.n14683 vss.n1429 759.029
R7592 vss.n14683 vss.n1430 759.029
R7593 vss.n2786 vss.n2751 759.029
R7594 vss.n2756 vss.n1529 759.029
R7595 vss.n2756 vss.n2755 759.029
R7596 vss.n2755 vss.n2750 759.029
R7597 vss.n14651 vss.n1533 759.029
R7598 vss.n14651 vss.n1534 759.029
R7599 vss.n2757 vss.n1534 759.029
R7600 vss.n2757 vss.n2751 759.029
R7601 vss.n1533 vss.n1523 759.029
R7602 vss.n1528 vss.n1524 759.029
R7603 vss.n14653 vss.n1528 759.029
R7604 vss.n14653 vss.n1529 759.029
R7605 vss.n14549 vss.n1637 759.029
R7606 vss.n14567 vss.n1582 759.029
R7607 vss.n14567 vss.n1640 759.029
R7608 vss.n14550 vss.n1640 759.029
R7609 vss.n14574 vss.n1632 759.029
R7610 vss.n14574 vss.n1633 759.029
R7611 vss.n14569 vss.n1633 759.029
R7612 vss.n14569 vss.n1637 759.029
R7613 vss.n1632 vss.n1576 759.029
R7614 vss.n1581 vss.n1577 759.029
R7615 vss.n14576 vss.n1581 759.029
R7616 vss.n14576 vss.n1582 759.029
R7617 vss.n2552 vss.n2517 759.029
R7618 vss.n2522 vss.n1687 759.029
R7619 vss.n2522 vss.n2521 759.029
R7620 vss.n2521 vss.n2516 759.029
R7621 vss.n14531 vss.n1691 759.029
R7622 vss.n14531 vss.n1692 759.029
R7623 vss.n2523 vss.n1692 759.029
R7624 vss.n2523 vss.n2517 759.029
R7625 vss.n1691 vss.n1681 759.029
R7626 vss.n1686 vss.n1682 759.029
R7627 vss.n14533 vss.n1686 759.029
R7628 vss.n14533 vss.n1687 759.029
R7629 vss.n1965 vss.n1871 759.029
R7630 vss.n1983 vss.n1862 759.029
R7631 vss.n1983 vss.n1874 759.029
R7632 vss.n1966 vss.n1874 759.029
R7633 vss.n14330 vss.n1866 759.029
R7634 vss.n14330 vss.n1867 759.029
R7635 vss.n1985 vss.n1867 759.029
R7636 vss.n1985 vss.n1871 759.029
R7637 vss.n1866 vss.n1856 759.029
R7638 vss.n1861 vss.n1857 759.029
R7639 vss.n14332 vss.n1861 759.029
R7640 vss.n14332 vss.n1862 759.029
R7641 vss.n1891 vss.n1890 759.029
R7642 vss.n1883 vss.n1878 759.029
R7643 vss.n1976 vss.n1878 759.029
R7644 vss.n1976 vss.n1879 759.029
R7645 vss.n1891 vss.n1877 759.029
R7646 vss.n1896 vss.n1877 759.029
R7647 vss.n1946 vss.n1896 759.029
R7648 vss.n1950 vss.n1946 759.029
R7649 vss.n1962 vss.n1879 759.029
R7650 vss.n1962 vss.n1961 759.029
R7651 vss.n1961 vss.n1960 759.029
R7652 vss.n1957 vss.n1950 759.029
R7653 vss.n2539 vss.n2527 759.029
R7654 vss.n2537 vss.n2525 759.029
R7655 vss.n2528 vss.n2525 759.029
R7656 vss.n2528 vss.n2509 759.029
R7657 vss.n2527 vss.n2526 759.029
R7658 vss.n2526 vss.n2514 759.029
R7659 vss.n2514 vss.n2508 759.029
R7660 vss.n2566 vss.n2508 759.029
R7661 vss.n2571 vss.n2509 759.029
R7662 vss.n2571 vss.n2510 759.029
R7663 vss.n2563 vss.n2510 759.029
R7664 vss.n2566 vss.n2565 759.029
R7665 vss.n1657 vss.n1656 759.029
R7666 vss.n1649 vss.n1644 759.029
R7667 vss.n14560 vss.n1644 759.029
R7668 vss.n14560 vss.n1645 759.029
R7669 vss.n1657 vss.n1643 759.029
R7670 vss.n1663 vss.n1643 759.029
R7671 vss.n1666 vss.n1663 759.029
R7672 vss.n1670 vss.n1666 759.029
R7673 vss.n14546 vss.n1645 759.029
R7674 vss.n14546 vss.n14545 759.029
R7675 vss.n14545 vss.n14544 759.029
R7676 vss.n1677 vss.n1670 759.029
R7677 vss.n2771 vss.n2761 759.029
R7678 vss.n2769 vss.n2760 759.029
R7679 vss.n2760 vss.n2759 759.029
R7680 vss.n2759 vss.n2745 759.029
R7681 vss.n2773 vss.n2761 759.029
R7682 vss.n2773 vss.n2748 759.029
R7683 vss.n2748 vss.n2744 759.029
R7684 vss.n2801 vss.n2744 759.029
R7685 vss.n2806 vss.n2745 759.029
R7686 vss.n2806 vss.n2746 759.029
R7687 vss.n2798 vss.n2746 759.029
R7688 vss.n2801 vss.n2800 759.029
R7689 vss.n7553 vss.n7543 759.029
R7690 vss.n7551 vss.n7542 759.029
R7691 vss.n7542 vss.n7541 759.029
R7692 vss.n7541 vss.n7527 759.029
R7693 vss.n7555 vss.n7543 759.029
R7694 vss.n7555 vss.n7530 759.029
R7695 vss.n7530 vss.n7526 759.029
R7696 vss.n7583 vss.n7526 759.029
R7697 vss.n7588 vss.n7527 759.029
R7698 vss.n7588 vss.n7528 759.029
R7699 vss.n7580 vss.n7528 759.029
R7700 vss.n7583 vss.n7582 759.029
R7701 vss.n1400 vss.n1399 759.029
R7702 vss.n1392 vss.n1387 759.029
R7703 vss.n14710 vss.n1387 759.029
R7704 vss.n14710 vss.n1388 759.029
R7705 vss.n1400 vss.n1386 759.029
R7706 vss.n1406 vss.n1386 759.029
R7707 vss.n1409 vss.n1406 759.029
R7708 vss.n1413 vss.n1409 759.029
R7709 vss.n14696 vss.n1388 759.029
R7710 vss.n14696 vss.n14695 759.029
R7711 vss.n14695 vss.n14694 759.029
R7712 vss.n1420 vss.n1413 759.029
R7713 vss.n2429 vss.n2422 759.029
R7714 vss.n8016 vss.n2424 759.029
R7715 vss.n2441 vss.n2424 759.029
R7716 vss.n2442 vss.n2441 759.029
R7717 vss.n2445 vss.n2429 759.029
R7718 vss.n2445 vss.n2443 759.029
R7719 vss.n6944 vss.n2443 759.029
R7720 vss.n6954 vss.n6944 759.029
R7721 vss.n6959 vss.n2442 759.029
R7722 vss.n6959 vss.n6945 759.029
R7723 vss.n6951 vss.n6945 759.029
R7724 vss.n6954 vss.n6953 759.029
R7725 vss.n3253 vss.n3252 759.029
R7726 vss.n3250 vss.n3238 759.029
R7727 vss.n3258 vss.n3238 759.029
R7728 vss.n3258 vss.n3188 759.029
R7729 vss.n3253 vss.n3237 759.029
R7730 vss.n3237 vss.n3189 759.029
R7731 vss.n3211 vss.n3189 759.029
R7732 vss.n3221 vss.n3211 759.029
R7733 vss.n3226 vss.n3188 759.029
R7734 vss.n3226 vss.n3212 759.029
R7735 vss.n3218 vss.n3212 759.029
R7736 vss.n3221 vss.n3220 759.029
R7737 vss.n12105 vss.n11873 759.029
R7738 vss.n12110 vss.n11878 759.029
R7739 vss.n12110 vss.n11879 759.029
R7740 vss.n11879 vss.n11874 759.029
R7741 vss.n12086 vss.n11937 759.029
R7742 vss.n12086 vss.n11882 759.029
R7743 vss.n12108 vss.n11882 759.029
R7744 vss.n12108 vss.n12105 759.029
R7745 vss.n12080 vss.n11939 759.029
R7746 vss.n12084 vss.n11939 759.029
R7747 vss.n12084 vss.n11878 759.029
R7748 vss.n12078 vss.n11937 759.029
R7749 vss.n10331 vss.n10274 759.029
R7750 vss.n10380 vss.n10279 759.029
R7751 vss.n10380 vss.n10280 759.029
R7752 vss.n10280 vss.n10275 759.029
R7753 vss.n10373 vss.n10334 759.029
R7754 vss.n10373 vss.n10329 759.029
R7755 vss.n10378 vss.n10329 759.029
R7756 vss.n10378 vss.n10331 759.029
R7757 vss.n10366 vss.n10338 759.029
R7758 vss.n10371 vss.n10338 759.029
R7759 vss.n10371 vss.n10279 759.029
R7760 vss.n10364 vss.n10334 759.029
R7761 vss.n8033 vss.n2358 709
R7762 vss.n8032 vss.n8031 709
R7763 vss.n14734 vss.n1315 709
R7764 vss.n14733 vss.n14732 709
R7765 vss.n14692 vss.n14691 709
R7766 vss.n14690 vss.n14689 709
R7767 vss.n14661 vss.n1520 709
R7768 vss.n14660 vss.n14659 709
R7769 vss.n14584 vss.n1573 709
R7770 vss.n14583 vss.n14582 709
R7771 vss.n14542 vss.n14541 709
R7772 vss.n14540 vss.n14539 709
R7773 vss.n14340 vss.n1853 709
R7774 vss.n14339 vss.n14338 709
R7775 vss.n4861 vss.n4860 709
R7776 vss.n4863 vss.n4862 709
R7777 vss.n15429 vss.n536 709
R7778 vss.n15428 vss.n15427 709
R7779 vss.n15387 vss.n15386 709
R7780 vss.n15385 vss.n15384 709
R7781 vss.n15356 vss.n741 709
R7782 vss.n15355 vss.n15354 709
R7783 vss.n15279 vss.n794 709
R7784 vss.n15278 vss.n15277 709
R7785 vss.n15237 vss.n15236 709
R7786 vss.n15235 vss.n15234 709
R7787 vss.n15035 vss.n1074 709
R7788 vss.n15034 vss.n15033 709
R7789 vss.n12829 vss.n12828 709
R7790 vss.n12827 vss.n12826 709
R7791 vss.n13163 vss.n8899 709
R7792 vss.n13162 vss.n13161 709
R7793 vss.n9172 vss.n9171 709
R7794 vss.n13003 vss.n13002 709
R7795 vss.n13306 vss.n13305 709
R7796 vss.n13304 vss.n13303 709
R7797 vss.n8571 vss.n8320 709
R7798 vss.n13715 vss.n13714 709
R7799 vss.n13686 vss.n8355 709
R7800 vss.n13685 vss.n13684 709
R7801 vss.n12074 vss.n12073 709
R7802 vss.n12076 vss.n12075 709
R7803 vss.n15527 vss.n15513 704.146
R7804 vss.n15527 vss.n15504 704.146
R7805 vss.n14826 vss.n14818 704.146
R7806 vss.n14832 vss.n14818 704.146
R7807 vss.n14174 vss.n14156 704.146
R7808 vss.n14167 vss.n14156 704.146
R7809 vss.n14167 vss.n14166 704.146
R7810 vss.n14166 vss.n1173 704.146
R7811 vss.n14800 vss.n1173 704.146
R7812 vss.n14800 vss.n1174 704.146
R7813 vss.n14794 vss.n1174 704.146
R7814 vss.n14794 vss.n14791 704.146
R7815 vss.n14868 vss.n14850 704.146
R7816 vss.n14861 vss.n14850 704.146
R7817 vss.n14861 vss.n14860 704.146
R7818 vss.n14860 vss.n394 704.146
R7819 vss.n15495 vss.n394 704.146
R7820 vss.n15495 vss.n395 704.146
R7821 vss.n15489 vss.n395 704.146
R7822 vss.n15489 vss.n15486 704.146
R7823 vss.n15551 vss.n15547 704.146
R7824 vss.n15551 vss.n372 704.146
R7825 vss.n15555 vss.n372 704.146
R7826 vss.n15555 vss.n365 704.146
R7827 vss.n15571 vss.n365 704.146
R7828 vss.n15571 vss.n366 704.146
R7829 vss.n15565 vss.n366 704.146
R7830 vss.n15565 vss.n303 704.146
R7831 vss.n12173 vss.n12143 704.146
R7832 vss.n12173 vss.n12144 704.146
R7833 vss.n13228 vss.n13225 704.146
R7834 vss.n13228 vss.n8828 704.146
R7835 vss.n13234 vss.n8828 704.146
R7836 vss.n13234 vss.n8819 704.146
R7837 vss.n13241 vss.n8819 704.146
R7838 vss.n13241 vss.n8820 704.146
R7839 vss.n8820 vss.n8811 704.146
R7840 vss.n13248 vss.n8811 704.146
R7841 vss.n8033 vss.n8032 704
R7842 vss.n14734 vss.n14733 704
R7843 vss.n14691 vss.n14690 704
R7844 vss.n14661 vss.n14660 704
R7845 vss.n14584 vss.n14583 704
R7846 vss.n14541 vss.n14540 704
R7847 vss.n14340 vss.n14339 704
R7848 vss.n4862 vss.n4861 704
R7849 vss.n15429 vss.n15428 704
R7850 vss.n15386 vss.n15385 704
R7851 vss.n15356 vss.n15355 704
R7852 vss.n15279 vss.n15278 704
R7853 vss.n15236 vss.n15235 704
R7854 vss.n15035 vss.n15034 704
R7855 vss.n12828 vss.n12827 704
R7856 vss.n13163 vss.n13162 704
R7857 vss.n13003 vss.n9172 704
R7858 vss.n13305 vss.n13304 704
R7859 vss.n13715 vss.n8320 704
R7860 vss.n13686 vss.n13685 704
R7861 vss.n12075 vss.n12074 704
R7862 vss.n11786 vss.n11763 700.481
R7863 vss.n11797 vss.n11763 700.481
R7864 vss.n15534 vss.n15504 694.048
R7865 vss.n12167 vss.n12144 694.048
R7866 vss.n12243 vss.n9744 691.532
R7867 vss.n12243 vss.n9737 691.532
R7868 vss.n12259 vss.n9737 691.532
R7869 vss.n12259 vss.n9738 691.532
R7870 vss.n12253 vss.n9738 691.532
R7871 vss.n12253 vss.n8687 691.532
R7872 vss.n12361 vss.n9614 691.532
R7873 vss.n12361 vss.n9607 691.532
R7874 vss.n12377 vss.n9607 691.532
R7875 vss.n12377 vss.n9608 691.532
R7876 vss.n12371 vss.n9608 691.532
R7877 vss.n12371 vss.n9207 691.532
R7878 vss.n12480 vss.n9485 691.532
R7879 vss.n12480 vss.n9478 691.532
R7880 vss.n12496 vss.n9478 691.532
R7881 vss.n12496 vss.n9479 691.532
R7882 vss.n12490 vss.n9479 691.532
R7883 vss.n12490 vss.n9280 691.532
R7884 vss.n11737 vss.n9873 691.532
R7885 vss.n11737 vss.n9866 691.532
R7886 vss.n11753 vss.n9866 691.532
R7887 vss.n11753 vss.n9867 691.532
R7888 vss.n11747 vss.n9867 691.532
R7889 vss.n11747 vss.n8806 691.532
R7890 vss.n5567 vss.n5553 691.532
R7891 vss.n5567 vss.n5546 691.532
R7892 vss.n5583 vss.n5546 691.532
R7893 vss.n5583 vss.n5547 691.532
R7894 vss.n5577 vss.n5547 691.532
R7895 vss.n5577 vss.n3730 691.532
R7896 vss.n5755 vss.n5741 691.532
R7897 vss.n5755 vss.n5734 691.532
R7898 vss.n5771 vss.n5734 691.532
R7899 vss.n5771 vss.n5735 691.532
R7900 vss.n5765 vss.n5735 691.532
R7901 vss.n5765 vss.n3849 691.532
R7902 vss.n5995 vss.n5981 691.532
R7903 vss.n5995 vss.n5974 691.532
R7904 vss.n6011 vss.n5974 691.532
R7905 vss.n6011 vss.n5975 691.532
R7906 vss.n6005 vss.n5975 691.532
R7907 vss.n6005 vss.n3968 691.532
R7908 vss.n6354 vss.n3334 691.532
R7909 vss.n6354 vss.n6344 691.532
R7910 vss.n6344 vss.n6340 691.532
R7911 vss.n6360 vss.n6340 691.532
R7912 vss.n6361 vss.n6360 691.532
R7913 vss.n6361 vss.n6335 691.532
R7914 vss.n4028 vss.n3326 691.532
R7915 vss.n4028 vss.n4020 691.532
R7916 vss.n4035 vss.n4020 691.532
R7917 vss.n4035 vss.n4014 691.532
R7918 vss.n5525 vss.n4014 691.532
R7919 vss.n5525 vss.n5524 691.532
R7920 vss.n4193 vss.n3318 691.532
R7921 vss.n4193 vss.n4184 691.532
R7922 vss.n4200 vss.n4184 691.532
R7923 vss.n4200 vss.n4199 691.532
R7924 vss.n4199 vss.n4180 691.532
R7925 vss.n4210 vss.n4180 691.532
R7926 vss.n4468 vss.n3310 691.532
R7927 vss.n4468 vss.n4459 691.532
R7928 vss.n4472 vss.n4459 691.532
R7929 vss.n4472 vss.n4452 691.532
R7930 vss.n4489 vss.n4452 691.532
R7931 vss.n4489 vss.n4453 691.532
R7932 vss.n14915 vss.n14900 691.532
R7933 vss.n14915 vss.n14893 691.532
R7934 vss.n14931 vss.n14893 691.532
R7935 vss.n14931 vss.n14894 691.532
R7936 vss.n14925 vss.n14894 691.532
R7937 vss.n14925 vss.n409 691.532
R7938 vss.n15135 vss.n15102 691.532
R7939 vss.n15135 vss.n15103 691.532
R7940 vss.n15129 vss.n15103 691.532
R7941 vss.n15129 vss.n15115 691.532
R7942 vss.n15123 vss.n15115 691.532
R7943 vss.n15123 vss.n417 691.532
R7944 vss.n3090 vss.n3076 691.532
R7945 vss.n3090 vss.n3069 691.532
R7946 vss.n3106 vss.n3069 691.532
R7947 vss.n3106 vss.n3070 691.532
R7948 vss.n3100 vss.n3070 691.532
R7949 vss.n3100 vss.n425 691.532
R7950 vss.n4681 vss.n4667 691.532
R7951 vss.n4681 vss.n4660 691.532
R7952 vss.n4697 vss.n4660 691.532
R7953 vss.n4697 vss.n4661 691.532
R7954 vss.n4691 vss.n4661 691.532
R7955 vss.n4691 vss.n433 691.532
R7956 vss.n7925 vss.n2643 691.532
R7957 vss.n2651 vss.n2643 691.532
R7958 vss.n7918 vss.n2651 691.532
R7959 vss.n7918 vss.n7917 691.532
R7960 vss.n7917 vss.n2655 691.532
R7961 vss.n2664 vss.n2655 691.532
R7962 vss.n2909 vss.n2477 691.532
R7963 vss.n2909 vss.n2899 691.532
R7964 vss.n2899 vss.n2895 691.532
R7965 vss.n2915 vss.n2895 691.532
R7966 vss.n2916 vss.n2915 691.532
R7967 vss.n2916 vss.n2890 691.532
R7968 vss.n7970 vss.n7959 691.532
R7969 vss.n7970 vss.n7960 691.532
R7970 vss.n7960 vss.n2465 691.532
R7971 vss.n7976 vss.n2465 691.532
R7972 vss.n7977 vss.n7976 691.532
R7973 vss.n7977 vss.n2460 691.532
R7974 vss.n6824 vss.n6805 691.532
R7975 vss.n6813 vss.n6805 691.532
R7976 vss.n6817 vss.n6813 691.532
R7977 vss.n6817 vss.n3144 691.532
R7978 vss.n7212 vss.n3144 691.532
R7979 vss.n7212 vss.n7211 691.532
R7980 vss.n14220 vss.n14205 691.532
R7981 vss.n14220 vss.n14198 691.532
R7982 vss.n14236 vss.n14198 691.532
R7983 vss.n14236 vss.n14199 691.532
R7984 vss.n14230 vss.n14199 691.532
R7985 vss.n14230 vss.n1188 691.532
R7986 vss.n14440 vss.n14407 691.532
R7987 vss.n14440 vss.n14408 691.532
R7988 vss.n14434 vss.n14408 691.532
R7989 vss.n14434 vss.n14420 691.532
R7990 vss.n14428 vss.n14420 691.532
R7991 vss.n14428 vss.n1196 691.532
R7992 vss.n13960 vss.n8164 691.532
R7993 vss.n13960 vss.n8157 691.532
R7994 vss.n13976 vss.n8157 691.532
R7995 vss.n13976 vss.n8158 691.532
R7996 vss.n13970 vss.n8158 691.532
R7997 vss.n13970 vss.n1204 691.532
R7998 vss.n2257 vss.n2243 691.532
R7999 vss.n2257 vss.n2236 691.532
R8000 vss.n2273 vss.n2236 691.532
R8001 vss.n2273 vss.n2237 691.532
R8002 vss.n2267 vss.n2237 691.532
R8003 vss.n2267 vss.n1212 691.532
R8004 vss.n13578 vss.n13574 691.532
R8005 vss.n13578 vss.n13568 691.532
R8006 vss.n13582 vss.n13568 691.532
R8007 vss.n13582 vss.n13561 691.532
R8008 vss.n13600 vss.n13561 691.532
R8009 vss.n13600 vss.n13562 691.532
R8010 vss.n13767 vss.n2107 691.532
R8011 vss.n13767 vss.n13758 691.532
R8012 vss.n13771 vss.n13758 691.532
R8013 vss.n13771 vss.n13751 691.532
R8014 vss.n13789 vss.n13751 691.532
R8015 vss.n13789 vss.n13752 691.532
R8016 vss.n13055 vss.n2115 691.532
R8017 vss.n13055 vss.n13046 691.532
R8018 vss.n13059 vss.n13046 691.532
R8019 vss.n13059 vss.n13039 691.532
R8020 vss.n13077 vss.n13039 691.532
R8021 vss.n13077 vss.n13040 691.532
R8022 vss.n2167 vss.n2123 691.532
R8023 vss.n2167 vss.n2158 691.532
R8024 vss.n2171 vss.n2158 691.532
R8025 vss.n2171 vss.n2151 691.532
R8026 vss.n14083 vss.n2151 691.532
R8027 vss.n14083 vss.n2152 691.532
R8028 vss.n3597 vss.n3581 691.532
R8029 vss.n3597 vss.n3572 691.532
R8030 vss.n3604 vss.n3572 691.532
R8031 vss.n3604 vss.n3573 691.532
R8032 vss.n3573 vss.n3564 691.532
R8033 vss.n3611 vss.n3564 691.532
R8034 vss.n11536 vss.n8837 691.532
R8035 vss.n11536 vss.n11527 691.532
R8036 vss.n11540 vss.n11527 691.532
R8037 vss.n11540 vss.n11520 691.532
R8038 vss.n11558 vss.n11520 691.532
R8039 vss.n11558 vss.n11521 691.532
R8040 vss.n11225 vss.n8845 691.532
R8041 vss.n11225 vss.n11216 691.532
R8042 vss.n11229 vss.n11216 691.532
R8043 vss.n11229 vss.n11209 691.532
R8044 vss.n11247 vss.n11209 691.532
R8045 vss.n11247 vss.n11210 691.532
R8046 vss.n10886 vss.n8853 691.532
R8047 vss.n10886 vss.n10877 691.532
R8048 vss.n10890 vss.n10877 691.532
R8049 vss.n10890 vss.n10870 691.532
R8050 vss.n10908 vss.n10870 691.532
R8051 vss.n10908 vss.n10871 691.532
R8052 vss.n10492 vss.n8861 691.532
R8053 vss.n10492 vss.n10483 691.532
R8054 vss.n10496 vss.n10483 691.532
R8055 vss.n10496 vss.n10476 691.532
R8056 vss.n10514 vss.n10476 691.532
R8057 vss.n10514 vss.n10477 691.532
R8058 vss.n10326 vss.n10281 669.716
R8059 vss.n10289 vss.n10281 669.716
R8060 vss.n10319 vss.n10289 669.716
R8061 vss.n10319 vss.n10318 669.716
R8062 vss.n10318 vss.n10293 669.716
R8063 vss.n10301 vss.n10293 669.716
R8064 vss.n10310 vss.n10301 669.716
R8065 vss.n10310 vss.n8864 669.716
R8066 vss.n11684 vss.n11680 669.716
R8067 vss.n11684 vss.n9923 669.716
R8068 vss.n11688 vss.n9923 669.716
R8069 vss.n11688 vss.n9916 669.716
R8070 vss.n11704 vss.n9916 669.716
R8071 vss.n11704 vss.n9917 669.716
R8072 vss.n11698 vss.n9917 669.716
R8073 vss.n11698 vss.n8839 669.716
R8074 vss.n11447 vss.n11443 669.716
R8075 vss.n11447 vss.n9978 669.716
R8076 vss.n11451 vss.n9978 669.716
R8077 vss.n11451 vss.n9971 669.716
R8078 vss.n11467 vss.n9971 669.716
R8079 vss.n11467 vss.n9972 669.716
R8080 vss.n11461 vss.n9972 669.716
R8081 vss.n11461 vss.n8843 669.716
R8082 vss.n11411 vss.n11366 669.716
R8083 vss.n11374 vss.n11366 669.716
R8084 vss.n11404 vss.n11374 669.716
R8085 vss.n11404 vss.n11375 669.716
R8086 vss.n11398 vss.n11375 669.716
R8087 vss.n11398 vss.n11384 669.716
R8088 vss.n11392 vss.n11384 669.716
R8089 vss.n11392 vss.n8840 669.716
R8090 vss.n11178 vss.n10055 669.716
R8091 vss.n11178 vss.n11169 669.716
R8092 vss.n11182 vss.n11169 669.716
R8093 vss.n11182 vss.n11162 669.716
R8094 vss.n11198 vss.n11162 669.716
R8095 vss.n11198 vss.n11163 669.716
R8096 vss.n11192 vss.n11163 669.716
R8097 vss.n11192 vss.n8847 669.716
R8098 vss.n11042 vss.n11038 669.716
R8099 vss.n11042 vss.n10138 669.716
R8100 vss.n11046 vss.n10138 669.716
R8101 vss.n11046 vss.n10131 669.716
R8102 vss.n11062 vss.n10131 669.716
R8103 vss.n11062 vss.n10132 669.716
R8104 vss.n11056 vss.n10132 669.716
R8105 vss.n11056 vss.n8851 669.716
R8106 vss.n10102 vss.n10098 669.716
R8107 vss.n10102 vss.n10092 669.716
R8108 vss.n10106 vss.n10092 669.716
R8109 vss.n10106 vss.n10085 669.716
R8110 vss.n10122 vss.n10085 669.716
R8111 vss.n10122 vss.n10086 669.716
R8112 vss.n10116 vss.n10086 669.716
R8113 vss.n10116 vss.n8848 669.716
R8114 vss.n10754 vss.n10710 669.716
R8115 vss.n10718 vss.n10710 669.716
R8116 vss.n10747 vss.n10718 669.716
R8117 vss.n10747 vss.n10719 669.716
R8118 vss.n10741 vss.n10719 669.716
R8119 vss.n10741 vss.n10726 669.716
R8120 vss.n10735 vss.n10726 669.716
R8121 vss.n10735 vss.n8855 669.716
R8122 vss.n10790 vss.n10786 669.716
R8123 vss.n10790 vss.n10225 669.716
R8124 vss.n10794 vss.n10225 669.716
R8125 vss.n10794 vss.n10218 669.716
R8126 vss.n10810 vss.n10218 669.716
R8127 vss.n10810 vss.n10219 669.716
R8128 vss.n10804 vss.n10219 669.716
R8129 vss.n10804 vss.n8859 669.716
R8130 vss.n10699 vss.n10654 669.716
R8131 vss.n10662 vss.n10654 669.716
R8132 vss.n10692 vss.n10662 669.716
R8133 vss.n10692 vss.n10663 669.716
R8134 vss.n10686 vss.n10663 669.716
R8135 vss.n10686 vss.n10672 669.716
R8136 vss.n10680 vss.n10672 669.716
R8137 vss.n10680 vss.n8856 669.716
R8138 vss.n10400 vss.n10396 669.716
R8139 vss.n10400 vss.n10267 669.716
R8140 vss.n10404 vss.n10267 669.716
R8141 vss.n10404 vss.n10260 669.716
R8142 vss.n10420 vss.n10260 669.716
R8143 vss.n10420 vss.n10261 669.716
R8144 vss.n10414 vss.n10261 669.716
R8145 vss.n10414 vss.n8863 669.716
R8146 vss.n11914 vss.n8808 669.716
R8147 vss.n11914 vss.n11906 669.716
R8148 vss.n11920 vss.n11906 669.716
R8149 vss.n11920 vss.n11897 669.716
R8150 vss.n11927 vss.n11897 669.716
R8151 vss.n11927 vss.n11898 669.716
R8152 vss.n11898 vss.n11889 669.716
R8153 vss.n11934 vss.n11889 669.716
R8154 vss.n9274 vss.n9273 669.716
R8155 vss.n9273 vss.n9257 669.716
R8156 vss.n9265 vss.n9257 669.716
R8157 vss.n9265 vss.n8889 669.716
R8158 vss.n13173 vss.n8889 669.716
R8159 vss.n13173 vss.n8890 669.716
R8160 vss.n13167 vss.n8890 669.716
R8161 vss.n13167 vss.n13164 669.716
R8162 vss.n12403 vss.n9205 669.716
R8163 vss.n12403 vss.n12394 669.716
R8164 vss.n12407 vss.n12394 669.716
R8165 vss.n12407 vss.n12387 669.716
R8166 vss.n12424 vss.n12387 669.716
R8167 vss.n12424 vss.n12388 669.716
R8168 vss.n12418 vss.n12388 669.716
R8169 vss.n12418 vss.n12415 669.716
R8170 vss.n13265 vss.n13261 669.716
R8171 vss.n13265 vss.n8631 669.716
R8172 vss.n13269 vss.n8631 669.716
R8173 vss.n13269 vss.n8624 669.716
R8174 vss.n13285 vss.n8624 669.716
R8175 vss.n13285 vss.n8625 669.716
R8176 vss.n13279 vss.n8625 669.716
R8177 vss.n13279 vss.n8440 669.716
R8178 vss.n12285 vss.n8688 669.716
R8179 vss.n12285 vss.n12276 669.716
R8180 vss.n12289 vss.n12276 669.716
R8181 vss.n12289 vss.n12269 669.716
R8182 vss.n12306 vss.n12269 669.716
R8183 vss.n12306 vss.n12270 669.716
R8184 vss.n12300 vss.n12270 669.716
R8185 vss.n12300 vss.n12297 669.716
R8186 vss.n8756 vss.n8755 669.716
R8187 vss.n8755 vss.n8739 669.716
R8188 vss.n8747 vss.n8739 669.716
R8189 vss.n8747 vss.n8345 669.716
R8190 vss.n13696 vss.n8345 669.716
R8191 vss.n13696 vss.n8346 669.716
R8192 vss.n13690 vss.n8346 669.716
R8193 vss.n13690 vss.n13687 669.716
R8194 vss.n11987 vss.n8807 669.716
R8195 vss.n11987 vss.n11979 669.716
R8196 vss.n11993 vss.n11979 669.716
R8197 vss.n11993 vss.n11970 669.716
R8198 vss.n12000 vss.n11970 669.716
R8199 vss.n12000 vss.n11971 669.716
R8200 vss.n11971 vss.n11963 669.716
R8201 vss.n12007 vss.n11963 669.716
R8202 vss.n8804 vss.n8803 669.716
R8203 vss.n8803 vss.n8758 669.716
R8204 vss.n8797 vss.n8758 669.716
R8205 vss.n8797 vss.n8766 669.716
R8206 vss.n8791 vss.n8766 669.716
R8207 vss.n8791 vss.n8776 669.716
R8208 vss.n8785 vss.n8776 669.716
R8209 vss.n8785 vss.n8782 669.716
R8210 vss.n8735 vss.n8734 669.716
R8211 vss.n8734 vss.n8690 669.716
R8212 vss.n8728 vss.n8690 669.716
R8213 vss.n8728 vss.n8697 669.716
R8214 vss.n8722 vss.n8697 669.716
R8215 vss.n8722 vss.n8707 669.716
R8216 vss.n8716 vss.n8707 669.716
R8217 vss.n8716 vss.n8713 669.716
R8218 vss.n9845 vss.n9813 669.716
R8219 vss.n9845 vss.n9814 669.716
R8220 vss.n9839 vss.n9814 669.716
R8221 vss.n9839 vss.n9825 669.716
R8222 vss.n9833 vss.n9825 669.716
R8223 vss.n9833 vss.n8737 669.716
R8224 vss.n8685 vss.n8684 669.716
R8225 vss.n8684 vss.n8639 669.716
R8226 vss.n8678 vss.n8639 669.716
R8227 vss.n8678 vss.n8647 669.716
R8228 vss.n8672 vss.n8647 669.716
R8229 vss.n8672 vss.n8657 669.716
R8230 vss.n8666 vss.n8657 669.716
R8231 vss.n8666 vss.n8663 669.716
R8232 vss.n12919 vss.n12916 669.716
R8233 vss.n12919 vss.n9199 669.716
R8234 vss.n12925 vss.n9199 669.716
R8235 vss.n12925 vss.n9190 669.716
R8236 vss.n12932 vss.n9190 669.716
R8237 vss.n12932 vss.n9191 669.716
R8238 vss.n9191 vss.n9182 669.716
R8239 vss.n12939 vss.n9182 669.716
R8240 vss.n9717 vss.n9684 669.716
R8241 vss.n9717 vss.n9685 669.716
R8242 vss.n9711 vss.n9685 669.716
R8243 vss.n9711 vss.n9696 669.716
R8244 vss.n9705 vss.n9696 669.716
R8245 vss.n9705 vss.n9702 669.716
R8246 vss.n9255 vss.n9254 669.716
R8247 vss.n9254 vss.n9209 669.716
R8248 vss.n9248 vss.n9209 669.716
R8249 vss.n9248 vss.n9217 669.716
R8250 vss.n9242 vss.n9217 669.716
R8251 vss.n9242 vss.n9227 669.716
R8252 vss.n9236 vss.n9227 669.716
R8253 vss.n9236 vss.n9233 669.716
R8254 vss.n9337 vss.n9281 669.716
R8255 vss.n9337 vss.n9329 669.716
R8256 vss.n9343 vss.n9329 669.716
R8257 vss.n9343 vss.n9320 669.716
R8258 vss.n9350 vss.n9320 669.716
R8259 vss.n9350 vss.n9321 669.716
R8260 vss.n9321 vss.n9311 669.716
R8261 vss.n9357 vss.n9311 669.716
R8262 vss.n12523 vss.n9278 669.716
R8263 vss.n12523 vss.n12515 669.716
R8264 vss.n12529 vss.n12515 669.716
R8265 vss.n12529 vss.n12506 669.716
R8266 vss.n12536 vss.n12506 669.716
R8267 vss.n12536 vss.n12507 669.716
R8268 vss.n12507 vss.n9418 669.716
R8269 vss.n12543 vss.n9418 669.716
R8270 vss.n12673 vss.n9277 669.716
R8271 vss.n12673 vss.n12665 669.716
R8272 vss.n12679 vss.n12665 669.716
R8273 vss.n12679 vss.n12656 669.716
R8274 vss.n12686 vss.n12656 669.716
R8275 vss.n12686 vss.n12657 669.716
R8276 vss.n12657 vss.n12648 669.716
R8277 vss.n12693 vss.n12648 669.716
R8278 vss.n9587 vss.n9555 669.716
R8279 vss.n9587 vss.n9556 669.716
R8280 vss.n9581 vss.n9556 669.716
R8281 vss.n9581 vss.n9567 669.716
R8282 vss.n9575 vss.n9567 669.716
R8283 vss.n9575 vss.n9276 669.716
R8284 vss.n3987 vss.n3969 669.716
R8285 vss.n3980 vss.n3969 669.716
R8286 vss.n3980 vss.n3979 669.716
R8287 vss.n3979 vss.n5 669.716
R8288 vss.n15900 vss.n5 669.716
R8289 vss.n15900 vss.n6 669.716
R8290 vss.n15894 vss.n6 669.716
R8291 vss.n15894 vss.n15891 669.716
R8292 vss.n5653 vss.n3660 669.716
R8293 vss.n5653 vss.n5644 669.716
R8294 vss.n5657 vss.n5644 669.716
R8295 vss.n5657 vss.n5637 669.716
R8296 vss.n5673 vss.n5637 669.716
R8297 vss.n5673 vss.n5638 669.716
R8298 vss.n5667 vss.n5638 669.716
R8299 vss.n5667 vss.n224 669.716
R8300 vss.n3728 vss.n3727 669.716
R8301 vss.n3727 vss.n3711 669.716
R8302 vss.n3719 vss.n3711 669.716
R8303 vss.n3719 vss.n170 669.716
R8304 vss.n15753 vss.n170 669.716
R8305 vss.n15753 vss.n171 669.716
R8306 vss.n15747 vss.n171 669.716
R8307 vss.n15747 vss.n15744 669.716
R8308 vss.n3709 vss.n3708 669.716
R8309 vss.n3708 vss.n3664 669.716
R8310 vss.n3702 vss.n3664 669.716
R8311 vss.n3702 vss.n3671 669.716
R8312 vss.n3696 vss.n3671 669.716
R8313 vss.n3696 vss.n3681 669.716
R8314 vss.n3690 vss.n3681 669.716
R8315 vss.n3690 vss.n3687 669.716
R8316 vss.n5845 vss.n3779 669.716
R8317 vss.n5845 vss.n5836 669.716
R8318 vss.n5849 vss.n5836 669.716
R8319 vss.n5849 vss.n5829 669.716
R8320 vss.n5865 vss.n5829 669.716
R8321 vss.n5865 vss.n5830 669.716
R8322 vss.n5859 vss.n5830 669.716
R8323 vss.n5859 vss.n146 669.716
R8324 vss.n3847 vss.n3846 669.716
R8325 vss.n3846 vss.n3830 669.716
R8326 vss.n3838 vss.n3830 669.716
R8327 vss.n3838 vss.n92 669.716
R8328 vss.n15809 vss.n92 669.716
R8329 vss.n15809 vss.n93 669.716
R8330 vss.n15803 vss.n93 669.716
R8331 vss.n15803 vss.n15800 669.716
R8332 vss.n3828 vss.n3827 669.716
R8333 vss.n3827 vss.n3783 669.716
R8334 vss.n3821 vss.n3783 669.716
R8335 vss.n3821 vss.n3790 669.716
R8336 vss.n3815 vss.n3790 669.716
R8337 vss.n3815 vss.n3800 669.716
R8338 vss.n3809 vss.n3800 669.716
R8339 vss.n3809 vss.n3806 669.716
R8340 vss.n3947 vss.n3946 669.716
R8341 vss.n3946 vss.n3902 669.716
R8342 vss.n3940 vss.n3902 669.716
R8343 vss.n3940 vss.n3909 669.716
R8344 vss.n3934 vss.n3909 669.716
R8345 vss.n3934 vss.n3919 669.716
R8346 vss.n3928 vss.n3919 669.716
R8347 vss.n3928 vss.n3925 669.716
R8348 vss.n6085 vss.n3898 669.716
R8349 vss.n6085 vss.n6076 669.716
R8350 vss.n6089 vss.n6076 669.716
R8351 vss.n6089 vss.n6069 669.716
R8352 vss.n6105 vss.n6069 669.716
R8353 vss.n6105 vss.n6070 669.716
R8354 vss.n6099 vss.n6070 669.716
R8355 vss.n6099 vss.n67 669.716
R8356 vss.n5612 vss.n5600 669.716
R8357 vss.n5612 vss.n5593 669.716
R8358 vss.n5628 vss.n5593 669.716
R8359 vss.n5628 vss.n5594 669.716
R8360 vss.n5622 vss.n5594 669.716
R8361 vss.n5622 vss.n3662 669.716
R8362 vss.n5906 vss.n5874 669.716
R8363 vss.n5906 vss.n5875 669.716
R8364 vss.n5900 vss.n5875 669.716
R8365 vss.n5900 vss.n5886 669.716
R8366 vss.n5894 vss.n5886 669.716
R8367 vss.n5894 vss.n3781 669.716
R8368 vss.n6145 vss.n6113 669.716
R8369 vss.n6145 vss.n6114 669.716
R8370 vss.n6139 vss.n6114 669.716
R8371 vss.n6139 vss.n6125 669.716
R8372 vss.n6133 vss.n6125 669.716
R8373 vss.n6133 vss.n3900 669.716
R8374 vss.n4553 vss.n4366 669.716
R8375 vss.n4374 vss.n4366 669.716
R8376 vss.n4546 vss.n4374 669.716
R8377 vss.n4546 vss.n4375 669.716
R8378 vss.n4398 vss.n4375 669.716
R8379 vss.n4398 vss.n4384 669.716
R8380 vss.n4392 vss.n4384 669.716
R8381 vss.n4392 vss.n3309 669.716
R8382 vss.n6636 vss.n1075 669.716
R8383 vss.n6636 vss.n6627 669.716
R8384 vss.n6640 vss.n6627 669.716
R8385 vss.n6640 vss.n6620 669.716
R8386 vss.n6656 vss.n6620 669.716
R8387 vss.n6656 vss.n6621 669.716
R8388 vss.n6650 vss.n6621 669.716
R8389 vss.n6650 vss.n3333 669.716
R8390 vss.n6587 vss.n6583 669.716
R8391 vss.n6587 vss.n6509 669.716
R8392 vss.n6591 vss.n6509 669.716
R8393 vss.n6591 vss.n6502 669.716
R8394 vss.n6608 vss.n6502 669.716
R8395 vss.n6608 vss.n6503 669.716
R8396 vss.n6602 vss.n6503 669.716
R8397 vss.n6602 vss.n6599 669.716
R8398 vss.n5234 vss.n795 669.716
R8399 vss.n5234 vss.n5225 669.716
R8400 vss.n5238 vss.n5225 669.716
R8401 vss.n5238 vss.n5218 669.716
R8402 vss.n5254 vss.n5218 669.716
R8403 vss.n5254 vss.n5219 669.716
R8404 vss.n5248 vss.n5219 669.716
R8405 vss.n5248 vss.n3325 669.716
R8406 vss.n5446 vss.n742 669.716
R8407 vss.n5446 vss.n5437 669.716
R8408 vss.n5450 vss.n5437 669.716
R8409 vss.n5450 vss.n5430 669.716
R8410 vss.n5466 vss.n5430 669.716
R8411 vss.n5466 vss.n5431 669.716
R8412 vss.n5460 vss.n5431 669.716
R8413 vss.n5460 vss.n3321 669.716
R8414 vss.n5399 vss.n5395 669.716
R8415 vss.n5399 vss.n5322 669.716
R8416 vss.n5403 vss.n5322 669.716
R8417 vss.n5403 vss.n5315 669.716
R8418 vss.n5419 vss.n5315 669.716
R8419 vss.n5419 vss.n5316 669.716
R8420 vss.n5413 vss.n5316 669.716
R8421 vss.n5413 vss.n3324 669.716
R8422 vss.n4149 vss.n643 669.716
R8423 vss.n4149 vss.n4140 669.716
R8424 vss.n4153 vss.n4140 669.716
R8425 vss.n4153 vss.n4133 669.716
R8426 vss.n4169 vss.n4133 669.716
R8427 vss.n4169 vss.n4134 669.716
R8428 vss.n4163 vss.n4134 669.716
R8429 vss.n4163 vss.n3317 669.716
R8430 vss.n4972 vss.n537 669.716
R8431 vss.n4972 vss.n4963 669.716
R8432 vss.n4976 vss.n4963 669.716
R8433 vss.n4976 vss.n4956 669.716
R8434 vss.n4992 vss.n4956 669.716
R8435 vss.n4992 vss.n4957 669.716
R8436 vss.n4986 vss.n4957 669.716
R8437 vss.n4986 vss.n3313 669.716
R8438 vss.n4103 vss.n628 669.716
R8439 vss.n4103 vss.n4094 669.716
R8440 vss.n4107 vss.n4094 669.716
R8441 vss.n4107 vss.n4087 669.716
R8442 vss.n4123 vss.n4087 669.716
R8443 vss.n4123 vss.n4088 669.716
R8444 vss.n4117 vss.n4088 669.716
R8445 vss.n4117 vss.n3316 669.716
R8446 vss.n4924 vss.n4920 669.716
R8447 vss.n4924 vss.n4277 669.716
R8448 vss.n4928 vss.n4277 669.716
R8449 vss.n4928 vss.n4270 669.716
R8450 vss.n4944 vss.n4270 669.716
R8451 vss.n4944 vss.n4271 669.716
R8452 vss.n4938 vss.n4271 669.716
R8453 vss.n4938 vss.n3312 669.716
R8454 vss.n5187 vss.n5183 669.716
R8455 vss.n5187 vss.n5110 669.716
R8456 vss.n5191 vss.n5110 669.716
R8457 vss.n5191 vss.n5103 669.716
R8458 vss.n5207 vss.n5103 669.716
R8459 vss.n5207 vss.n5104 669.716
R8460 vss.n5201 vss.n5104 669.716
R8461 vss.n5201 vss.n3320 669.716
R8462 vss.n3362 vss.n885 669.716
R8463 vss.n3362 vss.n3353 669.716
R8464 vss.n3366 vss.n3353 669.716
R8465 vss.n3366 vss.n3346 669.716
R8466 vss.n3382 vss.n3346 669.716
R8467 vss.n3382 vss.n3347 669.716
R8468 vss.n3376 vss.n3347 669.716
R8469 vss.n3376 vss.n3328 669.716
R8470 vss.n3409 vss.n900 669.716
R8471 vss.n3409 vss.n3400 669.716
R8472 vss.n3413 vss.n3400 669.716
R8473 vss.n3413 vss.n3393 669.716
R8474 vss.n3429 vss.n3393 669.716
R8475 vss.n3429 vss.n3394 669.716
R8476 vss.n3423 vss.n3394 669.716
R8477 vss.n3423 vss.n3329 669.716
R8478 vss.n6471 vss.n6467 669.716
R8479 vss.n6471 vss.n6394 669.716
R8480 vss.n6475 vss.n6394 669.716
R8481 vss.n6475 vss.n6387 669.716
R8482 vss.n6491 vss.n6387 669.716
R8483 vss.n6491 vss.n6388 669.716
R8484 vss.n6485 vss.n6388 669.716
R8485 vss.n6485 vss.n3332 669.716
R8486 vss.n3510 vss.n3330 669.716
R8487 vss.n3510 vss.n3502 669.716
R8488 vss.n3516 vss.n3502 669.716
R8489 vss.n3516 vss.n3496 669.716
R8490 vss.n3527 vss.n3496 669.716
R8491 vss.n3527 vss.n3526 669.716
R8492 vss.n4059 vss.n3322 669.716
R8493 vss.n4059 vss.n4050 669.716
R8494 vss.n4063 vss.n4050 669.716
R8495 vss.n4063 vss.n4043 669.716
R8496 vss.n4078 vss.n4043 669.716
R8497 vss.n4078 vss.n4044 669.716
R8498 vss.n4240 vss.n3314 669.716
R8499 vss.n4240 vss.n4231 669.716
R8500 vss.n4244 vss.n4231 669.716
R8501 vss.n4244 vss.n4224 669.716
R8502 vss.n4259 vss.n4224 669.716
R8503 vss.n4259 vss.n4225 669.716
R8504 vss.n4799 vss.n4753 669.716
R8505 vss.n4761 vss.n4753 669.716
R8506 vss.n4792 vss.n4761 669.716
R8507 vss.n4792 vss.n4762 669.716
R8508 vss.n4785 vss.n4762 669.716
R8509 vss.n4785 vss.n4771 669.716
R8510 vss.n4779 vss.n4771 669.716
R8511 vss.n4779 vss.n3308 669.716
R8512 vss.n1062 vss.n407 669.716
R8513 vss.n1062 vss.n1053 669.716
R8514 vss.n1066 vss.n1053 669.716
R8515 vss.n1066 vss.n1046 669.716
R8516 vss.n15045 vss.n1046 669.716
R8517 vss.n15045 vss.n1047 669.716
R8518 vss.n15039 vss.n1047 669.716
R8519 vss.n15039 vss.n15036 669.716
R8520 vss.n524 vss.n427 669.716
R8521 vss.n524 vss.n515 669.716
R8522 vss.n528 vss.n515 669.716
R8523 vss.n528 vss.n508 669.716
R8524 vss.n15439 vss.n508 669.716
R8525 vss.n15439 vss.n509 669.716
R8526 vss.n15433 vss.n509 669.716
R8527 vss.n15433 vss.n15430 669.716
R8528 vss.n7322 vss.n423 669.716
R8529 vss.n7322 vss.n7313 669.716
R8530 vss.n7326 vss.n7313 669.716
R8531 vss.n7326 vss.n7306 669.716
R8532 vss.n7342 vss.n7306 669.716
R8533 vss.n7342 vss.n7307 669.716
R8534 vss.n7336 vss.n7307 669.716
R8535 vss.n7336 vss.n642 669.716
R8536 vss.n729 vss.n419 669.716
R8537 vss.n729 vss.n720 669.716
R8538 vss.n733 vss.n720 669.716
R8539 vss.n733 vss.n713 669.716
R8540 vss.n15366 vss.n713 669.716
R8541 vss.n15366 vss.n714 669.716
R8542 vss.n15360 vss.n714 669.716
R8543 vss.n15360 vss.n15357 669.716
R8544 vss.n782 vss.n415 669.716
R8545 vss.n782 vss.n773 669.716
R8546 vss.n786 vss.n773 669.716
R8547 vss.n786 vss.n766 669.716
R8548 vss.n15289 vss.n766 669.716
R8549 vss.n15289 vss.n767 669.716
R8550 vss.n15283 vss.n767 669.716
R8551 vss.n15283 vss.n15280 669.716
R8552 vss.n15196 vss.n411 669.716
R8553 vss.n15196 vss.n15187 669.716
R8554 vss.n15200 vss.n15187 669.716
R8555 vss.n15200 vss.n15180 669.716
R8556 vss.n15216 vss.n15180 669.716
R8557 vss.n15216 vss.n15181 669.716
R8558 vss.n15210 vss.n15181 669.716
R8559 vss.n15210 vss.n899 669.716
R8560 vss.n939 vss.n410 669.716
R8561 vss.n939 vss.n930 669.716
R8562 vss.n943 vss.n930 669.716
R8563 vss.n943 vss.n923 669.716
R8564 vss.n960 vss.n923 669.716
R8565 vss.n960 vss.n924 669.716
R8566 vss.n954 vss.n924 669.716
R8567 vss.n954 vss.n951 669.716
R8568 vss.n830 vss.n414 669.716
R8569 vss.n830 vss.n822 669.716
R8570 vss.n836 vss.n822 669.716
R8571 vss.n836 vss.n813 669.716
R8572 vss.n843 vss.n813 669.716
R8573 vss.n843 vss.n814 669.716
R8574 vss.n814 vss.n805 669.716
R8575 vss.n850 vss.n805 669.716
R8576 vss.n15316 vss.n418 669.716
R8577 vss.n15316 vss.n15307 669.716
R8578 vss.n15320 vss.n15307 669.716
R8579 vss.n15320 vss.n15300 669.716
R8580 vss.n15337 vss.n15300 669.716
R8581 vss.n15337 vss.n15301 669.716
R8582 vss.n15331 vss.n15301 669.716
R8583 vss.n15331 vss.n15328 669.716
R8584 vss.n682 vss.n422 669.716
R8585 vss.n682 vss.n673 669.716
R8586 vss.n686 vss.n673 669.716
R8587 vss.n686 vss.n666 669.716
R8588 vss.n703 vss.n666 669.716
R8589 vss.n703 vss.n667 669.716
R8590 vss.n697 vss.n667 669.716
R8591 vss.n697 vss.n694 669.716
R8592 vss.n7433 vss.n7401 669.716
R8593 vss.n7433 vss.n7402 669.716
R8594 vss.n7427 vss.n7402 669.716
R8595 vss.n7427 vss.n7413 669.716
R8596 vss.n7421 vss.n7413 669.716
R8597 vss.n7421 vss.n421 669.716
R8598 vss.n573 vss.n426 669.716
R8599 vss.n573 vss.n565 669.716
R8600 vss.n579 vss.n565 669.716
R8601 vss.n579 vss.n556 669.716
R8602 vss.n586 vss.n556 669.716
R8603 vss.n586 vss.n557 669.716
R8604 vss.n557 vss.n547 669.716
R8605 vss.n593 vss.n547 669.716
R8606 vss.n474 vss.n434 669.716
R8607 vss.n474 vss.n465 669.716
R8608 vss.n478 vss.n465 669.716
R8609 vss.n478 vss.n458 669.716
R8610 vss.n495 vss.n458 669.716
R8611 vss.n495 vss.n459 669.716
R8612 vss.n489 vss.n459 669.716
R8613 vss.n489 vss.n486 669.716
R8614 vss.n4724 vss.n431 669.716
R8615 vss.n4724 vss.n4716 669.716
R8616 vss.n4730 vss.n4716 669.716
R8617 vss.n4730 vss.n4707 669.716
R8618 vss.n4737 vss.n4707 669.716
R8619 vss.n4737 vss.n4708 669.716
R8620 vss.n4708 vss.n4554 669.716
R8621 vss.n4744 vss.n4554 669.716
R8622 vss.n4339 vss.n430 669.716
R8623 vss.n4339 vss.n4331 669.716
R8624 vss.n4345 vss.n4331 669.716
R8625 vss.n4345 vss.n4322 669.716
R8626 vss.n4352 vss.n4322 669.716
R8627 vss.n4352 vss.n4323 669.716
R8628 vss.n4323 vss.n4314 669.716
R8629 vss.n4359 vss.n4314 669.716
R8630 vss.n7263 vss.n7231 669.716
R8631 vss.n7263 vss.n7232 669.716
R8632 vss.n7257 vss.n7232 669.716
R8633 vss.n7257 vss.n7243 669.716
R8634 vss.n7251 vss.n7243 669.716
R8635 vss.n7251 vss.n429 669.716
R8636 vss.n6852 vss.n2359 669.716
R8637 vss.n6852 vss.n6843 669.716
R8638 vss.n6856 vss.n6843 669.716
R8639 vss.n6856 vss.n6836 669.716
R8640 vss.n6872 vss.n6836 669.716
R8641 vss.n6872 vss.n6837 669.716
R8642 vss.n6866 vss.n6837 669.716
R8643 vss.n6866 vss.n6804 669.716
R8644 vss.n2621 vss.n1854 669.716
R8645 vss.n2621 vss.n2612 669.716
R8646 vss.n2627 vss.n2612 669.716
R8647 vss.n2627 vss.n2606 669.716
R8648 vss.n2635 vss.n2606 669.716
R8649 vss.n2635 vss.n2607 669.716
R8650 vss.n2607 vss.n2598 669.716
R8651 vss.n2642 vss.n2598 669.716
R8652 vss.n1944 vss.n1897 669.716
R8653 vss.n1905 vss.n1897 669.716
R8654 vss.n1937 vss.n1905 669.716
R8655 vss.n1937 vss.n1906 669.716
R8656 vss.n1930 vss.n1906 669.716
R8657 vss.n1930 vss.n1915 669.716
R8658 vss.n1924 vss.n1915 669.716
R8659 vss.n1924 vss.n1921 669.716
R8660 vss.n2859 vss.n1574 669.716
R8661 vss.n2859 vss.n2850 669.716
R8662 vss.n2863 vss.n2850 669.716
R8663 vss.n2863 vss.n2843 669.716
R8664 vss.n2879 vss.n2843 669.716
R8665 vss.n2879 vss.n2844 669.716
R8666 vss.n2873 vss.n2844 669.716
R8667 vss.n2873 vss.n2476 669.716
R8668 vss.n7643 vss.n1521 669.716
R8669 vss.n7643 vss.n7634 669.716
R8670 vss.n7647 vss.n7634 669.716
R8671 vss.n7647 vss.n7627 669.716
R8672 vss.n7663 vss.n7627 669.716
R8673 vss.n7663 vss.n7628 669.716
R8674 vss.n7657 vss.n7628 669.716
R8675 vss.n7657 vss.n2472 669.716
R8676 vss.n2813 vss.n2809 669.716
R8677 vss.n2813 vss.n2736 669.716
R8678 vss.n2817 vss.n2736 669.716
R8679 vss.n2817 vss.n2729 669.716
R8680 vss.n2833 vss.n2729 669.716
R8681 vss.n2833 vss.n2730 669.716
R8682 vss.n2827 vss.n2730 669.716
R8683 vss.n2827 vss.n2475 669.716
R8684 vss.n2951 vss.n1422 669.716
R8685 vss.n2951 vss.n2942 669.716
R8686 vss.n2955 vss.n2942 669.716
R8687 vss.n2955 vss.n2935 669.716
R8688 vss.n2972 vss.n2935 669.716
R8689 vss.n2972 vss.n2936 669.716
R8690 vss.n2966 vss.n2936 669.716
R8691 vss.n2966 vss.n2963 669.716
R8692 vss.n7010 vss.n1316 669.716
R8693 vss.n7010 vss.n7001 669.716
R8694 vss.n7016 vss.n7001 669.716
R8695 vss.n7016 vss.n6995 669.716
R8696 vss.n7024 vss.n6995 669.716
R8697 vss.n7024 vss.n6996 669.716
R8698 vss.n6996 vss.n6987 669.716
R8699 vss.n7031 vss.n6987 669.716
R8700 vss.n7149 vss.n1407 669.716
R8701 vss.n7149 vss.n7141 669.716
R8702 vss.n7155 vss.n7141 669.716
R8703 vss.n7155 vss.n7132 669.716
R8704 vss.n7162 vss.n7132 669.716
R8705 vss.n7162 vss.n7133 669.716
R8706 vss.n7133 vss.n7124 669.716
R8707 vss.n7169 vss.n7124 669.716
R8708 vss.n6965 vss.n6962 669.716
R8709 vss.n6965 vss.n6937 669.716
R8710 vss.n6971 vss.n6937 669.716
R8711 vss.n6971 vss.n6928 669.716
R8712 vss.n6979 vss.n6928 669.716
R8713 vss.n6979 vss.n6929 669.716
R8714 vss.n6929 vss.n6920 669.716
R8715 vss.n6986 vss.n6920 669.716
R8716 vss.n7595 vss.n7591 669.716
R8717 vss.n7595 vss.n7518 669.716
R8718 vss.n7599 vss.n7518 669.716
R8719 vss.n7599 vss.n7511 669.716
R8720 vss.n7615 vss.n7511 669.716
R8721 vss.n7615 vss.n7512 669.716
R8722 vss.n7609 vss.n7512 669.716
R8723 vss.n7609 vss.n2471 669.716
R8724 vss.n7790 vss.n1664 669.716
R8725 vss.n7790 vss.n7781 669.716
R8726 vss.n7794 vss.n7781 669.716
R8727 vss.n7794 vss.n7774 669.716
R8728 vss.n7810 vss.n7774 669.716
R8729 vss.n7810 vss.n7775 669.716
R8730 vss.n7804 vss.n7775 669.716
R8731 vss.n7804 vss.n2479 669.716
R8732 vss.n7838 vss.n1679 669.716
R8733 vss.n7838 vss.n7829 669.716
R8734 vss.n7842 vss.n7829 669.716
R8735 vss.n7842 vss.n7822 669.716
R8736 vss.n7858 vss.n7822 669.716
R8737 vss.n7858 vss.n7823 669.716
R8738 vss.n7852 vss.n7823 669.716
R8739 vss.n7852 vss.n2480 669.716
R8740 vss.n2577 vss.n2574 669.716
R8741 vss.n2577 vss.n2500 669.716
R8742 vss.n2583 vss.n2500 669.716
R8743 vss.n2583 vss.n2491 669.716
R8744 vss.n2590 vss.n2491 669.716
R8745 vss.n2590 vss.n2492 669.716
R8746 vss.n2492 vss.n2483 669.716
R8747 vss.n2597 vss.n2483 669.716
R8748 vss.n2700 vss.n2481 669.716
R8749 vss.n2700 vss.n2691 669.716
R8750 vss.n2704 vss.n2691 669.716
R8751 vss.n2704 vss.n2684 669.716
R8752 vss.n2719 vss.n2684 669.716
R8753 vss.n2719 vss.n2685 669.716
R8754 vss.n3034 vss.n2473 669.716
R8755 vss.n3034 vss.n3026 669.716
R8756 vss.n3040 vss.n3026 669.716
R8757 vss.n3040 vss.n3020 669.716
R8758 vss.n3051 vss.n3020 669.716
R8759 vss.n3051 vss.n3050 669.716
R8760 vss.n7076 vss.n7032 669.716
R8761 vss.n7040 vss.n7032 669.716
R8762 vss.n7069 vss.n7040 669.716
R8763 vss.n7069 vss.n7068 669.716
R8764 vss.n7068 vss.n7044 669.716
R8765 vss.n7060 vss.n7044 669.716
R8766 vss.n3209 vss.n3191 669.716
R8767 vss.n3198 vss.n3191 669.716
R8768 vss.n3202 vss.n3198 669.716
R8769 vss.n3202 vss.n3177 669.716
R8770 vss.n6796 vss.n3177 669.716
R8771 vss.n6796 vss.n3178 669.716
R8772 vss.n3178 vss.n3169 669.716
R8773 vss.n6803 vss.n3169 669.716
R8774 vss.n1841 vss.n1186 669.716
R8775 vss.n1841 vss.n1832 669.716
R8776 vss.n1845 vss.n1832 669.716
R8777 vss.n1845 vss.n1825 669.716
R8778 vss.n14350 vss.n1825 669.716
R8779 vss.n14350 vss.n1826 669.716
R8780 vss.n14344 vss.n1826 669.716
R8781 vss.n14344 vss.n14341 669.716
R8782 vss.n1303 vss.n1206 669.716
R8783 vss.n1303 vss.n1294 669.716
R8784 vss.n1307 vss.n1294 669.716
R8785 vss.n1307 vss.n1287 669.716
R8786 vss.n14744 vss.n1287 669.716
R8787 vss.n14744 vss.n1288 669.716
R8788 vss.n14738 vss.n1288 669.716
R8789 vss.n14738 vss.n14735 669.716
R8790 vss.n14002 vss.n1202 669.716
R8791 vss.n14002 vss.n13993 669.716
R8792 vss.n14006 vss.n13993 669.716
R8793 vss.n14006 vss.n13986 669.716
R8794 vss.n14022 vss.n13986 669.716
R8795 vss.n14022 vss.n13987 669.716
R8796 vss.n14016 vss.n13987 669.716
R8797 vss.n14016 vss.n1421 669.716
R8798 vss.n1508 vss.n1198 669.716
R8799 vss.n1508 vss.n1499 669.716
R8800 vss.n1512 vss.n1499 669.716
R8801 vss.n1512 vss.n1492 669.716
R8802 vss.n14671 vss.n1492 669.716
R8803 vss.n14671 vss.n1493 669.716
R8804 vss.n14665 vss.n1493 669.716
R8805 vss.n14665 vss.n14662 669.716
R8806 vss.n1561 vss.n1194 669.716
R8807 vss.n1561 vss.n1552 669.716
R8808 vss.n1565 vss.n1552 669.716
R8809 vss.n1565 vss.n1545 669.716
R8810 vss.n14594 vss.n1545 669.716
R8811 vss.n14594 vss.n1546 669.716
R8812 vss.n14588 vss.n1546 669.716
R8813 vss.n14588 vss.n14585 669.716
R8814 vss.n14501 vss.n1190 669.716
R8815 vss.n14501 vss.n14492 669.716
R8816 vss.n14505 vss.n14492 669.716
R8817 vss.n14505 vss.n14485 669.716
R8818 vss.n14521 vss.n14485 669.716
R8819 vss.n14521 vss.n14486 669.716
R8820 vss.n14515 vss.n14486 669.716
R8821 vss.n14515 vss.n1678 669.716
R8822 vss.n1718 vss.n1189 669.716
R8823 vss.n1718 vss.n1709 669.716
R8824 vss.n1722 vss.n1709 669.716
R8825 vss.n1722 vss.n1702 669.716
R8826 vss.n1739 vss.n1702 669.716
R8827 vss.n1739 vss.n1703 669.716
R8828 vss.n1733 vss.n1703 669.716
R8829 vss.n1733 vss.n1730 669.716
R8830 vss.n1609 vss.n1193 669.716
R8831 vss.n1609 vss.n1601 669.716
R8832 vss.n1615 vss.n1601 669.716
R8833 vss.n1615 vss.n1592 669.716
R8834 vss.n1622 vss.n1592 669.716
R8835 vss.n1622 vss.n1593 669.716
R8836 vss.n1593 vss.n1584 669.716
R8837 vss.n1629 vss.n1584 669.716
R8838 vss.n14621 vss.n1197 669.716
R8839 vss.n14621 vss.n14612 669.716
R8840 vss.n14625 vss.n14612 669.716
R8841 vss.n14625 vss.n14605 669.716
R8842 vss.n14642 vss.n14605 669.716
R8843 vss.n14642 vss.n14606 669.716
R8844 vss.n14636 vss.n14606 669.716
R8845 vss.n14636 vss.n14633 669.716
R8846 vss.n1461 vss.n1201 669.716
R8847 vss.n1461 vss.n1452 669.716
R8848 vss.n1465 vss.n1452 669.716
R8849 vss.n1465 vss.n1445 669.716
R8850 vss.n1482 vss.n1445 669.716
R8851 vss.n1482 vss.n1446 669.716
R8852 vss.n1476 vss.n1446 669.716
R8853 vss.n1476 vss.n1473 669.716
R8854 vss.n13898 vss.n13866 669.716
R8855 vss.n13898 vss.n13867 669.716
R8856 vss.n13892 vss.n13867 669.716
R8857 vss.n13892 vss.n13878 669.716
R8858 vss.n13886 vss.n13878 669.716
R8859 vss.n13886 vss.n1200 669.716
R8860 vss.n1352 vss.n1205 669.716
R8861 vss.n1352 vss.n1344 669.716
R8862 vss.n1358 vss.n1344 669.716
R8863 vss.n1358 vss.n1335 669.716
R8864 vss.n1365 vss.n1335 669.716
R8865 vss.n1365 vss.n1336 669.716
R8866 vss.n1336 vss.n1326 669.716
R8867 vss.n1372 vss.n1326 669.716
R8868 vss.n1253 vss.n1213 669.716
R8869 vss.n1253 vss.n1244 669.716
R8870 vss.n1257 vss.n1244 669.716
R8871 vss.n1257 vss.n1237 669.716
R8872 vss.n1274 vss.n1237 669.716
R8873 vss.n1274 vss.n1238 669.716
R8874 vss.n1268 vss.n1238 669.716
R8875 vss.n1268 vss.n1265 669.716
R8876 vss.n2346 vss.n1210 669.716
R8877 vss.n2346 vss.n2337 669.716
R8878 vss.n2350 vss.n2337 669.716
R8879 vss.n2350 vss.n2330 669.716
R8880 vss.n8043 vss.n2330 669.716
R8881 vss.n8043 vss.n2331 669.716
R8882 vss.n8037 vss.n2331 669.716
R8883 vss.n8037 vss.n8034 669.716
R8884 vss.n2394 vss.n1209 669.716
R8885 vss.n2394 vss.n2386 669.716
R8886 vss.n2400 vss.n2386 669.716
R8887 vss.n2400 vss.n2377 669.716
R8888 vss.n2407 vss.n2377 669.716
R8889 vss.n2407 vss.n2378 669.716
R8890 vss.n2378 vss.n2369 669.716
R8891 vss.n2414 vss.n2369 669.716
R8892 vss.n8137 vss.n8105 669.716
R8893 vss.n8137 vss.n8106 669.716
R8894 vss.n8131 vss.n8106 669.716
R8895 vss.n8131 vss.n8117 669.716
R8896 vss.n8125 vss.n8117 669.716
R8897 vss.n8125 vss.n1208 669.716
R8898 vss.n11962 vss.n11944 669.716
R8899 vss.n11951 vss.n11944 669.716
R8900 vss.n11955 vss.n11951 669.716
R8901 vss.n11955 vss.n2092 669.716
R8902 vss.n14134 vss.n2092 669.716
R8903 vss.n14134 vss.n2093 669.716
R8904 vss.n14128 vss.n2093 669.716
R8905 vss.n14128 vss.n14125 669.716
R8906 vss.n13488 vss.n8356 669.716
R8907 vss.n13488 vss.n13479 669.716
R8908 vss.n13492 vss.n13479 669.716
R8909 vss.n13492 vss.n13472 669.716
R8910 vss.n13508 vss.n13472 669.716
R8911 vss.n13508 vss.n13473 669.716
R8912 vss.n13502 vss.n13473 669.716
R8913 vss.n13502 vss.n2105 669.716
R8914 vss.n12060 vss.n12015 669.716
R8915 vss.n12023 vss.n12015 669.716
R8916 vss.n12053 vss.n12023 669.716
R8917 vss.n12053 vss.n12024 669.716
R8918 vss.n12047 vss.n12024 669.716
R8919 vss.n12047 vss.n12033 669.716
R8920 vss.n12041 vss.n12033 669.716
R8921 vss.n12041 vss.n2102 669.716
R8922 vss.n13720 vss.n13716 669.716
R8923 vss.n13720 vss.n8314 669.716
R8924 vss.n13724 vss.n8314 669.716
R8925 vss.n13724 vss.n8307 669.716
R8926 vss.n13740 vss.n8307 669.716
R8927 vss.n13740 vss.n8308 669.716
R8928 vss.n13734 vss.n8308 669.716
R8929 vss.n13734 vss.n2109 669.716
R8930 vss.n8486 vss.n8441 669.716
R8931 vss.n8449 vss.n8441 669.716
R8932 vss.n8479 vss.n8449 669.716
R8933 vss.n8479 vss.n8450 669.716
R8934 vss.n8473 vss.n8450 669.716
R8935 vss.n8473 vss.n8459 669.716
R8936 vss.n8467 vss.n8459 669.716
R8937 vss.n8467 vss.n2113 669.716
R8938 vss.n8563 vss.n8518 669.716
R8939 vss.n8526 vss.n8518 669.716
R8940 vss.n8556 vss.n8526 669.716
R8941 vss.n8556 vss.n8527 669.716
R8942 vss.n8550 vss.n8527 669.716
R8943 vss.n8550 vss.n8536 669.716
R8944 vss.n8544 vss.n8536 669.716
R8945 vss.n8544 vss.n2110 669.716
R8946 vss.n13008 vss.n13004 669.716
R8947 vss.n13008 vss.n9100 669.716
R8948 vss.n13012 vss.n9100 669.716
R8949 vss.n13012 vss.n9093 669.716
R8950 vss.n13028 vss.n9093 669.716
R8951 vss.n13028 vss.n9094 669.716
R8952 vss.n13022 vss.n9094 669.716
R8953 vss.n13022 vss.n2117 669.716
R8954 vss.n8973 vss.n8900 669.716
R8955 vss.n8973 vss.n8964 669.716
R8956 vss.n8977 vss.n8964 669.716
R8957 vss.n8977 vss.n8957 669.716
R8958 vss.n8993 vss.n8957 669.716
R8959 vss.n8993 vss.n8958 669.716
R8960 vss.n8987 vss.n8958 669.716
R8961 vss.n8987 vss.n2121 669.716
R8962 vss.n9158 vss.n9113 669.716
R8963 vss.n9121 vss.n9113 669.716
R8964 vss.n9151 vss.n9121 669.716
R8965 vss.n9151 vss.n9122 669.716
R8966 vss.n9145 vss.n9122 669.716
R8967 vss.n9145 vss.n9131 669.716
R8968 vss.n9139 vss.n9131 669.716
R8969 vss.n9139 vss.n2118 669.716
R8970 vss.n12638 vss.n12544 669.716
R8971 vss.n12552 vss.n12544 669.716
R8972 vss.n12631 vss.n12552 669.716
R8973 vss.n12631 vss.n12553 669.716
R8974 vss.n12576 vss.n12553 669.716
R8975 vss.n12576 vss.n12562 669.716
R8976 vss.n12570 vss.n12562 669.716
R8977 vss.n12570 vss.n2125 669.716
R8978 vss.n13533 vss.n2103 669.716
R8979 vss.n13533 vss.n13524 669.716
R8980 vss.n13537 vss.n13524 669.716
R8981 vss.n13537 vss.n13517 669.716
R8982 vss.n13552 vss.n13517 669.716
R8983 vss.n13552 vss.n13518 669.716
R8984 vss.n8245 vss.n2111 669.716
R8985 vss.n8245 vss.n8237 669.716
R8986 vss.n8251 vss.n8237 669.716
R8987 vss.n8251 vss.n8231 669.716
R8988 vss.n13852 vss.n8231 669.716
R8989 vss.n13852 vss.n13851 669.716
R8990 vss.n9018 vss.n2119 669.716
R8991 vss.n9018 vss.n9009 669.716
R8992 vss.n9022 vss.n9009 669.716
R8993 vss.n9022 vss.n9002 669.716
R8994 vss.n9037 vss.n9002 669.716
R8995 vss.n9037 vss.n9003 669.716
R8996 vss.n12845 vss.n12841 669.716
R8997 vss.n12845 vss.n9404 669.716
R8998 vss.n12849 vss.n9404 669.716
R8999 vss.n12849 vss.n9397 669.716
R9000 vss.n12865 vss.n9397 669.716
R9001 vss.n12865 vss.n9398 669.716
R9002 vss.n12859 vss.n9398 669.716
R9003 vss.n12859 vss.n2126 669.716
R9004 vss.n12774 vss.n12728 669.716
R9005 vss.n12736 vss.n12728 669.716
R9006 vss.n12767 vss.n12736 669.716
R9007 vss.n12767 vss.n12737 669.716
R9008 vss.n12760 vss.n12737 669.716
R9009 vss.n12760 vss.n12746 669.716
R9010 vss.n12754 vss.n12746 669.716
R9011 vss.n12754 vss.n2122 669.716
R9012 vss.n13322 vss.n13318 669.716
R9013 vss.n13322 vss.n8422 669.716
R9014 vss.n13326 vss.n8422 669.716
R9015 vss.n13326 vss.n8415 669.716
R9016 vss.n13342 vss.n8415 669.716
R9017 vss.n13342 vss.n8416 669.716
R9018 vss.n13336 vss.n8416 669.716
R9019 vss.n13336 vss.n2114 669.716
R9020 vss.n13441 vss.n13437 669.716
R9021 vss.n13441 vss.n13364 669.716
R9022 vss.n13445 vss.n13364 669.716
R9023 vss.n13445 vss.n13357 669.716
R9024 vss.n13461 vss.n13357 669.716
R9025 vss.n13461 vss.n13358 669.716
R9026 vss.n13455 vss.n13358 669.716
R9027 vss.n13455 vss.n2106 669.716
R9028 vss.n11865 vss.n11847 669.716
R9029 vss.n11854 vss.n11847 669.716
R9030 vss.n11858 vss.n11854 669.716
R9031 vss.n11858 vss.n2040 669.716
R9032 vss.n14186 vss.n2040 669.716
R9033 vss.n14186 vss.n2041 669.716
R9034 vss.n14180 vss.n2041 669.716
R9035 vss.n14180 vss.n14179 669.716
R9036 vss.n1807 vss.n1775 669.716
R9037 vss.n1807 vss.n1776 669.716
R9038 vss.n1801 vss.n1776 669.716
R9039 vss.n1801 vss.n1787 669.716
R9040 vss.n1795 vss.n1787 669.716
R9041 vss.n1795 vss.n1192 669.716
R9042 vss.n2008 vss.n1185 669.716
R9043 vss.n2008 vss.n1999 669.716
R9044 vss.n2012 vss.n1999 669.716
R9045 vss.n2012 vss.n1992 669.716
R9046 vss.n2029 vss.n1992 669.716
R9047 vss.n2029 vss.n1993 669.716
R9048 vss.n2023 vss.n1993 669.716
R9049 vss.n2023 vss.n2020 669.716
R9050 vss.n1028 vss.n996 669.716
R9051 vss.n1028 vss.n997 669.716
R9052 vss.n1022 vss.n997 669.716
R9053 vss.n1022 vss.n1008 669.716
R9054 vss.n1016 vss.n1008 669.716
R9055 vss.n1016 vss.n413 669.716
R9056 vss.n1113 vss.n406 669.716
R9057 vss.n1113 vss.n1104 669.716
R9058 vss.n1117 vss.n1104 669.716
R9059 vss.n1117 vss.n1097 669.716
R9060 vss.n1134 vss.n1097 669.716
R9061 vss.n1134 vss.n1098 669.716
R9062 vss.n1128 vss.n1098 669.716
R9063 vss.n1128 vss.n1125 669.716
R9064 vss.n3966 vss.n3965 669.716
R9065 vss.n3965 vss.n3949 669.716
R9066 vss.n3957 vss.n3949 669.716
R9067 vss.n3957 vss.n34 669.716
R9068 vss.n15865 vss.n34 669.716
R9069 vss.n15865 vss.n35 669.716
R9070 vss.n15859 vss.n35 669.716
R9071 vss.n15859 vss.n15856 669.716
R9072 vss.n3897 vss.n3896 669.716
R9073 vss.n3896 vss.n3851 669.716
R9074 vss.n3890 vss.n3851 669.716
R9075 vss.n3890 vss.n3859 669.716
R9076 vss.n3884 vss.n3859 669.716
R9077 vss.n3884 vss.n3869 669.716
R9078 vss.n3878 vss.n3869 669.716
R9079 vss.n3878 vss.n3875 669.716
R9080 vss.n3778 vss.n3777 669.716
R9081 vss.n3777 vss.n3732 669.716
R9082 vss.n3771 vss.n3732 669.716
R9083 vss.n3771 vss.n3740 669.716
R9084 vss.n3765 vss.n3740 669.716
R9085 vss.n3765 vss.n3750 669.716
R9086 vss.n3759 vss.n3750 669.716
R9087 vss.n3759 vss.n3756 669.716
R9088 vss.n3659 vss.n3658 669.716
R9089 vss.n3658 vss.n3613 669.716
R9090 vss.n3652 vss.n3613 669.716
R9091 vss.n3652 vss.n3621 669.716
R9092 vss.n3646 vss.n3621 669.716
R9093 vss.n3646 vss.n3631 669.716
R9094 vss.n3640 vss.n3631 669.716
R9095 vss.n3640 vss.n3637 669.716
R9096 vss.n6309 vss.n6291 669.716
R9097 vss.n6302 vss.n6291 669.716
R9098 vss.n6302 vss.n6301 669.716
R9099 vss.n6301 vss.n249 669.716
R9100 vss.n15697 vss.n249 669.716
R9101 vss.n15697 vss.n250 669.716
R9102 vss.n15691 vss.n250 669.716
R9103 vss.n15691 vss.n15688 669.716
R9104 vss.n350 vss.n349 669.716
R9105 vss.n349 vss.n305 669.716
R9106 vss.n343 vss.n305 669.716
R9107 vss.n343 vss.n312 669.716
R9108 vss.n337 vss.n312 669.716
R9109 vss.n337 vss.n322 669.716
R9110 vss.n331 vss.n322 669.716
R9111 vss.n331 vss.n328 669.716
R9112 vss.n11492 vss.n8841 669.716
R9113 vss.n11492 vss.n11483 669.716
R9114 vss.n11496 vss.n11483 669.716
R9115 vss.n11496 vss.n11476 669.716
R9116 vss.n11511 vss.n11476 669.716
R9117 vss.n11511 vss.n11477 669.716
R9118 vss.n11087 vss.n8849 669.716
R9119 vss.n11087 vss.n11078 669.716
R9120 vss.n11091 vss.n11078 669.716
R9121 vss.n11091 vss.n11071 669.716
R9122 vss.n11106 vss.n11071 669.716
R9123 vss.n11106 vss.n11072 669.716
R9124 vss.n10190 vss.n8857 669.716
R9125 vss.n10190 vss.n10181 669.716
R9126 vss.n10194 vss.n10181 669.716
R9127 vss.n10194 vss.n10174 669.716
R9128 vss.n10209 vss.n10174 669.716
R9129 vss.n10209 vss.n10175 669.716
R9130 vss.n10591 vss.n10587 669.716
R9131 vss.n10591 vss.n10581 669.716
R9132 vss.n10595 vss.n10581 669.716
R9133 vss.n10595 vss.n10574 669.716
R9134 vss.n10611 vss.n10574 669.716
R9135 vss.n10611 vss.n10575 669.716
R9136 vss.n10605 vss.n10575 669.716
R9137 vss.n10605 vss.n8860 669.716
R9138 vss.n10985 vss.n10981 669.716
R9139 vss.n10985 vss.n10975 669.716
R9140 vss.n10989 vss.n10975 669.716
R9141 vss.n10989 vss.n10968 669.716
R9142 vss.n11005 vss.n10968 669.716
R9143 vss.n11005 vss.n10969 669.716
R9144 vss.n10999 vss.n10969 669.716
R9145 vss.n10999 vss.n8852 669.716
R9146 vss.n10038 vss.n9992 669.716
R9147 vss.n10000 vss.n9992 669.716
R9148 vss.n10031 vss.n10000 669.716
R9149 vss.n10031 vss.n10001 669.716
R9150 vss.n10024 vss.n10001 669.716
R9151 vss.n10024 vss.n10010 669.716
R9152 vss.n10018 vss.n10010 669.716
R9153 vss.n10018 vss.n8844 669.716
R9154 vss.n11648 vss.n9948 669.716
R9155 vss.n9956 vss.n9948 669.716
R9156 vss.n11641 vss.n9956 669.716
R9157 vss.n11641 vss.n11640 669.716
R9158 vss.n11640 vss.n9960 669.716
R9159 vss.n11623 vss.n9960 669.716
R9160 vss.n11632 vss.n11623 669.716
R9161 vss.n11632 vss.n8836 669.716
R9162 vss.n14848 vss.n1159 641.981
R9163 vss.n15543 vss.n380 641.981
R9164 vss.n12183 vss.n12182 641.981
R9165 vss.n14832 vss.n14809 634.72
R9166 vss.n12182 vss.n12181 576.202
R9167 vss.n14848 vss.n14847 576.202
R9168 vss.n15543 vss.n15542 576.202
R9169 vss.n14826 vss.n1161 556.457
R9170 vss.n12239 vss.n9754 542.668
R9171 vss.n12357 vss.n9624 542.668
R9172 vss.n12476 vss.n9495 542.668
R9173 vss.n11733 vss.n11732 542.668
R9174 vss.n5556 vss.n5535 542.668
R9175 vss.n5744 vss.n3998 542.668
R9176 vss.n5984 vss.n3990 542.668
R9177 vss.n6369 vss.n6368 542.668
R9178 vss.n5534 vss.n4005 542.668
R9179 vss.n4211 vss.n3997 542.668
R9180 vss.n4479 vss.n3989 542.668
R9181 vss.n14911 vss.n14910 542.668
R9182 vss.n3079 vss.n3058 542.668
R9183 vss.n4670 vss.n3132 542.668
R9184 vss.n2674 vss.n2673 542.668
R9185 vss.n2924 vss.n2923 542.668
R9186 vss.n7985 vss.n7984 542.668
R9187 vss.n7221 vss.n3135 542.668
R9188 vss.n14216 vss.n14215 542.668
R9189 vss.n13956 vss.n8174 542.668
R9190 vss.n2246 vss.n2225 542.668
R9191 vss.n13591 vss.n13589 542.668
R9192 vss.n13780 vss.n13778 542.668
R9193 vss.n13068 vss.n13066 542.668
R9194 vss.n14074 vss.n2178 542.668
R9195 vss.n14446 vss.n14400 542.668
R9196 vss.n15141 vss.n15095 542.668
R9197 vss.n3591 vss.n3590 542.668
R9198 vss.n11549 vss.n11547 542.668
R9199 vss.n11238 vss.n11236 542.668
R9200 vss.n10899 vss.n10897 542.668
R9201 vss.n10505 vss.n10503 542.668
R9202 vss.n11832 vss.n11808 530.668
R9203 vss.n12184 vss.n11808 530.668
R9204 vss.n14271 vss.n14250 530.668
R9205 vss.n14250 vss.n1184 530.668
R9206 vss.n14312 vss.n14288 530.668
R9207 vss.n14320 vss.n14288 530.668
R9208 vss.n14966 vss.n14945 530.668
R9209 vss.n14945 vss.n405 530.668
R9210 vss.n15007 vss.n14983 530.668
R9211 vss.n15015 vss.n14983 530.668
R9212 vss.n15609 vss.n15588 530.668
R9213 vss.n15588 vss.n302 530.668
R9214 vss.n15648 vss.n353 530.668
R9215 vss.n15656 vss.n353 530.668
R9216 vss.n10361 vss.n10343 501.3
R9217 vss.n10350 vss.n10343 501.3
R9218 vss.n10354 vss.n10350 501.3
R9219 vss.n10354 vss.n8874 501.3
R9220 vss.n13192 vss.n8874 501.3
R9221 vss.n13192 vss.n13191 501.3
R9222 vss.n13191 vss.n8866 501.3
R9223 vss.n13199 vss.n8866 501.3
R9224 vss.n3295 vss.n436 501.3
R9225 vss.n3295 vss.n3286 501.3
R9226 vss.n3299 vss.n3286 501.3
R9227 vss.n3299 vss.n3279 501.3
R9228 vss.n6735 vss.n3279 501.3
R9229 vss.n6735 vss.n3280 501.3
R9230 vss.n6729 vss.n3280 501.3
R9231 vss.n6729 vss.n6726 501.3
R9232 vss.n6766 vss.n1215 501.3
R9233 vss.n6766 vss.n6757 501.3
R9234 vss.n6770 vss.n6757 501.3
R9235 vss.n6770 vss.n6750 501.3
R9236 vss.n6786 vss.n6750 501.3
R9237 vss.n6786 vss.n6751 501.3
R9238 vss.n6780 vss.n6751 501.3
R9239 vss.n6780 vss.n3168 501.3
R9240 vss.n9301 vss.n9283 501.3
R9241 vss.n9290 vss.n9283 501.3
R9242 vss.n9294 vss.n9290 501.3
R9243 vss.n9294 vss.n2136 501.3
R9244 vss.n14096 vss.n2136 501.3
R9245 vss.n14096 vss.n2137 501.3
R9246 vss.n2137 vss.n2128 501.3
R9247 vss.n14103 vss.n2128 501.3
R9248 vss.n9754 vss.n9744 498.046
R9249 vss.n9624 vss.n9614 498.046
R9250 vss.n9495 vss.n9485 498.046
R9251 vss.n11732 vss.n9873 498.046
R9252 vss.n5556 vss.n5553 498.046
R9253 vss.n5744 vss.n5741 498.046
R9254 vss.n5984 vss.n5981 498.046
R9255 vss.n6368 vss.n6335 498.046
R9256 vss.n5524 vss.n4005 498.046
R9257 vss.n4211 vss.n4210 498.046
R9258 vss.n4479 vss.n4453 498.046
R9259 vss.n14910 vss.n14900 498.046
R9260 vss.n15102 vss.n15095 498.046
R9261 vss.n3079 vss.n3076 498.046
R9262 vss.n4670 vss.n4667 498.046
R9263 vss.n2673 vss.n2664 498.046
R9264 vss.n2923 vss.n2890 498.046
R9265 vss.n7984 vss.n2460 498.046
R9266 vss.n7211 vss.n3135 498.046
R9267 vss.n14215 vss.n14205 498.046
R9268 vss.n14407 vss.n14400 498.046
R9269 vss.n8174 vss.n8164 498.046
R9270 vss.n2246 vss.n2243 498.046
R9271 vss.n13589 vss.n13562 498.046
R9272 vss.n13778 vss.n13752 498.046
R9273 vss.n13066 vss.n13040 498.046
R9274 vss.n2178 vss.n2152 498.046
R9275 vss.n3590 vss.n3581 498.046
R9276 vss.n11547 vss.n11521 498.046
R9277 vss.n11236 vss.n11210 498.046
R9278 vss.n10897 vss.n10871 498.046
R9279 vss.n10503 vss.n10477 498.046
R9280 vss.n15521 vss.n15513 497.128
R9281 vss.n12143 vss.n12133 497.128
R9282 vss.n9813 vss.n9807 482.334
R9283 vss.n9684 vss.n9678 482.334
R9284 vss.n9555 vss.n9549 482.334
R9285 vss.n5602 vss.n5600 482.334
R9286 vss.n5874 vss.n5725 482.334
R9287 vss.n6113 vss.n5965 482.334
R9288 vss.n3526 vss.n3523 482.334
R9289 vss.n4072 vss.n4044 482.334
R9290 vss.n4253 vss.n4225 482.334
R9291 vss.n7401 vss.n7395 482.334
R9292 vss.n7231 vss.n7225 482.334
R9293 vss.n2713 vss.n2685 482.334
R9294 vss.n3050 vss.n3047 482.334
R9295 vss.n7060 vss.n7059 482.334
R9296 vss.n13866 vss.n13860 482.334
R9297 vss.n8105 vss.n8099 482.334
R9298 vss.n13546 vss.n13518 482.334
R9299 vss.n13851 vss.n13848 482.334
R9300 vss.n9031 vss.n9003 482.334
R9301 vss.n1775 vss.n1769 482.334
R9302 vss.n996 vss.n990 482.334
R9303 vss.n11505 vss.n11477 482.334
R9304 vss.n11100 vss.n11072 482.334
R9305 vss.n10203 vss.n10175 482.334
R9306 vss.n12235 vss.n12234 475.476
R9307 vss.n12234 vss.n9853 475.476
R9308 vss.n12228 vss.n9853 475.476
R9309 vss.n12228 vss.n12197 475.476
R9310 vss.n12222 vss.n12197 475.476
R9311 vss.n12222 vss.n12207 475.476
R9312 vss.n9801 vss.n9755 475.476
R9313 vss.n9763 vss.n9755 475.476
R9314 vss.n9794 vss.n9763 475.476
R9315 vss.n9794 vss.n9764 475.476
R9316 vss.n9788 vss.n9764 475.476
R9317 vss.n9788 vss.n9773 475.476
R9318 vss.n12353 vss.n12352 475.476
R9319 vss.n12352 vss.n9725 475.476
R9320 vss.n12346 vss.n9725 475.476
R9321 vss.n12346 vss.n12315 475.476
R9322 vss.n12340 vss.n12315 475.476
R9323 vss.n12340 vss.n12325 475.476
R9324 vss.n9672 vss.n9625 475.476
R9325 vss.n9633 vss.n9625 475.476
R9326 vss.n9665 vss.n9633 475.476
R9327 vss.n9665 vss.n9634 475.476
R9328 vss.n9659 vss.n9634 475.476
R9329 vss.n9659 vss.n9643 475.476
R9330 vss.n12472 vss.n12471 475.476
R9331 vss.n12471 vss.n9595 475.476
R9332 vss.n12465 vss.n9595 475.476
R9333 vss.n12465 vss.n12434 475.476
R9334 vss.n12459 vss.n12434 475.476
R9335 vss.n12459 vss.n12444 475.476
R9336 vss.n9542 vss.n9496 475.476
R9337 vss.n9504 vss.n9496 475.476
R9338 vss.n9535 vss.n9504 475.476
R9339 vss.n9535 vss.n9505 475.476
R9340 vss.n9529 vss.n9505 475.476
R9341 vss.n9529 vss.n9514 475.476
R9342 vss.n9445 vss.n9441 475.476
R9343 vss.n9445 vss.n9435 475.476
R9344 vss.n9449 vss.n9435 475.476
R9345 vss.n9449 vss.n9428 475.476
R9346 vss.n9466 vss.n9428 475.476
R9347 vss.n9466 vss.n9429 475.476
R9348 vss.n6332 vss.n3536 475.476
R9349 vss.n3545 vss.n3536 475.476
R9350 vss.n6325 vss.n3545 475.476
R9351 vss.n6325 vss.n3546 475.476
R9352 vss.n6319 vss.n3546 475.476
R9353 vss.n6319 vss.n3555 475.476
R9354 vss.n5722 vss.n5536 475.476
R9355 vss.n5684 vss.n5536 475.476
R9356 vss.n5715 vss.n5684 475.476
R9357 vss.n5715 vss.n5685 475.476
R9358 vss.n5709 vss.n5685 475.476
R9359 vss.n5709 vss.n5694 475.476
R9360 vss.n5960 vss.n5913 475.476
R9361 vss.n5922 vss.n5913 475.476
R9362 vss.n5953 vss.n5922 475.476
R9363 vss.n5953 vss.n5923 475.476
R9364 vss.n5947 vss.n5923 475.476
R9365 vss.n5947 vss.n5932 475.476
R9366 vss.n5797 vss.n3999 475.476
R9367 vss.n5797 vss.n5788 475.476
R9368 vss.n5801 vss.n5788 475.476
R9369 vss.n5801 vss.n5781 475.476
R9370 vss.n5818 vss.n5781 475.476
R9371 vss.n5818 vss.n5782 475.476
R9372 vss.n6199 vss.n6152 475.476
R9373 vss.n6161 vss.n6152 475.476
R9374 vss.n6192 vss.n6161 475.476
R9375 vss.n6192 vss.n6162 475.476
R9376 vss.n6186 vss.n6162 475.476
R9377 vss.n6186 vss.n6171 475.476
R9378 vss.n6037 vss.n3991 475.476
R9379 vss.n6037 vss.n6028 475.476
R9380 vss.n6041 vss.n6028 475.476
R9381 vss.n6041 vss.n6021 475.476
R9382 vss.n6058 vss.n6021 475.476
R9383 vss.n6058 vss.n6022 475.476
R9384 vss.n6696 vss.n3335 475.476
R9385 vss.n6696 vss.n6665 475.476
R9386 vss.n6690 vss.n6665 475.476
R9387 vss.n6690 vss.n6689 475.476
R9388 vss.n6689 vss.n6677 475.476
R9389 vss.n6677 vss.n378 475.476
R9390 vss.n3470 vss.n3454 475.476
R9391 vss.n3470 vss.n3449 475.476
R9392 vss.n3479 vss.n3449 475.476
R9393 vss.n3479 vss.n3478 475.476
R9394 vss.n3478 vss.n3441 475.476
R9395 vss.n3486 vss.n3441 475.476
R9396 vss.n5284 vss.n5270 475.476
R9397 vss.n5284 vss.n5263 475.476
R9398 vss.n5301 vss.n5263 475.476
R9399 vss.n5301 vss.n5264 475.476
R9400 vss.n5295 vss.n5264 475.476
R9401 vss.n5295 vss.n5294 475.476
R9402 vss.n5499 vss.n5485 475.476
R9403 vss.n5499 vss.n5478 475.476
R9404 vss.n5515 vss.n5478 475.476
R9405 vss.n5515 vss.n5479 475.476
R9406 vss.n5509 vss.n5479 475.476
R9407 vss.n5509 vss.n4004 475.476
R9408 vss.n5073 vss.n5059 475.476
R9409 vss.n5073 vss.n5052 475.476
R9410 vss.n5089 vss.n5052 475.476
R9411 vss.n5089 vss.n5053 475.476
R9412 vss.n5083 vss.n5053 475.476
R9413 vss.n5083 vss.n4001 475.476
R9414 vss.n5025 vss.n5011 475.476
R9415 vss.n5025 vss.n5004 475.476
R9416 vss.n5041 vss.n5004 475.476
R9417 vss.n5041 vss.n5005 475.476
R9418 vss.n5035 vss.n5005 475.476
R9419 vss.n5035 vss.n3996 475.476
R9420 vss.n4520 vss.n4506 475.476
R9421 vss.n4520 vss.n4499 475.476
R9422 vss.n4536 vss.n4499 475.476
R9423 vss.n4536 vss.n4500 475.476
R9424 vss.n4530 vss.n4500 475.476
R9425 vss.n4530 vss.n3993 475.476
R9426 vss.n7487 vss.n7486 475.476
R9427 vss.n7486 vss.n7441 475.476
R9428 vss.n7480 vss.n7441 475.476
R9429 vss.n7480 vss.n7449 475.476
R9430 vss.n7474 vss.n7449 475.476
R9431 vss.n7474 vss.n7459 475.476
R9432 vss.n7392 vss.n3059 475.476
R9433 vss.n7354 vss.n3059 475.476
R9434 vss.n7385 vss.n7354 475.476
R9435 vss.n7385 vss.n7355 475.476
R9436 vss.n7379 vss.n7355 475.476
R9437 vss.n7379 vss.n7364 475.476
R9438 vss.n7275 vss.n7271 475.476
R9439 vss.n7275 vss.n3122 475.476
R9440 vss.n7279 vss.n3122 475.476
R9441 vss.n7279 vss.n3115 475.476
R9442 vss.n7296 vss.n3115 475.476
R9443 vss.n7296 vss.n3116 475.476
R9444 vss.n4628 vss.n3133 475.476
R9445 vss.n4628 vss.n4619 475.476
R9446 vss.n4632 vss.n4619 475.476
R9447 vss.n4632 vss.n4612 475.476
R9448 vss.n4649 vss.n4612 475.476
R9449 vss.n4649 vss.n4613 475.476
R9450 vss.n4581 vss.n4577 475.476
R9451 vss.n4581 vss.n4571 475.476
R9452 vss.n4585 vss.n4571 475.476
R9453 vss.n4585 vss.n4564 475.476
R9454 vss.n4602 vss.n4564 475.476
R9455 vss.n4602 vss.n4565 475.476
R9456 vss.n7936 vss.n7926 475.476
R9457 vss.n7936 vss.n1146 475.476
R9458 vss.n14878 vss.n1146 475.476
R9459 vss.n14878 vss.n1147 475.476
R9460 vss.n14872 vss.n1147 475.476
R9461 vss.n14872 vss.n14871 475.476
R9462 vss.n7891 vss.n7877 475.476
R9463 vss.n7891 vss.n7870 475.476
R9464 vss.n7908 vss.n7870 475.476
R9465 vss.n7908 vss.n7871 475.476
R9466 vss.n7902 vss.n7871 475.476
R9467 vss.n7902 vss.n7901 475.476
R9468 vss.n7745 vss.n7731 475.476
R9469 vss.n7745 vss.n7724 475.476
R9470 vss.n7761 vss.n7724 475.476
R9471 vss.n7761 vss.n7725 475.476
R9472 vss.n7755 vss.n7725 475.476
R9473 vss.n7755 vss.n986 475.476
R9474 vss.n7696 vss.n7682 475.476
R9475 vss.n7696 vss.n7675 475.476
R9476 vss.n7713 vss.n7675 475.476
R9477 vss.n7713 vss.n7676 475.476
R9478 vss.n7707 vss.n7676 475.476
R9479 vss.n7707 vss.n7706 475.476
R9480 vss.n3002 vss.n2988 475.476
R9481 vss.n3002 vss.n2981 475.476
R9482 vss.n7497 vss.n2981 475.476
R9483 vss.n7497 vss.n2982 475.476
R9484 vss.n7491 vss.n2982 475.476
R9485 vss.n7491 vss.n7490 475.476
R9486 vss.n7116 vss.n7077 475.476
R9487 vss.n7116 vss.n7084 475.476
R9488 vss.n7110 vss.n7084 475.476
R9489 vss.n7110 vss.n7109 475.476
R9490 vss.n7109 vss.n7096 475.476
R9491 vss.n7102 vss.n7096 475.476
R9492 vss.n6912 vss.n6825 475.476
R9493 vss.n6912 vss.n6881 475.476
R9494 vss.n6906 vss.n6881 475.476
R9495 vss.n6906 vss.n6905 475.476
R9496 vss.n6905 vss.n6893 475.476
R9497 vss.n6893 vss.n3130 475.476
R9498 vss.n13952 vss.n13951 475.476
R9499 vss.n13951 vss.n13906 475.476
R9500 vss.n13945 vss.n13906 475.476
R9501 vss.n13945 vss.n13914 475.476
R9502 vss.n13939 vss.n13914 475.476
R9503 vss.n13939 vss.n13924 475.476
R9504 vss.n8221 vss.n8175 475.476
R9505 vss.n8183 vss.n8175 475.476
R9506 vss.n8214 vss.n8183 475.476
R9507 vss.n8214 vss.n8184 475.476
R9508 vss.n8208 vss.n8184 475.476
R9509 vss.n8208 vss.n8193 475.476
R9510 vss.n14069 vss.n14068 475.476
R9511 vss.n14068 vss.n8145 475.476
R9512 vss.n14062 vss.n8145 475.476
R9513 vss.n14062 vss.n14031 475.476
R9514 vss.n14056 vss.n14031 475.476
R9515 vss.n14056 vss.n14041 475.476
R9516 vss.n8093 vss.n2226 475.476
R9517 vss.n8055 vss.n2226 475.476
R9518 vss.n8086 vss.n8055 475.476
R9519 vss.n8086 vss.n8056 475.476
R9520 vss.n8080 vss.n8056 475.476
R9521 vss.n8080 vss.n8065 475.476
R9522 vss.n2299 vss.n2295 475.476
R9523 vss.n2299 vss.n2289 475.476
R9524 vss.n2303 vss.n2289 475.476
R9525 vss.n2303 vss.n2282 475.476
R9526 vss.n2320 vss.n2282 475.476
R9527 vss.n2320 vss.n2283 475.476
R9528 vss.n2084 vss.n2068 475.476
R9529 vss.n2084 vss.n2062 475.476
R9530 vss.n14148 vss.n2062 475.476
R9531 vss.n14148 vss.n14147 475.476
R9532 vss.n14147 vss.n2054 475.476
R9533 vss.n14155 vss.n2054 475.476
R9534 vss.n13631 vss.n13617 475.476
R9535 vss.n13631 vss.n13610 475.476
R9536 vss.n13648 vss.n13610 475.476
R9537 vss.n13648 vss.n13611 475.476
R9538 vss.n13642 vss.n13611 475.476
R9539 vss.n13642 vss.n13641 475.476
R9540 vss.n8281 vss.n8267 475.476
R9541 vss.n8281 vss.n8260 475.476
R9542 vss.n8297 vss.n8260 475.476
R9543 vss.n8297 vss.n8261 475.476
R9544 vss.n8291 vss.n8261 475.476
R9545 vss.n8291 vss.n1765 475.476
R9546 vss.n13820 vss.n13806 475.476
R9547 vss.n13820 vss.n13799 475.476
R9548 vss.n13837 vss.n13799 475.476
R9549 vss.n13837 vss.n13800 475.476
R9550 vss.n13831 vss.n13800 475.476
R9551 vss.n13831 vss.n13830 475.476
R9552 vss.n9067 vss.n9053 475.476
R9553 vss.n9067 vss.n9046 475.476
R9554 vss.n9083 vss.n9046 475.476
R9555 vss.n9083 vss.n9047 475.476
R9556 vss.n9077 vss.n9047 475.476
R9557 vss.n9077 vss.n8223 475.476
R9558 vss.n13108 vss.n13094 475.476
R9559 vss.n13108 vss.n13087 475.476
R9560 vss.n13125 vss.n13087 475.476
R9561 vss.n13125 vss.n13088 475.476
R9562 vss.n13119 vss.n13088 475.476
R9563 vss.n13119 vss.n13118 475.476
R9564 vss.n12605 vss.n12591 475.476
R9565 vss.n12605 vss.n12584 475.476
R9566 vss.n12621 vss.n12584 475.476
R9567 vss.n12621 vss.n12585 475.476
R9568 vss.n12615 vss.n12585 475.476
R9569 vss.n12615 vss.n8095 475.476
R9570 vss.n14452 vss.n14448 475.476
R9571 vss.n14452 vss.n1757 475.476
R9572 vss.n14456 vss.n1757 475.476
R9573 vss.n14456 vss.n1750 475.476
R9574 vss.n14473 vss.n1750 475.476
R9575 vss.n14473 vss.n1751 475.476
R9576 vss.n14397 vss.n14396 475.476
R9577 vss.n14396 vss.n1815 475.476
R9578 vss.n14390 vss.n1815 475.476
R9579 vss.n14390 vss.n14359 475.476
R9580 vss.n14384 vss.n14359 475.476
R9581 vss.n14384 vss.n14369 475.476
R9582 vss.n15147 vss.n15143 475.476
R9583 vss.n15147 vss.n978 475.476
R9584 vss.n15151 vss.n978 475.476
R9585 vss.n15151 vss.n971 475.476
R9586 vss.n15168 vss.n971 475.476
R9587 vss.n15168 vss.n972 475.476
R9588 vss.n15092 vss.n15091 475.476
R9589 vss.n15091 vss.n1036 475.476
R9590 vss.n15085 vss.n1036 475.476
R9591 vss.n15085 vss.n15054 475.476
R9592 vss.n15079 vss.n15054 475.476
R9593 vss.n15079 vss.n15064 475.476
R9594 vss.n6251 vss.n6250 475.476
R9595 vss.n6250 vss.n6205 475.476
R9596 vss.n6244 vss.n6205 475.476
R9597 vss.n6244 vss.n6213 475.476
R9598 vss.n6238 vss.n6213 475.476
R9599 vss.n6238 vss.n6223 475.476
R9600 vss.n9908 vss.n9893 475.476
R9601 vss.n9908 vss.n9887 475.476
R9602 vss.n11718 vss.n9887 475.476
R9603 vss.n11718 vss.n11717 475.476
R9604 vss.n11717 vss.n9879 475.476
R9605 vss.n11725 vss.n9879 475.476
R9606 vss.n11589 vss.n11575 475.476
R9607 vss.n11589 vss.n11568 475.476
R9608 vss.n11606 vss.n11568 475.476
R9609 vss.n11606 vss.n11569 475.476
R9610 vss.n11600 vss.n11569 475.476
R9611 vss.n11600 vss.n11599 475.476
R9612 vss.n11136 vss.n11122 475.476
R9613 vss.n11136 vss.n11115 475.476
R9614 vss.n11152 vss.n11115 475.476
R9615 vss.n11152 vss.n11116 475.476
R9616 vss.n11146 vss.n11116 475.476
R9617 vss.n11146 vss.n9803 475.476
R9618 vss.n11278 vss.n11264 475.476
R9619 vss.n11278 vss.n11257 475.476
R9620 vss.n11295 vss.n11257 475.476
R9621 vss.n11295 vss.n11258 475.476
R9622 vss.n11289 vss.n11258 475.476
R9623 vss.n11289 vss.n11288 475.476
R9624 vss.n10939 vss.n10925 475.476
R9625 vss.n10939 vss.n10918 475.476
R9626 vss.n10955 vss.n10918 475.476
R9627 vss.n10955 vss.n10919 475.476
R9628 vss.n10949 vss.n10919 475.476
R9629 vss.n10949 vss.n9674 475.476
R9630 vss.n10843 vss.n10829 475.476
R9631 vss.n10843 vss.n10822 475.476
R9632 vss.n10860 vss.n10822 475.476
R9633 vss.n10860 vss.n10823 475.476
R9634 vss.n10854 vss.n10823 475.476
R9635 vss.n10854 vss.n10853 475.476
R9636 vss.n10545 vss.n10531 475.476
R9637 vss.n10545 vss.n10524 475.476
R9638 vss.n10561 vss.n10524 475.476
R9639 vss.n10561 vss.n10525 475.476
R9640 vss.n10555 vss.n10525 475.476
R9641 vss.n10555 vss.n9545 475.476
R9642 vss.n15521 vss.n382 460.522
R9643 vss.n14839 vss.n14809 460.522
R9644 vss.n14839 vss.n14810 460.522
R9645 vss.n14810 vss.n1162 460.522
R9646 vss.n14846 vss.n1162 460.522
R9647 vss.n15534 vss.n15505 460.522
R9648 vss.n15505 vss.n383 460.522
R9649 vss.n15541 vss.n383 460.522
R9650 vss.n12167 vss.n12153 460.522
R9651 vss.n12161 vss.n12153 460.522
R9652 vss.n12161 vss.n12132 460.522
R9653 vss.n12180 vss.n12133 460.522
R9654 vss.n12908 vss.n12907 376
R9655 vss.n12911 vss.n12910 376
R9656 vss.n12914 vss.n12913 376
R9657 vss.n13260 vss.n8637 376
R9658 vss.n13258 vss.n13257 376
R9659 vss.n13255 vss.n13254 376
R9660 vss.n13252 vss.n13251 376
R9661 vss.n14107 vss.n14106 376
R9662 vss.n14110 vss.n14109 376
R9663 vss.n14113 vss.n14112 376
R9664 vss.n14116 vss.n14115 376
R9665 vss.n14119 vss.n14118 376
R9666 vss.n14122 vss.n14121 376
R9667 vss.n14124 vss.n2053 376
R9668 vss.n14769 vss.n14768 376
R9669 vss.n14772 vss.n14771 376
R9670 vss.n14775 vss.n14774 376
R9671 vss.n14778 vss.n14777 376
R9672 vss.n14781 vss.n14780 376
R9673 vss.n14784 vss.n14783 376
R9674 vss.n14787 vss.n14786 376
R9675 vss.n7175 vss.n7174 376
R9676 vss.n7172 vss.n7171 376
R9677 vss.n7958 vss.n2470 376
R9678 vss.n7956 vss.n7955 376
R9679 vss.n7953 vss.n7952 376
R9680 vss.n7950 vss.n7949 376
R9681 vss.n7947 vss.n7946 376
R9682 vss.n15464 vss.n15463 376
R9683 vss.n15467 vss.n15466 376
R9684 vss.n15470 vss.n15469 376
R9685 vss.n15473 vss.n15472 376
R9686 vss.n15476 vss.n15475 376
R9687 vss.n15479 vss.n15478 376
R9688 vss.n15482 vss.n15481 376
R9689 vss.n6723 vss.n6722 376
R9690 vss.n6720 vss.n6719 376
R9691 vss.n6717 vss.n6716 376
R9692 vss.n6714 vss.n6713 376
R9693 vss.n6711 vss.n6710 376
R9694 vss.n6708 vss.n6707 376
R9695 vss.n6705 vss.n6704 376
R9696 vss.n6274 vss.n6273 376
R9697 vss.n6277 vss.n6276 376
R9698 vss.n6280 vss.n6279 376
R9699 vss.n6283 vss.n6282 376
R9700 vss.n6286 vss.n6285 376
R9701 vss.n6289 vss.n6288 376
R9702 vss.n6311 vss.n6310 376
R9703 vss.n13203 vss.n13202 376
R9704 vss.n13206 vss.n13205 376
R9705 vss.n13209 vss.n13208 376
R9706 vss.n13212 vss.n13211 376
R9707 vss.n13215 vss.n13214 376
R9708 vss.n13218 vss.n13217 376
R9709 vss.n13221 vss.n13220 376
R9710 vss.n6270 vss.n6253 342.738
R9711 vss.n6263 vss.n6253 342.738
R9712 vss.n6263 vss.n15 342.738
R9713 vss.n15889 vss.n16 342.738
R9714 vss.n15881 vss.n16 342.738
R9715 vss.n15881 vss.n15880 342.738
R9716 vss.n15880 vss.n25 342.738
R9717 vss.n15854 vss.n44 342.738
R9718 vss.n52 vss.n44 342.738
R9719 vss.n15847 vss.n52 342.738
R9720 vss.n15840 vss.n62 342.738
R9721 vss.n15840 vss.n63 342.738
R9722 vss.n15832 vss.n63 342.738
R9723 vss.n15832 vss.n15829 342.738
R9724 vss.n15827 vss.n68 342.738
R9725 vss.n76 vss.n68 342.738
R9726 vss.n15820 vss.n76 342.738
R9727 vss.n114 vss.n111 342.738
R9728 vss.n115 vss.n114 342.738
R9729 vss.n115 vss.n102 342.738
R9730 vss.n122 vss.n102 342.738
R9731 vss.n15798 vss.n123 342.738
R9732 vss.n131 vss.n123 342.738
R9733 vss.n15791 vss.n131 342.738
R9734 vss.n15784 vss.n141 342.738
R9735 vss.n15784 vss.n142 342.738
R9736 vss.n15776 vss.n142 342.738
R9737 vss.n15776 vss.n15773 342.738
R9738 vss.n15771 vss.n147 342.738
R9739 vss.n155 vss.n147 342.738
R9740 vss.n15764 vss.n155 342.738
R9741 vss.n192 vss.n189 342.738
R9742 vss.n193 vss.n192 342.738
R9743 vss.n193 vss.n180 342.738
R9744 vss.n200 vss.n180 342.738
R9745 vss.n15742 vss.n201 342.738
R9746 vss.n209 vss.n201 342.738
R9747 vss.n15735 vss.n209 342.738
R9748 vss.n15728 vss.n219 342.738
R9749 vss.n15728 vss.n220 342.738
R9750 vss.n15720 vss.n220 342.738
R9751 vss.n15720 vss.n15717 342.738
R9752 vss.n15715 vss.n225 342.738
R9753 vss.n233 vss.n225 342.738
R9754 vss.n15708 vss.n233 342.738
R9755 vss.n271 vss.n268 342.738
R9756 vss.n272 vss.n271 342.738
R9757 vss.n272 vss.n259 342.738
R9758 vss.n279 vss.n259 342.738
R9759 vss.n15686 vss.n280 342.738
R9760 vss.n15679 vss.n280 342.738
R9761 vss.n15679 vss.n15678 342.738
R9762 vss.n15671 vss.n294 342.738
R9763 vss.n15671 vss.n295 342.738
R9764 vss.n15663 vss.n295 342.738
R9765 vss.n15663 vss.n15660 342.738
R9766 vss.n10365 vss.n10362 342.738
R9767 vss.n10365 vss.n10335 342.738
R9768 vss.n10372 vss.n10335 342.738
R9769 vss.n10372 vss.n10337 342.738
R9770 vss.n10379 vss.n10328 342.738
R9771 vss.n10328 vss.n10273 342.738
R9772 vss.n10386 vss.n10273 342.738
R9773 vss.n10394 vss.n10387 342.738
R9774 vss.n10387 vss.n10247 342.738
R9775 vss.n10621 vss.n10247 342.738
R9776 vss.n10621 vss.n10249 342.738
R9777 vss.n10628 vss.n10240 342.738
R9778 vss.n10240 vss.n10231 342.738
R9779 vss.n10635 vss.n10231 342.738
R9780 vss.n10784 vss.n10636 342.738
R9781 vss.n10644 vss.n10636 342.738
R9782 vss.n10777 vss.n10644 342.738
R9783 vss.n10777 vss.n10645 342.738
R9784 vss.n10771 vss.n10701 342.738
R9785 vss.n10709 vss.n10701 342.738
R9786 vss.n10764 vss.n10709 342.738
R9787 vss.n10762 vss.n10755 342.738
R9788 vss.n10755 vss.n10160 342.738
R9789 vss.n11014 vss.n10160 342.738
R9790 vss.n11014 vss.n10162 342.738
R9791 vss.n11021 vss.n10153 342.738
R9792 vss.n10153 vss.n10144 342.738
R9793 vss.n11028 vss.n10144 342.738
R9794 vss.n11036 vss.n11029 342.738
R9795 vss.n11029 vss.n10072 342.738
R9796 vss.n11308 vss.n10072 342.738
R9797 vss.n11308 vss.n10074 342.738
R9798 vss.n11315 vss.n10065 342.738
R9799 vss.n10065 vss.n10056 342.738
R9800 vss.n11322 vss.n10056 342.738
R9801 vss.n11327 vss.n11324 342.738
R9802 vss.n11327 vss.n10047 342.738
R9803 vss.n11334 vss.n10047 342.738
R9804 vss.n11334 vss.n10049 342.738
R9805 vss.n11341 vss.n10040 342.738
R9806 vss.n10040 vss.n9984 342.738
R9807 vss.n11348 vss.n9984 342.738
R9808 vss.n11441 vss.n11349 342.738
R9809 vss.n11356 vss.n11349 342.738
R9810 vss.n11434 vss.n11356 342.738
R9811 vss.n11434 vss.n11357 342.738
R9812 vss.n11428 vss.n11413 342.738
R9813 vss.n11420 vss.n11413 342.738
R9814 vss.n11420 vss.n9929 342.738
R9815 vss.n11678 vss.n9930 342.738
R9816 vss.n9938 vss.n9930 342.738
R9817 vss.n11671 vss.n9938 342.738
R9818 vss.n11671 vss.n9939 342.738
R9819 vss.n11665 vss.n11650 342.738
R9820 vss.n11657 vss.n11650 342.738
R9821 vss.n11657 vss.n8834 342.738
R9822 vss.n12207 vss.n8805 342.442
R9823 vss.n9773 vss.n8736 342.442
R9824 vss.n12325 vss.n8686 342.442
R9825 vss.n9650 vss.n9643 342.442
R9826 vss.n12444 vss.n9206 342.442
R9827 vss.n9514 vss.n9275 342.442
R9828 vss.n9429 vss.n9279 342.442
R9829 vss.n6312 vss.n3555 342.442
R9830 vss.n5694 vss.n3661 342.442
R9831 vss.n5932 vss.n3729 342.442
R9832 vss.n5782 vss.n3780 342.442
R9833 vss.n6171 vss.n3848 342.442
R9834 vss.n6022 vss.n3899 342.442
R9835 vss.n6703 vss.n3335 342.442
R9836 vss.n3454 vss.n3331 342.442
R9837 vss.n5270 vss.n3327 342.442
R9838 vss.n5485 vss.n3323 342.442
R9839 vss.n5059 vss.n3319 342.442
R9840 vss.n5011 vss.n3315 342.442
R9841 vss.n4506 vss.n3311 342.442
R9842 vss.n7459 vss.n416 342.442
R9843 vss.n7364 vss.n420 342.442
R9844 vss.n3116 vss.n424 342.442
R9845 vss.n4613 vss.n428 342.442
R9846 vss.n4565 vss.n432 342.442
R9847 vss.n7945 vss.n7926 342.442
R9848 vss.n7877 vss.n2482 342.442
R9849 vss.n7731 vss.n2478 342.442
R9850 vss.n7682 vss.n2474 342.442
R9851 vss.n2988 vss.n2469 342.442
R9852 vss.n7123 vss.n7077 342.442
R9853 vss.n6919 vss.n6825 342.442
R9854 vss.n13924 vss.n1195 342.442
R9855 vss.n8193 vss.n1199 342.442
R9856 vss.n14041 vss.n1203 342.442
R9857 vss.n8065 vss.n1207 342.442
R9858 vss.n2283 vss.n1211 342.442
R9859 vss.n2074 vss.n2068 342.442
R9860 vss.n13617 vss.n2104 342.442
R9861 vss.n8267 vss.n2108 342.442
R9862 vss.n13806 vss.n2112 342.442
R9863 vss.n9053 vss.n2116 342.442
R9864 vss.n13094 vss.n2120 342.442
R9865 vss.n12591 vss.n2124 342.442
R9866 vss.n1751 vss.n1191 342.442
R9867 vss.n14369 vss.n1187 342.442
R9868 vss.n972 vss.n412 342.442
R9869 vss.n15064 vss.n408 342.442
R9870 vss.n6223 vss.n3967 342.442
R9871 vss.n9893 vss.n8838 342.442
R9872 vss.n11575 vss.n8842 342.442
R9873 vss.n11122 vss.n8846 342.442
R9874 vss.n11264 vss.n8850 342.442
R9875 vss.n10925 vss.n8854 342.442
R9876 vss.n10829 vss.n8858 342.442
R9877 vss.n10531 vss.n8862 342.442
R9878 vss.n4422 vss.n3307 315.219
R9879 vss.n4422 vss.n4413 315.219
R9880 vss.n4426 vss.n4413 315.219
R9881 vss.n4426 vss.n4406 315.219
R9882 vss.n4442 vss.n4406 315.219
R9883 vss.n4442 vss.n4407 315.219
R9884 vss.n4436 vss.n4407 315.219
R9885 vss.n4436 vss.n3988 315.219
R9886 vss.n7182 vss.n7178 315.219
R9887 vss.n7182 vss.n3162 315.219
R9888 vss.n7186 vss.n3162 315.219
R9889 vss.n7186 vss.n3155 315.219
R9890 vss.n7202 vss.n3155 315.219
R9891 vss.n7202 vss.n3156 315.219
R9892 vss.n7196 vss.n3156 315.219
R9893 vss.n7196 vss.n3134 315.219
R9894 vss.n2203 vss.n2127 315.219
R9895 vss.n2203 vss.n2194 315.219
R9896 vss.n2209 vss.n2194 315.219
R9897 vss.n2209 vss.n2188 315.219
R9898 vss.n2217 vss.n2188 315.219
R9899 vss.n2217 vss.n2189 315.219
R9900 vss.n2189 vss.n2180 315.219
R9901 vss.n2224 vss.n2180 315.219
R9902 vss.n10445 vss.n8865 315.219
R9903 vss.n10445 vss.n10436 315.219
R9904 vss.n10449 vss.n10436 315.219
R9905 vss.n10449 vss.n10429 315.219
R9906 vss.n10466 vss.n10429 315.219
R9907 vss.n10466 vss.n10430 315.219
R9908 vss.n10460 vss.n10430 315.219
R9909 vss.n10460 vss.n10457 315.219
R9910 vss.n14847 vss.n14846 293.493
R9911 vss.n15667 vss.n292 263.154
R9912 vss.n15875 vss.n24 263.154
R9913 vss.n15724 vss.n216 263.154
R9914 vss.n15780 vss.n138 263.154
R9915 vss.n15836 vss.n59 263.154
R9916 vss.n6577 vss.n6567 263.154
R9917 vss.n6549 vss.n6548 263.154
R9918 vss.n6563 vss.n6496 263.154
R9919 vss.n5389 vss.n5380 263.154
R9920 vss.n5362 vss.n5361 263.154
R9921 vss.n5376 vss.n5309 263.154
R9922 vss.n638 vss.n636 263.154
R9923 vss.n624 vss.n623 263.154
R9924 vss.n15402 vss.n626 263.154
R9925 vss.n4914 vss.n4905 263.154
R9926 vss.n4887 vss.n4886 263.154
R9927 vss.n4901 vss.n4264 263.154
R9928 vss.n5177 vss.n5168 263.154
R9929 vss.n5150 vss.n5149 263.154
R9930 vss.n5164 vss.n5097 263.154
R9931 vss.n895 vss.n893 263.154
R9932 vss.n881 vss.n880 263.154
R9933 vss.n15252 vss.n883 263.154
R9934 vss.n6461 vss.n6452 263.154
R9935 vss.n6434 vss.n6433 263.154
R9936 vss.n6448 vss.n6381 263.154
R9937 vss.n4856 vss.n4749 263.154
R9938 vss.n4833 vss.n4832 263.154
R9939 vss.n4848 vss.n4750 263.154
R9940 vss.n6439 vss.n6411 263.154
R9941 vss.n15259 vss.n857 263.154
R9942 vss.n5367 vss.n5339 263.154
R9943 vss.n5155 vss.n5127 263.154
R9944 vss.n15409 vss.n600 263.154
R9945 vss.n4840 vss.n4811 263.154
R9946 vss.n4892 vss.n4294 263.154
R9947 vss.n1954 vss.n1952 263.154
R9948 vss.n1893 vss.n1882 263.154
R9949 vss.n1973 vss.n1138 263.154
R9950 vss.n2803 vss.n2794 263.154
R9951 vss.n2776 vss.n2775 263.154
R9952 vss.n2790 vss.n2723 263.154
R9953 vss.n1417 vss.n1415 263.154
R9954 vss.n1403 vss.n1402 263.154
R9955 vss.n14707 vss.n1405 263.154
R9956 vss.n6956 vss.n6947 263.154
R9957 vss.n8013 vss.n2428 263.154
R9958 vss.n7999 vss.n7998 263.154
R9959 vss.n7585 vss.n7576 263.154
R9960 vss.n7558 vss.n7557 263.154
R9961 vss.n7572 vss.n7505 263.154
R9962 vss.n1674 vss.n1672 263.154
R9963 vss.n1660 vss.n1659 263.154
R9964 vss.n14557 vss.n1662 263.154
R9965 vss.n2568 vss.n2559 263.154
R9966 vss.n2542 vss.n2541 263.154
R9967 vss.n2557 vss.n2556 263.154
R9968 vss.n3223 vss.n3214 263.154
R9969 vss.n3255 vss.n3240 263.154
R9970 vss.n3271 vss.n3270 263.154
R9971 vss.n2547 vss.n2519 263.154
R9972 vss.n14564 vss.n1636 263.154
R9973 vss.n2781 vss.n2753 263.154
R9974 vss.n7563 vss.n7535 263.154
R9975 vss.n14714 vss.n1379 263.154
R9976 vss.n3262 vss.n3233 263.154
R9977 vss.n8008 vss.n2435 263.154
R9978 vss.n12127 vss.n11844 263.154
R9979 vss.n12098 vss.n12097 263.154
R9980 vss.n12119 vss.n2034 263.154
R9981 vss.n12069 vss.n12068 263.154
R9982 vss.n8401 vss.n8387 263.154
R9983 vss.n13659 vss.n13658 263.154
R9984 vss.n8577 vss.n8576 263.154
R9985 vss.n8597 vss.n8596 263.154
R9986 vss.n8603 vss.n8407 263.154
R9987 vss.n9167 vss.n9166 263.154
R9988 vss.n8945 vss.n8931 263.154
R9989 vss.n13136 vss.n13135 263.154
R9990 vss.n12835 vss.n9414 263.154
R9991 vss.n12885 vss.n9371 263.154
R9992 vss.n12871 vss.n12870 263.154
R9993 vss.n12786 vss.n12726 263.154
R9994 vss.n12808 vss.n12707 263.154
R9995 vss.n12794 vss.n12793 263.154
R9996 vss.n13312 vss.n8436 263.154
R9997 vss.n12973 vss.n12972 263.154
R9998 vss.n12977 vss.n8409 263.154
R9999 vss.n13431 vss.n13422 263.154
R10000 vss.n13403 vss.n13402 263.154
R10001 vss.n13418 vss.n13351 263.154
R10002 vss.n1980 vss.n1870 263.154
R10003 vss.n6554 vss.n6526 263.154
R10004 vss.n117 vss.n107 263.154
R10005 vss.n195 vss.n185 263.154
R10006 vss.n274 vss.n264 263.154
R10007 vss.n6578 vss.n6577 252.988
R10008 vss.n6549 vss.n6535 252.988
R10009 vss.n6564 vss.n6563 252.988
R10010 vss.n5390 vss.n5389 252.988
R10011 vss.n5362 vss.n5348 252.988
R10012 vss.n5377 vss.n5376 252.988
R10013 vss.n636 vss.n635 252.988
R10014 vss.n623 vss.n610 252.988
R10015 vss.n15403 vss.n15402 252.988
R10016 vss.n4915 vss.n4914 252.988
R10017 vss.n4887 vss.n4301 252.988
R10018 vss.n4902 vss.n4901 252.988
R10019 vss.n5178 vss.n5177 252.988
R10020 vss.n5150 vss.n5136 252.988
R10021 vss.n5165 vss.n5164 252.988
R10022 vss.n893 vss.n892 252.988
R10023 vss.n880 vss.n867 252.988
R10024 vss.n15253 vss.n15252 252.988
R10025 vss.n6462 vss.n6461 252.988
R10026 vss.n6434 vss.n6420 252.988
R10027 vss.n6449 vss.n6448 252.988
R10028 vss.n4850 vss.n4749 252.988
R10029 vss.n4833 vss.n4818 252.988
R10030 vss.n4849 vss.n4848 252.988
R10031 vss.n1952 vss.n1951 252.988
R10032 vss.n1894 vss.n1893 252.988
R10033 vss.n1974 vss.n1973 252.988
R10034 vss.n2804 vss.n2803 252.988
R10035 vss.n2776 vss.n2762 252.988
R10036 vss.n2791 vss.n2790 252.988
R10037 vss.n1415 vss.n1414 252.988
R10038 vss.n1402 vss.n1389 252.988
R10039 vss.n14708 vss.n14707 252.988
R10040 vss.n6957 vss.n6956 252.988
R10041 vss.n8014 vss.n8013 252.988
R10042 vss.n7999 vss.n2444 252.988
R10043 vss.n7586 vss.n7585 252.988
R10044 vss.n7558 vss.n7544 252.988
R10045 vss.n7573 vss.n7572 252.988
R10046 vss.n1672 vss.n1671 252.988
R10047 vss.n1659 vss.n1646 252.988
R10048 vss.n14558 vss.n14557 252.988
R10049 vss.n2569 vss.n2568 252.988
R10050 vss.n2542 vss.n2530 252.988
R10051 vss.n2556 vss.n2511 252.988
R10052 vss.n3224 vss.n3223 252.988
R10053 vss.n3256 vss.n3255 252.988
R10054 vss.n3270 vss.n3187 252.988
R10055 vss.n12121 vss.n11844 252.988
R10056 vss.n12098 vss.n11886 252.988
R10057 vss.n12120 vss.n12119 252.988
R10058 vss.n12068 vss.n12012 252.988
R10059 vss.n8401 vss.n8400 252.988
R10060 vss.n13659 vss.n8386 252.988
R10061 vss.n8576 vss.n8516 252.988
R10062 vss.n8597 vss.n8583 252.988
R10063 vss.n8603 vss.n8602 252.988
R10064 vss.n9166 vss.n9110 252.988
R10065 vss.n8945 vss.n8944 252.988
R10066 vss.n13136 vss.n8930 252.988
R10067 vss.n12836 vss.n12835 252.988
R10068 vss.n12886 vss.n12885 252.988
R10069 vss.n12871 vss.n9387 252.988
R10070 vss.n12787 vss.n12786 252.988
R10071 vss.n12809 vss.n12808 252.988
R10072 vss.n12794 vss.n12723 252.988
R10073 vss.n13313 vss.n13312 252.988
R10074 vss.n12972 vss.n12959 252.988
R10075 vss.n12977 vss.n8433 252.988
R10076 vss.n13432 vss.n13431 252.988
R10077 vss.n13403 vss.n13390 252.988
R10078 vss.n13419 vss.n13418 252.988
R10079 vss.n10340 vss.n10333 239.812
R10080 vss.n10368 vss.n10340 239.812
R10081 vss.n10375 vss.n10332 239.812
R10082 vss.n10332 vss.n10278 239.812
R10083 vss.n11654 vss.n9946 239.812
R10084 vss.n11662 vss.n11654 239.812
R10085 vss.n11668 vss.n9945 239.812
R10086 vss.n11652 vss.n9945 239.812
R10087 vss.n9943 vss.n9934 239.812
R10088 vss.n11674 vss.n9934 239.812
R10089 vss.n11417 vss.n11364 239.812
R10090 vss.n11425 vss.n11417 239.812
R10091 vss.n11431 vss.n11363 239.812
R10092 vss.n11415 vss.n11363 239.812
R10093 vss.n11361 vss.n11353 239.812
R10094 vss.n11437 vss.n11353 239.812
R10095 vss.n11312 vss.n10060 239.812
R10096 vss.n11318 vss.n10060 239.812
R10097 vss.n11311 vss.n10069 239.812
R10098 vss.n10069 vss.n10061 239.812
R10099 vss.n10077 vss.n10070 239.812
R10100 vss.n10078 vss.n10077 239.812
R10101 vss.n10705 vss.n10652 239.812
R10102 vss.n10768 vss.n10705 239.812
R10103 vss.n10774 vss.n10651 239.812
R10104 vss.n10703 vss.n10651 239.812
R10105 vss.n10649 vss.n10640 239.812
R10106 vss.n10780 vss.n10640 239.812
R10107 vss.n11941 vss.n11936 239.812
R10108 vss.n12082 vss.n11941 239.812
R10109 vss.n12089 vss.n12088 239.812
R10110 vss.n12089 vss.n11877 239.812
R10111 vss.n8370 vss.n8361 239.812
R10112 vss.n13680 vss.n8361 239.812
R10113 vss.n13674 vss.n8371 239.812
R10114 vss.n8371 vss.n8362 239.812
R10115 vss.n8377 vss.n8372 239.812
R10116 vss.n13667 vss.n8377 239.812
R10117 vss.n8334 vss.n8325 239.812
R10118 vss.n13710 vss.n8325 239.812
R10119 vss.n13704 vss.n8335 239.812
R10120 vss.n8335 vss.n8326 239.812
R10121 vss.n13382 vss.n13381 239.812
R10122 vss.n13410 vss.n13382 239.812
R10123 vss.n8500 vss.n8491 239.812
R10124 vss.n13299 vss.n8491 239.812
R10125 vss.n13293 vss.n8501 239.812
R10126 vss.n8501 vss.n8492 239.812
R10127 vss.n8507 vss.n8502 239.812
R10128 vss.n8611 vss.n8507 239.812
R10129 vss.n12944 vss.n9177 239.812
R10130 vss.n12998 vss.n9177 239.812
R10131 vss.n12992 vss.n12945 239.812
R10132 vss.n12945 vss.n9178 239.812
R10133 vss.n12951 vss.n12946 239.812
R10134 vss.n12985 vss.n12951 239.812
R10135 vss.n8914 vss.n8905 239.812
R10136 vss.n13157 vss.n8905 239.812
R10137 vss.n13151 vss.n8915 239.812
R10138 vss.n8915 vss.n8906 239.812
R10139 vss.n8921 vss.n8916 239.812
R10140 vss.n13144 vss.n8921 239.812
R10141 vss.n9362 vss.n9306 239.812
R10142 vss.n12899 vss.n9306 239.812
R10143 vss.n12893 vss.n12892 239.812
R10144 vss.n12892 vss.n9307 239.812
R10145 vss.n12880 vss.n9378 239.812
R10146 vss.n12880 vss.n12879 239.812
R10147 vss.n12698 vss.n12643 239.812
R10148 vss.n12822 vss.n12643 239.812
R10149 vss.n12816 vss.n12815 239.812
R10150 vss.n12815 vss.n12644 239.812
R10151 vss.n12803 vss.n12714 239.812
R10152 vss.n12803 vss.n12802 239.812
R10153 vss.n15675 vss.n291 239.812
R10154 vss.n299 vss.n291 239.812
R10155 vss.n15668 vss.n15667 239.812
R10156 vss.n15681 vss.n285 239.812
R10157 vss.n15682 vss.n15681 239.812
R10158 vss.n15887 vss.n19 239.812
R10159 vss.n15887 vss.n15886 239.812
R10160 vss.n24 vss.n21 239.812
R10161 vss.n6265 vss.n6257 239.812
R10162 vss.n6266 vss.n6265 239.812
R10163 vss.n214 vss.n205 239.812
R10164 vss.n15738 vss.n205 239.812
R10165 vss.n15732 vss.n215 239.812
R10166 vss.n215 vss.n206 239.812
R10167 vss.n15725 vss.n15724 239.812
R10168 vss.n136 vss.n127 239.812
R10169 vss.n15794 vss.n127 239.812
R10170 vss.n15788 vss.n137 239.812
R10171 vss.n137 vss.n128 239.812
R10172 vss.n15781 vss.n15780 239.812
R10173 vss.n57 vss.n48 239.812
R10174 vss.n15850 vss.n48 239.812
R10175 vss.n15844 vss.n58 239.812
R10176 vss.n58 vss.n49 239.812
R10177 vss.n15837 vss.n15836 239.812
R10178 vss.n914 vss.n905 239.812
R10179 vss.n15230 vss.n905 239.812
R10180 vss.n15224 vss.n915 239.812
R10181 vss.n915 vss.n906 239.812
R10182 vss.n6440 vss.n6439 239.812
R10183 vss.n855 vss.n800 239.812
R10184 vss.n15273 vss.n800 239.812
R10185 vss.n15267 vss.n856 239.812
R10186 vss.n856 vss.n801 239.812
R10187 vss.n15260 vss.n15259 239.812
R10188 vss.n756 vss.n747 239.812
R10189 vss.n15350 vss.n747 239.812
R10190 vss.n15344 vss.n757 239.812
R10191 vss.n757 vss.n748 239.812
R10192 vss.n5368 vss.n5367 239.812
R10193 vss.n657 vss.n648 239.812
R10194 vss.n15380 vss.n648 239.812
R10195 vss.n15374 vss.n658 239.812
R10196 vss.n658 vss.n649 239.812
R10197 vss.n5156 vss.n5155 239.812
R10198 vss.n598 vss.n542 239.812
R10199 vss.n15423 vss.n542 239.812
R10200 vss.n15417 vss.n599 239.812
R10201 vss.n599 vss.n543 239.812
R10202 vss.n15410 vss.n15409 239.812
R10203 vss.n450 vss.n441 239.812
R10204 vss.n15455 vss.n441 239.812
R10205 vss.n15449 vss.n451 239.812
R10206 vss.n451 vss.n442 239.812
R10207 vss.n4841 vss.n4840 239.812
R10208 vss.n4869 vss.n4363 239.812
R10209 vss.n4363 vss.n4311 239.812
R10210 vss.n4876 vss.n4310 239.812
R10211 vss.n4876 vss.n4875 239.812
R10212 vss.n4893 vss.n4892 239.812
R10213 vss.n1693 vss.n1684 239.812
R10214 vss.n14535 vss.n1684 239.812
R10215 vss.n14529 vss.n1694 239.812
R10216 vss.n1694 vss.n1685 239.812
R10217 vss.n2548 vss.n2547 239.812
R10218 vss.n1634 vss.n1579 239.812
R10219 vss.n14578 vss.n1579 239.812
R10220 vss.n14572 vss.n1635 239.812
R10221 vss.n1635 vss.n1580 239.812
R10222 vss.n14565 vss.n14564 239.812
R10223 vss.n1535 vss.n1526 239.812
R10224 vss.n14655 vss.n1526 239.812
R10225 vss.n14649 vss.n1536 239.812
R10226 vss.n1536 vss.n1527 239.812
R10227 vss.n2782 vss.n2781 239.812
R10228 vss.n1436 vss.n1427 239.812
R10229 vss.n14685 vss.n1427 239.812
R10230 vss.n14679 vss.n1437 239.812
R10231 vss.n1437 vss.n1428 239.812
R10232 vss.n7564 vss.n7563 239.812
R10233 vss.n1377 vss.n1321 239.812
R10234 vss.n14728 vss.n1321 239.812
R10235 vss.n14722 vss.n1378 239.812
R10236 vss.n1378 vss.n1322 239.812
R10237 vss.n14715 vss.n14714 239.812
R10238 vss.n1229 vss.n1220 239.812
R10239 vss.n14760 vss.n1220 239.812
R10240 vss.n14754 vss.n1230 239.812
R10241 vss.n1230 vss.n1221 239.812
R10242 vss.n3263 vss.n3262 239.812
R10243 vss.n2419 vss.n2364 239.812
R10244 vss.n8027 vss.n2364 239.812
R10245 vss.n8021 vss.n8020 239.812
R10246 vss.n8020 vss.n2365 239.812
R10247 vss.n8008 vss.n8007 239.812
R10248 vss.n1868 vss.n1859 239.812
R10249 vss.n14334 vss.n1859 239.812
R10250 vss.n14328 vss.n1869 239.812
R10251 vss.n1869 vss.n1860 239.812
R10252 vss.n1981 vss.n1980 239.812
R10253 vss.n1089 vss.n1080 239.812
R10254 vss.n15029 vss.n1080 239.812
R10255 vss.n15023 vss.n1090 239.812
R10256 vss.n1090 vss.n1081 239.812
R10257 vss.n6555 vss.n6554 239.812
R10258 vss.n81 vss.n72 239.812
R10259 vss.n15823 vss.n72 239.812
R10260 vss.n15817 vss.n82 239.812
R10261 vss.n82 vss.n73 239.812
R10262 vss.n118 vss.n117 239.812
R10263 vss.n160 vss.n151 239.812
R10264 vss.n15767 vss.n151 239.812
R10265 vss.n15761 vss.n161 239.812
R10266 vss.n161 vss.n152 239.812
R10267 vss.n196 vss.n195 239.812
R10268 vss.n238 vss.n229 239.812
R10269 vss.n15711 vss.n229 239.812
R10270 vss.n15705 vss.n239 239.812
R10271 vss.n239 vss.n230 239.812
R10272 vss.n275 vss.n274 239.812
R10273 vss.n12106 vss.n11876 239.812
R10274 vss.n12112 vss.n11876 239.812
R10275 vss.n10625 vss.n10235 239.812
R10276 vss.n10631 vss.n10235 239.812
R10277 vss.n10624 vss.n10244 239.812
R10278 vss.n10244 vss.n10236 239.812
R10279 vss.n10252 vss.n10245 239.812
R10280 vss.n10253 vss.n10252 239.812
R10281 vss.n11018 vss.n10148 239.812
R10282 vss.n11024 vss.n10148 239.812
R10283 vss.n11017 vss.n10157 239.812
R10284 vss.n10157 vss.n10149 239.812
R10285 vss.n10165 vss.n10158 239.812
R10286 vss.n10166 vss.n10165 239.812
R10287 vss.n11338 vss.n9988 239.812
R10288 vss.n11344 vss.n9988 239.812
R10289 vss.n11337 vss.n10044 239.812
R10290 vss.n10044 vss.n9989 239.812
R10291 vss.n10052 vss.n10045 239.812
R10292 vss.n11330 vss.n10052 239.812
R10293 vss.n10376 vss.n10277 239.812
R10294 vss.n10382 vss.n10277 239.812
R10295 vss.n15890 vss.n15889 229.263
R10296 vss.n62 vss.n53 229.263
R10297 vss.n111 vss.n77 229.263
R10298 vss.n141 vss.n132 229.263
R10299 vss.n189 vss.n156 229.263
R10300 vss.n219 vss.n210 229.263
R10301 vss.n268 vss.n234 229.263
R10302 vss.n294 vss.n288 229.263
R10303 vss.n10337 vss.n10327 229.263
R10304 vss.n10249 vss.n10239 229.263
R10305 vss.n10700 vss.n10645 229.263
R10306 vss.n10162 vss.n10152 229.263
R10307 vss.n10074 vss.n10064 229.263
R10308 vss.n10049 vss.n10039 229.263
R10309 vss.n11412 vss.n11357 229.263
R10310 vss.n11649 vss.n9939 229.263
R10311 vss.n10327 vss.n10326 183.912
R10312 vss.n13201 vss.n8864 183.912
R10313 vss.n11680 vss.n11679 183.912
R10314 vss.n13220 vss.n8839 183.912
R10315 vss.n11443 vss.n11442 183.912
R10316 vss.n13217 vss.n8843 183.912
R10317 vss.n11412 vss.n11411 183.912
R10318 vss.n13219 vss.n8840 183.912
R10319 vss.n11323 vss.n10055 183.912
R10320 vss.n13214 vss.n8847 183.912
R10321 vss.n11038 vss.n11037 183.912
R10322 vss.n13211 vss.n8851 183.912
R10323 vss.n10098 vss.n10064 183.912
R10324 vss.n13213 vss.n8848 183.912
R10325 vss.n10763 vss.n10754 183.912
R10326 vss.n13208 vss.n8855 183.912
R10327 vss.n10786 vss.n10785 183.912
R10328 vss.n13205 vss.n8859 183.912
R10329 vss.n10700 vss.n10699 183.912
R10330 vss.n13207 vss.n8856 183.912
R10331 vss.n10396 vss.n10395 183.912
R10332 vss.n13202 vss.n8863 183.912
R10333 vss.n13250 vss.n8808 183.912
R10334 vss.n11935 vss.n11934 183.912
R10335 vss.n12911 vss.n9274 183.912
R10336 vss.n13164 vss.n13163 183.912
R10337 vss.n12914 vss.n9205 183.912
R10338 vss.n12415 vss.n9172 183.912
R10339 vss.n13261 vss.n13260 183.912
R10340 vss.n13305 vss.n8440 183.912
R10341 vss.n13257 vss.n8688 183.912
R10342 vss.n12297 vss.n8320 183.912
R10343 vss.n13254 vss.n8756 183.912
R10344 vss.n13687 vss.n13686 183.912
R10345 vss.n13251 vss.n8807 183.912
R10346 vss.n12074 vss.n12007 183.912
R10347 vss.n13253 vss.n8804 183.912
R10348 vss.n8782 vss.n8366 183.912
R10349 vss.n13256 vss.n8735 183.912
R10350 vss.n8713 vss.n8330 183.912
R10351 vss.n13259 vss.n8685 183.912
R10352 vss.n8663 vss.n8496 183.912
R10353 vss.n12916 vss.n12915 183.912
R10354 vss.n12940 vss.n12939 183.912
R10355 vss.n12912 vss.n9255 183.912
R10356 vss.n9233 vss.n8910 183.912
R10357 vss.n12906 vss.n9281 183.912
R10358 vss.n9358 vss.n9357 183.912
R10359 vss.n12908 vss.n9278 183.912
R10360 vss.n12828 vss.n12543 183.912
R10361 vss.n12909 vss.n9277 183.912
R10362 vss.n12694 vss.n12693 183.912
R10363 vss.n6272 vss.n3987 183.912
R10364 vss.n15891 vss.n15890 183.912
R10365 vss.n6289 vss.n3660 183.912
R10366 vss.n15716 vss.n224 183.912
R10367 vss.n6286 vss.n3728 183.912
R10368 vss.n15744 vss.n15743 183.912
R10369 vss.n6287 vss.n3709 183.912
R10370 vss.n3687 vss.n210 183.912
R10371 vss.n6283 vss.n3779 183.912
R10372 vss.n15772 vss.n146 183.912
R10373 vss.n6280 vss.n3847 183.912
R10374 vss.n15800 vss.n15799 183.912
R10375 vss.n6281 vss.n3828 183.912
R10376 vss.n3806 vss.n132 183.912
R10377 vss.n6275 vss.n3947 183.912
R10378 vss.n3925 vss.n53 183.912
R10379 vss.n6277 vss.n3898 183.912
R10380 vss.n15828 vss.n67 183.912
R10381 vss.n4862 vss.n4553 183.912
R10382 vss.n6723 vss.n3309 183.912
R10383 vss.n15034 vss.n1075 183.912
R10384 vss.n6705 vss.n3333 183.912
R10385 vss.n6583 vss.n6582 183.912
R10386 vss.n6599 vss.n379 183.912
R10387 vss.n15278 vss.n795 183.912
R10388 vss.n6711 vss.n3325 183.912
R10389 vss.n15355 vss.n742 183.912
R10390 vss.n6714 vss.n3321 183.912
R10391 vss.n5395 vss.n5394 183.912
R10392 vss.n6712 vss.n3324 183.912
R10393 vss.n15385 vss.n643 183.912
R10394 vss.n6717 vss.n3317 183.912
R10395 vss.n15428 vss.n537 183.912
R10396 vss.n6720 vss.n3313 183.912
R10397 vss.n15393 vss.n628 183.912
R10398 vss.n6718 vss.n3316 183.912
R10399 vss.n4920 vss.n4919 183.912
R10400 vss.n6721 vss.n3312 183.912
R10401 vss.n5183 vss.n5182 183.912
R10402 vss.n6715 vss.n3320 183.912
R10403 vss.n15243 vss.n885 183.912
R10404 vss.n6709 vss.n3328 183.912
R10405 vss.n15235 vss.n900 183.912
R10406 vss.n6708 vss.n3329 183.912
R10407 vss.n6467 vss.n6466 183.912
R10408 vss.n6706 vss.n3332 183.912
R10409 vss.n4800 vss.n4799 183.912
R10410 vss.n6724 vss.n3308 183.912
R10411 vss.n15482 vss.n407 183.912
R10412 vss.n15036 vss.n15035 183.912
R10413 vss.n15467 vss.n427 183.912
R10414 vss.n15430 vss.n15429 183.912
R10415 vss.n15470 vss.n423 183.912
R10416 vss.n15386 vss.n642 183.912
R10417 vss.n15473 vss.n419 183.912
R10418 vss.n15357 vss.n15356 183.912
R10419 vss.n15476 vss.n415 183.912
R10420 vss.n15280 vss.n15279 183.912
R10421 vss.n15479 vss.n411 183.912
R10422 vss.n15236 vss.n899 183.912
R10423 vss.n15480 vss.n410 183.912
R10424 vss.n951 vss.n910 183.912
R10425 vss.n15477 vss.n414 183.912
R10426 vss.n851 vss.n850 183.912
R10427 vss.n15474 vss.n418 183.912
R10428 vss.n15328 vss.n752 183.912
R10429 vss.n15471 vss.n422 183.912
R10430 vss.n694 vss.n653 183.912
R10431 vss.n15468 vss.n426 183.912
R10432 vss.n594 vss.n593 183.912
R10433 vss.n15462 vss.n434 183.912
R10434 vss.n486 vss.n446 183.912
R10435 vss.n15464 vss.n431 183.912
R10436 vss.n4861 vss.n4744 183.912
R10437 vss.n15465 vss.n430 183.912
R10438 vss.n4360 vss.n4359 183.912
R10439 vss.n8032 vss.n2359 183.912
R10440 vss.n7175 vss.n6804 183.912
R10441 vss.n14339 vss.n1854 183.912
R10442 vss.n7947 vss.n2642 183.912
R10443 vss.n1964 vss.n1944 183.912
R10444 vss.n1921 vss.n1158 183.912
R10445 vss.n14583 vss.n1574 183.912
R10446 vss.n7953 vss.n2476 183.912
R10447 vss.n14660 vss.n1521 183.912
R10448 vss.n7956 vss.n2472 183.912
R10449 vss.n2809 vss.n2808 183.912
R10450 vss.n7954 vss.n2475 183.912
R10451 vss.n14690 vss.n1422 183.912
R10452 vss.n2963 vss.n2470 183.912
R10453 vss.n14733 vss.n1316 183.912
R10454 vss.n7172 vss.n7031 183.912
R10455 vss.n14698 vss.n1407 183.912
R10456 vss.n7170 vss.n7169 183.912
R10457 vss.n6962 vss.n6961 183.912
R10458 vss.n7173 vss.n6986 183.912
R10459 vss.n7591 vss.n7590 183.912
R10460 vss.n7957 vss.n2471 183.912
R10461 vss.n14548 vss.n1664 183.912
R10462 vss.n7951 vss.n2479 183.912
R10463 vss.n14540 vss.n1679 183.912
R10464 vss.n7950 vss.n2480 183.912
R10465 vss.n2574 vss.n2573 183.912
R10466 vss.n7948 vss.n2597 183.912
R10467 vss.n3228 vss.n3209 183.912
R10468 vss.n7176 vss.n6803 183.912
R10469 vss.n14787 vss.n1186 183.912
R10470 vss.n14341 vss.n14340 183.912
R10471 vss.n14772 vss.n1206 183.912
R10472 vss.n14735 vss.n14734 183.912
R10473 vss.n14775 vss.n1202 183.912
R10474 vss.n14691 vss.n1421 183.912
R10475 vss.n14778 vss.n1198 183.912
R10476 vss.n14662 vss.n14661 183.912
R10477 vss.n14781 vss.n1194 183.912
R10478 vss.n14585 vss.n14584 183.912
R10479 vss.n14784 vss.n1190 183.912
R10480 vss.n14541 vss.n1678 183.912
R10481 vss.n14785 vss.n1189 183.912
R10482 vss.n1730 vss.n1689 183.912
R10483 vss.n14782 vss.n1193 183.912
R10484 vss.n1630 vss.n1629 183.912
R10485 vss.n14779 vss.n1197 183.912
R10486 vss.n14633 vss.n1531 183.912
R10487 vss.n14776 vss.n1201 183.912
R10488 vss.n1473 vss.n1432 183.912
R10489 vss.n14773 vss.n1205 183.912
R10490 vss.n1373 vss.n1372 183.912
R10491 vss.n14767 vss.n1213 183.912
R10492 vss.n1265 vss.n1225 183.912
R10493 vss.n14769 vss.n1210 183.912
R10494 vss.n8034 vss.n8033 183.912
R10495 vss.n14770 vss.n1209 183.912
R10496 vss.n2415 vss.n2414 183.912
R10497 vss.n12075 vss.n11962 183.912
R10498 vss.n14125 vss.n14124 183.912
R10499 vss.n13685 vss.n8356 183.912
R10500 vss.n14121 vss.n2105 183.912
R10501 vss.n12061 vss.n12060 183.912
R10502 vss.n14123 vss.n2102 183.912
R10503 vss.n13716 vss.n13715 183.912
R10504 vss.n14118 vss.n2109 183.912
R10505 vss.n13304 vss.n8486 183.912
R10506 vss.n14115 vss.n2113 183.912
R10507 vss.n8564 vss.n8563 183.912
R10508 vss.n14117 vss.n2110 183.912
R10509 vss.n13004 vss.n13003 183.912
R10510 vss.n14112 vss.n2117 183.912
R10511 vss.n13162 vss.n8900 183.912
R10512 vss.n14109 vss.n2121 183.912
R10513 vss.n9159 vss.n9158 183.912
R10514 vss.n14111 vss.n2118 183.912
R10515 vss.n12827 vss.n12638 183.912
R10516 vss.n14106 vss.n2125 183.912
R10517 vss.n12841 vss.n12840 183.912
R10518 vss.n14105 vss.n2126 183.912
R10519 vss.n12775 vss.n12774 183.912
R10520 vss.n14108 vss.n2122 183.912
R10521 vss.n13318 vss.n13317 183.912
R10522 vss.n14114 vss.n2114 183.912
R10523 vss.n13437 vss.n13436 183.912
R10524 vss.n14120 vss.n2106 183.912
R10525 vss.n11866 vss.n11865 183.912
R10526 vss.n14179 vss.n14178 183.912
R10527 vss.n14788 vss.n1185 183.912
R10528 vss.n2020 vss.n1864 183.912
R10529 vss.n15483 vss.n406 183.912
R10530 vss.n1125 vss.n1085 183.912
R10531 vss.n6274 vss.n3966 183.912
R10532 vss.n15856 vss.n15855 183.912
R10533 vss.n6278 vss.n3897 183.912
R10534 vss.n3875 vss.n77 183.912
R10535 vss.n6284 vss.n3778 183.912
R10536 vss.n3756 vss.n156 183.912
R10537 vss.n6290 vss.n3659 183.912
R10538 vss.n3637 vss.n234 183.912
R10539 vss.n6310 vss.n6309 183.912
R10540 vss.n15688 vss.n15687 183.912
R10541 vss.n351 vss.n350 183.912
R10542 vss.n328 vss.n288 183.912
R10543 vss.n10587 vss.n10239 183.912
R10544 vss.n13204 vss.n8860 183.912
R10545 vss.n10981 vss.n10152 183.912
R10546 vss.n13210 vss.n8852 183.912
R10547 vss.n10039 vss.n10038 183.912
R10548 vss.n13216 vss.n8844 183.912
R10549 vss.n11649 vss.n11648 183.912
R10550 vss.n13222 vss.n8836 183.912
R10551 vss.n14764 vss.n1216 148
R10552 vss.n1224 vss.n1216 148
R10553 vss.n14757 vss.n1224 148
R10554 vss.n3227 vss.n3210 148
R10555 vss.n3219 vss.n3210 148
R10556 vss.n3219 vss.n2358 148
R10557 vss.n8031 vss.n2360 148
R10558 vss.n2368 vss.n2360 148
R10559 vss.n8024 vss.n2368 148
R10560 vss.n6960 vss.n6943 148
R10561 vss.n6952 vss.n6943 148
R10562 vss.n6952 vss.n1315 148
R10563 vss.n14732 vss.n1317 148
R10564 vss.n1325 vss.n1317 148
R10565 vss.n14725 vss.n1325 148
R10566 vss.n14697 vss.n1408 148
R10567 vss.n14693 vss.n1408 148
R10568 vss.n14693 vss.n14692 148
R10569 vss.n14689 vss.n1423 148
R10570 vss.n1431 vss.n1423 148
R10571 vss.n14682 vss.n1431 148
R10572 vss.n7589 vss.n7525 148
R10573 vss.n7581 vss.n7525 148
R10574 vss.n7581 vss.n1520 148
R10575 vss.n14659 vss.n1522 148
R10576 vss.n1530 vss.n1522 148
R10577 vss.n14652 vss.n1530 148
R10578 vss.n2807 vss.n2743 148
R10579 vss.n2799 vss.n2743 148
R10580 vss.n2799 vss.n1573 148
R10581 vss.n14582 vss.n1575 148
R10582 vss.n1583 vss.n1575 148
R10583 vss.n14575 vss.n1583 148
R10584 vss.n14547 vss.n1665 148
R10585 vss.n14543 vss.n1665 148
R10586 vss.n14543 vss.n14542 148
R10587 vss.n14539 vss.n1680 148
R10588 vss.n1688 vss.n1680 148
R10589 vss.n14532 vss.n1688 148
R10590 vss.n2572 vss.n2507 148
R10591 vss.n2564 vss.n2507 148
R10592 vss.n2564 vss.n1853 148
R10593 vss.n14338 vss.n1855 148
R10594 vss.n1863 vss.n1855 148
R10595 vss.n14331 vss.n1863 148
R10596 vss.n1963 vss.n1945 148
R10597 vss.n1959 vss.n1945 148
R10598 vss.n1959 vss.n1958 148
R10599 vss.n15459 vss.n437 148
R10600 vss.n445 vss.n437 148
R10601 vss.n15452 vss.n445 148
R10602 vss.n4853 vss.n4801 148
R10603 vss.n4801 vss.n4745 148
R10604 vss.n4860 vss.n4745 148
R10605 vss.n4866 vss.n4863 148
R10606 vss.n4866 vss.n4313 148
R10607 vss.n4872 vss.n4313 148
R10608 vss.n4918 vss.n4284 148
R10609 vss.n4910 vss.n4284 148
R10610 vss.n4910 vss.n536 148
R10611 vss.n15427 vss.n538 148
R10612 vss.n546 vss.n538 148
R10613 vss.n15420 vss.n546 148
R10614 vss.n15392 vss.n629 148
R10615 vss.n15388 vss.n629 148
R10616 vss.n15388 vss.n15387 148
R10617 vss.n15384 vss.n644 148
R10618 vss.n652 vss.n644 148
R10619 vss.n15377 vss.n652 148
R10620 vss.n5181 vss.n5117 148
R10621 vss.n5173 vss.n5117 148
R10622 vss.n5173 vss.n741 148
R10623 vss.n15354 vss.n743 148
R10624 vss.n751 vss.n743 148
R10625 vss.n15347 vss.n751 148
R10626 vss.n5393 vss.n5329 148
R10627 vss.n5385 vss.n5329 148
R10628 vss.n5385 vss.n794 148
R10629 vss.n15277 vss.n796 148
R10630 vss.n804 vss.n796 148
R10631 vss.n15270 vss.n804 148
R10632 vss.n15242 vss.n886 148
R10633 vss.n15238 vss.n886 148
R10634 vss.n15238 vss.n15237 148
R10635 vss.n15234 vss.n901 148
R10636 vss.n909 vss.n901 148
R10637 vss.n15227 vss.n909 148
R10638 vss.n6465 vss.n6401 148
R10639 vss.n6457 vss.n6401 148
R10640 vss.n6457 vss.n1074 148
R10641 vss.n15033 vss.n1076 148
R10642 vss.n1084 vss.n1076 148
R10643 vss.n15026 vss.n1084 148
R10644 vss.n6581 vss.n6516 148
R10645 vss.n6573 vss.n6516 148
R10646 vss.n6573 vss.n6571 148
R10647 vss.n12903 vss.n9302 148
R10648 vss.n9310 vss.n9302 148
R10649 vss.n12896 vss.n9310 148
R10650 vss.n12839 vss.n9410 148
R10651 vss.n12831 vss.n9410 148
R10652 vss.n12831 vss.n12829 148
R10653 vss.n12826 vss.n12639 148
R10654 vss.n12647 vss.n12639 148
R10655 vss.n12819 vss.n12647 148
R10656 vss.n12790 vss.n12776 148
R10657 vss.n12782 vss.n12776 148
R10658 vss.n12782 vss.n8899 148
R10659 vss.n13161 vss.n8901 148
R10660 vss.n8909 vss.n8901 148
R10661 vss.n13154 vss.n8909 148
R10662 vss.n9164 vss.n9163 148
R10663 vss.n9164 vss.n9106 148
R10664 vss.n9171 vss.n9106 148
R10665 vss.n13002 vss.n9173 148
R10666 vss.n9181 vss.n9173 148
R10667 vss.n12995 vss.n9181 148
R10668 vss.n13316 vss.n8429 148
R10669 vss.n13308 vss.n8429 148
R10670 vss.n13308 vss.n13306 148
R10671 vss.n13303 vss.n8487 148
R10672 vss.n8495 vss.n8487 148
R10673 vss.n13296 vss.n8495 148
R10674 vss.n8580 vss.n8565 148
R10675 vss.n8570 vss.n8565 148
R10676 vss.n8571 vss.n8570 148
R10677 vss.n13714 vss.n8321 148
R10678 vss.n8329 vss.n8321 148
R10679 vss.n13707 vss.n8329 148
R10680 vss.n13435 vss.n13371 148
R10681 vss.n13427 vss.n13371 148
R10682 vss.n13427 vss.n8355 148
R10683 vss.n13684 vss.n8357 148
R10684 vss.n8365 vss.n8357 148
R10685 vss.n13677 vss.n8365 148
R10686 vss.n12066 vss.n12065 148
R10687 vss.n12066 vss.n12008 148
R10688 vss.n12073 vss.n12008 148
R10689 vss.n12079 vss.n12076 148
R10690 vss.n12079 vss.n11938 148
R10691 vss.n12085 vss.n11938 148
R10692 vss.n12124 vss.n11867 148
R10693 vss.n11867 vss.n11840 148
R10694 vss.n12131 vss.n11840 148
R10695 vss.n11676 vss.n9933 146.834
R10696 vss.n11660 vss.n11656 146.834
R10697 vss.n11439 vss.n11352 146.834
R10698 vss.n11423 vss.n11419 146.834
R10699 vss.n11034 vss.n11032 146.834
R10700 vss.n11320 vss.n10059 146.834
R10701 vss.n10782 vss.n10639 146.834
R10702 vss.n10766 vss.n10707 146.834
R10703 vss.n13682 vss.n13681 146.834
R10704 vss.n13666 vss.n8378 146.834
R10705 vss.n13712 vss.n13711 146.834
R10706 vss.n13412 vss.n13411 146.834
R10707 vss.n13301 vss.n13300 146.834
R10708 vss.n8610 vss.n8508 146.834
R10709 vss.n13000 vss.n12999 146.834
R10710 vss.n12984 vss.n12952 146.834
R10711 vss.n13159 vss.n13158 146.834
R10712 vss.n13143 vss.n8922 146.834
R10713 vss.n12901 vss.n12900 146.834
R10714 vss.n12878 vss.n9381 146.834
R10715 vss.n12824 vss.n12823 146.834
R10716 vss.n12801 vss.n12717 146.834
R10717 vss.n15665 vss.n300 146.834
R10718 vss.n15684 vss.n15683 146.834
R10719 vss.n15877 vss.n15876 146.834
R10720 vss.n6268 vss.n6267 146.834
R10721 vss.n15722 vss.n222 146.834
R10722 vss.n15740 vss.n15739 146.834
R10723 vss.n15778 vss.n144 146.834
R10724 vss.n15796 vss.n15795 146.834
R10725 vss.n15834 vss.n65 146.834
R10726 vss.n15852 vss.n15851 146.834
R10727 vss.n6569 vss.n6565 146.834
R10728 vss.n6541 vss.n6536 146.834
R10729 vss.n5382 vss.n5378 146.834
R10730 vss.n5354 vss.n5349 146.834
R10731 vss.n639 vss.n633 146.834
R10732 vss.n615 vss.n614 146.834
R10733 vss.n4907 vss.n4903 146.834
R10734 vss.n4879 vss.n4302 146.834
R10735 vss.n5170 vss.n5166 146.834
R10736 vss.n5142 vss.n5137 146.834
R10737 vss.n896 vss.n890 146.834
R10738 vss.n872 vss.n871 146.834
R10739 vss.n6454 vss.n6450 146.834
R10740 vss.n6426 vss.n6421 146.834
R10741 vss.n4858 vss.n4748 146.834
R10742 vss.n4820 vss.n4819 146.834
R10743 vss.n6442 vss.n6441 146.834
R10744 vss.n15232 vss.n15231 146.834
R10745 vss.n15247 vss.n862 146.834
R10746 vss.n15275 vss.n15274 146.834
R10747 vss.n5370 vss.n5369 146.834
R10748 vss.n15352 vss.n15351 146.834
R10749 vss.n5158 vss.n5157 146.834
R10750 vss.n15382 vss.n15381 146.834
R10751 vss.n15397 vss.n605 146.834
R10752 vss.n15425 vss.n15424 146.834
R10753 vss.n4843 vss.n4842 146.834
R10754 vss.n15457 vss.n15456 146.834
R10755 vss.n4895 vss.n4894 146.834
R10756 vss.n4864 vss.n4364 146.834
R10757 vss.n1955 vss.n1949 146.834
R10758 vss.n1888 vss.n1880 146.834
R10759 vss.n2796 vss.n2792 146.834
R10760 vss.n2768 vss.n2763 146.834
R10761 vss.n1418 vss.n1412 146.834
R10762 vss.n1394 vss.n1393 146.834
R10763 vss.n6949 vss.n6946 146.834
R10764 vss.n8015 vss.n2425 146.834
R10765 vss.n7578 vss.n7574 146.834
R10766 vss.n7550 vss.n7545 146.834
R10767 vss.n1675 vss.n1669 146.834
R10768 vss.n1651 vss.n1650 146.834
R10769 vss.n2561 vss.n2512 146.834
R10770 vss.n2536 vss.n2531 146.834
R10771 vss.n3216 vss.n3213 146.834
R10772 vss.n3242 vss.n3239 146.834
R10773 vss.n2550 vss.n2549 146.834
R10774 vss.n14537 vss.n14536 146.834
R10775 vss.n14552 vss.n1641 146.834
R10776 vss.n14580 vss.n14579 146.834
R10777 vss.n2784 vss.n2783 146.834
R10778 vss.n14657 vss.n14656 146.834
R10779 vss.n7566 vss.n7565 146.834
R10780 vss.n14687 vss.n14686 146.834
R10781 vss.n14702 vss.n1384 146.834
R10782 vss.n14730 vss.n14729 146.834
R10783 vss.n3265 vss.n3264 146.834
R10784 vss.n14762 vss.n14761 146.834
R10785 vss.n8006 vss.n2438 146.834
R10786 vss.n8029 vss.n8028 146.834
R10787 vss.n12129 vss.n11843 146.834
R10788 vss.n11888 vss.n11887 146.834
R10789 vss.n12071 vss.n12011 146.834
R10790 vss.n8397 vss.n8391 146.834
R10791 vss.n8573 vss.n8568 146.834
R10792 vss.n8587 vss.n8586 146.834
R10793 vss.n9169 vss.n9109 146.834
R10794 vss.n8941 vss.n8935 146.834
R10795 vss.n9416 vss.n9413 146.834
R10796 vss.n12887 vss.n9368 146.834
R10797 vss.n12784 vss.n12778 146.834
R10798 vss.n12810 vss.n12704 146.834
R10799 vss.n8438 vss.n8434 146.834
R10800 vss.n12966 vss.n12965 146.834
R10801 vss.n13424 vss.n13420 146.834
R10802 vss.n13392 vss.n13391 146.834
R10803 vss.n1968 vss.n1875 146.834
R10804 vss.n14336 vss.n14335 146.834
R10805 vss.n6557 vss.n6556 146.834
R10806 vss.n15031 vss.n15030 146.834
R10807 vss.n120 vss.n119 146.834
R10808 vss.n15825 vss.n15824 146.834
R10809 vss.n198 vss.n197 146.834
R10810 vss.n15769 vss.n15768 146.834
R10811 vss.n277 vss.n276 146.834
R10812 vss.n15713 vss.n15712 146.834
R10813 vss.n12081 vss.n11942 146.834
R10814 vss.n12114 vss.n12113 146.834
R10815 vss.n10392 vss.n10390 146.834
R10816 vss.n10633 vss.n10234 146.834
R10817 vss.n10760 vss.n10758 146.834
R10818 vss.n11026 vss.n10147 146.834
R10819 vss.n11325 vss.n10053 146.834
R10820 vss.n11346 vss.n9987 146.834
R10821 vss.n10363 vss.n10341 146.834
R10822 vss.n10384 vss.n10276 146.834
R10823 vss.n13662 vss.n8378 141.34
R10824 vss.n13413 vss.n13412 141.34
R10825 vss.n8606 vss.n8508 141.34
R10826 vss.n12980 vss.n12952 141.34
R10827 vss.n13139 vss.n8922 141.34
R10828 vss.n12874 vss.n9381 141.34
R10829 vss.n12797 vss.n12717 141.34
R10830 vss.n15661 vss.n300 141.34
R10831 vss.n15878 vss.n15877 141.34
R10832 vss.n15718 vss.n222 141.34
R10833 vss.n15774 vss.n144 141.34
R10834 vss.n15830 vss.n65 141.34
R10835 vss.n6570 vss.n6569 141.34
R10836 vss.n6545 vss.n6536 141.34
R10837 vss.n5383 vss.n5382 141.34
R10838 vss.n5358 vss.n5349 141.34
R10839 vss.n640 vss.n639 141.34
R10840 vss.n615 vss.n612 141.34
R10841 vss.n4908 vss.n4907 141.34
R10842 vss.n4883 vss.n4302 141.34
R10843 vss.n5171 vss.n5170 141.34
R10844 vss.n5146 vss.n5137 141.34
R10845 vss.n897 vss.n896 141.34
R10846 vss.n872 vss.n869 141.34
R10847 vss.n6455 vss.n6454 141.34
R10848 vss.n6430 vss.n6421 141.34
R10849 vss.n4858 vss.n4857 141.34
R10850 vss.n4830 vss.n4820 141.34
R10851 vss.n6443 vss.n6442 141.34
R10852 vss.n15247 vss.n15246 141.34
R10853 vss.n5371 vss.n5370 141.34
R10854 vss.n5159 vss.n5158 141.34
R10855 vss.n15397 vss.n15396 141.34
R10856 vss.n4843 vss.n4809 141.34
R10857 vss.n4896 vss.n4895 141.34
R10858 vss.n1956 vss.n1955 141.34
R10859 vss.n1889 vss.n1888 141.34
R10860 vss.n2797 vss.n2796 141.34
R10861 vss.n2772 vss.n2763 141.34
R10862 vss.n1419 vss.n1418 141.34
R10863 vss.n1394 vss.n1391 141.34
R10864 vss.n6950 vss.n6949 141.34
R10865 vss.n2427 vss.n2425 141.34
R10866 vss.n7579 vss.n7578 141.34
R10867 vss.n7554 vss.n7545 141.34
R10868 vss.n1676 vss.n1675 141.34
R10869 vss.n1651 vss.n1648 141.34
R10870 vss.n2562 vss.n2561 141.34
R10871 vss.n2540 vss.n2531 141.34
R10872 vss.n3217 vss.n3216 141.34
R10873 vss.n3243 vss.n3242 141.34
R10874 vss.n2551 vss.n2550 141.34
R10875 vss.n14552 vss.n14551 141.34
R10876 vss.n2785 vss.n2784 141.34
R10877 vss.n7567 vss.n7566 141.34
R10878 vss.n14702 vss.n14701 141.34
R10879 vss.n3265 vss.n3231 141.34
R10880 vss.n8002 vss.n2438 141.34
R10881 vss.n12129 vss.n12128 141.34
R10882 vss.n12095 vss.n11888 141.34
R10883 vss.n12071 vss.n12070 141.34
R10884 vss.n8391 vss.n8390 141.34
R10885 vss.n8574 vss.n8573 141.34
R10886 vss.n8593 vss.n8587 141.34
R10887 vss.n9169 vss.n9168 141.34
R10888 vss.n8935 vss.n8934 141.34
R10889 vss.n9417 vss.n9416 141.34
R10890 vss.n9370 vss.n9368 141.34
R10891 vss.n12780 vss.n12778 141.34
R10892 vss.n12706 vss.n12704 141.34
R10893 vss.n8439 vss.n8438 141.34
R10894 vss.n12965 vss.n12958 141.34
R10895 vss.n13425 vss.n13424 141.34
R10896 vss.n13399 vss.n13391 141.34
R10897 vss.n1968 vss.n1967 141.34
R10898 vss.n6558 vss.n6557 141.34
R10899 vss.n120 vss.n105 141.34
R10900 vss.n198 vss.n183 141.34
R10901 vss.n277 vss.n262 141.34
R10902 vss.n12114 vss.n11875 141.34
R10903 vss.n15460 vss.n436 137.662
R10904 vss.n14765 vss.n1215 137.662
R10905 vss.n12904 vss.n9301 137.662
R10906 vss.n11676 vss.n11675 133.615
R10907 vss.n11661 vss.n11660 133.615
R10908 vss.n11439 vss.n11438 133.615
R10909 vss.n11424 vss.n11423 133.615
R10910 vss.n11034 vss.n11033 133.615
R10911 vss.n11320 vss.n11319 133.615
R10912 vss.n10782 vss.n10781 133.615
R10913 vss.n10767 vss.n10766 133.615
R10914 vss.n13682 vss.n8360 133.615
R10915 vss.n13712 vss.n8324 133.615
R10916 vss.n13301 vss.n8490 133.615
R10917 vss.n13000 vss.n9176 133.615
R10918 vss.n13159 vss.n8904 133.615
R10919 vss.n12901 vss.n9305 133.615
R10920 vss.n12824 vss.n12642 133.615
R10921 vss.n15684 vss.n283 133.615
R10922 vss.n6268 vss.n6256 133.615
R10923 vss.n15740 vss.n204 133.615
R10924 vss.n15796 vss.n126 133.615
R10925 vss.n15852 vss.n47 133.615
R10926 vss.n15232 vss.n904 133.615
R10927 vss.n15275 vss.n799 133.615
R10928 vss.n15352 vss.n746 133.615
R10929 vss.n15382 vss.n647 133.615
R10930 vss.n15425 vss.n541 133.615
R10931 vss.n15457 vss.n440 133.615
R10932 vss.n4868 vss.n4364 133.615
R10933 vss.n14537 vss.n1683 133.615
R10934 vss.n14580 vss.n1578 133.615
R10935 vss.n14657 vss.n1525 133.615
R10936 vss.n14687 vss.n1426 133.615
R10937 vss.n14730 vss.n1320 133.615
R10938 vss.n14762 vss.n1219 133.615
R10939 vss.n8029 vss.n2363 133.615
R10940 vss.n14336 vss.n1858 133.615
R10941 vss.n15031 vss.n1079 133.615
R10942 vss.n15825 vss.n71 133.615
R10943 vss.n15769 vss.n150 133.615
R10944 vss.n15713 vss.n228 133.615
R10945 vss.n12077 vss.n11942 133.615
R10946 vss.n10392 vss.n10391 133.615
R10947 vss.n10633 vss.n10632 133.615
R10948 vss.n10760 vss.n10759 133.615
R10949 vss.n11026 vss.n11025 133.615
R10950 vss.n11329 vss.n10053 133.615
R10951 vss.n11346 vss.n11345 133.615
R10952 vss.n10367 vss.n10341 133.615
R10953 vss.n10384 vss.n10383 133.615
R10954 vss.n11726 vss.n11725 130.571
R10955 vss.n15890 vss.n15 113.475
R10956 vss.n15847 vss.n53 113.475
R10957 vss.n15820 vss.n77 113.475
R10958 vss.n15791 vss.n132 113.475
R10959 vss.n15764 vss.n156 113.475
R10960 vss.n15735 vss.n210 113.475
R10961 vss.n15708 vss.n234 113.475
R10962 vss.n15678 vss.n288 113.475
R10963 vss.n10379 vss.n10327 113.475
R10964 vss.n10628 vss.n10239 113.475
R10965 vss.n10771 vss.n10700 113.475
R10966 vss.n11021 vss.n10152 113.475
R10967 vss.n11315 vss.n10064 113.475
R10968 vss.n11341 vss.n10039 113.475
R10969 vss.n11428 vss.n11412 113.475
R10970 vss.n11665 vss.n11649 113.475
R10971 vss.n6725 vss.n3307 86.5632
R10972 vss.n7178 vss.n7177 86.5632
R10973 vss.n14104 vss.n2127 86.5632
R10974 vss.n13200 vss.n8865 86.5632
R10975 vss.n3246 vss.n3244 86.0005
R10976 vss.n3251 vss.n3249 86.0005
R10977 vss.n3260 vss.n3236 86.0005
R10978 vss.n3259 vss.n3190 86.0005
R10979 vss.n3268 vss.n3267 86.0005
R10980 vss.n8018 vss.n2420 86.0005
R10981 vss.n8017 vss.n2421 86.0005
R10982 vss.n8011 vss.n8010 86.0005
R10983 vss.n8004 vss.n2430 86.0005
R10984 vss.n8001 vss.n2440 86.0005
R10985 vss.n1397 vss.n1396 86.0005
R10986 vss.n14718 vss.n1381 86.0005
R10987 vss.n14712 vss.n1382 86.0005
R10988 vss.n14711 vss.n1385 86.0005
R10989 vss.n14705 vss.n14704 86.0005
R10990 vss.n7549 vss.n7547 86.0005
R10991 vss.n7552 vss.n7540 86.0005
R10992 vss.n7561 vss.n7560 86.0005
R10993 vss.n7569 vss.n7531 86.0005
R10994 vss.n7570 vss.n7524 86.0005
R10995 vss.n2767 vss.n2765 86.0005
R10996 vss.n2770 vss.n2758 86.0005
R10997 vss.n2779 vss.n2778 86.0005
R10998 vss.n2787 vss.n2749 86.0005
R10999 vss.n2788 vss.n2742 86.0005
R11000 vss.n1654 vss.n1653 86.0005
R11001 vss.n14568 vss.n1638 86.0005
R11002 vss.n14562 vss.n1639 86.0005
R11003 vss.n14561 vss.n1642 86.0005
R11004 vss.n14555 vss.n14554 86.0005
R11005 vss.n2535 vss.n2533 86.0005
R11006 vss.n2538 vss.n2524 86.0005
R11007 vss.n2545 vss.n2544 86.0005
R11008 vss.n2553 vss.n2515 86.0005
R11009 vss.n2554 vss.n2506 86.0005
R11010 vss.n1886 vss.n1885 86.0005
R11011 vss.n1984 vss.n1872 86.0005
R11012 vss.n1978 vss.n1873 86.0005
R11013 vss.n1977 vss.n1876 86.0005
R11014 vss.n1971 vss.n1970 86.0005
R11015 vss.n4824 vss.n4822 86.0005
R11016 vss.n4828 vss.n4827 86.0005
R11017 vss.n4838 vss.n4814 86.0005
R11018 vss.n4837 vss.n4806 86.0005
R11019 vss.n4846 vss.n4845 86.0005
R11020 vss.n4878 vss.n4304 86.0005
R11021 vss.n4881 vss.n4297 86.0005
R11022 vss.n4890 vss.n4889 86.0005
R11023 vss.n4898 vss.n4290 86.0005
R11024 vss.n4899 vss.n4283 86.0005
R11025 vss.n618 vss.n617 86.0005
R11026 vss.n15413 vss.n602 86.0005
R11027 vss.n15407 vss.n603 86.0005
R11028 vss.n15406 vss.n606 86.0005
R11029 vss.n15400 vss.n15399 86.0005
R11030 vss.n5141 vss.n5139 86.0005
R11031 vss.n5144 vss.n5132 86.0005
R11032 vss.n5153 vss.n5152 86.0005
R11033 vss.n5161 vss.n5123 86.0005
R11034 vss.n5162 vss.n5116 86.0005
R11035 vss.n5353 vss.n5351 86.0005
R11036 vss.n5356 vss.n5344 86.0005
R11037 vss.n5365 vss.n5364 86.0005
R11038 vss.n5373 vss.n5335 86.0005
R11039 vss.n5374 vss.n5328 86.0005
R11040 vss.n875 vss.n874 86.0005
R11041 vss.n15263 vss.n859 86.0005
R11042 vss.n15257 vss.n860 86.0005
R11043 vss.n15256 vss.n863 86.0005
R11044 vss.n15250 vss.n15249 86.0005
R11045 vss.n6425 vss.n6423 86.0005
R11046 vss.n6428 vss.n6416 86.0005
R11047 vss.n6437 vss.n6436 86.0005
R11048 vss.n6445 vss.n6407 86.0005
R11049 vss.n6446 vss.n6400 86.0005
R11050 vss.n6540 vss.n6538 86.0005
R11051 vss.n6543 vss.n6531 86.0005
R11052 vss.n6552 vss.n6551 86.0005
R11053 vss.n6560 vss.n6522 86.0005
R11054 vss.n6561 vss.n6515 86.0005
R11055 vss.n12890 vss.n9363 86.0005
R11056 vss.n12889 vss.n9364 86.0005
R11057 vss.n12883 vss.n12882 86.0005
R11058 vss.n12876 vss.n9373 86.0005
R11059 vss.n12873 vss.n9383 86.0005
R11060 vss.n12813 vss.n12699 86.0005
R11061 vss.n12812 vss.n12700 86.0005
R11062 vss.n12806 vss.n12805 86.0005
R11063 vss.n12799 vss.n12709 86.0005
R11064 vss.n12796 vss.n12719 86.0005
R11065 vss.n8938 vss.n8937 86.0005
R11066 vss.n13147 vss.n8918 86.0005
R11067 vss.n8925 vss.n8919 86.0005
R11068 vss.n13141 vss.n8926 86.0005
R11069 vss.n13138 vss.n8927 86.0005
R11070 vss.n12963 vss.n12962 86.0005
R11071 vss.n12988 vss.n12948 86.0005
R11072 vss.n12955 vss.n12949 86.0005
R11073 vss.n12982 vss.n12956 86.0005
R11074 vss.n12979 vss.n8428 86.0005
R11075 vss.n8590 vss.n8589 86.0005
R11076 vss.n8614 vss.n8504 86.0005
R11077 vss.n8511 vss.n8505 86.0005
R11078 vss.n8608 vss.n8512 86.0005
R11079 vss.n8605 vss.n8513 86.0005
R11080 vss.n13396 vss.n13395 86.0005
R11081 vss.n13407 vss.n13384 86.0005
R11082 vss.n13405 vss.n13386 86.0005
R11083 vss.n13415 vss.n13377 86.0005
R11084 vss.n13416 vss.n13370 86.0005
R11085 vss.n8394 vss.n8393 86.0005
R11086 vss.n13670 vss.n8374 86.0005
R11087 vss.n8381 vss.n8375 86.0005
R11088 vss.n13664 vss.n8382 86.0005
R11089 vss.n13661 vss.n8383 86.0005
R11090 vss.n12092 vss.n12091 86.0005
R11091 vss.n12109 vss.n11880 86.0005
R11092 vss.n12103 vss.n11881 86.0005
R11093 vss.n12102 vss.n11872 86.0005
R11094 vss.n12117 vss.n12116 86.0005
R11095 vss.n13197 vss.n13196 71.8634
R11096 vss.n10359 vss.n10358 71.8634
R11097 vss.n10308 vss.n10307 71.8634
R11098 vss.n10324 vss.n10323 71.8634
R11099 vss.n11700 vss.n11694 71.8634
R11100 vss.n11682 vss.n11681 71.8634
R11101 vss.n11463 vss.n11457 71.8634
R11102 vss.n11445 vss.n11444 71.8634
R11103 vss.n11394 vss.n11388 71.8634
R11104 vss.n11409 vss.n11408 71.8634
R11105 vss.n11194 vss.n11188 71.8634
R11106 vss.n11176 vss.n11175 71.8634
R11107 vss.n11058 vss.n11052 71.8634
R11108 vss.n11040 vss.n11039 71.8634
R11109 vss.n10118 vss.n10112 71.8634
R11110 vss.n10100 vss.n10099 71.8634
R11111 vss.n10737 vss.n10730 71.8634
R11112 vss.n10752 vss.n10751 71.8634
R11113 vss.n10806 vss.n10800 71.8634
R11114 vss.n10788 vss.n10787 71.8634
R11115 vss.n10682 vss.n10676 71.8634
R11116 vss.n10697 vss.n10696 71.8634
R11117 vss.n10416 vss.n10410 71.8634
R11118 vss.n10398 vss.n10397 71.8634
R11119 vss.n10510 vss.n10502 71.8634
R11120 vss.n10490 vss.n10489 71.8634
R11121 vss.n10557 vss.n10551 71.8634
R11122 vss.n10538 vss.n10537 71.8634
R11123 vss.n10856 vss.n10849 71.8634
R11124 vss.n10836 vss.n10835 71.8634
R11125 vss.n10904 vss.n10896 71.8634
R11126 vss.n10884 vss.n10883 71.8634
R11127 vss.n10951 vss.n10945 71.8634
R11128 vss.n10932 vss.n10931 71.8634
R11129 vss.n11291 vss.n11284 71.8634
R11130 vss.n11271 vss.n11270 71.8634
R11131 vss.n11243 vss.n11235 71.8634
R11132 vss.n11223 vss.n11222 71.8634
R11133 vss.n11148 vss.n11142 71.8634
R11134 vss.n11129 vss.n11128 71.8634
R11135 vss.n11602 vss.n11595 71.8634
R11136 vss.n11582 vss.n11581 71.8634
R11137 vss.n11554 vss.n11546 71.8634
R11138 vss.n11534 vss.n11533 71.8634
R11139 vss.n11723 vss.n11722 71.8634
R11140 vss.n9904 vss.n9897 71.8634
R11141 vss.n11815 vss.n11813 71.8634
R11142 vss.n11830 vss.n11829 71.8634
R11143 vss.n11912 vss.n11910 71.8634
R11144 vss.n11932 vss.n11892 71.8634
R11145 vss.n9261 vss.n9260 71.8634
R11146 vss.n13169 vss.n8897 71.8634
R11147 vss.n12401 vss.n12400 71.8634
R11148 vss.n12420 vss.n12413 71.8634
R11149 vss.n9670 vss.n9628 71.8634
R11150 vss.n9654 vss.n9648 71.8634
R11151 vss.n9621 vss.n9620 71.8634
R11152 vss.n12373 vss.n12367 71.8634
R11153 vss.n13263 vss.n13262 71.8634
R11154 vss.n13281 vss.n13275 71.8634
R11155 vss.n12283 vss.n12282 71.8634
R11156 vss.n12302 vss.n12295 71.8634
R11157 vss.n9799 vss.n9758 71.8634
R11158 vss.n9783 vss.n9778 71.8634
R11159 vss.n9751 vss.n9750 71.8634
R11160 vss.n12255 vss.n12249 71.8634
R11161 vss.n8743 vss.n8742 71.8634
R11162 vss.n13692 vss.n8353 71.8634
R11163 vss.n11985 vss.n11983 71.8634
R11164 vss.n12005 vss.n11966 71.8634
R11165 vss.n11728 vss.n11727 71.8634
R11166 vss.n11749 vss.n11743 71.8634
R11167 vss.n12201 vss.n9856 71.8634
R11168 vss.n12213 vss.n12211 71.8634
R11169 vss.n8770 vss.n8761 71.8634
R11170 vss.n8783 vss.n8780 71.8634
R11171 vss.n8701 vss.n8693 71.8634
R11172 vss.n8714 vss.n8711 71.8634
R11173 vss.n9819 vss.n9809 71.8634
R11174 vss.n9831 vss.n9829 71.8634
R11175 vss.n12319 vss.n9728 71.8634
R11176 vss.n12331 vss.n12329 71.8634
R11177 vss.n8651 vss.n8642 71.8634
R11178 vss.n8664 vss.n8661 71.8634
R11179 vss.n12917 vss.n9203 71.8634
R11180 vss.n12937 vss.n9185 71.8634
R11181 vss.n9690 vss.n9680 71.8634
R11182 vss.n9703 vss.n9700 71.8634
R11183 vss.n12438 vss.n9598 71.8634
R11184 vss.n12450 vss.n12448 71.8634
R11185 vss.n9221 vss.n9212 71.8634
R11186 vss.n9234 vss.n9231 71.8634
R11187 vss.n9335 vss.n9333 71.8634
R11188 vss.n9355 vss.n9314 71.8634
R11189 vss.n12521 vss.n12519 71.8634
R11190 vss.n12541 vss.n9421 71.8634
R11191 vss.n9492 vss.n9491 71.8634
R11192 vss.n12492 vss.n12486 71.8634
R11193 vss.n9540 vss.n9499 71.8634
R11194 vss.n9524 vss.n9519 71.8634
R11195 vss.n9443 vss.n9442 71.8634
R11196 vss.n9462 vss.n9455 71.8634
R11197 vss.n12671 vss.n12669 71.8634
R11198 vss.n12691 vss.n12651 71.8634
R11199 vss.n9561 vss.n9551 71.8634
R11200 vss.n9573 vss.n9571 71.8634
R11201 vss.n10188 vss.n10187 71.8634
R11202 vss.n10205 vss.n10202 71.8634
R11203 vss.n11085 vss.n11084 71.8634
R11204 vss.n11102 vss.n11099 71.8634
R11205 vss.n11490 vss.n11489 71.8634
R11206 vss.n11507 vss.n11504 71.8634
R11207 vss.n13226 vss.n8832 71.8634
R11208 vss.n13246 vss.n8814 71.8634
R11209 vss.n15641 vss.n15640 71.8634
R11210 vss.n15651 vss.n15624 71.8634
R11211 vss.n3985 vss.n3972 71.8634
R11212 vss.n15896 vss.n13 71.8634
R11213 vss.n5651 vss.n5650 71.8634
R11214 vss.n5669 vss.n5663 71.8634
R11215 vss.n3715 vss.n3714 71.8634
R11216 vss.n15749 vss.n178 71.8634
R11217 vss.n3675 vss.n3667 71.8634
R11218 vss.n3688 vss.n3685 71.8634
R11219 vss.n5843 vss.n5842 71.8634
R11220 vss.n5861 vss.n5855 71.8634
R11221 vss.n3834 vss.n3833 71.8634
R11222 vss.n15805 vss.n100 71.8634
R11223 vss.n3794 vss.n3786 71.8634
R11224 vss.n3807 vss.n3804 71.8634
R11225 vss.n3913 vss.n3905 71.8634
R11226 vss.n3926 vss.n3923 71.8634
R11227 vss.n6083 vss.n6082 71.8634
R11228 vss.n6101 vss.n6095 71.8634
R11229 vss.n6035 vss.n6034 71.8634
R11230 vss.n6054 vss.n6047 71.8634
R11231 vss.n6197 vss.n6155 71.8634
R11232 vss.n6177 vss.n6175 71.8634
R11233 vss.n5748 vss.n5747 71.8634
R11234 vss.n5767 vss.n5761 71.8634
R11235 vss.n5795 vss.n5794 71.8634
R11236 vss.n5814 vss.n5807 71.8634
R11237 vss.n5958 vss.n5916 71.8634
R11238 vss.n5938 vss.n5936 71.8634
R11239 vss.n5560 vss.n5559 71.8634
R11240 vss.n5579 vss.n5573 71.8634
R11241 vss.n5720 vss.n5539 71.8634
R11242 vss.n5700 vss.n5698 71.8634
R11243 vss.n6330 vss.n3539 71.8634
R11244 vss.n3561 vss.n3559 71.8634
R11245 vss.n5605 vss.n5604 71.8634
R11246 vss.n5624 vss.n5618 71.8634
R11247 vss.n5880 vss.n5727 71.8634
R11248 vss.n5892 vss.n5890 71.8634
R11249 vss.n6119 vss.n5967 71.8634
R11250 vss.n6131 vss.n6129 71.8634
R11251 vss.n5988 vss.n5987 71.8634
R11252 vss.n6007 vss.n6001 71.8634
R11253 vss.n4394 vss.n4388 71.8634
R11254 vss.n4551 vss.n4550 71.8634
R11255 vss.n4485 vss.n4478 71.8634
R11256 vss.n4466 vss.n4465 71.8634
R11257 vss.n4532 vss.n4526 71.8634
R11258 vss.n4513 vss.n4512 71.8634
R11259 vss.n6652 vss.n6646 71.8634
R11260 vss.n6634 vss.n6633 71.8634
R11261 vss.n6604 vss.n6597 71.8634
R11262 vss.n6585 vss.n6584 71.8634
R11263 vss.n5250 vss.n5244 71.8634
R11264 vss.n5232 vss.n5231 71.8634
R11265 vss.n5297 vss.n5290 71.8634
R11266 vss.n5277 vss.n5276 71.8634
R11267 vss.n5531 vss.n5530 71.8634
R11268 vss.n4030 vss.n4024 71.8634
R11269 vss.n5511 vss.n5505 71.8634
R11270 vss.n5492 vss.n5491 71.8634
R11271 vss.n4074 vss.n4071 71.8634
R11272 vss.n4057 vss.n4056 71.8634
R11273 vss.n5462 vss.n5456 71.8634
R11274 vss.n5444 vss.n5443 71.8634
R11275 vss.n5415 vss.n5409 71.8634
R11276 vss.n5397 vss.n5396 71.8634
R11277 vss.n4165 vss.n4159 71.8634
R11278 vss.n4147 vss.n4146 71.8634
R11279 vss.n5085 vss.n5079 71.8634
R11280 vss.n5066 vss.n5065 71.8634
R11281 vss.n4204 vss.n4177 71.8634
R11282 vss.n4191 vss.n4190 71.8634
R11283 vss.n5037 vss.n5031 71.8634
R11284 vss.n5018 vss.n5017 71.8634
R11285 vss.n4255 vss.n4252 71.8634
R11286 vss.n4238 vss.n4237 71.8634
R11287 vss.n4988 vss.n4982 71.8634
R11288 vss.n4970 vss.n4969 71.8634
R11289 vss.n4119 vss.n4113 71.8634
R11290 vss.n4101 vss.n4100 71.8634
R11291 vss.n4940 vss.n4934 71.8634
R11292 vss.n4922 vss.n4921 71.8634
R11293 vss.n5203 vss.n5197 71.8634
R11294 vss.n5185 vss.n5184 71.8634
R11295 vss.n3378 vss.n3372 71.8634
R11296 vss.n3360 vss.n3359 71.8634
R11297 vss.n3425 vss.n3419 71.8634
R11298 vss.n3407 vss.n3406 71.8634
R11299 vss.n3484 vss.n3483 71.8634
R11300 vss.n3466 vss.n3458 71.8634
R11301 vss.n6365 vss.n3438 71.8634
R11302 vss.n6352 vss.n6346 71.8634
R11303 vss.n3532 vss.n3531 71.8634
R11304 vss.n3512 vss.n3506 71.8634
R11305 vss.n6487 vss.n6481 71.8634
R11306 vss.n6469 vss.n6468 71.8634
R11307 vss.n6681 vss.n6680 71.8634
R11308 vss.n6670 vss.n3339 71.8634
R11309 vss.n4438 vss.n4432 71.8634
R11310 vss.n4420 vss.n4419 71.8634
R11311 vss.n4781 vss.n4775 71.8634
R11312 vss.n4797 vss.n4796 71.8634
R11313 vss.n3293 vss.n3292 71.8634
R11314 vss.n6731 vss.n3305 71.8634
R11315 vss.n15519 vss.n15517 71.8634
R11316 vss.n15539 vss.n386 71.8634
R11317 vss.n14866 vss.n14853 71.8634
R11318 vss.n15491 vss.n402 71.8634
R11319 vss.n14990 vss.n14988 71.8634
R11320 vss.n15005 vss.n15004 71.8634
R11321 vss.n1060 vss.n1059 71.8634
R11322 vss.n15041 vss.n1072 71.8634
R11323 vss.n14907 vss.n14906 71.8634
R11324 vss.n14927 vss.n14921 71.8634
R11325 vss.n522 vss.n521 71.8634
R11326 vss.n15435 vss.n534 71.8634
R11327 vss.n7320 vss.n7319 71.8634
R11328 vss.n7338 vss.n7332 71.8634
R11329 vss.n7390 vss.n3062 71.8634
R11330 vss.n7374 vss.n7369 71.8634
R11331 vss.n3083 vss.n3082 71.8634
R11332 vss.n3102 vss.n3096 71.8634
R11333 vss.n727 vss.n726 71.8634
R11334 vss.n15362 vss.n739 71.8634
R11335 vss.n780 vss.n779 71.8634
R11336 vss.n15285 vss.n792 71.8634
R11337 vss.n15145 vss.n15144 71.8634
R11338 vss.n15164 vss.n15157 71.8634
R11339 vss.n15194 vss.n15193 71.8634
R11340 vss.n15212 vss.n15206 71.8634
R11341 vss.n937 vss.n936 71.8634
R11342 vss.n956 vss.n949 71.8634
R11343 vss.n828 vss.n826 71.8634
R11344 vss.n848 vss.n808 71.8634
R11345 vss.n15109 vss.n15098 71.8634
R11346 vss.n15121 vss.n15119 71.8634
R11347 vss.n7453 vss.n7444 71.8634
R11348 vss.n7465 vss.n7463 71.8634
R11349 vss.n15314 vss.n15313 71.8634
R11350 vss.n15333 vss.n15326 71.8634
R11351 vss.n680 vss.n679 71.8634
R11352 vss.n699 vss.n692 71.8634
R11353 vss.n7407 vss.n7397 71.8634
R11354 vss.n7419 vss.n7417 71.8634
R11355 vss.n7273 vss.n7272 71.8634
R11356 vss.n7292 vss.n7285 71.8634
R11357 vss.n571 vss.n569 71.8634
R11358 vss.n591 vss.n550 71.8634
R11359 vss.n472 vss.n471 71.8634
R11360 vss.n491 vss.n484 71.8634
R11361 vss.n4722 vss.n4720 71.8634
R11362 vss.n4742 vss.n4557 71.8634
R11363 vss.n4674 vss.n4673 71.8634
R11364 vss.n4693 vss.n4687 71.8634
R11365 vss.n4626 vss.n4625 71.8634
R11366 vss.n4645 vss.n4638 71.8634
R11367 vss.n4579 vss.n4578 71.8634
R11368 vss.n4598 vss.n4591 71.8634
R11369 vss.n4337 vss.n4335 71.8634
R11370 vss.n4357 vss.n4317 71.8634
R11371 vss.n7237 vss.n7227 71.8634
R11372 vss.n7249 vss.n7247 71.8634
R11373 vss.n6868 vss.n6862 71.8634
R11374 vss.n6850 vss.n6849 71.8634
R11375 vss.n7218 vss.n7217 71.8634
R11376 vss.n6822 vss.n6821 71.8634
R11377 vss.n6897 vss.n6896 71.8634
R11378 vss.n6886 vss.n6829 71.8634
R11379 vss.n2640 vss.n2639 71.8634
R11380 vss.n2623 vss.n2616 71.8634
R11381 vss.n1926 vss.n1919 71.8634
R11382 vss.n1942 vss.n1941 71.8634
R11383 vss.n2875 vss.n2869 71.8634
R11384 vss.n2857 vss.n2856 71.8634
R11385 vss.n7757 vss.n7751 71.8634
R11386 vss.n7738 vss.n7737 71.8634
R11387 vss.n2920 vss.n2887 71.8634
R11388 vss.n2907 vss.n2901 71.8634
R11389 vss.n7709 vss.n7702 71.8634
R11390 vss.n7689 vss.n7688 71.8634
R11391 vss.n3056 vss.n3055 71.8634
R11392 vss.n3036 vss.n3030 71.8634
R11393 vss.n7659 vss.n7653 71.8634
R11394 vss.n7641 vss.n7640 71.8634
R11395 vss.n2829 vss.n2823 71.8634
R11396 vss.n2811 vss.n2810 71.8634
R11397 vss.n2968 vss.n2961 71.8634
R11398 vss.n2949 vss.n2948 71.8634
R11399 vss.n7493 vss.n3008 71.8634
R11400 vss.n2995 vss.n2994 71.8634
R11401 vss.n7981 vss.n2456 71.8634
R11402 vss.n7968 vss.n7962 71.8634
R11403 vss.n7104 vss.n7100 71.8634
R11404 vss.n7089 vss.n7081 71.8634
R11405 vss.n7057 vss.n7056 71.8634
R11406 vss.n7074 vss.n7073 71.8634
R11407 vss.n7029 vss.n7028 71.8634
R11408 vss.n7012 vss.n7005 71.8634
R11409 vss.n7167 vss.n7166 71.8634
R11410 vss.n7151 vss.n7145 71.8634
R11411 vss.n6984 vss.n6983 71.8634
R11412 vss.n6967 vss.n6941 71.8634
R11413 vss.n7611 vss.n7605 71.8634
R11414 vss.n7593 vss.n7592 71.8634
R11415 vss.n7806 vss.n7800 71.8634
R11416 vss.n7788 vss.n7787 71.8634
R11417 vss.n7854 vss.n7848 71.8634
R11418 vss.n7836 vss.n7835 71.8634
R11419 vss.n7904 vss.n7897 71.8634
R11420 vss.n7884 vss.n7883 71.8634
R11421 vss.n2670 vss.n2661 71.8634
R11422 vss.n7923 vss.n7922 71.8634
R11423 vss.n2715 vss.n2712 71.8634
R11424 vss.n2698 vss.n2697 71.8634
R11425 vss.n2595 vss.n2594 71.8634
R11426 vss.n2579 vss.n2504 71.8634
R11427 vss.n14874 vss.n1154 71.8634
R11428 vss.n7932 vss.n7930 71.8634
R11429 vss.n7198 vss.n7192 71.8634
R11430 vss.n7180 vss.n7179 71.8634
R11431 vss.n6801 vss.n6800 71.8634
R11432 vss.n3207 vss.n3206 71.8634
R11433 vss.n6782 vss.n6776 71.8634
R11434 vss.n6764 vss.n6763 71.8634
R11435 vss.n14824 vss.n14822 71.8634
R11436 vss.n14844 vss.n1165 71.8634
R11437 vss.n14172 vss.n14159 71.8634
R11438 vss.n14796 vss.n1181 71.8634
R11439 vss.n14295 vss.n14293 71.8634
R11440 vss.n14310 vss.n14309 71.8634
R11441 vss.n1839 vss.n1838 71.8634
R11442 vss.n14346 vss.n1851 71.8634
R11443 vss.n14212 vss.n14211 71.8634
R11444 vss.n14232 vss.n14226 71.8634
R11445 vss.n1301 vss.n1300 71.8634
R11446 vss.n14740 vss.n1313 71.8634
R11447 vss.n14000 vss.n13999 71.8634
R11448 vss.n14018 vss.n14012 71.8634
R11449 vss.n8219 vss.n8178 71.8634
R11450 vss.n8203 vss.n8198 71.8634
R11451 vss.n8171 vss.n8170 71.8634
R11452 vss.n13972 vss.n13966 71.8634
R11453 vss.n1506 vss.n1505 71.8634
R11454 vss.n14667 vss.n1518 71.8634
R11455 vss.n1559 vss.n1558 71.8634
R11456 vss.n14590 vss.n1571 71.8634
R11457 vss.n14450 vss.n14449 71.8634
R11458 vss.n14469 vss.n14462 71.8634
R11459 vss.n14499 vss.n14498 71.8634
R11460 vss.n14517 vss.n14511 71.8634
R11461 vss.n1716 vss.n1715 71.8634
R11462 vss.n1735 vss.n1728 71.8634
R11463 vss.n1607 vss.n1605 71.8634
R11464 vss.n1627 vss.n1587 71.8634
R11465 vss.n14414 vss.n14403 71.8634
R11466 vss.n14426 vss.n14424 71.8634
R11467 vss.n13918 vss.n13909 71.8634
R11468 vss.n13930 vss.n13928 71.8634
R11469 vss.n14619 vss.n14618 71.8634
R11470 vss.n14638 vss.n14631 71.8634
R11471 vss.n1459 vss.n1458 71.8634
R11472 vss.n1478 vss.n1471 71.8634
R11473 vss.n13872 vss.n13862 71.8634
R11474 vss.n13884 vss.n13882 71.8634
R11475 vss.n14035 vss.n8148 71.8634
R11476 vss.n14047 vss.n14045 71.8634
R11477 vss.n1350 vss.n1348 71.8634
R11478 vss.n1370 vss.n1329 71.8634
R11479 vss.n1251 vss.n1250 71.8634
R11480 vss.n1270 vss.n1263 71.8634
R11481 vss.n2344 vss.n2343 71.8634
R11482 vss.n8039 vss.n2356 71.8634
R11483 vss.n2250 vss.n2249 71.8634
R11484 vss.n2269 vss.n2263 71.8634
R11485 vss.n8091 vss.n2229 71.8634
R11486 vss.n8075 vss.n8070 71.8634
R11487 vss.n2297 vss.n2296 71.8634
R11488 vss.n2316 vss.n2309 71.8634
R11489 vss.n2392 vss.n2390 71.8634
R11490 vss.n2412 vss.n2372 71.8634
R11491 vss.n8111 vss.n8101 71.8634
R11492 vss.n8123 vss.n8121 71.8634
R11493 vss.n14130 vss.n2100 71.8634
R11494 vss.n11960 vss.n11959 71.8634
R11495 vss.n13504 vss.n13498 71.8634
R11496 vss.n13486 vss.n13485 71.8634
R11497 vss.n12043 vss.n12037 71.8634
R11498 vss.n12058 vss.n12057 71.8634
R11499 vss.n13736 vss.n13730 71.8634
R11500 vss.n13718 vss.n13717 71.8634
R11501 vss.n8469 vss.n8463 71.8634
R11502 vss.n8484 vss.n8483 71.8634
R11503 vss.n8546 vss.n8540 71.8634
R11504 vss.n8561 vss.n8560 71.8634
R11505 vss.n13024 vss.n13018 71.8634
R11506 vss.n13006 vss.n13005 71.8634
R11507 vss.n8989 vss.n8983 71.8634
R11508 vss.n8971 vss.n8970 71.8634
R11509 vss.n9141 vss.n9135 71.8634
R11510 vss.n9156 vss.n9155 71.8634
R11511 vss.n12572 vss.n12566 71.8634
R11512 vss.n12636 vss.n12635 71.8634
R11513 vss.n14079 vss.n2177 71.8634
R11514 vss.n2165 vss.n2164 71.8634
R11515 vss.n12617 vss.n12611 71.8634
R11516 vss.n12598 vss.n12597 71.8634
R11517 vss.n9033 vss.n9030 71.8634
R11518 vss.n9016 vss.n9015 71.8634
R11519 vss.n13121 vss.n13114 71.8634
R11520 vss.n13101 vss.n13100 71.8634
R11521 vss.n13073 vss.n13065 71.8634
R11522 vss.n13053 vss.n13052 71.8634
R11523 vss.n9079 vss.n9073 71.8634
R11524 vss.n9060 vss.n9059 71.8634
R11525 vss.n13857 vss.n13856 71.8634
R11526 vss.n8247 vss.n8241 71.8634
R11527 vss.n13833 vss.n13826 71.8634
R11528 vss.n13813 vss.n13812 71.8634
R11529 vss.n13785 vss.n13777 71.8634
R11530 vss.n13765 vss.n13764 71.8634
R11531 vss.n8293 vss.n8287 71.8634
R11532 vss.n8274 vss.n8273 71.8634
R11533 vss.n13548 vss.n13545 71.8634
R11534 vss.n13531 vss.n13530 71.8634
R11535 vss.n13644 vss.n13637 71.8634
R11536 vss.n13624 vss.n13623 71.8634
R11537 vss.n13596 vss.n13588 71.8634
R11538 vss.n13576 vss.n13575 71.8634
R11539 vss.n14153 vss.n14152 71.8634
R11540 vss.n2080 vss.n2072 71.8634
R11541 vss.n2222 vss.n2221 71.8634
R11542 vss.n2205 vss.n2198 71.8634
R11543 vss.n14101 vss.n14100 71.8634
R11544 vss.n9299 vss.n9298 71.8634
R11545 vss.n12861 vss.n12855 71.8634
R11546 vss.n12843 vss.n12842 71.8634
R11547 vss.n12756 vss.n12750 71.8634
R11548 vss.n12772 vss.n12771 71.8634
R11549 vss.n13338 vss.n13332 71.8634
R11550 vss.n13320 vss.n13319 71.8634
R11551 vss.n13457 vss.n13451 71.8634
R11552 vss.n13439 vss.n13438 71.8634
R11553 vss.n14182 vss.n2048 71.8634
R11554 vss.n11863 vss.n11862 71.8634
R11555 vss.n1781 vss.n1771 71.8634
R11556 vss.n1793 vss.n1791 71.8634
R11557 vss.n14363 vss.n1818 71.8634
R11558 vss.n14375 vss.n14373 71.8634
R11559 vss.n2006 vss.n2005 71.8634
R11560 vss.n2025 vss.n2018 71.8634
R11561 vss.n14265 vss.n14264 71.8634
R11562 vss.n14274 vss.n14273 71.8634
R11563 vss.n1002 vss.n992 71.8634
R11564 vss.n1014 vss.n1012 71.8634
R11565 vss.n15058 vss.n1039 71.8634
R11566 vss.n15070 vss.n15068 71.8634
R11567 vss.n1111 vss.n1110 71.8634
R11568 vss.n1130 vss.n1123 71.8634
R11569 vss.n14960 vss.n14959 71.8634
R11570 vss.n14969 vss.n14968 71.8634
R11571 vss.n6217 vss.n6208 71.8634
R11572 vss.n6229 vss.n6227 71.8634
R11573 vss.n3953 vss.n3952 71.8634
R11574 vss.n15861 vss.n42 71.8634
R11575 vss.n3863 vss.n3854 71.8634
R11576 vss.n3876 vss.n3873 71.8634
R11577 vss.n3744 vss.n3735 71.8634
R11578 vss.n3757 vss.n3754 71.8634
R11579 vss.n3625 vss.n3616 71.8634
R11580 vss.n3638 vss.n3635 71.8634
R11581 vss.n6307 vss.n6294 71.8634
R11582 vss.n15693 vss.n257 71.8634
R11583 vss.n15603 vss.n15602 71.8634
R11584 vss.n15612 vss.n15611 71.8634
R11585 vss.n316 vss.n308 71.8634
R11586 vss.n329 vss.n326 71.8634
R11587 vss.n3587 vss.n3585 71.8634
R11588 vss.n3609 vss.n3567 71.8634
R11589 vss.n15549 vss.n15548 71.8634
R11590 vss.n15567 vss.n15561 71.8634
R11591 vss.n12178 vss.n12136 71.8634
R11592 vss.n12159 vss.n12157 71.8634
R11593 vss.n11790 vss.n11769 71.8634
R11594 vss.n11784 vss.n11783 71.8634
R11595 vss.n10462 vss.n10455 71.8634
R11596 vss.n10443 vss.n10442 71.8634
R11597 vss.n10607 vss.n10601 71.8634
R11598 vss.n10589 vss.n10588 71.8634
R11599 vss.n11001 vss.n10995 71.8634
R11600 vss.n10983 vss.n10982 71.8634
R11601 vss.n10020 vss.n10014 71.8634
R11602 vss.n10036 vss.n10035 71.8634
R11603 vss.n11630 vss.n11629 71.8634
R11604 vss.n11646 vss.n11645 71.8634
R11605 vss.n10348 vss.n10347 68.5181
R11606 vss.n10357 vss.n10348 68.5181
R11607 vss.n13185 vss.n8877 68.5181
R11608 vss.n8877 vss.n8871 68.5181
R11609 vss.n13186 vss.n8870 68.5181
R11610 vss.n13195 vss.n8870 68.5181
R11611 vss.n10295 vss.n10285 68.5181
R11612 vss.n10322 vss.n10285 68.5181
R11613 vss.n10316 vss.n10315 68.5181
R11614 vss.n10316 vss.n10286 68.5181
R11615 vss.n10303 vss.n10297 68.5181
R11616 vss.n10306 vss.n10303 68.5181
R11617 vss.n11693 vss.n9913 68.5181
R11618 vss.n11701 vss.n11693 68.5181
R11619 vss.n11707 vss.n9911 68.5181
R11620 vss.n11691 vss.n9911 68.5181
R11621 vss.n9927 vss.n9926 68.5181
R11622 vss.n9926 vss.n9921 68.5181
R11623 vss.n11456 vss.n9968 68.5181
R11624 vss.n11464 vss.n11456 68.5181
R11625 vss.n11470 vss.n9966 68.5181
R11626 vss.n11454 vss.n9966 68.5181
R11627 vss.n9982 vss.n9981 68.5181
R11628 vss.n9981 vss.n9976 68.5181
R11629 vss.n11387 vss.n11382 68.5181
R11630 vss.n11395 vss.n11387 68.5181
R11631 vss.n11401 vss.n11381 68.5181
R11632 vss.n11381 vss.n11371 68.5181
R11633 vss.n11379 vss.n11370 68.5181
R11634 vss.n11407 vss.n11370 68.5181
R11635 vss.n11187 vss.n11159 68.5181
R11636 vss.n11195 vss.n11187 68.5181
R11637 vss.n11201 vss.n11157 68.5181
R11638 vss.n11185 vss.n11157 68.5181
R11639 vss.n11173 vss.n11172 68.5181
R11640 vss.n11172 vss.n11167 68.5181
R11641 vss.n11051 vss.n10128 68.5181
R11642 vss.n11059 vss.n11051 68.5181
R11643 vss.n11065 vss.n10126 68.5181
R11644 vss.n11049 vss.n10126 68.5181
R11645 vss.n10142 vss.n10141 68.5181
R11646 vss.n10141 vss.n10136 68.5181
R11647 vss.n10111 vss.n10082 68.5181
R11648 vss.n10119 vss.n10111 68.5181
R11649 vss.n10125 vss.n10080 68.5181
R11650 vss.n10109 vss.n10080 68.5181
R11651 vss.n10096 vss.n10095 68.5181
R11652 vss.n10095 vss.n10090 68.5181
R11653 vss.n10732 vss.n10729 68.5181
R11654 vss.n10738 vss.n10729 68.5181
R11655 vss.n10722 vss.n10168 68.5181
R11656 vss.n10722 vss.n10715 68.5181
R11657 vss.n10744 vss.n10714 68.5181
R11658 vss.n10750 vss.n10714 68.5181
R11659 vss.n10799 vss.n10215 68.5181
R11660 vss.n10807 vss.n10799 68.5181
R11661 vss.n10813 vss.n10213 68.5181
R11662 vss.n10797 vss.n10213 68.5181
R11663 vss.n10229 vss.n10228 68.5181
R11664 vss.n10228 vss.n10223 68.5181
R11665 vss.n10675 vss.n10670 68.5181
R11666 vss.n10683 vss.n10675 68.5181
R11667 vss.n10689 vss.n10669 68.5181
R11668 vss.n10669 vss.n10659 68.5181
R11669 vss.n10667 vss.n10658 68.5181
R11670 vss.n10695 vss.n10658 68.5181
R11671 vss.n10409 vss.n10257 68.5181
R11672 vss.n10417 vss.n10409 68.5181
R11673 vss.n10423 vss.n10255 68.5181
R11674 vss.n10407 vss.n10255 68.5181
R11675 vss.n10271 vss.n10270 68.5181
R11676 vss.n10270 vss.n10265 68.5181
R11677 vss.n10454 vss.n10426 68.5181
R11678 vss.n10463 vss.n10454 68.5181
R11679 vss.n10469 vss.n10424 68.5181
R11680 vss.n10452 vss.n10424 68.5181
R11681 vss.n10487 vss.n10486 68.5181
R11682 vss.n10486 vss.n10481 68.5181
R11683 vss.n10517 vss.n10471 68.5181
R11684 vss.n10499 vss.n10471 68.5181
R11685 vss.n10501 vss.n10473 68.5181
R11686 vss.n10511 vss.n10501 68.5181
R11687 vss.n10535 vss.n10534 68.5181
R11688 vss.n10534 vss.n10529 68.5181
R11689 vss.n10564 vss.n10519 68.5181
R11690 vss.n10548 vss.n10519 68.5181
R11691 vss.n10550 vss.n10521 68.5181
R11692 vss.n10558 vss.n10550 68.5181
R11693 vss.n10833 vss.n10832 68.5181
R11694 vss.n10832 vss.n10827 68.5181
R11695 vss.n10863 vss.n10817 68.5181
R11696 vss.n10846 vss.n10817 68.5181
R11697 vss.n10848 vss.n10819 68.5181
R11698 vss.n10857 vss.n10848 68.5181
R11699 vss.n10881 vss.n10880 68.5181
R11700 vss.n10880 vss.n10875 68.5181
R11701 vss.n10911 vss.n10865 68.5181
R11702 vss.n10893 vss.n10865 68.5181
R11703 vss.n10895 vss.n10867 68.5181
R11704 vss.n10905 vss.n10895 68.5181
R11705 vss.n10929 vss.n10928 68.5181
R11706 vss.n10928 vss.n10923 68.5181
R11707 vss.n10958 vss.n10913 68.5181
R11708 vss.n10942 vss.n10913 68.5181
R11709 vss.n10944 vss.n10915 68.5181
R11710 vss.n10952 vss.n10944 68.5181
R11711 vss.n11268 vss.n11267 68.5181
R11712 vss.n11267 vss.n11262 68.5181
R11713 vss.n11298 vss.n11252 68.5181
R11714 vss.n11281 vss.n11252 68.5181
R11715 vss.n11283 vss.n11254 68.5181
R11716 vss.n11292 vss.n11283 68.5181
R11717 vss.n11220 vss.n11219 68.5181
R11718 vss.n11219 vss.n11214 68.5181
R11719 vss.n11250 vss.n11204 68.5181
R11720 vss.n11232 vss.n11204 68.5181
R11721 vss.n11234 vss.n11206 68.5181
R11722 vss.n11244 vss.n11234 68.5181
R11723 vss.n11126 vss.n11125 68.5181
R11724 vss.n11125 vss.n11120 68.5181
R11725 vss.n11155 vss.n11110 68.5181
R11726 vss.n11139 vss.n11110 68.5181
R11727 vss.n11141 vss.n11112 68.5181
R11728 vss.n11149 vss.n11141 68.5181
R11729 vss.n11579 vss.n11578 68.5181
R11730 vss.n11578 vss.n11573 68.5181
R11731 vss.n11609 vss.n11563 68.5181
R11732 vss.n11592 vss.n11563 68.5181
R11733 vss.n11594 vss.n11565 68.5181
R11734 vss.n11603 vss.n11594 68.5181
R11735 vss.n11531 vss.n11530 68.5181
R11736 vss.n11530 vss.n11525 68.5181
R11737 vss.n11561 vss.n11515 68.5181
R11738 vss.n11543 vss.n11515 68.5181
R11739 vss.n11545 vss.n11517 68.5181
R11740 vss.n11555 vss.n11545 68.5181
R11741 vss.n9896 vss.n9891 68.5181
R11742 vss.n9905 vss.n9896 68.5181
R11743 vss.n11711 vss.n9890 68.5181
R11744 vss.n9890 vss.n9884 68.5181
R11745 vss.n11712 vss.n9883 68.5181
R11746 vss.n11721 vss.n9883 68.5181
R11747 vss.n11827 vss.n11824 68.5181
R11748 vss.n11824 vss.n11805 68.5181
R11749 vss.n11825 vss.n11803 68.5181
R11750 vss.n12187 vss.n11803 68.5181
R11751 vss.n11836 vss.n11814 68.5181
R11752 vss.n11837 vss.n11836 68.5181
R11753 vss.n11924 vss.n11893 68.5181
R11754 vss.n11930 vss.n11893 68.5181
R11755 vss.n11923 vss.n11903 68.5181
R11756 vss.n11903 vss.n11894 68.5181
R11757 vss.n11909 vss.n11904 68.5181
R11758 vss.n11917 vss.n11909 68.5181
R11759 vss.n13170 vss.n8896 68.5181
R11760 vss.n8896 vss.n8886 68.5181
R11761 vss.n8894 vss.n8884 68.5181
R11762 vss.n13176 vss.n8884 68.5181
R11763 vss.n9269 vss.n9262 68.5181
R11764 vss.n9270 vss.n9269 68.5181
R11765 vss.n12421 vss.n12412 68.5181
R11766 vss.n12412 vss.n12384 68.5181
R11767 vss.n12410 vss.n12382 68.5181
R11768 vss.n12427 vss.n12382 68.5181
R11769 vss.n12397 vss.n12392 68.5181
R11770 vss.n12398 vss.n12397 68.5181
R11771 vss.n12447 vss.n12442 68.5181
R11772 vss.n12456 vss.n12447 68.5181
R11773 vss.n12462 vss.n12441 68.5181
R11774 vss.n12441 vss.n12432 68.5181
R11775 vss.n9646 vss.n9641 68.5181
R11776 vss.n9656 vss.n9646 68.5181
R11777 vss.n9662 vss.n9640 68.5181
R11778 vss.n9640 vss.n9630 68.5181
R11779 vss.n9638 vss.n9629 68.5181
R11780 vss.n9668 vss.n9629 68.5181
R11781 vss.n12374 vss.n12366 68.5181
R11782 vss.n12366 vss.n9604 68.5181
R11783 vss.n12364 vss.n9602 68.5181
R11784 vss.n12380 vss.n9602 68.5181
R11785 vss.n9617 vss.n9612 68.5181
R11786 vss.n9618 vss.n9617 68.5181
R11787 vss.n13282 vss.n13274 68.5181
R11788 vss.n13274 vss.n8621 68.5181
R11789 vss.n13272 vss.n8619 68.5181
R11790 vss.n13288 vss.n8619 68.5181
R11791 vss.n8634 vss.n8629 68.5181
R11792 vss.n8635 vss.n8634 68.5181
R11793 vss.n12303 vss.n12294 68.5181
R11794 vss.n12294 vss.n12266 68.5181
R11795 vss.n12292 vss.n12264 68.5181
R11796 vss.n12309 vss.n12264 68.5181
R11797 vss.n12279 vss.n12274 68.5181
R11798 vss.n12280 vss.n12279 68.5181
R11799 vss.n12328 vss.n12323 68.5181
R11800 vss.n12337 vss.n12328 68.5181
R11801 vss.n12343 vss.n12322 68.5181
R11802 vss.n12322 vss.n12313 68.5181
R11803 vss.n9776 vss.n9771 68.5181
R11804 vss.n9785 vss.n9776 68.5181
R11805 vss.n9791 vss.n9770 68.5181
R11806 vss.n9770 vss.n9760 68.5181
R11807 vss.n9768 vss.n9759 68.5181
R11808 vss.n9797 vss.n9759 68.5181
R11809 vss.n12256 vss.n12248 68.5181
R11810 vss.n12248 vss.n9734 68.5181
R11811 vss.n12246 vss.n9732 68.5181
R11812 vss.n12262 vss.n9732 68.5181
R11813 vss.n9747 vss.n9742 68.5181
R11814 vss.n9748 vss.n9747 68.5181
R11815 vss.n13693 vss.n8352 68.5181
R11816 vss.n8352 vss.n8342 68.5181
R11817 vss.n8350 vss.n8340 68.5181
R11818 vss.n13699 vss.n8340 68.5181
R11819 vss.n8751 vss.n8744 68.5181
R11820 vss.n8752 vss.n8751 68.5181
R11821 vss.n11997 vss.n11967 68.5181
R11822 vss.n12003 vss.n11967 68.5181
R11823 vss.n11996 vss.n11976 68.5181
R11824 vss.n11976 vss.n9858 68.5181
R11825 vss.n11982 vss.n11977 68.5181
R11826 vss.n11990 vss.n11982 68.5181
R11827 vss.n11750 vss.n11742 68.5181
R11828 vss.n11742 vss.n9863 68.5181
R11829 vss.n11740 vss.n9861 68.5181
R11830 vss.n11756 vss.n9861 68.5181
R11831 vss.n9876 vss.n9871 68.5181
R11832 vss.n9877 vss.n9876 68.5181
R11833 vss.n12210 vss.n12205 68.5181
R11834 vss.n12219 vss.n12210 68.5181
R11835 vss.n12225 vss.n12204 68.5181
R11836 vss.n12204 vss.n12195 68.5181
R11837 vss.n12202 vss.n9857 68.5181
R11838 vss.n12231 vss.n9857 68.5181
R11839 vss.n8779 vss.n8774 68.5181
R11840 vss.n8788 vss.n8779 68.5181
R11841 vss.n8794 vss.n8773 68.5181
R11842 vss.n8773 vss.n8764 68.5181
R11843 vss.n8771 vss.n8762 68.5181
R11844 vss.n8800 vss.n8762 68.5181
R11845 vss.n8710 vss.n8705 68.5181
R11846 vss.n8719 vss.n8710 68.5181
R11847 vss.n8725 vss.n8704 68.5181
R11848 vss.n8704 vss.n8695 68.5181
R11849 vss.n8702 vss.n8694 68.5181
R11850 vss.n8731 vss.n8694 68.5181
R11851 vss.n9828 vss.n9823 68.5181
R11852 vss.n9836 vss.n9828 68.5181
R11853 vss.n9842 vss.n9822 68.5181
R11854 vss.n9822 vss.n9811 68.5181
R11855 vss.n9820 vss.n9810 68.5181
R11856 vss.n9848 vss.n9810 68.5181
R11857 vss.n12320 vss.n9729 68.5181
R11858 vss.n12349 vss.n9729 68.5181
R11859 vss.n8660 vss.n8655 68.5181
R11860 vss.n8669 vss.n8660 68.5181
R11861 vss.n8675 vss.n8654 68.5181
R11862 vss.n8654 vss.n8645 68.5181
R11863 vss.n8652 vss.n8643 68.5181
R11864 vss.n8681 vss.n8643 68.5181
R11865 vss.n12929 vss.n9186 68.5181
R11866 vss.n12935 vss.n9186 68.5181
R11867 vss.n12928 vss.n9196 68.5181
R11868 vss.n9196 vss.n9187 68.5181
R11869 vss.n9202 vss.n9197 68.5181
R11870 vss.n12922 vss.n9202 68.5181
R11871 vss.n9699 vss.n9694 68.5181
R11872 vss.n9708 vss.n9699 68.5181
R11873 vss.n9714 vss.n9693 68.5181
R11874 vss.n9693 vss.n9682 68.5181
R11875 vss.n9691 vss.n9681 68.5181
R11876 vss.n9720 vss.n9681 68.5181
R11877 vss.n12439 vss.n9599 68.5181
R11878 vss.n12468 vss.n9599 68.5181
R11879 vss.n9230 vss.n9225 68.5181
R11880 vss.n9239 vss.n9230 68.5181
R11881 vss.n9245 vss.n9224 68.5181
R11882 vss.n9224 vss.n9215 68.5181
R11883 vss.n9222 vss.n9213 68.5181
R11884 vss.n9251 vss.n9213 68.5181
R11885 vss.n9347 vss.n9315 68.5181
R11886 vss.n9353 vss.n9315 68.5181
R11887 vss.n9346 vss.n9326 68.5181
R11888 vss.n9326 vss.n9317 68.5181
R11889 vss.n9332 vss.n9327 68.5181
R11890 vss.n9340 vss.n9332 68.5181
R11891 vss.n12533 vss.n9422 68.5181
R11892 vss.n12539 vss.n9422 68.5181
R11893 vss.n12532 vss.n12512 68.5181
R11894 vss.n12512 vss.n12503 68.5181
R11895 vss.n12518 vss.n12513 68.5181
R11896 vss.n12526 vss.n12518 68.5181
R11897 vss.n12493 vss.n12485 68.5181
R11898 vss.n12485 vss.n9475 68.5181
R11899 vss.n12483 vss.n9473 68.5181
R11900 vss.n12499 vss.n9473 68.5181
R11901 vss.n9488 vss.n9483 68.5181
R11902 vss.n9489 vss.n9488 68.5181
R11903 vss.n9517 vss.n9512 68.5181
R11904 vss.n9526 vss.n9517 68.5181
R11905 vss.n9532 vss.n9511 68.5181
R11906 vss.n9511 vss.n9501 68.5181
R11907 vss.n9509 vss.n9500 68.5181
R11908 vss.n9538 vss.n9500 68.5181
R11909 vss.n9463 vss.n9454 68.5181
R11910 vss.n9454 vss.n9425 68.5181
R11911 vss.n9452 vss.n9423 68.5181
R11912 vss.n9469 vss.n9423 68.5181
R11913 vss.n9438 vss.n9433 68.5181
R11914 vss.n9439 vss.n9438 68.5181
R11915 vss.n12683 vss.n12652 68.5181
R11916 vss.n12689 vss.n12652 68.5181
R11917 vss.n12682 vss.n12662 68.5181
R11918 vss.n12662 vss.n12653 68.5181
R11919 vss.n12668 vss.n12663 68.5181
R11920 vss.n12676 vss.n12668 68.5181
R11921 vss.n9570 vss.n9565 68.5181
R11922 vss.n9578 vss.n9570 68.5181
R11923 vss.n9584 vss.n9564 68.5181
R11924 vss.n9564 vss.n9553 68.5181
R11925 vss.n9562 vss.n9552 68.5181
R11926 vss.n9590 vss.n9552 68.5181
R11927 vss.n10212 vss.n10169 68.5181
R11928 vss.n10197 vss.n10169 68.5181
R11929 vss.n10185 vss.n10184 68.5181
R11930 vss.n10184 vss.n10179 68.5181
R11931 vss.n10199 vss.n10171 68.5181
R11932 vss.n10206 vss.n10199 68.5181
R11933 vss.n11109 vss.n11066 68.5181
R11934 vss.n11094 vss.n11066 68.5181
R11935 vss.n11082 vss.n11081 68.5181
R11936 vss.n11081 vss.n11076 68.5181
R11937 vss.n11096 vss.n11068 68.5181
R11938 vss.n11103 vss.n11096 68.5181
R11939 vss.n11514 vss.n11471 68.5181
R11940 vss.n11499 vss.n11471 68.5181
R11941 vss.n11487 vss.n11486 68.5181
R11942 vss.n11486 vss.n11481 68.5181
R11943 vss.n11501 vss.n11473 68.5181
R11944 vss.n11508 vss.n11501 68.5181
R11945 vss.n13238 vss.n8815 68.5181
R11946 vss.n13244 vss.n8815 68.5181
R11947 vss.n13237 vss.n8825 68.5181
R11948 vss.n8825 vss.n8816 68.5181
R11949 vss.n8831 vss.n8826 68.5181
R11950 vss.n13231 vss.n8831 68.5181
R11951 vss.n15568 vss.n15560 68.5181
R11952 vss.n15560 vss.n362 68.5181
R11953 vss.n15558 vss.n360 68.5181
R11954 vss.n15574 vss.n360 68.5181
R11955 vss.n15645 vss.n15623 68.5181
R11956 vss.n15653 vss.n15623 68.5181
R11957 vss.n15644 vss.n15631 68.5181
R11958 vss.n15631 vss.n15622 68.5181
R11959 vss.n15642 vss.n15635 68.5181
R11960 vss.n15637 vss.n15635 68.5181
R11961 vss.n325 vss.n320 68.5181
R11962 vss.n334 vss.n325 68.5181
R11963 vss.n340 vss.n319 68.5181
R11964 vss.n319 vss.n310 68.5181
R11965 vss.n15897 vss.n12 68.5181
R11966 vss.n12 vss.n2 68.5181
R11967 vss.n10 vss.n0 68.5181
R11968 vss.n15903 vss.n0 68.5181
R11969 vss.n3982 vss.n3973 68.5181
R11970 vss.n3983 vss.n3982 68.5181
R11971 vss.n5670 vss.n5662 68.5181
R11972 vss.n5662 vss.n5634 68.5181
R11973 vss.n5660 vss.n5632 68.5181
R11974 vss.n5676 vss.n5632 68.5181
R11975 vss.n5647 vss.n5642 68.5181
R11976 vss.n5648 vss.n5647 68.5181
R11977 vss.n15750 vss.n177 68.5181
R11978 vss.n177 vss.n167 68.5181
R11979 vss.n175 vss.n165 68.5181
R11980 vss.n15756 vss.n165 68.5181
R11981 vss.n3723 vss.n3716 68.5181
R11982 vss.n3724 vss.n3723 68.5181
R11983 vss.n3684 vss.n3679 68.5181
R11984 vss.n3693 vss.n3684 68.5181
R11985 vss.n3699 vss.n3678 68.5181
R11986 vss.n3678 vss.n3669 68.5181
R11987 vss.n3676 vss.n3668 68.5181
R11988 vss.n3705 vss.n3668 68.5181
R11989 vss.n5862 vss.n5854 68.5181
R11990 vss.n5854 vss.n5826 68.5181
R11991 vss.n5852 vss.n5824 68.5181
R11992 vss.n5868 vss.n5824 68.5181
R11993 vss.n5839 vss.n5834 68.5181
R11994 vss.n5840 vss.n5839 68.5181
R11995 vss.n15806 vss.n99 68.5181
R11996 vss.n99 vss.n89 68.5181
R11997 vss.n97 vss.n87 68.5181
R11998 vss.n15812 vss.n87 68.5181
R11999 vss.n3842 vss.n3835 68.5181
R12000 vss.n3843 vss.n3842 68.5181
R12001 vss.n3803 vss.n3798 68.5181
R12002 vss.n3812 vss.n3803 68.5181
R12003 vss.n3818 vss.n3797 68.5181
R12004 vss.n3797 vss.n3788 68.5181
R12005 vss.n3795 vss.n3787 68.5181
R12006 vss.n3824 vss.n3787 68.5181
R12007 vss.n3922 vss.n3917 68.5181
R12008 vss.n3931 vss.n3922 68.5181
R12009 vss.n3937 vss.n3916 68.5181
R12010 vss.n3916 vss.n3907 68.5181
R12011 vss.n3914 vss.n3906 68.5181
R12012 vss.n3943 vss.n3906 68.5181
R12013 vss.n6102 vss.n6094 68.5181
R12014 vss.n6094 vss.n6066 68.5181
R12015 vss.n6092 vss.n6064 68.5181
R12016 vss.n6108 vss.n6064 68.5181
R12017 vss.n6079 vss.n6074 68.5181
R12018 vss.n6080 vss.n6079 68.5181
R12019 vss.n6226 vss.n6221 68.5181
R12020 vss.n6235 vss.n6226 68.5181
R12021 vss.n6241 vss.n6220 68.5181
R12022 vss.n6220 vss.n6211 68.5181
R12023 vss.n6055 vss.n6046 68.5181
R12024 vss.n6046 vss.n6018 68.5181
R12025 vss.n6044 vss.n6016 68.5181
R12026 vss.n6061 vss.n6016 68.5181
R12027 vss.n6031 vss.n6026 68.5181
R12028 vss.n6032 vss.n6031 68.5181
R12029 vss.n6174 vss.n6169 68.5181
R12030 vss.n6183 vss.n6174 68.5181
R12031 vss.n6189 vss.n6168 68.5181
R12032 vss.n6168 vss.n6158 68.5181
R12033 vss.n6166 vss.n6156 68.5181
R12034 vss.n6195 vss.n6156 68.5181
R12035 vss.n5768 vss.n5760 68.5181
R12036 vss.n5760 vss.n5731 68.5181
R12037 vss.n5758 vss.n5729 68.5181
R12038 vss.n5774 vss.n5729 68.5181
R12039 vss.n5749 vss.n5739 68.5181
R12040 vss.n5750 vss.n5749 68.5181
R12041 vss.n5815 vss.n5806 68.5181
R12042 vss.n5806 vss.n5778 68.5181
R12043 vss.n5804 vss.n5776 68.5181
R12044 vss.n5821 vss.n5776 68.5181
R12045 vss.n5791 vss.n5786 68.5181
R12046 vss.n5792 vss.n5791 68.5181
R12047 vss.n5935 vss.n5930 68.5181
R12048 vss.n5944 vss.n5935 68.5181
R12049 vss.n5950 vss.n5929 68.5181
R12050 vss.n5929 vss.n5919 68.5181
R12051 vss.n5927 vss.n5917 68.5181
R12052 vss.n5956 vss.n5917 68.5181
R12053 vss.n5580 vss.n5572 68.5181
R12054 vss.n5572 vss.n5543 68.5181
R12055 vss.n5570 vss.n5541 68.5181
R12056 vss.n5586 vss.n5541 68.5181
R12057 vss.n5561 vss.n5551 68.5181
R12058 vss.n5562 vss.n5561 68.5181
R12059 vss.n5697 vss.n5692 68.5181
R12060 vss.n5706 vss.n5697 68.5181
R12061 vss.n5712 vss.n5691 68.5181
R12062 vss.n5691 vss.n5681 68.5181
R12063 vss.n5689 vss.n5540 68.5181
R12064 vss.n5718 vss.n5540 68.5181
R12065 vss.n3558 vss.n3553 68.5181
R12066 vss.n6316 vss.n3558 68.5181
R12067 vss.n6322 vss.n3552 68.5181
R12068 vss.n3552 vss.n3542 68.5181
R12069 vss.n3550 vss.n3540 68.5181
R12070 vss.n6328 vss.n3540 68.5181
R12071 vss.n5625 vss.n5617 68.5181
R12072 vss.n5617 vss.n5590 68.5181
R12073 vss.n5615 vss.n5588 68.5181
R12074 vss.n5631 vss.n5588 68.5181
R12075 vss.n5606 vss.n5598 68.5181
R12076 vss.n5607 vss.n5606 68.5181
R12077 vss.n5889 vss.n5884 68.5181
R12078 vss.n5897 vss.n5889 68.5181
R12079 vss.n5903 vss.n5883 68.5181
R12080 vss.n5883 vss.n5872 68.5181
R12081 vss.n5881 vss.n5728 68.5181
R12082 vss.n5909 vss.n5728 68.5181
R12083 vss.n6128 vss.n6123 68.5181
R12084 vss.n6136 vss.n6128 68.5181
R12085 vss.n6142 vss.n6122 68.5181
R12086 vss.n6122 vss.n6111 68.5181
R12087 vss.n6120 vss.n5968 68.5181
R12088 vss.n6148 vss.n5968 68.5181
R12089 vss.n6008 vss.n6000 68.5181
R12090 vss.n6000 vss.n5971 68.5181
R12091 vss.n5998 vss.n5969 68.5181
R12092 vss.n6014 vss.n5969 68.5181
R12093 vss.n5989 vss.n5979 68.5181
R12094 vss.n5990 vss.n5989 68.5181
R12095 vss.n6738 vss.n3274 68.5181
R12096 vss.n3302 vss.n3274 68.5181
R12097 vss.n4387 vss.n4382 68.5181
R12098 vss.n4395 vss.n4387 68.5181
R12099 vss.n4543 vss.n4381 68.5181
R12100 vss.n4381 vss.n4371 68.5181
R12101 vss.n4379 vss.n4370 68.5181
R12102 vss.n4549 vss.n4370 68.5181
R12103 vss.n4431 vss.n4403 68.5181
R12104 vss.n4439 vss.n4431 68.5181
R12105 vss.n4445 vss.n4401 68.5181
R12106 vss.n4429 vss.n4401 68.5181
R12107 vss.n4463 vss.n4462 68.5181
R12108 vss.n4462 vss.n4457 68.5181
R12109 vss.n4492 vss.n4447 68.5181
R12110 vss.n4475 vss.n4447 68.5181
R12111 vss.n4477 vss.n4449 68.5181
R12112 vss.n4486 vss.n4477 68.5181
R12113 vss.n4510 vss.n4509 68.5181
R12114 vss.n4509 vss.n4504 68.5181
R12115 vss.n4539 vss.n4494 68.5181
R12116 vss.n4523 vss.n4494 68.5181
R12117 vss.n4525 vss.n4496 68.5181
R12118 vss.n4533 vss.n4525 68.5181
R12119 vss.n6645 vss.n6617 68.5181
R12120 vss.n6653 vss.n6645 68.5181
R12121 vss.n6659 vss.n6615 68.5181
R12122 vss.n6643 vss.n6615 68.5181
R12123 vss.n6631 vss.n6630 68.5181
R12124 vss.n6630 vss.n6625 68.5181
R12125 vss.n6596 vss.n6499 68.5181
R12126 vss.n6605 vss.n6596 68.5181
R12127 vss.n6611 vss.n6497 68.5181
R12128 vss.n6594 vss.n6497 68.5181
R12129 vss.n6513 vss.n6512 68.5181
R12130 vss.n6512 vss.n6507 68.5181
R12131 vss.n5243 vss.n5215 68.5181
R12132 vss.n5251 vss.n5243 68.5181
R12133 vss.n5257 vss.n5213 68.5181
R12134 vss.n5241 vss.n5213 68.5181
R12135 vss.n5229 vss.n5228 68.5181
R12136 vss.n5228 vss.n5223 68.5181
R12137 vss.n5274 vss.n5273 68.5181
R12138 vss.n5273 vss.n5268 68.5181
R12139 vss.n5304 vss.n5258 68.5181
R12140 vss.n5287 vss.n5258 68.5181
R12141 vss.n5289 vss.n5260 68.5181
R12142 vss.n5298 vss.n5289 68.5181
R12143 vss.n4023 vss.n4018 68.5181
R12144 vss.n4031 vss.n4023 68.5181
R12145 vss.n5521 vss.n4017 68.5181
R12146 vss.n4032 vss.n4017 68.5181
R12147 vss.n4010 vss.n4008 68.5181
R12148 vss.n4010 vss.n4009 68.5181
R12149 vss.n5489 vss.n5488 68.5181
R12150 vss.n5488 vss.n5483 68.5181
R12151 vss.n5518 vss.n5473 68.5181
R12152 vss.n5502 vss.n5473 68.5181
R12153 vss.n5504 vss.n5475 68.5181
R12154 vss.n5512 vss.n5504 68.5181
R12155 vss.n4054 vss.n4053 68.5181
R12156 vss.n4053 vss.n4048 68.5181
R12157 vss.n4081 vss.n4038 68.5181
R12158 vss.n4066 vss.n4038 68.5181
R12159 vss.n4068 vss.n4040 68.5181
R12160 vss.n4075 vss.n4068 68.5181
R12161 vss.n5455 vss.n5427 68.5181
R12162 vss.n5463 vss.n5455 68.5181
R12163 vss.n5469 vss.n5425 68.5181
R12164 vss.n5453 vss.n5425 68.5181
R12165 vss.n5441 vss.n5440 68.5181
R12166 vss.n5440 vss.n5435 68.5181
R12167 vss.n5408 vss.n5312 68.5181
R12168 vss.n5416 vss.n5408 68.5181
R12169 vss.n5422 vss.n5310 68.5181
R12170 vss.n5406 vss.n5310 68.5181
R12171 vss.n5326 vss.n5325 68.5181
R12172 vss.n5325 vss.n5320 68.5181
R12173 vss.n4158 vss.n4130 68.5181
R12174 vss.n4166 vss.n4158 68.5181
R12175 vss.n4172 vss.n4128 68.5181
R12176 vss.n4156 vss.n4128 68.5181
R12177 vss.n4144 vss.n4143 68.5181
R12178 vss.n4143 vss.n4138 68.5181
R12179 vss.n5063 vss.n5062 68.5181
R12180 vss.n5062 vss.n5057 68.5181
R12181 vss.n5092 vss.n5047 68.5181
R12182 vss.n5076 vss.n5047 68.5181
R12183 vss.n5078 vss.n5049 68.5181
R12184 vss.n5086 vss.n5078 68.5181
R12185 vss.n4188 vss.n4187 68.5181
R12186 vss.n4187 vss.n4182 68.5181
R12187 vss.n4218 vss.n4173 68.5181
R12188 vss.n4203 vss.n4173 68.5181
R12189 vss.n4216 vss.n4176 68.5181
R12190 vss.n4205 vss.n4176 68.5181
R12191 vss.n5015 vss.n5014 68.5181
R12192 vss.n5014 vss.n5009 68.5181
R12193 vss.n5044 vss.n4999 68.5181
R12194 vss.n5028 vss.n4999 68.5181
R12195 vss.n5030 vss.n5001 68.5181
R12196 vss.n5038 vss.n5030 68.5181
R12197 vss.n4235 vss.n4234 68.5181
R12198 vss.n4234 vss.n4229 68.5181
R12199 vss.n4262 vss.n4219 68.5181
R12200 vss.n4247 vss.n4219 68.5181
R12201 vss.n4249 vss.n4221 68.5181
R12202 vss.n4256 vss.n4249 68.5181
R12203 vss.n4981 vss.n4953 68.5181
R12204 vss.n4989 vss.n4981 68.5181
R12205 vss.n4995 vss.n4951 68.5181
R12206 vss.n4979 vss.n4951 68.5181
R12207 vss.n4967 vss.n4966 68.5181
R12208 vss.n4966 vss.n4961 68.5181
R12209 vss.n4112 vss.n4084 68.5181
R12210 vss.n4120 vss.n4112 68.5181
R12211 vss.n4126 vss.n4082 68.5181
R12212 vss.n4110 vss.n4082 68.5181
R12213 vss.n4098 vss.n4097 68.5181
R12214 vss.n4097 vss.n4092 68.5181
R12215 vss.n4933 vss.n4267 68.5181
R12216 vss.n4941 vss.n4933 68.5181
R12217 vss.n4947 vss.n4265 68.5181
R12218 vss.n4931 vss.n4265 68.5181
R12219 vss.n4281 vss.n4280 68.5181
R12220 vss.n4280 vss.n4275 68.5181
R12221 vss.n5196 vss.n5100 68.5181
R12222 vss.n5204 vss.n5196 68.5181
R12223 vss.n5210 vss.n5098 68.5181
R12224 vss.n5194 vss.n5098 68.5181
R12225 vss.n5114 vss.n5113 68.5181
R12226 vss.n5113 vss.n5108 68.5181
R12227 vss.n3371 vss.n3343 68.5181
R12228 vss.n3379 vss.n3371 68.5181
R12229 vss.n3385 vss.n3341 68.5181
R12230 vss.n3369 vss.n3341 68.5181
R12231 vss.n3357 vss.n3356 68.5181
R12232 vss.n3356 vss.n3351 68.5181
R12233 vss.n3418 vss.n3390 68.5181
R12234 vss.n3426 vss.n3418 68.5181
R12235 vss.n3432 vss.n3388 68.5181
R12236 vss.n3416 vss.n3388 68.5181
R12237 vss.n3404 vss.n3403 68.5181
R12238 vss.n3403 vss.n3398 68.5181
R12239 vss.n3460 vss.n3457 68.5181
R12240 vss.n3467 vss.n3457 68.5181
R12241 vss.n3450 vss.n3433 68.5181
R12242 vss.n3450 vss.n3446 68.5181
R12243 vss.n3473 vss.n3445 68.5181
R12244 vss.n3482 vss.n3445 68.5181
R12245 vss.n6348 vss.n6347 68.5181
R12246 vss.n6351 vss.n6348 68.5181
R12247 vss.n6374 vss.n3434 68.5181
R12248 vss.n6338 vss.n3434 68.5181
R12249 vss.n6372 vss.n3437 68.5181
R12250 vss.n6364 vss.n3437 68.5181
R12251 vss.n3505 vss.n3500 68.5181
R12252 vss.n3513 vss.n3505 68.5181
R12253 vss.n3519 vss.n3499 68.5181
R12254 vss.n3499 vss.n3493 68.5181
R12255 vss.n3520 vss.n3492 68.5181
R12256 vss.n3530 vss.n3492 68.5181
R12257 vss.n6480 vss.n6384 68.5181
R12258 vss.n6488 vss.n6480 68.5181
R12259 vss.n6494 vss.n6382 68.5181
R12260 vss.n6478 vss.n6382 68.5181
R12261 vss.n6398 vss.n6397 68.5181
R12262 vss.n6397 vss.n6392 68.5181
R12263 vss.n6699 vss.n3340 68.5181
R12264 vss.n6671 vss.n3340 68.5181
R12265 vss.n6673 vss.n6663 68.5181
R12266 vss.n6693 vss.n6673 68.5181
R12267 vss.n6687 vss.n6686 68.5181
R12268 vss.n6687 vss.n6674 68.5181
R12269 vss.n4417 vss.n4416 68.5181
R12270 vss.n4416 vss.n4411 68.5181
R12271 vss.n4774 vss.n4769 68.5181
R12272 vss.n4782 vss.n4774 68.5181
R12273 vss.n4789 vss.n4768 68.5181
R12274 vss.n4768 vss.n4758 68.5181
R12275 vss.n4766 vss.n4757 68.5181
R12276 vss.n4795 vss.n4757 68.5181
R12277 vss.n3304 vss.n3276 68.5181
R12278 vss.n6732 vss.n3304 68.5181
R12279 vss.n3290 vss.n3289 68.5181
R12280 vss.n3289 vss.n3284 68.5181
R12281 vss.n15531 vss.n387 68.5181
R12282 vss.n15537 vss.n387 68.5181
R12283 vss.n15530 vss.n15510 68.5181
R12284 vss.n15510 vss.n15501 68.5181
R12285 vss.n15516 vss.n15511 68.5181
R12286 vss.n15524 vss.n15516 68.5181
R12287 vss.n15492 vss.n401 68.5181
R12288 vss.n401 vss.n391 68.5181
R12289 vss.n399 vss.n389 68.5181
R12290 vss.n15498 vss.n389 68.5181
R12291 vss.n14863 vss.n14854 68.5181
R12292 vss.n14864 vss.n14863 68.5181
R12293 vss.n15002 vss.n14999 68.5181
R12294 vss.n14999 vss.n14980 68.5181
R12295 vss.n15000 vss.n14978 68.5181
R12296 vss.n15018 vss.n14978 68.5181
R12297 vss.n15011 vss.n14989 68.5181
R12298 vss.n15012 vss.n15011 68.5181
R12299 vss.n15042 vss.n1071 68.5181
R12300 vss.n1071 vss.n1043 68.5181
R12301 vss.n1069 vss.n1041 68.5181
R12302 vss.n15048 vss.n1041 68.5181
R12303 vss.n1056 vss.n1051 68.5181
R12304 vss.n1057 vss.n1056 68.5181
R12305 vss.n15067 vss.n15062 68.5181
R12306 vss.n15076 vss.n15067 68.5181
R12307 vss.n15082 vss.n15061 68.5181
R12308 vss.n15061 vss.n15052 68.5181
R12309 vss.n1011 vss.n1006 68.5181
R12310 vss.n1019 vss.n1011 68.5181
R12311 vss.n14928 vss.n14920 68.5181
R12312 vss.n14920 vss.n14890 68.5181
R12313 vss.n14918 vss.n14888 68.5181
R12314 vss.n14934 vss.n14888 68.5181
R12315 vss.n14903 vss.n14898 68.5181
R12316 vss.n14904 vss.n14903 68.5181
R12317 vss.n15436 vss.n533 68.5181
R12318 vss.n533 vss.n505 68.5181
R12319 vss.n531 vss.n503 68.5181
R12320 vss.n15442 vss.n503 68.5181
R12321 vss.n518 vss.n513 68.5181
R12322 vss.n519 vss.n518 68.5181
R12323 vss.n7339 vss.n7331 68.5181
R12324 vss.n7331 vss.n7303 68.5181
R12325 vss.n7329 vss.n7301 68.5181
R12326 vss.n7345 vss.n7301 68.5181
R12327 vss.n7316 vss.n7311 68.5181
R12328 vss.n7317 vss.n7316 68.5181
R12329 vss.n7293 vss.n7284 68.5181
R12330 vss.n7284 vss.n3112 68.5181
R12331 vss.n7282 vss.n3110 68.5181
R12332 vss.n7299 vss.n3110 68.5181
R12333 vss.n7367 vss.n7362 68.5181
R12334 vss.n7376 vss.n7367 68.5181
R12335 vss.n7382 vss.n7361 68.5181
R12336 vss.n7361 vss.n7351 68.5181
R12337 vss.n7359 vss.n3063 68.5181
R12338 vss.n7388 vss.n3063 68.5181
R12339 vss.n3103 vss.n3095 68.5181
R12340 vss.n3095 vss.n3066 68.5181
R12341 vss.n3093 vss.n3064 68.5181
R12342 vss.n3109 vss.n3064 68.5181
R12343 vss.n3084 vss.n3074 68.5181
R12344 vss.n3085 vss.n3084 68.5181
R12345 vss.n15363 vss.n738 68.5181
R12346 vss.n738 vss.n710 68.5181
R12347 vss.n736 vss.n708 68.5181
R12348 vss.n15369 vss.n708 68.5181
R12349 vss.n723 vss.n718 68.5181
R12350 vss.n724 vss.n723 68.5181
R12351 vss.n15286 vss.n791 68.5181
R12352 vss.n791 vss.n763 68.5181
R12353 vss.n789 vss.n761 68.5181
R12354 vss.n15292 vss.n761 68.5181
R12355 vss.n776 vss.n771 68.5181
R12356 vss.n777 vss.n776 68.5181
R12357 vss.n7462 vss.n7457 68.5181
R12358 vss.n7471 vss.n7462 68.5181
R12359 vss.n7477 vss.n7456 68.5181
R12360 vss.n7456 vss.n7447 68.5181
R12361 vss.n15165 vss.n15156 68.5181
R12362 vss.n15156 vss.n968 68.5181
R12363 vss.n15154 vss.n966 68.5181
R12364 vss.n15171 vss.n966 68.5181
R12365 vss.n981 vss.n976 68.5181
R12366 vss.n982 vss.n981 68.5181
R12367 vss.n15213 vss.n15205 68.5181
R12368 vss.n15205 vss.n15177 68.5181
R12369 vss.n15203 vss.n15175 68.5181
R12370 vss.n15219 vss.n15175 68.5181
R12371 vss.n15190 vss.n15185 68.5181
R12372 vss.n15191 vss.n15190 68.5181
R12373 vss.n957 vss.n948 68.5181
R12374 vss.n948 vss.n920 68.5181
R12375 vss.n946 vss.n918 68.5181
R12376 vss.n963 vss.n918 68.5181
R12377 vss.n933 vss.n928 68.5181
R12378 vss.n934 vss.n933 68.5181
R12379 vss.n840 vss.n809 68.5181
R12380 vss.n846 vss.n809 68.5181
R12381 vss.n839 vss.n819 68.5181
R12382 vss.n819 vss.n810 68.5181
R12383 vss.n825 vss.n820 68.5181
R12384 vss.n833 vss.n825 68.5181
R12385 vss.n15118 vss.n15113 68.5181
R12386 vss.n15126 vss.n15118 68.5181
R12387 vss.n15132 vss.n15112 68.5181
R12388 vss.n15112 vss.n15100 68.5181
R12389 vss.n15110 vss.n15099 68.5181
R12390 vss.n15138 vss.n15099 68.5181
R12391 vss.n7454 vss.n7445 68.5181
R12392 vss.n7483 vss.n7445 68.5181
R12393 vss.n15334 vss.n15325 68.5181
R12394 vss.n15325 vss.n15297 68.5181
R12395 vss.n15323 vss.n15295 68.5181
R12396 vss.n15340 vss.n15295 68.5181
R12397 vss.n15310 vss.n15305 68.5181
R12398 vss.n15311 vss.n15310 68.5181
R12399 vss.n700 vss.n691 68.5181
R12400 vss.n691 vss.n663 68.5181
R12401 vss.n689 vss.n661 68.5181
R12402 vss.n706 vss.n661 68.5181
R12403 vss.n676 vss.n671 68.5181
R12404 vss.n677 vss.n676 68.5181
R12405 vss.n7416 vss.n7411 68.5181
R12406 vss.n7424 vss.n7416 68.5181
R12407 vss.n7430 vss.n7410 68.5181
R12408 vss.n7410 vss.n7399 68.5181
R12409 vss.n7408 vss.n7398 68.5181
R12410 vss.n7436 vss.n7398 68.5181
R12411 vss.n3125 vss.n3120 68.5181
R12412 vss.n3126 vss.n3125 68.5181
R12413 vss.n583 vss.n551 68.5181
R12414 vss.n589 vss.n551 68.5181
R12415 vss.n582 vss.n562 68.5181
R12416 vss.n562 vss.n553 68.5181
R12417 vss.n568 vss.n563 68.5181
R12418 vss.n576 vss.n568 68.5181
R12419 vss.n492 vss.n483 68.5181
R12420 vss.n483 vss.n455 68.5181
R12421 vss.n481 vss.n453 68.5181
R12422 vss.n498 vss.n453 68.5181
R12423 vss.n468 vss.n463 68.5181
R12424 vss.n469 vss.n468 68.5181
R12425 vss.n4734 vss.n4558 68.5181
R12426 vss.n4740 vss.n4558 68.5181
R12427 vss.n4733 vss.n4713 68.5181
R12428 vss.n4713 vss.n4704 68.5181
R12429 vss.n4719 vss.n4714 68.5181
R12430 vss.n4727 vss.n4719 68.5181
R12431 vss.n4694 vss.n4686 68.5181
R12432 vss.n4686 vss.n4657 68.5181
R12433 vss.n4684 vss.n4655 68.5181
R12434 vss.n4700 vss.n4655 68.5181
R12435 vss.n4675 vss.n4665 68.5181
R12436 vss.n4676 vss.n4675 68.5181
R12437 vss.n4646 vss.n4637 68.5181
R12438 vss.n4637 vss.n4609 68.5181
R12439 vss.n4635 vss.n4607 68.5181
R12440 vss.n4652 vss.n4607 68.5181
R12441 vss.n4622 vss.n4617 68.5181
R12442 vss.n4623 vss.n4622 68.5181
R12443 vss.n4599 vss.n4590 68.5181
R12444 vss.n4590 vss.n4561 68.5181
R12445 vss.n4588 vss.n4559 68.5181
R12446 vss.n4605 vss.n4559 68.5181
R12447 vss.n4574 vss.n4569 68.5181
R12448 vss.n4575 vss.n4574 68.5181
R12449 vss.n4349 vss.n4318 68.5181
R12450 vss.n4355 vss.n4318 68.5181
R12451 vss.n4348 vss.n4328 68.5181
R12452 vss.n4328 vss.n4319 68.5181
R12453 vss.n4334 vss.n4329 68.5181
R12454 vss.n4342 vss.n4334 68.5181
R12455 vss.n7246 vss.n7241 68.5181
R12456 vss.n7254 vss.n7246 68.5181
R12457 vss.n7260 vss.n7240 68.5181
R12458 vss.n7240 vss.n7229 68.5181
R12459 vss.n7238 vss.n7228 68.5181
R12460 vss.n7266 vss.n7228 68.5181
R12461 vss.n6861 vss.n6833 68.5181
R12462 vss.n6869 vss.n6861 68.5181
R12463 vss.n6875 vss.n6831 68.5181
R12464 vss.n6859 vss.n6831 68.5181
R12465 vss.n6847 vss.n6846 68.5181
R12466 vss.n6846 vss.n6841 68.5181
R12467 vss.n7191 vss.n3152 68.5181
R12468 vss.n7199 vss.n7191 68.5181
R12469 vss.n7205 vss.n3150 68.5181
R12470 vss.n7189 vss.n3150 68.5181
R12471 vss.n6810 vss.n6809 68.5181
R12472 vss.n6820 vss.n6810 68.5181
R12473 vss.n7208 vss.n3147 68.5181
R12474 vss.n6811 vss.n3147 68.5181
R12475 vss.n3140 vss.n3138 68.5181
R12476 vss.n3140 vss.n3139 68.5181
R12477 vss.n6915 vss.n6830 68.5181
R12478 vss.n6887 vss.n6830 68.5181
R12479 vss.n6889 vss.n6879 68.5181
R12480 vss.n6909 vss.n6889 68.5181
R12481 vss.n6903 vss.n6902 68.5181
R12482 vss.n6903 vss.n6890 68.5181
R12483 vss.n2632 vss.n2602 68.5181
R12484 vss.n2638 vss.n2602 68.5181
R12485 vss.n2608 vss.n1140 68.5181
R12486 vss.n2608 vss.n2603 68.5181
R12487 vss.n2618 vss.n2615 68.5181
R12488 vss.n2624 vss.n2615 68.5181
R12489 vss.n1918 vss.n1913 68.5181
R12490 vss.n1927 vss.n1918 68.5181
R12491 vss.n1934 vss.n1912 68.5181
R12492 vss.n1912 vss.n1902 68.5181
R12493 vss.n1910 vss.n1901 68.5181
R12494 vss.n1940 vss.n1901 68.5181
R12495 vss.n2868 vss.n2840 68.5181
R12496 vss.n2876 vss.n2868 68.5181
R12497 vss.n2882 vss.n2838 68.5181
R12498 vss.n2866 vss.n2838 68.5181
R12499 vss.n2854 vss.n2853 68.5181
R12500 vss.n2853 vss.n2848 68.5181
R12501 vss.n7735 vss.n7734 68.5181
R12502 vss.n7734 vss.n7729 68.5181
R12503 vss.n7764 vss.n7719 68.5181
R12504 vss.n7748 vss.n7719 68.5181
R12505 vss.n7750 vss.n7721 68.5181
R12506 vss.n7758 vss.n7750 68.5181
R12507 vss.n2903 vss.n2902 68.5181
R12508 vss.n2906 vss.n2903 68.5181
R12509 vss.n2929 vss.n2883 68.5181
R12510 vss.n2893 vss.n2883 68.5181
R12511 vss.n2927 vss.n2886 68.5181
R12512 vss.n2919 vss.n2886 68.5181
R12513 vss.n7686 vss.n7685 68.5181
R12514 vss.n7685 vss.n7680 68.5181
R12515 vss.n7716 vss.n7670 68.5181
R12516 vss.n7699 vss.n7670 68.5181
R12517 vss.n7701 vss.n7672 68.5181
R12518 vss.n7710 vss.n7701 68.5181
R12519 vss.n3029 vss.n3024 68.5181
R12520 vss.n3037 vss.n3029 68.5181
R12521 vss.n3043 vss.n3023 68.5181
R12522 vss.n3023 vss.n3017 68.5181
R12523 vss.n3044 vss.n3016 68.5181
R12524 vss.n3054 vss.n3016 68.5181
R12525 vss.n7652 vss.n7624 68.5181
R12526 vss.n7660 vss.n7652 68.5181
R12527 vss.n7666 vss.n7622 68.5181
R12528 vss.n7650 vss.n7622 68.5181
R12529 vss.n7638 vss.n7637 68.5181
R12530 vss.n7637 vss.n7632 68.5181
R12531 vss.n2822 vss.n2726 68.5181
R12532 vss.n2830 vss.n2822 68.5181
R12533 vss.n2836 vss.n2724 68.5181
R12534 vss.n2820 vss.n2724 68.5181
R12535 vss.n2740 vss.n2739 68.5181
R12536 vss.n2739 vss.n2734 68.5181
R12537 vss.n2960 vss.n2932 68.5181
R12538 vss.n2969 vss.n2960 68.5181
R12539 vss.n2975 vss.n2930 68.5181
R12540 vss.n2958 vss.n2930 68.5181
R12541 vss.n2946 vss.n2945 68.5181
R12542 vss.n2945 vss.n2940 68.5181
R12543 vss.n2992 vss.n2991 68.5181
R12544 vss.n2991 vss.n2986 68.5181
R12545 vss.n7500 vss.n2976 68.5181
R12546 vss.n3005 vss.n2976 68.5181
R12547 vss.n3007 vss.n2978 68.5181
R12548 vss.n7494 vss.n3007 68.5181
R12549 vss.n7964 vss.n7963 68.5181
R12550 vss.n7967 vss.n7964 68.5181
R12551 vss.n7990 vss.n2452 68.5181
R12552 vss.n2463 vss.n2452 68.5181
R12553 vss.n7988 vss.n2455 68.5181
R12554 vss.n7980 vss.n2455 68.5181
R12555 vss.n7119 vss.n7082 68.5181
R12556 vss.n7090 vss.n7082 68.5181
R12557 vss.n7092 vss.n2451 68.5181
R12558 vss.n7113 vss.n7092 68.5181
R12559 vss.n7107 vss.n7106 68.5181
R12560 vss.n7107 vss.n7093 68.5181
R12561 vss.n7046 vss.n7036 68.5181
R12562 vss.n7072 vss.n7036 68.5181
R12563 vss.n7066 vss.n7065 68.5181
R12564 vss.n7066 vss.n7037 68.5181
R12565 vss.n7051 vss.n7048 68.5181
R12566 vss.n7054 vss.n7051 68.5181
R12567 vss.n7021 vss.n6991 68.5181
R12568 vss.n7027 vss.n6991 68.5181
R12569 vss.n6997 vss.n2450 68.5181
R12570 vss.n6997 vss.n6992 68.5181
R12571 vss.n7007 vss.n7004 68.5181
R12572 vss.n7013 vss.n7004 68.5181
R12573 vss.n7159 vss.n7128 68.5181
R12574 vss.n7165 vss.n7128 68.5181
R12575 vss.n7158 vss.n7138 68.5181
R12576 vss.n7138 vss.n7129 68.5181
R12577 vss.n7144 vss.n7139 68.5181
R12578 vss.n7152 vss.n7144 68.5181
R12579 vss.n6976 vss.n6924 68.5181
R12580 vss.n6982 vss.n6924 68.5181
R12581 vss.n6975 vss.n6934 68.5181
R12582 vss.n6934 vss.n6925 68.5181
R12583 vss.n6940 vss.n6935 68.5181
R12584 vss.n6968 vss.n6940 68.5181
R12585 vss.n7604 vss.n7508 68.5181
R12586 vss.n7612 vss.n7604 68.5181
R12587 vss.n7618 vss.n7506 68.5181
R12588 vss.n7602 vss.n7506 68.5181
R12589 vss.n7522 vss.n7521 68.5181
R12590 vss.n7521 vss.n7516 68.5181
R12591 vss.n7799 vss.n7771 68.5181
R12592 vss.n7807 vss.n7799 68.5181
R12593 vss.n7813 vss.n7769 68.5181
R12594 vss.n7797 vss.n7769 68.5181
R12595 vss.n7785 vss.n7784 68.5181
R12596 vss.n7784 vss.n7779 68.5181
R12597 vss.n7847 vss.n7819 68.5181
R12598 vss.n7855 vss.n7847 68.5181
R12599 vss.n7861 vss.n7817 68.5181
R12600 vss.n7845 vss.n7817 68.5181
R12601 vss.n7833 vss.n7832 68.5181
R12602 vss.n7832 vss.n7827 68.5181
R12603 vss.n7881 vss.n7880 68.5181
R12604 vss.n7880 vss.n7875 68.5181
R12605 vss.n7911 vss.n7865 68.5181
R12606 vss.n7894 vss.n7865 68.5181
R12607 vss.n7896 vss.n7867 68.5181
R12608 vss.n7905 vss.n7896 68.5181
R12609 vss.n2657 vss.n2647 68.5181
R12610 vss.n7921 vss.n2647 68.5181
R12611 vss.n7915 vss.n7914 68.5181
R12612 vss.n7915 vss.n2648 68.5181
R12613 vss.n2677 vss.n2660 68.5181
R12614 vss.n2669 vss.n2660 68.5181
R12615 vss.n2695 vss.n2694 68.5181
R12616 vss.n2694 vss.n2689 68.5181
R12617 vss.n2722 vss.n2679 68.5181
R12618 vss.n2707 vss.n2679 68.5181
R12619 vss.n2709 vss.n2681 68.5181
R12620 vss.n2716 vss.n2709 68.5181
R12621 vss.n2587 vss.n2487 68.5181
R12622 vss.n2593 vss.n2487 68.5181
R12623 vss.n2586 vss.n2497 68.5181
R12624 vss.n2497 vss.n2488 68.5181
R12625 vss.n2503 vss.n2498 68.5181
R12626 vss.n2580 vss.n2503 68.5181
R12627 vss.n7941 vss.n7940 68.5181
R12628 vss.n7940 vss.n7931 68.5181
R12629 vss.n14881 vss.n1141 68.5181
R12630 vss.n1151 vss.n1141 68.5181
R12631 vss.n1153 vss.n1143 68.5181
R12632 vss.n14875 vss.n1153 68.5181
R12633 vss.n3166 vss.n3165 68.5181
R12634 vss.n3165 vss.n3160 68.5181
R12635 vss.n6793 vss.n3173 68.5181
R12636 vss.n6799 vss.n3173 68.5181
R12637 vss.n6792 vss.n3183 68.5181
R12638 vss.n3183 vss.n3174 68.5181
R12639 vss.n3196 vss.n3195 68.5181
R12640 vss.n3205 vss.n3196 68.5181
R12641 vss.n6761 vss.n6760 68.5181
R12642 vss.n6760 vss.n6755 68.5181
R12643 vss.n6789 vss.n6745 68.5181
R12644 vss.n6773 vss.n6745 68.5181
R12645 vss.n6775 vss.n6747 68.5181
R12646 vss.n6783 vss.n6775 68.5181
R12647 vss.n14836 vss.n1166 68.5181
R12648 vss.n14842 vss.n1166 68.5181
R12649 vss.n14835 vss.n14815 68.5181
R12650 vss.n14815 vss.n14806 68.5181
R12651 vss.n14821 vss.n14816 68.5181
R12652 vss.n14829 vss.n14821 68.5181
R12653 vss.n14797 vss.n1180 68.5181
R12654 vss.n1180 vss.n1170 68.5181
R12655 vss.n1178 vss.n1168 68.5181
R12656 vss.n14803 vss.n1168 68.5181
R12657 vss.n14169 vss.n14160 68.5181
R12658 vss.n14170 vss.n14169 68.5181
R12659 vss.n14307 vss.n14304 68.5181
R12660 vss.n14304 vss.n14285 68.5181
R12661 vss.n14305 vss.n14283 68.5181
R12662 vss.n14323 vss.n14283 68.5181
R12663 vss.n14316 vss.n14294 68.5181
R12664 vss.n14317 vss.n14316 68.5181
R12665 vss.n14347 vss.n1850 68.5181
R12666 vss.n1850 vss.n1822 68.5181
R12667 vss.n1848 vss.n1820 68.5181
R12668 vss.n14353 vss.n1820 68.5181
R12669 vss.n1835 vss.n1830 68.5181
R12670 vss.n1836 vss.n1835 68.5181
R12671 vss.n14372 vss.n14367 68.5181
R12672 vss.n14381 vss.n14372 68.5181
R12673 vss.n14387 vss.n14366 68.5181
R12674 vss.n14366 vss.n14357 68.5181
R12675 vss.n1790 vss.n1785 68.5181
R12676 vss.n1798 vss.n1790 68.5181
R12677 vss.n14233 vss.n14225 68.5181
R12678 vss.n14225 vss.n14195 68.5181
R12679 vss.n14223 vss.n14193 68.5181
R12680 vss.n14239 vss.n14193 68.5181
R12681 vss.n14208 vss.n14203 68.5181
R12682 vss.n14209 vss.n14208 68.5181
R12683 vss.n14741 vss.n1312 68.5181
R12684 vss.n1312 vss.n1284 68.5181
R12685 vss.n1310 vss.n1282 68.5181
R12686 vss.n14747 vss.n1282 68.5181
R12687 vss.n1297 vss.n1292 68.5181
R12688 vss.n1298 vss.n1297 68.5181
R12689 vss.n14019 vss.n14011 68.5181
R12690 vss.n14011 vss.n13983 68.5181
R12691 vss.n14009 vss.n13981 68.5181
R12692 vss.n14025 vss.n13981 68.5181
R12693 vss.n13996 vss.n13991 68.5181
R12694 vss.n13997 vss.n13996 68.5181
R12695 vss.n14044 vss.n14039 68.5181
R12696 vss.n14053 vss.n14044 68.5181
R12697 vss.n14059 vss.n14038 68.5181
R12698 vss.n14038 vss.n14029 68.5181
R12699 vss.n8196 vss.n8191 68.5181
R12700 vss.n8205 vss.n8196 68.5181
R12701 vss.n8211 vss.n8190 68.5181
R12702 vss.n8190 vss.n8180 68.5181
R12703 vss.n8188 vss.n8179 68.5181
R12704 vss.n8217 vss.n8179 68.5181
R12705 vss.n13973 vss.n13965 68.5181
R12706 vss.n13965 vss.n8154 68.5181
R12707 vss.n13963 vss.n8152 68.5181
R12708 vss.n13979 vss.n8152 68.5181
R12709 vss.n8167 vss.n8162 68.5181
R12710 vss.n8168 vss.n8167 68.5181
R12711 vss.n14668 vss.n1517 68.5181
R12712 vss.n1517 vss.n1489 68.5181
R12713 vss.n1515 vss.n1487 68.5181
R12714 vss.n14674 vss.n1487 68.5181
R12715 vss.n1502 vss.n1497 68.5181
R12716 vss.n1503 vss.n1502 68.5181
R12717 vss.n14591 vss.n1570 68.5181
R12718 vss.n1570 vss.n1542 68.5181
R12719 vss.n1568 vss.n1540 68.5181
R12720 vss.n14597 vss.n1540 68.5181
R12721 vss.n1555 vss.n1550 68.5181
R12722 vss.n1556 vss.n1555 68.5181
R12723 vss.n13927 vss.n13922 68.5181
R12724 vss.n13936 vss.n13927 68.5181
R12725 vss.n13942 vss.n13921 68.5181
R12726 vss.n13921 vss.n13912 68.5181
R12727 vss.n14470 vss.n14461 68.5181
R12728 vss.n14461 vss.n1747 68.5181
R12729 vss.n14459 vss.n1745 68.5181
R12730 vss.n14476 vss.n1745 68.5181
R12731 vss.n1760 vss.n1755 68.5181
R12732 vss.n1761 vss.n1760 68.5181
R12733 vss.n14518 vss.n14510 68.5181
R12734 vss.n14510 vss.n14482 68.5181
R12735 vss.n14508 vss.n14480 68.5181
R12736 vss.n14524 vss.n14480 68.5181
R12737 vss.n14495 vss.n14490 68.5181
R12738 vss.n14496 vss.n14495 68.5181
R12739 vss.n1736 vss.n1727 68.5181
R12740 vss.n1727 vss.n1699 68.5181
R12741 vss.n1725 vss.n1697 68.5181
R12742 vss.n1742 vss.n1697 68.5181
R12743 vss.n1712 vss.n1707 68.5181
R12744 vss.n1713 vss.n1712 68.5181
R12745 vss.n1619 vss.n1588 68.5181
R12746 vss.n1625 vss.n1588 68.5181
R12747 vss.n1618 vss.n1598 68.5181
R12748 vss.n1598 vss.n1589 68.5181
R12749 vss.n1604 vss.n1599 68.5181
R12750 vss.n1612 vss.n1604 68.5181
R12751 vss.n14423 vss.n14418 68.5181
R12752 vss.n14431 vss.n14423 68.5181
R12753 vss.n14437 vss.n14417 68.5181
R12754 vss.n14417 vss.n14405 68.5181
R12755 vss.n14415 vss.n14404 68.5181
R12756 vss.n14443 vss.n14404 68.5181
R12757 vss.n13919 vss.n13910 68.5181
R12758 vss.n13948 vss.n13910 68.5181
R12759 vss.n14639 vss.n14630 68.5181
R12760 vss.n14630 vss.n14602 68.5181
R12761 vss.n14628 vss.n14600 68.5181
R12762 vss.n14645 vss.n14600 68.5181
R12763 vss.n14615 vss.n14610 68.5181
R12764 vss.n14616 vss.n14615 68.5181
R12765 vss.n1479 vss.n1470 68.5181
R12766 vss.n1470 vss.n1442 68.5181
R12767 vss.n1468 vss.n1440 68.5181
R12768 vss.n1485 vss.n1440 68.5181
R12769 vss.n1455 vss.n1450 68.5181
R12770 vss.n1456 vss.n1455 68.5181
R12771 vss.n13881 vss.n13876 68.5181
R12772 vss.n13889 vss.n13881 68.5181
R12773 vss.n13895 vss.n13875 68.5181
R12774 vss.n13875 vss.n13864 68.5181
R12775 vss.n13873 vss.n13863 68.5181
R12776 vss.n13901 vss.n13863 68.5181
R12777 vss.n14036 vss.n8149 68.5181
R12778 vss.n14065 vss.n8149 68.5181
R12779 vss.n1362 vss.n1330 68.5181
R12780 vss.n1368 vss.n1330 68.5181
R12781 vss.n1361 vss.n1341 68.5181
R12782 vss.n1341 vss.n1332 68.5181
R12783 vss.n1347 vss.n1342 68.5181
R12784 vss.n1355 vss.n1347 68.5181
R12785 vss.n1271 vss.n1262 68.5181
R12786 vss.n1262 vss.n1234 68.5181
R12787 vss.n1260 vss.n1232 68.5181
R12788 vss.n1277 vss.n1232 68.5181
R12789 vss.n1247 vss.n1242 68.5181
R12790 vss.n1248 vss.n1247 68.5181
R12791 vss.n8040 vss.n2355 68.5181
R12792 vss.n2355 vss.n2327 68.5181
R12793 vss.n2353 vss.n2325 68.5181
R12794 vss.n8046 vss.n2325 68.5181
R12795 vss.n2340 vss.n2335 68.5181
R12796 vss.n2341 vss.n2340 68.5181
R12797 vss.n2270 vss.n2262 68.5181
R12798 vss.n2262 vss.n2233 68.5181
R12799 vss.n2260 vss.n2231 68.5181
R12800 vss.n2276 vss.n2231 68.5181
R12801 vss.n2251 vss.n2241 68.5181
R12802 vss.n2252 vss.n2251 68.5181
R12803 vss.n8068 vss.n8063 68.5181
R12804 vss.n8077 vss.n8068 68.5181
R12805 vss.n8083 vss.n8062 68.5181
R12806 vss.n8062 vss.n8052 68.5181
R12807 vss.n8060 vss.n2230 68.5181
R12808 vss.n8089 vss.n2230 68.5181
R12809 vss.n2317 vss.n2308 68.5181
R12810 vss.n2308 vss.n2279 68.5181
R12811 vss.n2306 vss.n2277 68.5181
R12812 vss.n2323 vss.n2277 68.5181
R12813 vss.n2292 vss.n2287 68.5181
R12814 vss.n2293 vss.n2292 68.5181
R12815 vss.n2404 vss.n2373 68.5181
R12816 vss.n2410 vss.n2373 68.5181
R12817 vss.n2403 vss.n2383 68.5181
R12818 vss.n2383 vss.n2374 68.5181
R12819 vss.n2389 vss.n2384 68.5181
R12820 vss.n2397 vss.n2389 68.5181
R12821 vss.n8120 vss.n8115 68.5181
R12822 vss.n8128 vss.n8120 68.5181
R12823 vss.n8134 vss.n8114 68.5181
R12824 vss.n8114 vss.n8103 68.5181
R12825 vss.n8112 vss.n8102 68.5181
R12826 vss.n8140 vss.n8102 68.5181
R12827 vss.n2099 vss.n2089 68.5181
R12828 vss.n14131 vss.n2099 68.5181
R12829 vss.n14137 vss.n2087 68.5181
R12830 vss.n2097 vss.n2087 68.5181
R12831 vss.n11949 vss.n11948 68.5181
R12832 vss.n11958 vss.n11949 68.5181
R12833 vss.n13497 vss.n13469 68.5181
R12834 vss.n13505 vss.n13497 68.5181
R12835 vss.n13511 vss.n13467 68.5181
R12836 vss.n13495 vss.n13467 68.5181
R12837 vss.n13483 vss.n13482 68.5181
R12838 vss.n13482 vss.n13477 68.5181
R12839 vss.n12036 vss.n12031 68.5181
R12840 vss.n12044 vss.n12036 68.5181
R12841 vss.n12050 vss.n12030 68.5181
R12842 vss.n12030 vss.n12020 68.5181
R12843 vss.n12028 vss.n12019 68.5181
R12844 vss.n12056 vss.n12019 68.5181
R12845 vss.n13729 vss.n8304 68.5181
R12846 vss.n13737 vss.n13729 68.5181
R12847 vss.n13743 vss.n8302 68.5181
R12848 vss.n13727 vss.n8302 68.5181
R12849 vss.n8318 vss.n8317 68.5181
R12850 vss.n8317 vss.n8312 68.5181
R12851 vss.n8462 vss.n8457 68.5181
R12852 vss.n8470 vss.n8462 68.5181
R12853 vss.n8476 vss.n8456 68.5181
R12854 vss.n8456 vss.n8446 68.5181
R12855 vss.n8454 vss.n8445 68.5181
R12856 vss.n8482 vss.n8445 68.5181
R12857 vss.n8539 vss.n8534 68.5181
R12858 vss.n8547 vss.n8539 68.5181
R12859 vss.n8553 vss.n8533 68.5181
R12860 vss.n8533 vss.n8523 68.5181
R12861 vss.n8531 vss.n8522 68.5181
R12862 vss.n8559 vss.n8522 68.5181
R12863 vss.n13017 vss.n9090 68.5181
R12864 vss.n13025 vss.n13017 68.5181
R12865 vss.n13031 vss.n9088 68.5181
R12866 vss.n13015 vss.n9088 68.5181
R12867 vss.n9104 vss.n9103 68.5181
R12868 vss.n9103 vss.n9098 68.5181
R12869 vss.n8982 vss.n8954 68.5181
R12870 vss.n8990 vss.n8982 68.5181
R12871 vss.n8996 vss.n8952 68.5181
R12872 vss.n8980 vss.n8952 68.5181
R12873 vss.n8968 vss.n8967 68.5181
R12874 vss.n8967 vss.n8962 68.5181
R12875 vss.n9134 vss.n9129 68.5181
R12876 vss.n9142 vss.n9134 68.5181
R12877 vss.n9148 vss.n9128 68.5181
R12878 vss.n9128 vss.n9118 68.5181
R12879 vss.n9126 vss.n9117 68.5181
R12880 vss.n9154 vss.n9117 68.5181
R12881 vss.n12565 vss.n12560 68.5181
R12882 vss.n12573 vss.n12565 68.5181
R12883 vss.n12628 vss.n12559 68.5181
R12884 vss.n12559 vss.n12549 68.5181
R12885 vss.n12557 vss.n12548 68.5181
R12886 vss.n12634 vss.n12548 68.5181
R12887 vss.n2214 vss.n2184 68.5181
R12888 vss.n2220 vss.n2184 68.5181
R12889 vss.n2190 vss.n2145 68.5181
R12890 vss.n2190 vss.n2185 68.5181
R12891 vss.n2162 vss.n2161 68.5181
R12892 vss.n2161 vss.n2156 68.5181
R12893 vss.n14086 vss.n2146 68.5181
R12894 vss.n2174 vss.n2146 68.5181
R12895 vss.n2176 vss.n2148 68.5181
R12896 vss.n14080 vss.n2176 68.5181
R12897 vss.n12595 vss.n12594 68.5181
R12898 vss.n12594 vss.n12589 68.5181
R12899 vss.n12624 vss.n12579 68.5181
R12900 vss.n12608 vss.n12579 68.5181
R12901 vss.n12610 vss.n12581 68.5181
R12902 vss.n12618 vss.n12610 68.5181
R12903 vss.n9013 vss.n9012 68.5181
R12904 vss.n9012 vss.n9007 68.5181
R12905 vss.n9040 vss.n8997 68.5181
R12906 vss.n9025 vss.n8997 68.5181
R12907 vss.n9027 vss.n8999 68.5181
R12908 vss.n9034 vss.n9027 68.5181
R12909 vss.n13098 vss.n13097 68.5181
R12910 vss.n13097 vss.n13092 68.5181
R12911 vss.n13128 vss.n13082 68.5181
R12912 vss.n13111 vss.n13082 68.5181
R12913 vss.n13113 vss.n13084 68.5181
R12914 vss.n13122 vss.n13113 68.5181
R12915 vss.n13050 vss.n13049 68.5181
R12916 vss.n13049 vss.n13044 68.5181
R12917 vss.n13080 vss.n13034 68.5181
R12918 vss.n13062 vss.n13034 68.5181
R12919 vss.n13064 vss.n13036 68.5181
R12920 vss.n13074 vss.n13064 68.5181
R12921 vss.n9057 vss.n9056 68.5181
R12922 vss.n9056 vss.n9051 68.5181
R12923 vss.n9086 vss.n9041 68.5181
R12924 vss.n9070 vss.n9041 68.5181
R12925 vss.n9072 vss.n9043 68.5181
R12926 vss.n9080 vss.n9072 68.5181
R12927 vss.n8240 vss.n8235 68.5181
R12928 vss.n8248 vss.n8240 68.5181
R12929 vss.n13844 vss.n8234 68.5181
R12930 vss.n8234 vss.n8228 68.5181
R12931 vss.n13845 vss.n8227 68.5181
R12932 vss.n13855 vss.n8227 68.5181
R12933 vss.n13810 vss.n13809 68.5181
R12934 vss.n13809 vss.n13804 68.5181
R12935 vss.n13840 vss.n13794 68.5181
R12936 vss.n13823 vss.n13794 68.5181
R12937 vss.n13825 vss.n13796 68.5181
R12938 vss.n13834 vss.n13825 68.5181
R12939 vss.n13762 vss.n13761 68.5181
R12940 vss.n13761 vss.n13756 68.5181
R12941 vss.n13792 vss.n13746 68.5181
R12942 vss.n13774 vss.n13746 68.5181
R12943 vss.n13776 vss.n13748 68.5181
R12944 vss.n13786 vss.n13776 68.5181
R12945 vss.n8271 vss.n8270 68.5181
R12946 vss.n8270 vss.n8265 68.5181
R12947 vss.n8300 vss.n8255 68.5181
R12948 vss.n8284 vss.n8255 68.5181
R12949 vss.n8286 vss.n8257 68.5181
R12950 vss.n8294 vss.n8286 68.5181
R12951 vss.n13528 vss.n13527 68.5181
R12952 vss.n13527 vss.n13522 68.5181
R12953 vss.n13555 vss.n13512 68.5181
R12954 vss.n13540 vss.n13512 68.5181
R12955 vss.n13542 vss.n13514 68.5181
R12956 vss.n13549 vss.n13542 68.5181
R12957 vss.n13621 vss.n13620 68.5181
R12958 vss.n13620 vss.n13615 68.5181
R12959 vss.n13651 vss.n13605 68.5181
R12960 vss.n13634 vss.n13605 68.5181
R12961 vss.n13636 vss.n13607 68.5181
R12962 vss.n13645 vss.n13636 68.5181
R12963 vss.n13572 vss.n13571 68.5181
R12964 vss.n13571 vss.n13566 68.5181
R12965 vss.n13603 vss.n13556 68.5181
R12966 vss.n13585 vss.n13556 68.5181
R12967 vss.n13587 vss.n13558 68.5181
R12968 vss.n13597 vss.n13587 68.5181
R12969 vss.n2071 vss.n2066 68.5181
R12970 vss.n2081 vss.n2071 68.5181
R12971 vss.n14141 vss.n2065 68.5181
R12972 vss.n2065 vss.n2059 68.5181
R12973 vss.n14142 vss.n2058 68.5181
R12974 vss.n14151 vss.n2058 68.5181
R12975 vss.n2200 vss.n2197 68.5181
R12976 vss.n2206 vss.n2197 68.5181
R12977 vss.n14093 vss.n2132 68.5181
R12978 vss.n14099 vss.n2132 68.5181
R12979 vss.n14092 vss.n2142 68.5181
R12980 vss.n2142 vss.n2133 68.5181
R12981 vss.n9288 vss.n9287 68.5181
R12982 vss.n9297 vss.n9288 68.5181
R12983 vss.n12854 vss.n9394 68.5181
R12984 vss.n12862 vss.n12854 68.5181
R12985 vss.n12868 vss.n9392 68.5181
R12986 vss.n12852 vss.n9392 68.5181
R12987 vss.n9408 vss.n9407 68.5181
R12988 vss.n9407 vss.n9402 68.5181
R12989 vss.n12749 vss.n12744 68.5181
R12990 vss.n12757 vss.n12749 68.5181
R12991 vss.n12764 vss.n12743 68.5181
R12992 vss.n12743 vss.n12733 68.5181
R12993 vss.n12741 vss.n12732 68.5181
R12994 vss.n12770 vss.n12732 68.5181
R12995 vss.n13331 vss.n8412 68.5181
R12996 vss.n13339 vss.n13331 68.5181
R12997 vss.n13345 vss.n8410 68.5181
R12998 vss.n13329 vss.n8410 68.5181
R12999 vss.n8426 vss.n8425 68.5181
R13000 vss.n8425 vss.n8420 68.5181
R13001 vss.n13450 vss.n13354 68.5181
R13002 vss.n13458 vss.n13450 68.5181
R13003 vss.n13464 vss.n13352 68.5181
R13004 vss.n13448 vss.n13352 68.5181
R13005 vss.n13368 vss.n13367 68.5181
R13006 vss.n13367 vss.n13362 68.5181
R13007 vss.n11852 vss.n11851 68.5181
R13008 vss.n11861 vss.n11852 68.5181
R13009 vss.n14189 vss.n2035 68.5181
R13010 vss.n2045 vss.n2035 68.5181
R13011 vss.n2047 vss.n2037 68.5181
R13012 vss.n14183 vss.n2047 68.5181
R13013 vss.n1804 vss.n1784 68.5181
R13014 vss.n1784 vss.n1773 68.5181
R13015 vss.n1782 vss.n1772 68.5181
R13016 vss.n1810 vss.n1772 68.5181
R13017 vss.n14364 vss.n1819 68.5181
R13018 vss.n14393 vss.n1819 68.5181
R13019 vss.n2026 vss.n2017 68.5181
R13020 vss.n2017 vss.n1989 68.5181
R13021 vss.n2015 vss.n1987 68.5181
R13022 vss.n2032 vss.n1987 68.5181
R13023 vss.n2002 vss.n1997 68.5181
R13024 vss.n2003 vss.n2002 68.5181
R13025 vss.n14248 vss.n14247 68.5181
R13026 vss.n14247 vss.n14243 68.5181
R13027 vss.n14268 vss.n14241 68.5181
R13028 vss.n14280 vss.n14241 68.5181
R13029 vss.n14266 vss.n14255 68.5181
R13030 vss.n14256 vss.n14255 68.5181
R13031 vss.n1025 vss.n1005 68.5181
R13032 vss.n1005 vss.n994 68.5181
R13033 vss.n1003 vss.n993 68.5181
R13034 vss.n1031 vss.n993 68.5181
R13035 vss.n15059 vss.n1040 68.5181
R13036 vss.n15088 vss.n1040 68.5181
R13037 vss.n1131 vss.n1122 68.5181
R13038 vss.n1122 vss.n1094 68.5181
R13039 vss.n1120 vss.n1092 68.5181
R13040 vss.n1137 vss.n1092 68.5181
R13041 vss.n1107 vss.n1102 68.5181
R13042 vss.n1108 vss.n1107 68.5181
R13043 vss.n14943 vss.n14942 68.5181
R13044 vss.n14942 vss.n14938 68.5181
R13045 vss.n14963 vss.n14936 68.5181
R13046 vss.n14975 vss.n14936 68.5181
R13047 vss.n14961 vss.n14950 68.5181
R13048 vss.n14951 vss.n14950 68.5181
R13049 vss.n6218 vss.n6209 68.5181
R13050 vss.n6247 vss.n6209 68.5181
R13051 vss.n15862 vss.n41 68.5181
R13052 vss.n41 vss.n31 68.5181
R13053 vss.n39 vss.n29 68.5181
R13054 vss.n15868 vss.n29 68.5181
R13055 vss.n3961 vss.n3954 68.5181
R13056 vss.n3962 vss.n3961 68.5181
R13057 vss.n3872 vss.n3867 68.5181
R13058 vss.n3881 vss.n3872 68.5181
R13059 vss.n3887 vss.n3866 68.5181
R13060 vss.n3866 vss.n3857 68.5181
R13061 vss.n3864 vss.n3855 68.5181
R13062 vss.n3893 vss.n3855 68.5181
R13063 vss.n3753 vss.n3748 68.5181
R13064 vss.n3762 vss.n3753 68.5181
R13065 vss.n3768 vss.n3747 68.5181
R13066 vss.n3747 vss.n3738 68.5181
R13067 vss.n3745 vss.n3736 68.5181
R13068 vss.n3774 vss.n3736 68.5181
R13069 vss.n3634 vss.n3629 68.5181
R13070 vss.n3643 vss.n3634 68.5181
R13071 vss.n3649 vss.n3628 68.5181
R13072 vss.n3628 vss.n3619 68.5181
R13073 vss.n3626 vss.n3617 68.5181
R13074 vss.n3655 vss.n3617 68.5181
R13075 vss.n15694 vss.n256 68.5181
R13076 vss.n256 vss.n246 68.5181
R13077 vss.n254 vss.n244 68.5181
R13078 vss.n15700 vss.n244 68.5181
R13079 vss.n6304 vss.n6295 68.5181
R13080 vss.n6305 vss.n6304 68.5181
R13081 vss.n15586 vss.n15585 68.5181
R13082 vss.n15585 vss.n15581 68.5181
R13083 vss.n15606 vss.n15579 68.5181
R13084 vss.n15618 vss.n15579 68.5181
R13085 vss.n15604 vss.n15593 68.5181
R13086 vss.n15594 vss.n15593 68.5181
R13087 vss.n317 vss.n309 68.5181
R13088 vss.n346 vss.n309 68.5181
R13089 vss.n3601 vss.n3568 68.5181
R13090 vss.n3607 vss.n3568 68.5181
R13091 vss.n3600 vss.n3578 68.5181
R13092 vss.n3578 vss.n3569 68.5181
R13093 vss.n3584 vss.n3579 68.5181
R13094 vss.n3594 vss.n3584 68.5181
R13095 vss.n375 vss.n370 68.5181
R13096 vss.n376 vss.n375 68.5181
R13097 vss.n12156 vss.n12151 68.5181
R13098 vss.n12164 vss.n12156 68.5181
R13099 vss.n12170 vss.n12150 68.5181
R13100 vss.n12150 vss.n12140 68.5181
R13101 vss.n12148 vss.n12137 68.5181
R13102 vss.n12176 vss.n12137 68.5181
R13103 vss.n11781 vss.n11779 68.5181
R13104 vss.n11779 vss.n11760 68.5181
R13105 vss.n11772 vss.n11758 68.5181
R13106 vss.n11800 vss.n11758 68.5181
R13107 vss.n11789 vss.n11771 68.5181
R13108 vss.n11771 vss.n11770 68.5181
R13109 vss.n10440 vss.n10439 68.5181
R13110 vss.n10439 vss.n10434 68.5181
R13111 vss.n10600 vss.n10571 68.5181
R13112 vss.n10608 vss.n10600 68.5181
R13113 vss.n10614 vss.n10569 68.5181
R13114 vss.n10598 vss.n10569 68.5181
R13115 vss.n10585 vss.n10584 68.5181
R13116 vss.n10584 vss.n10579 68.5181
R13117 vss.n10994 vss.n10965 68.5181
R13118 vss.n11002 vss.n10994 68.5181
R13119 vss.n11008 vss.n10963 68.5181
R13120 vss.n10992 vss.n10963 68.5181
R13121 vss.n10979 vss.n10978 68.5181
R13122 vss.n10978 vss.n10973 68.5181
R13123 vss.n10013 vss.n10008 68.5181
R13124 vss.n10021 vss.n10013 68.5181
R13125 vss.n10028 vss.n10007 68.5181
R13126 vss.n10007 vss.n9997 68.5181
R13127 vss.n10005 vss.n9996 68.5181
R13128 vss.n10034 vss.n9996 68.5181
R13129 vss.n9962 vss.n9952 68.5181
R13130 vss.n11644 vss.n9952 68.5181
R13131 vss.n11638 vss.n11637 68.5181
R13132 vss.n11638 vss.n9953 68.5181
R13133 vss.n11625 vss.n11619 68.5181
R13134 vss.n11628 vss.n11625 68.5181
R13135 vss.n3251 vss.n3246 62.0005
R13136 vss.n3249 vss.n3236 62.0005
R13137 vss.n3260 vss.n3259 62.0005
R13138 vss.n3268 vss.n3190 62.0005
R13139 vss.n8018 vss.n8017 62.0005
R13140 vss.n8011 vss.n2421 62.0005
R13141 vss.n8010 vss.n2430 62.0005
R13142 vss.n8004 vss.n8001 62.0005
R13143 vss.n1396 vss.n1381 62.0005
R13144 vss.n14718 vss.n1382 62.0005
R13145 vss.n14712 vss.n14711 62.0005
R13146 vss.n14705 vss.n1385 62.0005
R13147 vss.n7552 vss.n7549 62.0005
R13148 vss.n7560 vss.n7540 62.0005
R13149 vss.n7561 vss.n7531 62.0005
R13150 vss.n7570 vss.n7569 62.0005
R13151 vss.n2770 vss.n2767 62.0005
R13152 vss.n2778 vss.n2758 62.0005
R13153 vss.n2779 vss.n2749 62.0005
R13154 vss.n2788 vss.n2787 62.0005
R13155 vss.n1653 vss.n1638 62.0005
R13156 vss.n14568 vss.n1639 62.0005
R13157 vss.n14562 vss.n14561 62.0005
R13158 vss.n14555 vss.n1642 62.0005
R13159 vss.n2538 vss.n2535 62.0005
R13160 vss.n2544 vss.n2524 62.0005
R13161 vss.n2545 vss.n2515 62.0005
R13162 vss.n2554 vss.n2553 62.0005
R13163 vss.n1885 vss.n1872 62.0005
R13164 vss.n1984 vss.n1873 62.0005
R13165 vss.n1978 vss.n1977 62.0005
R13166 vss.n1971 vss.n1876 62.0005
R13167 vss.n4828 vss.n4824 62.0005
R13168 vss.n4827 vss.n4814 62.0005
R13169 vss.n4838 vss.n4837 62.0005
R13170 vss.n4846 vss.n4806 62.0005
R13171 vss.n4881 vss.n4878 62.0005
R13172 vss.n4889 vss.n4297 62.0005
R13173 vss.n4890 vss.n4290 62.0005
R13174 vss.n4899 vss.n4898 62.0005
R13175 vss.n617 vss.n602 62.0005
R13176 vss.n15413 vss.n603 62.0005
R13177 vss.n15407 vss.n15406 62.0005
R13178 vss.n15400 vss.n606 62.0005
R13179 vss.n5144 vss.n5141 62.0005
R13180 vss.n5152 vss.n5132 62.0005
R13181 vss.n5153 vss.n5123 62.0005
R13182 vss.n5162 vss.n5161 62.0005
R13183 vss.n5356 vss.n5353 62.0005
R13184 vss.n5364 vss.n5344 62.0005
R13185 vss.n5365 vss.n5335 62.0005
R13186 vss.n5374 vss.n5373 62.0005
R13187 vss.n874 vss.n859 62.0005
R13188 vss.n15263 vss.n860 62.0005
R13189 vss.n15257 vss.n15256 62.0005
R13190 vss.n15250 vss.n863 62.0005
R13191 vss.n6428 vss.n6425 62.0005
R13192 vss.n6436 vss.n6416 62.0005
R13193 vss.n6437 vss.n6407 62.0005
R13194 vss.n6446 vss.n6445 62.0005
R13195 vss.n6543 vss.n6540 62.0005
R13196 vss.n6551 vss.n6531 62.0005
R13197 vss.n6552 vss.n6522 62.0005
R13198 vss.n6561 vss.n6560 62.0005
R13199 vss.n12890 vss.n12889 62.0005
R13200 vss.n12883 vss.n9364 62.0005
R13201 vss.n12882 vss.n9373 62.0005
R13202 vss.n12876 vss.n12873 62.0005
R13203 vss.n12813 vss.n12812 62.0005
R13204 vss.n12806 vss.n12700 62.0005
R13205 vss.n12805 vss.n12709 62.0005
R13206 vss.n12799 vss.n12796 62.0005
R13207 vss.n8937 vss.n8918 62.0005
R13208 vss.n13147 vss.n8919 62.0005
R13209 vss.n8926 vss.n8925 62.0005
R13210 vss.n13141 vss.n13138 62.0005
R13211 vss.n12962 vss.n12948 62.0005
R13212 vss.n12988 vss.n12949 62.0005
R13213 vss.n12956 vss.n12955 62.0005
R13214 vss.n12982 vss.n12979 62.0005
R13215 vss.n8589 vss.n8504 62.0005
R13216 vss.n8614 vss.n8505 62.0005
R13217 vss.n8512 vss.n8511 62.0005
R13218 vss.n8608 vss.n8605 62.0005
R13219 vss.n13395 vss.n13384 62.0005
R13220 vss.n13407 vss.n13405 62.0005
R13221 vss.n13386 vss.n13377 62.0005
R13222 vss.n13416 vss.n13415 62.0005
R13223 vss.n8393 vss.n8374 62.0005
R13224 vss.n13670 vss.n8375 62.0005
R13225 vss.n8382 vss.n8381 62.0005
R13226 vss.n13664 vss.n13661 62.0005
R13227 vss.n12091 vss.n11880 62.0005
R13228 vss.n12109 vss.n11881 62.0005
R13229 vss.n12103 vss.n12102 62.0005
R13230 vss.n12117 vss.n11872 62.0005
R13231 vss.n13197 vss.n8869 51.0489
R13232 vss.n10359 vss.n10346 51.0489
R13233 vss.n10307 vss.n10300 51.0489
R13234 vss.n10324 vss.n10284 51.0489
R13235 vss.n11696 vss.n11694 51.0489
R13236 vss.n11681 vss.n9928 51.0489
R13237 vss.n11459 vss.n11457 51.0489
R13238 vss.n11444 vss.n9983 51.0489
R13239 vss.n11390 vss.n11388 51.0489
R13240 vss.n11409 vss.n11369 51.0489
R13241 vss.n11190 vss.n11188 51.0489
R13242 vss.n11175 vss.n11174 51.0489
R13243 vss.n11054 vss.n11052 51.0489
R13244 vss.n11039 vss.n10143 51.0489
R13245 vss.n10114 vss.n10112 51.0489
R13246 vss.n10099 vss.n10097 51.0489
R13247 vss.n10733 vss.n10730 51.0489
R13248 vss.n10752 vss.n10713 51.0489
R13249 vss.n10802 vss.n10800 51.0489
R13250 vss.n10787 vss.n10230 51.0489
R13251 vss.n10678 vss.n10676 51.0489
R13252 vss.n10697 vss.n10657 51.0489
R13253 vss.n10412 vss.n10410 51.0489
R13254 vss.n10397 vss.n10272 51.0489
R13255 vss.n10504 vss.n10502 51.0489
R13256 vss.n10489 vss.n10488 51.0489
R13257 vss.n10553 vss.n10551 51.0489
R13258 vss.n10537 vss.n10536 51.0489
R13259 vss.n10851 vss.n10849 51.0489
R13260 vss.n10835 vss.n10834 51.0489
R13261 vss.n10898 vss.n10896 51.0489
R13262 vss.n10883 vss.n10882 51.0489
R13263 vss.n10947 vss.n10945 51.0489
R13264 vss.n10931 vss.n10930 51.0489
R13265 vss.n11286 vss.n11284 51.0489
R13266 vss.n11270 vss.n11269 51.0489
R13267 vss.n11237 vss.n11235 51.0489
R13268 vss.n11222 vss.n11221 51.0489
R13269 vss.n11144 vss.n11142 51.0489
R13270 vss.n11128 vss.n11127 51.0489
R13271 vss.n11597 vss.n11595 51.0489
R13272 vss.n11581 vss.n11580 51.0489
R13273 vss.n11548 vss.n11546 51.0489
R13274 vss.n11533 vss.n11532 51.0489
R13275 vss.n11723 vss.n9882 51.0489
R13276 vss.n9899 vss.n9897 51.0489
R13277 vss.n11838 vss.n11813 51.0489
R13278 vss.n11829 vss.n11828 51.0489
R13279 vss.n11916 vss.n11910 51.0489
R13280 vss.n11932 vss.n11931 51.0489
R13281 vss.n9271 vss.n9260 51.0489
R13282 vss.n13165 vss.n8897 51.0489
R13283 vss.n12400 vss.n12399 51.0489
R13284 vss.n12416 vss.n12413 51.0489
R13285 vss.n9670 vss.n9669 51.0489
R13286 vss.n9655 vss.n9654 51.0489
R13287 vss.n9620 vss.n9619 51.0489
R13288 vss.n12369 vss.n12367 51.0489
R13289 vss.n13262 vss.n8636 51.0489
R13290 vss.n13277 vss.n13275 51.0489
R13291 vss.n12282 vss.n12281 51.0489
R13292 vss.n12298 vss.n12295 51.0489
R13293 vss.n9799 vss.n9798 51.0489
R13294 vss.n9784 vss.n9783 51.0489
R13295 vss.n9750 vss.n9749 51.0489
R13296 vss.n12251 vss.n12249 51.0489
R13297 vss.n8753 vss.n8742 51.0489
R13298 vss.n13688 vss.n8353 51.0489
R13299 vss.n11989 vss.n11983 51.0489
R13300 vss.n12005 vss.n12004 51.0489
R13301 vss.n11727 vss.n9878 51.0489
R13302 vss.n11745 vss.n11743 51.0489
R13303 vss.n12232 vss.n9856 51.0489
R13304 vss.n12218 vss.n12211 51.0489
R13305 vss.n8801 vss.n8761 51.0489
R13306 vss.n8787 vss.n8780 51.0489
R13307 vss.n8732 vss.n8693 51.0489
R13308 vss.n8718 vss.n8711 51.0489
R13309 vss.n9835 vss.n9829 51.0489
R13310 vss.n9849 vss.n9809 51.0489
R13311 vss.n12350 vss.n9728 51.0489
R13312 vss.n12336 vss.n12329 51.0489
R13313 vss.n8682 vss.n8642 51.0489
R13314 vss.n8668 vss.n8661 51.0489
R13315 vss.n12921 vss.n9203 51.0489
R13316 vss.n12937 vss.n12936 51.0489
R13317 vss.n9707 vss.n9700 51.0489
R13318 vss.n9721 vss.n9680 51.0489
R13319 vss.n12469 vss.n9598 51.0489
R13320 vss.n12455 vss.n12448 51.0489
R13321 vss.n9252 vss.n9212 51.0489
R13322 vss.n9238 vss.n9231 51.0489
R13323 vss.n9339 vss.n9333 51.0489
R13324 vss.n9355 vss.n9354 51.0489
R13325 vss.n12525 vss.n12519 51.0489
R13326 vss.n12541 vss.n12540 51.0489
R13327 vss.n9491 vss.n9490 51.0489
R13328 vss.n12488 vss.n12486 51.0489
R13329 vss.n9540 vss.n9539 51.0489
R13330 vss.n9525 vss.n9524 51.0489
R13331 vss.n9442 vss.n9440 51.0489
R13332 vss.n9457 vss.n9455 51.0489
R13333 vss.n12675 vss.n12669 51.0489
R13334 vss.n12691 vss.n12690 51.0489
R13335 vss.n9577 vss.n9571 51.0489
R13336 vss.n9591 vss.n9551 51.0489
R13337 vss.n10187 vss.n10186 51.0489
R13338 vss.n10202 vss.n10201 51.0489
R13339 vss.n11084 vss.n11083 51.0489
R13340 vss.n11099 vss.n11098 51.0489
R13341 vss.n11489 vss.n11488 51.0489
R13342 vss.n11504 vss.n11503 51.0489
R13343 vss.n13230 vss.n8832 51.0489
R13344 vss.n13246 vss.n13245 51.0489
R13345 vss.n15640 vss.n15638 51.0489
R13346 vss.n15652 vss.n15651 51.0489
R13347 vss.n3985 vss.n3984 51.0489
R13348 vss.n15892 vss.n13 51.0489
R13349 vss.n5650 vss.n5649 51.0489
R13350 vss.n5665 vss.n5663 51.0489
R13351 vss.n3725 vss.n3714 51.0489
R13352 vss.n15745 vss.n178 51.0489
R13353 vss.n3706 vss.n3667 51.0489
R13354 vss.n3692 vss.n3685 51.0489
R13355 vss.n5842 vss.n5841 51.0489
R13356 vss.n5857 vss.n5855 51.0489
R13357 vss.n3844 vss.n3833 51.0489
R13358 vss.n15801 vss.n100 51.0489
R13359 vss.n3825 vss.n3786 51.0489
R13360 vss.n3811 vss.n3804 51.0489
R13361 vss.n3944 vss.n3905 51.0489
R13362 vss.n3930 vss.n3923 51.0489
R13363 vss.n6082 vss.n6081 51.0489
R13364 vss.n6097 vss.n6095 51.0489
R13365 vss.n6034 vss.n6033 51.0489
R13366 vss.n6049 vss.n6047 51.0489
R13367 vss.n6197 vss.n6196 51.0489
R13368 vss.n6182 vss.n6175 51.0489
R13369 vss.n5751 vss.n5748 51.0489
R13370 vss.n5763 vss.n5761 51.0489
R13371 vss.n5794 vss.n5793 51.0489
R13372 vss.n5809 vss.n5807 51.0489
R13373 vss.n5958 vss.n5957 51.0489
R13374 vss.n5943 vss.n5936 51.0489
R13375 vss.n5563 vss.n5560 51.0489
R13376 vss.n5575 vss.n5573 51.0489
R13377 vss.n5720 vss.n5719 51.0489
R13378 vss.n5705 vss.n5698 51.0489
R13379 vss.n6330 vss.n6329 51.0489
R13380 vss.n6315 vss.n3559 51.0489
R13381 vss.n5620 vss.n5618 51.0489
R13382 vss.n5608 vss.n5605 51.0489
R13383 vss.n5896 vss.n5890 51.0489
R13384 vss.n5910 vss.n5727 51.0489
R13385 vss.n6135 vss.n6129 51.0489
R13386 vss.n6149 vss.n5967 51.0489
R13387 vss.n5991 vss.n5988 51.0489
R13388 vss.n6003 vss.n6001 51.0489
R13389 vss.n4390 vss.n4388 51.0489
R13390 vss.n4551 vss.n4369 51.0489
R13391 vss.n4480 vss.n4478 51.0489
R13392 vss.n4465 vss.n4464 51.0489
R13393 vss.n4528 vss.n4526 51.0489
R13394 vss.n4512 vss.n4511 51.0489
R13395 vss.n6648 vss.n6646 51.0489
R13396 vss.n6633 vss.n6632 51.0489
R13397 vss.n6600 vss.n6597 51.0489
R13398 vss.n6584 vss.n6514 51.0489
R13399 vss.n5246 vss.n5244 51.0489
R13400 vss.n5231 vss.n5230 51.0489
R13401 vss.n5292 vss.n5290 51.0489
R13402 vss.n5276 vss.n5275 51.0489
R13403 vss.n5532 vss.n5531 51.0489
R13404 vss.n4026 vss.n4024 51.0489
R13405 vss.n5507 vss.n5505 51.0489
R13406 vss.n5491 vss.n5490 51.0489
R13407 vss.n4071 vss.n4070 51.0489
R13408 vss.n4056 vss.n4055 51.0489
R13409 vss.n5458 vss.n5456 51.0489
R13410 vss.n5443 vss.n5442 51.0489
R13411 vss.n5411 vss.n5409 51.0489
R13412 vss.n5396 vss.n5327 51.0489
R13413 vss.n4161 vss.n4159 51.0489
R13414 vss.n4146 vss.n4145 51.0489
R13415 vss.n5081 vss.n5079 51.0489
R13416 vss.n5065 vss.n5064 51.0489
R13417 vss.n4215 vss.n4177 51.0489
R13418 vss.n4190 vss.n4189 51.0489
R13419 vss.n5033 vss.n5031 51.0489
R13420 vss.n5017 vss.n5016 51.0489
R13421 vss.n4252 vss.n4251 51.0489
R13422 vss.n4237 vss.n4236 51.0489
R13423 vss.n4984 vss.n4982 51.0489
R13424 vss.n4969 vss.n4968 51.0489
R13425 vss.n4115 vss.n4113 51.0489
R13426 vss.n4100 vss.n4099 51.0489
R13427 vss.n4936 vss.n4934 51.0489
R13428 vss.n4921 vss.n4282 51.0489
R13429 vss.n5199 vss.n5197 51.0489
R13430 vss.n5184 vss.n5115 51.0489
R13431 vss.n3374 vss.n3372 51.0489
R13432 vss.n3359 vss.n3358 51.0489
R13433 vss.n3421 vss.n3419 51.0489
R13434 vss.n3406 vss.n3405 51.0489
R13435 vss.n3484 vss.n3444 51.0489
R13436 vss.n3461 vss.n3458 51.0489
R13437 vss.n6371 vss.n3438 51.0489
R13438 vss.n6346 vss.n6343 51.0489
R13439 vss.n3532 vss.n3491 51.0489
R13440 vss.n3508 vss.n3506 51.0489
R13441 vss.n6483 vss.n6481 51.0489
R13442 vss.n6468 vss.n6399 51.0489
R13443 vss.n6685 vss.n6680 51.0489
R13444 vss.n6700 vss.n3339 51.0489
R13445 vss.n4434 vss.n4432 51.0489
R13446 vss.n4419 vss.n4418 51.0489
R13447 vss.n4777 vss.n4775 51.0489
R13448 vss.n4797 vss.n4756 51.0489
R13449 vss.n3292 vss.n3291 51.0489
R13450 vss.n6727 vss.n3305 51.0489
R13451 vss.n15523 vss.n15517 51.0489
R13452 vss.n15539 vss.n15538 51.0489
R13453 vss.n14866 vss.n14865 51.0489
R13454 vss.n15487 vss.n402 51.0489
R13455 vss.n15013 vss.n14988 51.0489
R13456 vss.n15004 vss.n15003 51.0489
R13457 vss.n1059 vss.n1058 51.0489
R13458 vss.n15037 vss.n1072 51.0489
R13459 vss.n14906 vss.n14905 51.0489
R13460 vss.n14923 vss.n14921 51.0489
R13461 vss.n521 vss.n520 51.0489
R13462 vss.n15431 vss.n534 51.0489
R13463 vss.n7319 vss.n7318 51.0489
R13464 vss.n7334 vss.n7332 51.0489
R13465 vss.n7390 vss.n7389 51.0489
R13466 vss.n7375 vss.n7374 51.0489
R13467 vss.n3086 vss.n3083 51.0489
R13468 vss.n3098 vss.n3096 51.0489
R13469 vss.n726 vss.n725 51.0489
R13470 vss.n15358 vss.n739 51.0489
R13471 vss.n779 vss.n778 51.0489
R13472 vss.n15281 vss.n792 51.0489
R13473 vss.n15144 vss.n983 51.0489
R13474 vss.n15159 vss.n15157 51.0489
R13475 vss.n15193 vss.n15192 51.0489
R13476 vss.n15208 vss.n15206 51.0489
R13477 vss.n936 vss.n935 51.0489
R13478 vss.n952 vss.n949 51.0489
R13479 vss.n832 vss.n826 51.0489
R13480 vss.n848 vss.n847 51.0489
R13481 vss.n15139 vss.n15098 51.0489
R13482 vss.n15125 vss.n15119 51.0489
R13483 vss.n7484 vss.n7444 51.0489
R13484 vss.n7470 vss.n7463 51.0489
R13485 vss.n15313 vss.n15312 51.0489
R13486 vss.n15329 vss.n15326 51.0489
R13487 vss.n679 vss.n678 51.0489
R13488 vss.n695 vss.n692 51.0489
R13489 vss.n7423 vss.n7417 51.0489
R13490 vss.n7437 vss.n7397 51.0489
R13491 vss.n7272 vss.n3127 51.0489
R13492 vss.n7287 vss.n7285 51.0489
R13493 vss.n575 vss.n569 51.0489
R13494 vss.n591 vss.n590 51.0489
R13495 vss.n471 vss.n470 51.0489
R13496 vss.n487 vss.n484 51.0489
R13497 vss.n4726 vss.n4720 51.0489
R13498 vss.n4742 vss.n4741 51.0489
R13499 vss.n4677 vss.n4674 51.0489
R13500 vss.n4689 vss.n4687 51.0489
R13501 vss.n4625 vss.n4624 51.0489
R13502 vss.n4640 vss.n4638 51.0489
R13503 vss.n4578 vss.n4576 51.0489
R13504 vss.n4593 vss.n4591 51.0489
R13505 vss.n4341 vss.n4335 51.0489
R13506 vss.n4357 vss.n4356 51.0489
R13507 vss.n7253 vss.n7247 51.0489
R13508 vss.n7267 vss.n7227 51.0489
R13509 vss.n6864 vss.n6862 51.0489
R13510 vss.n6849 vss.n6848 51.0489
R13511 vss.n7219 vss.n7218 51.0489
R13512 vss.n6822 vss.n6808 51.0489
R13513 vss.n6901 vss.n6896 51.0489
R13514 vss.n6916 vss.n6829 51.0489
R13515 vss.n2640 vss.n2601 51.0489
R13516 vss.n2619 vss.n2616 51.0489
R13517 vss.n1922 vss.n1919 51.0489
R13518 vss.n1942 vss.n1900 51.0489
R13519 vss.n2871 vss.n2869 51.0489
R13520 vss.n2856 vss.n2855 51.0489
R13521 vss.n7753 vss.n7751 51.0489
R13522 vss.n7737 vss.n7736 51.0489
R13523 vss.n2926 vss.n2887 51.0489
R13524 vss.n2901 vss.n2898 51.0489
R13525 vss.n7704 vss.n7702 51.0489
R13526 vss.n7688 vss.n7687 51.0489
R13527 vss.n3056 vss.n3015 51.0489
R13528 vss.n3032 vss.n3030 51.0489
R13529 vss.n7655 vss.n7653 51.0489
R13530 vss.n7640 vss.n7639 51.0489
R13531 vss.n2825 vss.n2823 51.0489
R13532 vss.n2810 vss.n2741 51.0489
R13533 vss.n2964 vss.n2961 51.0489
R13534 vss.n2948 vss.n2947 51.0489
R13535 vss.n3010 vss.n3008 51.0489
R13536 vss.n2994 vss.n2993 51.0489
R13537 vss.n7987 vss.n2456 51.0489
R13538 vss.n7962 vss.n2468 51.0489
R13539 vss.n7105 vss.n7104 51.0489
R13540 vss.n7120 vss.n7081 51.0489
R13541 vss.n7056 vss.n7055 51.0489
R13542 vss.n7074 vss.n7035 51.0489
R13543 vss.n7029 vss.n6990 51.0489
R13544 vss.n7008 vss.n7005 51.0489
R13545 vss.n7167 vss.n7127 51.0489
R13546 vss.n7147 vss.n7145 51.0489
R13547 vss.n6984 vss.n6923 51.0489
R13548 vss.n6963 vss.n6941 51.0489
R13549 vss.n7607 vss.n7605 51.0489
R13550 vss.n7592 vss.n7523 51.0489
R13551 vss.n7802 vss.n7800 51.0489
R13552 vss.n7787 vss.n7786 51.0489
R13553 vss.n7850 vss.n7848 51.0489
R13554 vss.n7835 vss.n7834 51.0489
R13555 vss.n7899 vss.n7897 51.0489
R13556 vss.n7883 vss.n7882 51.0489
R13557 vss.n2676 vss.n2661 51.0489
R13558 vss.n7923 vss.n2646 51.0489
R13559 vss.n2712 vss.n2711 51.0489
R13560 vss.n2697 vss.n2696 51.0489
R13561 vss.n2595 vss.n2486 51.0489
R13562 vss.n2575 vss.n2504 51.0489
R13563 vss.n1156 vss.n1154 51.0489
R13564 vss.n7942 vss.n7930 51.0489
R13565 vss.n7194 vss.n7192 51.0489
R13566 vss.n7179 vss.n3167 51.0489
R13567 vss.n6801 vss.n3172 51.0489
R13568 vss.n3207 vss.n3194 51.0489
R13569 vss.n6778 vss.n6776 51.0489
R13570 vss.n6763 vss.n6762 51.0489
R13571 vss.n14828 vss.n14822 51.0489
R13572 vss.n14844 vss.n14843 51.0489
R13573 vss.n14172 vss.n14171 51.0489
R13574 vss.n14792 vss.n1181 51.0489
R13575 vss.n14318 vss.n14293 51.0489
R13576 vss.n14309 vss.n14308 51.0489
R13577 vss.n1838 vss.n1837 51.0489
R13578 vss.n14342 vss.n1851 51.0489
R13579 vss.n14211 vss.n14210 51.0489
R13580 vss.n14228 vss.n14226 51.0489
R13581 vss.n1300 vss.n1299 51.0489
R13582 vss.n14736 vss.n1313 51.0489
R13583 vss.n13999 vss.n13998 51.0489
R13584 vss.n14014 vss.n14012 51.0489
R13585 vss.n8219 vss.n8218 51.0489
R13586 vss.n8204 vss.n8203 51.0489
R13587 vss.n8170 vss.n8169 51.0489
R13588 vss.n13968 vss.n13966 51.0489
R13589 vss.n1505 vss.n1504 51.0489
R13590 vss.n14663 vss.n1518 51.0489
R13591 vss.n1558 vss.n1557 51.0489
R13592 vss.n14586 vss.n1571 51.0489
R13593 vss.n14449 vss.n1762 51.0489
R13594 vss.n14464 vss.n14462 51.0489
R13595 vss.n14498 vss.n14497 51.0489
R13596 vss.n14513 vss.n14511 51.0489
R13597 vss.n1715 vss.n1714 51.0489
R13598 vss.n1731 vss.n1728 51.0489
R13599 vss.n1611 vss.n1605 51.0489
R13600 vss.n1627 vss.n1626 51.0489
R13601 vss.n14444 vss.n14403 51.0489
R13602 vss.n14430 vss.n14424 51.0489
R13603 vss.n13949 vss.n13909 51.0489
R13604 vss.n13935 vss.n13928 51.0489
R13605 vss.n14618 vss.n14617 51.0489
R13606 vss.n14634 vss.n14631 51.0489
R13607 vss.n1458 vss.n1457 51.0489
R13608 vss.n1474 vss.n1471 51.0489
R13609 vss.n13888 vss.n13882 51.0489
R13610 vss.n13902 vss.n13862 51.0489
R13611 vss.n14066 vss.n8148 51.0489
R13612 vss.n14052 vss.n14045 51.0489
R13613 vss.n1354 vss.n1348 51.0489
R13614 vss.n1370 vss.n1369 51.0489
R13615 vss.n1250 vss.n1249 51.0489
R13616 vss.n1266 vss.n1263 51.0489
R13617 vss.n2343 vss.n2342 51.0489
R13618 vss.n8035 vss.n2356 51.0489
R13619 vss.n2253 vss.n2250 51.0489
R13620 vss.n2265 vss.n2263 51.0489
R13621 vss.n8091 vss.n8090 51.0489
R13622 vss.n8076 vss.n8075 51.0489
R13623 vss.n2296 vss.n2294 51.0489
R13624 vss.n2311 vss.n2309 51.0489
R13625 vss.n2396 vss.n2390 51.0489
R13626 vss.n2412 vss.n2411 51.0489
R13627 vss.n8127 vss.n8121 51.0489
R13628 vss.n8141 vss.n8101 51.0489
R13629 vss.n14126 vss.n2100 51.0489
R13630 vss.n11960 vss.n11947 51.0489
R13631 vss.n13500 vss.n13498 51.0489
R13632 vss.n13485 vss.n13484 51.0489
R13633 vss.n12039 vss.n12037 51.0489
R13634 vss.n12058 vss.n12018 51.0489
R13635 vss.n13732 vss.n13730 51.0489
R13636 vss.n13717 vss.n8319 51.0489
R13637 vss.n8465 vss.n8463 51.0489
R13638 vss.n8484 vss.n8444 51.0489
R13639 vss.n8542 vss.n8540 51.0489
R13640 vss.n8561 vss.n8521 51.0489
R13641 vss.n13020 vss.n13018 51.0489
R13642 vss.n13005 vss.n9105 51.0489
R13643 vss.n8985 vss.n8983 51.0489
R13644 vss.n8970 vss.n8969 51.0489
R13645 vss.n9137 vss.n9135 51.0489
R13646 vss.n9156 vss.n9116 51.0489
R13647 vss.n12568 vss.n12566 51.0489
R13648 vss.n12636 vss.n12547 51.0489
R13649 vss.n2179 vss.n2177 51.0489
R13650 vss.n2164 vss.n2163 51.0489
R13651 vss.n12613 vss.n12611 51.0489
R13652 vss.n12597 vss.n12596 51.0489
R13653 vss.n9030 vss.n9029 51.0489
R13654 vss.n9015 vss.n9014 51.0489
R13655 vss.n13116 vss.n13114 51.0489
R13656 vss.n13100 vss.n13099 51.0489
R13657 vss.n13067 vss.n13065 51.0489
R13658 vss.n13052 vss.n13051 51.0489
R13659 vss.n9075 vss.n9073 51.0489
R13660 vss.n9059 vss.n9058 51.0489
R13661 vss.n13857 vss.n8226 51.0489
R13662 vss.n8243 vss.n8241 51.0489
R13663 vss.n13828 vss.n13826 51.0489
R13664 vss.n13812 vss.n13811 51.0489
R13665 vss.n13779 vss.n13777 51.0489
R13666 vss.n13764 vss.n13763 51.0489
R13667 vss.n8289 vss.n8287 51.0489
R13668 vss.n8273 vss.n8272 51.0489
R13669 vss.n13545 vss.n13544 51.0489
R13670 vss.n13530 vss.n13529 51.0489
R13671 vss.n13639 vss.n13637 51.0489
R13672 vss.n13623 vss.n13622 51.0489
R13673 vss.n13590 vss.n13588 51.0489
R13674 vss.n13575 vss.n13573 51.0489
R13675 vss.n14153 vss.n2057 51.0489
R13676 vss.n2075 vss.n2072 51.0489
R13677 vss.n2222 vss.n2183 51.0489
R13678 vss.n2201 vss.n2198 51.0489
R13679 vss.n14101 vss.n2131 51.0489
R13680 vss.n9299 vss.n9286 51.0489
R13681 vss.n12857 vss.n12855 51.0489
R13682 vss.n12842 vss.n9409 51.0489
R13683 vss.n12752 vss.n12750 51.0489
R13684 vss.n12772 vss.n12731 51.0489
R13685 vss.n13334 vss.n13332 51.0489
R13686 vss.n13319 vss.n8427 51.0489
R13687 vss.n13453 vss.n13451 51.0489
R13688 vss.n13438 vss.n13369 51.0489
R13689 vss.n2050 vss.n2048 51.0489
R13690 vss.n11863 vss.n11850 51.0489
R13691 vss.n1797 vss.n1791 51.0489
R13692 vss.n1811 vss.n1771 51.0489
R13693 vss.n14394 vss.n1818 51.0489
R13694 vss.n14380 vss.n14373 51.0489
R13695 vss.n2005 vss.n2004 51.0489
R13696 vss.n2021 vss.n2018 51.0489
R13697 vss.n14264 vss.n14257 51.0489
R13698 vss.n14275 vss.n14274 51.0489
R13699 vss.n1018 vss.n1012 51.0489
R13700 vss.n1032 vss.n992 51.0489
R13701 vss.n15089 vss.n1039 51.0489
R13702 vss.n15075 vss.n15068 51.0489
R13703 vss.n1110 vss.n1109 51.0489
R13704 vss.n1126 vss.n1123 51.0489
R13705 vss.n14959 vss.n14952 51.0489
R13706 vss.n14970 vss.n14969 51.0489
R13707 vss.n6248 vss.n6208 51.0489
R13708 vss.n6234 vss.n6227 51.0489
R13709 vss.n3963 vss.n3952 51.0489
R13710 vss.n15857 vss.n42 51.0489
R13711 vss.n3894 vss.n3854 51.0489
R13712 vss.n3880 vss.n3873 51.0489
R13713 vss.n3775 vss.n3735 51.0489
R13714 vss.n3761 vss.n3754 51.0489
R13715 vss.n3656 vss.n3616 51.0489
R13716 vss.n3642 vss.n3635 51.0489
R13717 vss.n6307 vss.n6306 51.0489
R13718 vss.n15689 vss.n257 51.0489
R13719 vss.n15602 vss.n15595 51.0489
R13720 vss.n15613 vss.n15612 51.0489
R13721 vss.n347 vss.n308 51.0489
R13722 vss.n333 vss.n326 51.0489
R13723 vss.n3593 vss.n3585 51.0489
R13724 vss.n3609 vss.n3608 51.0489
R13725 vss.n15548 vss.n377 51.0489
R13726 vss.n15563 vss.n15561 51.0489
R13727 vss.n12178 vss.n12177 51.0489
R13728 vss.n12163 vss.n12157 51.0489
R13729 vss.n11769 vss.n11767 51.0489
R13730 vss.n11783 vss.n11782 51.0489
R13731 vss.n10458 vss.n10455 51.0489
R13732 vss.n10442 vss.n10441 51.0489
R13733 vss.n10603 vss.n10601 51.0489
R13734 vss.n10588 vss.n10586 51.0489
R13735 vss.n10997 vss.n10995 51.0489
R13736 vss.n10982 vss.n10980 51.0489
R13737 vss.n10016 vss.n10014 51.0489
R13738 vss.n10036 vss.n9995 51.0489
R13739 vss.n11629 vss.n11622 51.0489
R13740 vss.n11646 vss.n9951 51.0489
R13741 vss.n14757 vss.n1225 49.0005
R13742 vss.n3228 vss.n3227 49.0005
R13743 vss.n8024 vss.n2415 49.0005
R13744 vss.n6961 vss.n6960 49.0005
R13745 vss.n14725 vss.n1373 49.0005
R13746 vss.n14698 vss.n14697 49.0005
R13747 vss.n14682 vss.n1432 49.0005
R13748 vss.n7590 vss.n7589 49.0005
R13749 vss.n14652 vss.n1531 49.0005
R13750 vss.n2808 vss.n2807 49.0005
R13751 vss.n14575 vss.n1630 49.0005
R13752 vss.n14548 vss.n14547 49.0005
R13753 vss.n14532 vss.n1689 49.0005
R13754 vss.n2573 vss.n2572 49.0005
R13755 vss.n14331 vss.n1864 49.0005
R13756 vss.n1964 vss.n1963 49.0005
R13757 vss.n15452 vss.n446 49.0005
R13758 vss.n4853 vss.n4800 49.0005
R13759 vss.n4872 vss.n4360 49.0005
R13760 vss.n4919 vss.n4918 49.0005
R13761 vss.n15420 vss.n594 49.0005
R13762 vss.n15393 vss.n15392 49.0005
R13763 vss.n15377 vss.n653 49.0005
R13764 vss.n5182 vss.n5181 49.0005
R13765 vss.n15347 vss.n752 49.0005
R13766 vss.n5394 vss.n5393 49.0005
R13767 vss.n15270 vss.n851 49.0005
R13768 vss.n15243 vss.n15242 49.0005
R13769 vss.n15227 vss.n910 49.0005
R13770 vss.n6466 vss.n6465 49.0005
R13771 vss.n15026 vss.n1085 49.0005
R13772 vss.n6582 vss.n6581 49.0005
R13773 vss.n12896 vss.n9358 49.0005
R13774 vss.n12840 vss.n12839 49.0005
R13775 vss.n12819 vss.n12694 49.0005
R13776 vss.n12790 vss.n12775 49.0005
R13777 vss.n13154 vss.n8910 49.0005
R13778 vss.n9163 vss.n9159 49.0005
R13779 vss.n12995 vss.n12940 49.0005
R13780 vss.n13317 vss.n13316 49.0005
R13781 vss.n13296 vss.n8496 49.0005
R13782 vss.n8580 vss.n8564 49.0005
R13783 vss.n13707 vss.n8330 49.0005
R13784 vss.n13436 vss.n13435 49.0005
R13785 vss.n13677 vss.n8366 49.0005
R13786 vss.n12065 vss.n12061 49.0005
R13787 vss.n12085 vss.n11935 49.0005
R13788 vss.n12124 vss.n11866 49.0005
R13789 vss.n10358 vss.n10357 35.2919
R13790 vss.n10357 vss.n10356 35.2919
R13791 vss.n10356 vss.n8871 35.2919
R13792 vss.n13194 vss.n8871 35.2919
R13793 vss.n13195 vss.n13194 35.2919
R13794 vss.n13196 vss.n13195 35.2919
R13795 vss.n10323 vss.n10322 35.2919
R13796 vss.n10322 vss.n10321 35.2919
R13797 vss.n10321 vss.n10286 35.2919
R13798 vss.n10305 vss.n10286 35.2919
R13799 vss.n10306 vss.n10305 35.2919
R13800 vss.n10308 vss.n10306 35.2919
R13801 vss.n11682 vss.n9921 35.2919
R13802 vss.n11690 vss.n9921 35.2919
R13803 vss.n11691 vss.n11690 35.2919
R13804 vss.n11702 vss.n11691 35.2919
R13805 vss.n11702 vss.n11701 35.2919
R13806 vss.n11701 vss.n11700 35.2919
R13807 vss.n11445 vss.n9976 35.2919
R13808 vss.n11453 vss.n9976 35.2919
R13809 vss.n11454 vss.n11453 35.2919
R13810 vss.n11465 vss.n11454 35.2919
R13811 vss.n11465 vss.n11464 35.2919
R13812 vss.n11464 vss.n11463 35.2919
R13813 vss.n11408 vss.n11407 35.2919
R13814 vss.n11407 vss.n11406 35.2919
R13815 vss.n11406 vss.n11371 35.2919
R13816 vss.n11396 vss.n11371 35.2919
R13817 vss.n11396 vss.n11395 35.2919
R13818 vss.n11395 vss.n11394 35.2919
R13819 vss.n11176 vss.n11167 35.2919
R13820 vss.n11184 vss.n11167 35.2919
R13821 vss.n11185 vss.n11184 35.2919
R13822 vss.n11196 vss.n11185 35.2919
R13823 vss.n11196 vss.n11195 35.2919
R13824 vss.n11195 vss.n11194 35.2919
R13825 vss.n11040 vss.n10136 35.2919
R13826 vss.n11048 vss.n10136 35.2919
R13827 vss.n11049 vss.n11048 35.2919
R13828 vss.n11060 vss.n11049 35.2919
R13829 vss.n11060 vss.n11059 35.2919
R13830 vss.n11059 vss.n11058 35.2919
R13831 vss.n10100 vss.n10090 35.2919
R13832 vss.n10108 vss.n10090 35.2919
R13833 vss.n10109 vss.n10108 35.2919
R13834 vss.n10120 vss.n10109 35.2919
R13835 vss.n10120 vss.n10119 35.2919
R13836 vss.n10119 vss.n10118 35.2919
R13837 vss.n10751 vss.n10750 35.2919
R13838 vss.n10750 vss.n10749 35.2919
R13839 vss.n10749 vss.n10715 35.2919
R13840 vss.n10739 vss.n10715 35.2919
R13841 vss.n10739 vss.n10738 35.2919
R13842 vss.n10738 vss.n10737 35.2919
R13843 vss.n10788 vss.n10223 35.2919
R13844 vss.n10796 vss.n10223 35.2919
R13845 vss.n10797 vss.n10796 35.2919
R13846 vss.n10808 vss.n10797 35.2919
R13847 vss.n10808 vss.n10807 35.2919
R13848 vss.n10807 vss.n10806 35.2919
R13849 vss.n10696 vss.n10695 35.2919
R13850 vss.n10695 vss.n10694 35.2919
R13851 vss.n10694 vss.n10659 35.2919
R13852 vss.n10684 vss.n10659 35.2919
R13853 vss.n10684 vss.n10683 35.2919
R13854 vss.n10683 vss.n10682 35.2919
R13855 vss.n10398 vss.n10265 35.2919
R13856 vss.n10406 vss.n10265 35.2919
R13857 vss.n10407 vss.n10406 35.2919
R13858 vss.n10418 vss.n10407 35.2919
R13859 vss.n10418 vss.n10417 35.2919
R13860 vss.n10417 vss.n10416 35.2919
R13861 vss.n10490 vss.n10481 35.2919
R13862 vss.n10498 vss.n10481 35.2919
R13863 vss.n10499 vss.n10498 35.2919
R13864 vss.n10512 vss.n10499 35.2919
R13865 vss.n10512 vss.n10511 35.2919
R13866 vss.n10511 vss.n10510 35.2919
R13867 vss.n10538 vss.n10529 35.2919
R13868 vss.n10547 vss.n10529 35.2919
R13869 vss.n10548 vss.n10547 35.2919
R13870 vss.n10559 vss.n10548 35.2919
R13871 vss.n10559 vss.n10558 35.2919
R13872 vss.n10558 vss.n10557 35.2919
R13873 vss.n10836 vss.n10827 35.2919
R13874 vss.n10845 vss.n10827 35.2919
R13875 vss.n10846 vss.n10845 35.2919
R13876 vss.n10858 vss.n10846 35.2919
R13877 vss.n10858 vss.n10857 35.2919
R13878 vss.n10857 vss.n10856 35.2919
R13879 vss.n10884 vss.n10875 35.2919
R13880 vss.n10892 vss.n10875 35.2919
R13881 vss.n10893 vss.n10892 35.2919
R13882 vss.n10906 vss.n10893 35.2919
R13883 vss.n10906 vss.n10905 35.2919
R13884 vss.n10905 vss.n10904 35.2919
R13885 vss.n10932 vss.n10923 35.2919
R13886 vss.n10941 vss.n10923 35.2919
R13887 vss.n10942 vss.n10941 35.2919
R13888 vss.n10953 vss.n10942 35.2919
R13889 vss.n10953 vss.n10952 35.2919
R13890 vss.n10952 vss.n10951 35.2919
R13891 vss.n11271 vss.n11262 35.2919
R13892 vss.n11280 vss.n11262 35.2919
R13893 vss.n11281 vss.n11280 35.2919
R13894 vss.n11293 vss.n11281 35.2919
R13895 vss.n11293 vss.n11292 35.2919
R13896 vss.n11292 vss.n11291 35.2919
R13897 vss.n11223 vss.n11214 35.2919
R13898 vss.n11231 vss.n11214 35.2919
R13899 vss.n11232 vss.n11231 35.2919
R13900 vss.n11245 vss.n11232 35.2919
R13901 vss.n11245 vss.n11244 35.2919
R13902 vss.n11244 vss.n11243 35.2919
R13903 vss.n11129 vss.n11120 35.2919
R13904 vss.n11138 vss.n11120 35.2919
R13905 vss.n11139 vss.n11138 35.2919
R13906 vss.n11150 vss.n11139 35.2919
R13907 vss.n11150 vss.n11149 35.2919
R13908 vss.n11149 vss.n11148 35.2919
R13909 vss.n11582 vss.n11573 35.2919
R13910 vss.n11591 vss.n11573 35.2919
R13911 vss.n11592 vss.n11591 35.2919
R13912 vss.n11604 vss.n11592 35.2919
R13913 vss.n11604 vss.n11603 35.2919
R13914 vss.n11603 vss.n11602 35.2919
R13915 vss.n11534 vss.n11525 35.2919
R13916 vss.n11542 vss.n11525 35.2919
R13917 vss.n11543 vss.n11542 35.2919
R13918 vss.n11556 vss.n11543 35.2919
R13919 vss.n11556 vss.n11555 35.2919
R13920 vss.n11555 vss.n11554 35.2919
R13921 vss.n9905 vss.n9904 35.2919
R13922 vss.n9906 vss.n9905 35.2919
R13923 vss.n9906 vss.n9884 35.2919
R13924 vss.n11720 vss.n9884 35.2919
R13925 vss.n11721 vss.n11720 35.2919
R13926 vss.n11722 vss.n11721 35.2919
R13927 vss.n11815 vss.n11814 35.2919
R13928 vss.n11819 vss.n11814 35.2919
R13929 vss.n11825 vss.n11819 35.2919
R13930 vss.n11826 vss.n11825 35.2919
R13931 vss.n11827 vss.n11826 35.2919
R13932 vss.n11830 vss.n11827 35.2919
R13933 vss.n11912 vss.n11904 35.2919
R13934 vss.n11922 vss.n11904 35.2919
R13935 vss.n11923 vss.n11922 35.2919
R13936 vss.n11925 vss.n11923 35.2919
R13937 vss.n11925 vss.n11924 35.2919
R13938 vss.n11924 vss.n11892 35.2919
R13939 vss.n9262 vss.n9261 35.2919
R13940 vss.n9263 vss.n9262 35.2919
R13941 vss.n9263 vss.n8894 35.2919
R13942 vss.n13171 vss.n8894 35.2919
R13943 vss.n13171 vss.n13170 35.2919
R13944 vss.n13170 vss.n13169 35.2919
R13945 vss.n12401 vss.n12392 35.2919
R13946 vss.n12409 vss.n12392 35.2919
R13947 vss.n12410 vss.n12409 35.2919
R13948 vss.n12422 vss.n12410 35.2919
R13949 vss.n12422 vss.n12421 35.2919
R13950 vss.n12421 vss.n12420 35.2919
R13951 vss.n9638 vss.n9628 35.2919
R13952 vss.n9663 vss.n9638 35.2919
R13953 vss.n9663 vss.n9662 35.2919
R13954 vss.n9662 vss.n9661 35.2919
R13955 vss.n9661 vss.n9641 35.2919
R13956 vss.n9648 vss.n9641 35.2919
R13957 vss.n9621 vss.n9612 35.2919
R13958 vss.n12363 vss.n9612 35.2919
R13959 vss.n12364 vss.n12363 35.2919
R13960 vss.n12375 vss.n12364 35.2919
R13961 vss.n12375 vss.n12374 35.2919
R13962 vss.n12374 vss.n12373 35.2919
R13963 vss.n13263 vss.n8629 35.2919
R13964 vss.n13271 vss.n8629 35.2919
R13965 vss.n13272 vss.n13271 35.2919
R13966 vss.n13283 vss.n13272 35.2919
R13967 vss.n13283 vss.n13282 35.2919
R13968 vss.n13282 vss.n13281 35.2919
R13969 vss.n12283 vss.n12274 35.2919
R13970 vss.n12291 vss.n12274 35.2919
R13971 vss.n12292 vss.n12291 35.2919
R13972 vss.n12304 vss.n12292 35.2919
R13973 vss.n12304 vss.n12303 35.2919
R13974 vss.n12303 vss.n12302 35.2919
R13975 vss.n9768 vss.n9758 35.2919
R13976 vss.n9792 vss.n9768 35.2919
R13977 vss.n9792 vss.n9791 35.2919
R13978 vss.n9791 vss.n9790 35.2919
R13979 vss.n9790 vss.n9771 35.2919
R13980 vss.n9778 vss.n9771 35.2919
R13981 vss.n9751 vss.n9742 35.2919
R13982 vss.n12245 vss.n9742 35.2919
R13983 vss.n12246 vss.n12245 35.2919
R13984 vss.n12257 vss.n12246 35.2919
R13985 vss.n12257 vss.n12256 35.2919
R13986 vss.n12256 vss.n12255 35.2919
R13987 vss.n8744 vss.n8743 35.2919
R13988 vss.n8745 vss.n8744 35.2919
R13989 vss.n8745 vss.n8350 35.2919
R13990 vss.n13694 vss.n8350 35.2919
R13991 vss.n13694 vss.n13693 35.2919
R13992 vss.n13693 vss.n13692 35.2919
R13993 vss.n11985 vss.n11977 35.2919
R13994 vss.n11995 vss.n11977 35.2919
R13995 vss.n11996 vss.n11995 35.2919
R13996 vss.n11998 vss.n11996 35.2919
R13997 vss.n11998 vss.n11997 35.2919
R13998 vss.n11997 vss.n11966 35.2919
R13999 vss.n11728 vss.n9871 35.2919
R14000 vss.n11739 vss.n9871 35.2919
R14001 vss.n11740 vss.n11739 35.2919
R14002 vss.n11751 vss.n11740 35.2919
R14003 vss.n11751 vss.n11750 35.2919
R14004 vss.n11750 vss.n11749 35.2919
R14005 vss.n12202 vss.n12201 35.2919
R14006 vss.n12226 vss.n12202 35.2919
R14007 vss.n12226 vss.n12225 35.2919
R14008 vss.n12225 vss.n12224 35.2919
R14009 vss.n12224 vss.n12205 35.2919
R14010 vss.n12213 vss.n12205 35.2919
R14011 vss.n8771 vss.n8770 35.2919
R14012 vss.n8795 vss.n8771 35.2919
R14013 vss.n8795 vss.n8794 35.2919
R14014 vss.n8794 vss.n8793 35.2919
R14015 vss.n8793 vss.n8774 35.2919
R14016 vss.n8783 vss.n8774 35.2919
R14017 vss.n8702 vss.n8701 35.2919
R14018 vss.n8726 vss.n8702 35.2919
R14019 vss.n8726 vss.n8725 35.2919
R14020 vss.n8725 vss.n8724 35.2919
R14021 vss.n8724 vss.n8705 35.2919
R14022 vss.n8714 vss.n8705 35.2919
R14023 vss.n9820 vss.n9819 35.2919
R14024 vss.n9843 vss.n9820 35.2919
R14025 vss.n9843 vss.n9842 35.2919
R14026 vss.n9842 vss.n9841 35.2919
R14027 vss.n9841 vss.n9823 35.2919
R14028 vss.n9831 vss.n9823 35.2919
R14029 vss.n12320 vss.n12319 35.2919
R14030 vss.n12344 vss.n12320 35.2919
R14031 vss.n12344 vss.n12343 35.2919
R14032 vss.n12343 vss.n12342 35.2919
R14033 vss.n12342 vss.n12323 35.2919
R14034 vss.n12331 vss.n12323 35.2919
R14035 vss.n8652 vss.n8651 35.2919
R14036 vss.n8676 vss.n8652 35.2919
R14037 vss.n8676 vss.n8675 35.2919
R14038 vss.n8675 vss.n8674 35.2919
R14039 vss.n8674 vss.n8655 35.2919
R14040 vss.n8664 vss.n8655 35.2919
R14041 vss.n12917 vss.n9197 35.2919
R14042 vss.n12927 vss.n9197 35.2919
R14043 vss.n12928 vss.n12927 35.2919
R14044 vss.n12930 vss.n12928 35.2919
R14045 vss.n12930 vss.n12929 35.2919
R14046 vss.n12929 vss.n9185 35.2919
R14047 vss.n9691 vss.n9690 35.2919
R14048 vss.n9715 vss.n9691 35.2919
R14049 vss.n9715 vss.n9714 35.2919
R14050 vss.n9714 vss.n9713 35.2919
R14051 vss.n9713 vss.n9694 35.2919
R14052 vss.n9703 vss.n9694 35.2919
R14053 vss.n12439 vss.n12438 35.2919
R14054 vss.n12463 vss.n12439 35.2919
R14055 vss.n12463 vss.n12462 35.2919
R14056 vss.n12462 vss.n12461 35.2919
R14057 vss.n12461 vss.n12442 35.2919
R14058 vss.n12450 vss.n12442 35.2919
R14059 vss.n9222 vss.n9221 35.2919
R14060 vss.n9246 vss.n9222 35.2919
R14061 vss.n9246 vss.n9245 35.2919
R14062 vss.n9245 vss.n9244 35.2919
R14063 vss.n9244 vss.n9225 35.2919
R14064 vss.n9234 vss.n9225 35.2919
R14065 vss.n9335 vss.n9327 35.2919
R14066 vss.n9345 vss.n9327 35.2919
R14067 vss.n9346 vss.n9345 35.2919
R14068 vss.n9348 vss.n9346 35.2919
R14069 vss.n9348 vss.n9347 35.2919
R14070 vss.n9347 vss.n9314 35.2919
R14071 vss.n12521 vss.n12513 35.2919
R14072 vss.n12531 vss.n12513 35.2919
R14073 vss.n12532 vss.n12531 35.2919
R14074 vss.n12534 vss.n12532 35.2919
R14075 vss.n12534 vss.n12533 35.2919
R14076 vss.n12533 vss.n9421 35.2919
R14077 vss.n9492 vss.n9483 35.2919
R14078 vss.n12482 vss.n9483 35.2919
R14079 vss.n12483 vss.n12482 35.2919
R14080 vss.n12494 vss.n12483 35.2919
R14081 vss.n12494 vss.n12493 35.2919
R14082 vss.n12493 vss.n12492 35.2919
R14083 vss.n9509 vss.n9499 35.2919
R14084 vss.n9533 vss.n9509 35.2919
R14085 vss.n9533 vss.n9532 35.2919
R14086 vss.n9532 vss.n9531 35.2919
R14087 vss.n9531 vss.n9512 35.2919
R14088 vss.n9519 vss.n9512 35.2919
R14089 vss.n9443 vss.n9433 35.2919
R14090 vss.n9451 vss.n9433 35.2919
R14091 vss.n9452 vss.n9451 35.2919
R14092 vss.n9464 vss.n9452 35.2919
R14093 vss.n9464 vss.n9463 35.2919
R14094 vss.n9463 vss.n9462 35.2919
R14095 vss.n12671 vss.n12663 35.2919
R14096 vss.n12681 vss.n12663 35.2919
R14097 vss.n12682 vss.n12681 35.2919
R14098 vss.n12684 vss.n12682 35.2919
R14099 vss.n12684 vss.n12683 35.2919
R14100 vss.n12683 vss.n12651 35.2919
R14101 vss.n9562 vss.n9561 35.2919
R14102 vss.n9585 vss.n9562 35.2919
R14103 vss.n9585 vss.n9584 35.2919
R14104 vss.n9584 vss.n9583 35.2919
R14105 vss.n9583 vss.n9565 35.2919
R14106 vss.n9573 vss.n9565 35.2919
R14107 vss.n10188 vss.n10179 35.2919
R14108 vss.n10196 vss.n10179 35.2919
R14109 vss.n10197 vss.n10196 35.2919
R14110 vss.n10207 vss.n10197 35.2919
R14111 vss.n10207 vss.n10206 35.2919
R14112 vss.n10206 vss.n10205 35.2919
R14113 vss.n11085 vss.n11076 35.2919
R14114 vss.n11093 vss.n11076 35.2919
R14115 vss.n11094 vss.n11093 35.2919
R14116 vss.n11104 vss.n11094 35.2919
R14117 vss.n11104 vss.n11103 35.2919
R14118 vss.n11103 vss.n11102 35.2919
R14119 vss.n11490 vss.n11481 35.2919
R14120 vss.n11498 vss.n11481 35.2919
R14121 vss.n11499 vss.n11498 35.2919
R14122 vss.n11509 vss.n11499 35.2919
R14123 vss.n11509 vss.n11508 35.2919
R14124 vss.n11508 vss.n11507 35.2919
R14125 vss.n13226 vss.n8826 35.2919
R14126 vss.n13236 vss.n8826 35.2919
R14127 vss.n13237 vss.n13236 35.2919
R14128 vss.n13239 vss.n13237 35.2919
R14129 vss.n13239 vss.n13238 35.2919
R14130 vss.n13238 vss.n8814 35.2919
R14131 vss.n15642 vss.n15641 35.2919
R14132 vss.n15643 vss.n15642 35.2919
R14133 vss.n15644 vss.n15643 35.2919
R14134 vss.n15646 vss.n15644 35.2919
R14135 vss.n15646 vss.n15645 35.2919
R14136 vss.n15645 vss.n15624 35.2919
R14137 vss.n3973 vss.n3972 35.2919
R14138 vss.n3977 vss.n3973 35.2919
R14139 vss.n3977 vss.n10 35.2919
R14140 vss.n15898 vss.n10 35.2919
R14141 vss.n15898 vss.n15897 35.2919
R14142 vss.n15897 vss.n15896 35.2919
R14143 vss.n5651 vss.n5642 35.2919
R14144 vss.n5659 vss.n5642 35.2919
R14145 vss.n5660 vss.n5659 35.2919
R14146 vss.n5671 vss.n5660 35.2919
R14147 vss.n5671 vss.n5670 35.2919
R14148 vss.n5670 vss.n5669 35.2919
R14149 vss.n3716 vss.n3715 35.2919
R14150 vss.n3717 vss.n3716 35.2919
R14151 vss.n3717 vss.n175 35.2919
R14152 vss.n15751 vss.n175 35.2919
R14153 vss.n15751 vss.n15750 35.2919
R14154 vss.n15750 vss.n15749 35.2919
R14155 vss.n3676 vss.n3675 35.2919
R14156 vss.n3700 vss.n3676 35.2919
R14157 vss.n3700 vss.n3699 35.2919
R14158 vss.n3699 vss.n3698 35.2919
R14159 vss.n3698 vss.n3679 35.2919
R14160 vss.n3688 vss.n3679 35.2919
R14161 vss.n5843 vss.n5834 35.2919
R14162 vss.n5851 vss.n5834 35.2919
R14163 vss.n5852 vss.n5851 35.2919
R14164 vss.n5863 vss.n5852 35.2919
R14165 vss.n5863 vss.n5862 35.2919
R14166 vss.n5862 vss.n5861 35.2919
R14167 vss.n3835 vss.n3834 35.2919
R14168 vss.n3836 vss.n3835 35.2919
R14169 vss.n3836 vss.n97 35.2919
R14170 vss.n15807 vss.n97 35.2919
R14171 vss.n15807 vss.n15806 35.2919
R14172 vss.n15806 vss.n15805 35.2919
R14173 vss.n3795 vss.n3794 35.2919
R14174 vss.n3819 vss.n3795 35.2919
R14175 vss.n3819 vss.n3818 35.2919
R14176 vss.n3818 vss.n3817 35.2919
R14177 vss.n3817 vss.n3798 35.2919
R14178 vss.n3807 vss.n3798 35.2919
R14179 vss.n3914 vss.n3913 35.2919
R14180 vss.n3938 vss.n3914 35.2919
R14181 vss.n3938 vss.n3937 35.2919
R14182 vss.n3937 vss.n3936 35.2919
R14183 vss.n3936 vss.n3917 35.2919
R14184 vss.n3926 vss.n3917 35.2919
R14185 vss.n6083 vss.n6074 35.2919
R14186 vss.n6091 vss.n6074 35.2919
R14187 vss.n6092 vss.n6091 35.2919
R14188 vss.n6103 vss.n6092 35.2919
R14189 vss.n6103 vss.n6102 35.2919
R14190 vss.n6102 vss.n6101 35.2919
R14191 vss.n6035 vss.n6026 35.2919
R14192 vss.n6043 vss.n6026 35.2919
R14193 vss.n6044 vss.n6043 35.2919
R14194 vss.n6056 vss.n6044 35.2919
R14195 vss.n6056 vss.n6055 35.2919
R14196 vss.n6055 vss.n6054 35.2919
R14197 vss.n6166 vss.n6155 35.2919
R14198 vss.n6190 vss.n6166 35.2919
R14199 vss.n6190 vss.n6189 35.2919
R14200 vss.n6189 vss.n6188 35.2919
R14201 vss.n6188 vss.n6169 35.2919
R14202 vss.n6177 vss.n6169 35.2919
R14203 vss.n5747 vss.n5739 35.2919
R14204 vss.n5757 vss.n5739 35.2919
R14205 vss.n5758 vss.n5757 35.2919
R14206 vss.n5769 vss.n5758 35.2919
R14207 vss.n5769 vss.n5768 35.2919
R14208 vss.n5768 vss.n5767 35.2919
R14209 vss.n5795 vss.n5786 35.2919
R14210 vss.n5803 vss.n5786 35.2919
R14211 vss.n5804 vss.n5803 35.2919
R14212 vss.n5816 vss.n5804 35.2919
R14213 vss.n5816 vss.n5815 35.2919
R14214 vss.n5815 vss.n5814 35.2919
R14215 vss.n5927 vss.n5916 35.2919
R14216 vss.n5951 vss.n5927 35.2919
R14217 vss.n5951 vss.n5950 35.2919
R14218 vss.n5950 vss.n5949 35.2919
R14219 vss.n5949 vss.n5930 35.2919
R14220 vss.n5938 vss.n5930 35.2919
R14221 vss.n5559 vss.n5551 35.2919
R14222 vss.n5569 vss.n5551 35.2919
R14223 vss.n5570 vss.n5569 35.2919
R14224 vss.n5581 vss.n5570 35.2919
R14225 vss.n5581 vss.n5580 35.2919
R14226 vss.n5580 vss.n5579 35.2919
R14227 vss.n5689 vss.n5539 35.2919
R14228 vss.n5713 vss.n5689 35.2919
R14229 vss.n5713 vss.n5712 35.2919
R14230 vss.n5712 vss.n5711 35.2919
R14231 vss.n5711 vss.n5692 35.2919
R14232 vss.n5700 vss.n5692 35.2919
R14233 vss.n3550 vss.n3539 35.2919
R14234 vss.n6323 vss.n3550 35.2919
R14235 vss.n6323 vss.n6322 35.2919
R14236 vss.n6322 vss.n6321 35.2919
R14237 vss.n6321 vss.n3553 35.2919
R14238 vss.n3561 vss.n3553 35.2919
R14239 vss.n5604 vss.n5598 35.2919
R14240 vss.n5614 vss.n5598 35.2919
R14241 vss.n5615 vss.n5614 35.2919
R14242 vss.n5626 vss.n5615 35.2919
R14243 vss.n5626 vss.n5625 35.2919
R14244 vss.n5625 vss.n5624 35.2919
R14245 vss.n5881 vss.n5880 35.2919
R14246 vss.n5904 vss.n5881 35.2919
R14247 vss.n5904 vss.n5903 35.2919
R14248 vss.n5903 vss.n5902 35.2919
R14249 vss.n5902 vss.n5884 35.2919
R14250 vss.n5892 vss.n5884 35.2919
R14251 vss.n6120 vss.n6119 35.2919
R14252 vss.n6143 vss.n6120 35.2919
R14253 vss.n6143 vss.n6142 35.2919
R14254 vss.n6142 vss.n6141 35.2919
R14255 vss.n6141 vss.n6123 35.2919
R14256 vss.n6131 vss.n6123 35.2919
R14257 vss.n5987 vss.n5979 35.2919
R14258 vss.n5997 vss.n5979 35.2919
R14259 vss.n5998 vss.n5997 35.2919
R14260 vss.n6009 vss.n5998 35.2919
R14261 vss.n6009 vss.n6008 35.2919
R14262 vss.n6008 vss.n6007 35.2919
R14263 vss.n4550 vss.n4549 35.2919
R14264 vss.n4549 vss.n4548 35.2919
R14265 vss.n4548 vss.n4371 35.2919
R14266 vss.n4396 vss.n4371 35.2919
R14267 vss.n4396 vss.n4395 35.2919
R14268 vss.n4395 vss.n4394 35.2919
R14269 vss.n4466 vss.n4457 35.2919
R14270 vss.n4474 vss.n4457 35.2919
R14271 vss.n4475 vss.n4474 35.2919
R14272 vss.n4487 vss.n4475 35.2919
R14273 vss.n4487 vss.n4486 35.2919
R14274 vss.n4486 vss.n4485 35.2919
R14275 vss.n4513 vss.n4504 35.2919
R14276 vss.n4522 vss.n4504 35.2919
R14277 vss.n4523 vss.n4522 35.2919
R14278 vss.n4534 vss.n4523 35.2919
R14279 vss.n4534 vss.n4533 35.2919
R14280 vss.n4533 vss.n4532 35.2919
R14281 vss.n6634 vss.n6625 35.2919
R14282 vss.n6642 vss.n6625 35.2919
R14283 vss.n6643 vss.n6642 35.2919
R14284 vss.n6654 vss.n6643 35.2919
R14285 vss.n6654 vss.n6653 35.2919
R14286 vss.n6653 vss.n6652 35.2919
R14287 vss.n6585 vss.n6507 35.2919
R14288 vss.n6593 vss.n6507 35.2919
R14289 vss.n6594 vss.n6593 35.2919
R14290 vss.n6606 vss.n6594 35.2919
R14291 vss.n6606 vss.n6605 35.2919
R14292 vss.n6605 vss.n6604 35.2919
R14293 vss.n5232 vss.n5223 35.2919
R14294 vss.n5240 vss.n5223 35.2919
R14295 vss.n5241 vss.n5240 35.2919
R14296 vss.n5252 vss.n5241 35.2919
R14297 vss.n5252 vss.n5251 35.2919
R14298 vss.n5251 vss.n5250 35.2919
R14299 vss.n5277 vss.n5268 35.2919
R14300 vss.n5286 vss.n5268 35.2919
R14301 vss.n5287 vss.n5286 35.2919
R14302 vss.n5299 vss.n5287 35.2919
R14303 vss.n5299 vss.n5298 35.2919
R14304 vss.n5298 vss.n5297 35.2919
R14305 vss.n4031 vss.n4030 35.2919
R14306 vss.n4033 vss.n4031 35.2919
R14307 vss.n4033 vss.n4032 35.2919
R14308 vss.n4032 vss.n4013 35.2919
R14309 vss.n4013 vss.n4009 35.2919
R14310 vss.n5530 vss.n4009 35.2919
R14311 vss.n5492 vss.n5483 35.2919
R14312 vss.n5501 vss.n5483 35.2919
R14313 vss.n5502 vss.n5501 35.2919
R14314 vss.n5513 vss.n5502 35.2919
R14315 vss.n5513 vss.n5512 35.2919
R14316 vss.n5512 vss.n5511 35.2919
R14317 vss.n4057 vss.n4048 35.2919
R14318 vss.n4065 vss.n4048 35.2919
R14319 vss.n4066 vss.n4065 35.2919
R14320 vss.n4076 vss.n4066 35.2919
R14321 vss.n4076 vss.n4075 35.2919
R14322 vss.n4075 vss.n4074 35.2919
R14323 vss.n5444 vss.n5435 35.2919
R14324 vss.n5452 vss.n5435 35.2919
R14325 vss.n5453 vss.n5452 35.2919
R14326 vss.n5464 vss.n5453 35.2919
R14327 vss.n5464 vss.n5463 35.2919
R14328 vss.n5463 vss.n5462 35.2919
R14329 vss.n5397 vss.n5320 35.2919
R14330 vss.n5405 vss.n5320 35.2919
R14331 vss.n5406 vss.n5405 35.2919
R14332 vss.n5417 vss.n5406 35.2919
R14333 vss.n5417 vss.n5416 35.2919
R14334 vss.n5416 vss.n5415 35.2919
R14335 vss.n4147 vss.n4138 35.2919
R14336 vss.n4155 vss.n4138 35.2919
R14337 vss.n4156 vss.n4155 35.2919
R14338 vss.n4167 vss.n4156 35.2919
R14339 vss.n4167 vss.n4166 35.2919
R14340 vss.n4166 vss.n4165 35.2919
R14341 vss.n5066 vss.n5057 35.2919
R14342 vss.n5075 vss.n5057 35.2919
R14343 vss.n5076 vss.n5075 35.2919
R14344 vss.n5087 vss.n5076 35.2919
R14345 vss.n5087 vss.n5086 35.2919
R14346 vss.n5086 vss.n5085 35.2919
R14347 vss.n4191 vss.n4182 35.2919
R14348 vss.n4202 vss.n4182 35.2919
R14349 vss.n4203 vss.n4202 35.2919
R14350 vss.n4206 vss.n4203 35.2919
R14351 vss.n4206 vss.n4205 35.2919
R14352 vss.n4205 vss.n4204 35.2919
R14353 vss.n5018 vss.n5009 35.2919
R14354 vss.n5027 vss.n5009 35.2919
R14355 vss.n5028 vss.n5027 35.2919
R14356 vss.n5039 vss.n5028 35.2919
R14357 vss.n5039 vss.n5038 35.2919
R14358 vss.n5038 vss.n5037 35.2919
R14359 vss.n4238 vss.n4229 35.2919
R14360 vss.n4246 vss.n4229 35.2919
R14361 vss.n4247 vss.n4246 35.2919
R14362 vss.n4257 vss.n4247 35.2919
R14363 vss.n4257 vss.n4256 35.2919
R14364 vss.n4256 vss.n4255 35.2919
R14365 vss.n4970 vss.n4961 35.2919
R14366 vss.n4978 vss.n4961 35.2919
R14367 vss.n4979 vss.n4978 35.2919
R14368 vss.n4990 vss.n4979 35.2919
R14369 vss.n4990 vss.n4989 35.2919
R14370 vss.n4989 vss.n4988 35.2919
R14371 vss.n4101 vss.n4092 35.2919
R14372 vss.n4109 vss.n4092 35.2919
R14373 vss.n4110 vss.n4109 35.2919
R14374 vss.n4121 vss.n4110 35.2919
R14375 vss.n4121 vss.n4120 35.2919
R14376 vss.n4120 vss.n4119 35.2919
R14377 vss.n4922 vss.n4275 35.2919
R14378 vss.n4930 vss.n4275 35.2919
R14379 vss.n4931 vss.n4930 35.2919
R14380 vss.n4942 vss.n4931 35.2919
R14381 vss.n4942 vss.n4941 35.2919
R14382 vss.n4941 vss.n4940 35.2919
R14383 vss.n5185 vss.n5108 35.2919
R14384 vss.n5193 vss.n5108 35.2919
R14385 vss.n5194 vss.n5193 35.2919
R14386 vss.n5205 vss.n5194 35.2919
R14387 vss.n5205 vss.n5204 35.2919
R14388 vss.n5204 vss.n5203 35.2919
R14389 vss.n3360 vss.n3351 35.2919
R14390 vss.n3368 vss.n3351 35.2919
R14391 vss.n3369 vss.n3368 35.2919
R14392 vss.n3380 vss.n3369 35.2919
R14393 vss.n3380 vss.n3379 35.2919
R14394 vss.n3379 vss.n3378 35.2919
R14395 vss.n3407 vss.n3398 35.2919
R14396 vss.n3415 vss.n3398 35.2919
R14397 vss.n3416 vss.n3415 35.2919
R14398 vss.n3427 vss.n3416 35.2919
R14399 vss.n3427 vss.n3426 35.2919
R14400 vss.n3426 vss.n3425 35.2919
R14401 vss.n3467 vss.n3466 35.2919
R14402 vss.n3468 vss.n3467 35.2919
R14403 vss.n3468 vss.n3446 35.2919
R14404 vss.n3481 vss.n3446 35.2919
R14405 vss.n3482 vss.n3481 35.2919
R14406 vss.n3483 vss.n3482 35.2919
R14407 vss.n6352 vss.n6351 35.2919
R14408 vss.n6351 vss.n6350 35.2919
R14409 vss.n6350 vss.n6338 35.2919
R14410 vss.n6363 vss.n6338 35.2919
R14411 vss.n6364 vss.n6363 35.2919
R14412 vss.n6365 vss.n6364 35.2919
R14413 vss.n3513 vss.n3512 35.2919
R14414 vss.n3514 vss.n3513 35.2919
R14415 vss.n3514 vss.n3493 35.2919
R14416 vss.n3529 vss.n3493 35.2919
R14417 vss.n3530 vss.n3529 35.2919
R14418 vss.n3531 vss.n3530 35.2919
R14419 vss.n6469 vss.n6392 35.2919
R14420 vss.n6477 vss.n6392 35.2919
R14421 vss.n6478 vss.n6477 35.2919
R14422 vss.n6489 vss.n6478 35.2919
R14423 vss.n6489 vss.n6488 35.2919
R14424 vss.n6488 vss.n6487 35.2919
R14425 vss.n6671 vss.n6670 35.2919
R14426 vss.n6694 vss.n6671 35.2919
R14427 vss.n6694 vss.n6693 35.2919
R14428 vss.n6693 vss.n6692 35.2919
R14429 vss.n6692 vss.n6674 35.2919
R14430 vss.n6681 vss.n6674 35.2919
R14431 vss.n4420 vss.n4411 35.2919
R14432 vss.n4428 vss.n4411 35.2919
R14433 vss.n4429 vss.n4428 35.2919
R14434 vss.n4440 vss.n4429 35.2919
R14435 vss.n4440 vss.n4439 35.2919
R14436 vss.n4439 vss.n4438 35.2919
R14437 vss.n4796 vss.n4795 35.2919
R14438 vss.n4795 vss.n4794 35.2919
R14439 vss.n4794 vss.n4758 35.2919
R14440 vss.n4783 vss.n4758 35.2919
R14441 vss.n4783 vss.n4782 35.2919
R14442 vss.n4782 vss.n4781 35.2919
R14443 vss.n3293 vss.n3284 35.2919
R14444 vss.n3301 vss.n3284 35.2919
R14445 vss.n3302 vss.n3301 35.2919
R14446 vss.n6733 vss.n3302 35.2919
R14447 vss.n6733 vss.n6732 35.2919
R14448 vss.n6732 vss.n6731 35.2919
R14449 vss.n15519 vss.n15511 35.2919
R14450 vss.n15529 vss.n15511 35.2919
R14451 vss.n15530 vss.n15529 35.2919
R14452 vss.n15532 vss.n15530 35.2919
R14453 vss.n15532 vss.n15531 35.2919
R14454 vss.n15531 vss.n386 35.2919
R14455 vss.n14854 vss.n14853 35.2919
R14456 vss.n14858 vss.n14854 35.2919
R14457 vss.n14858 vss.n399 35.2919
R14458 vss.n15493 vss.n399 35.2919
R14459 vss.n15493 vss.n15492 35.2919
R14460 vss.n15492 vss.n15491 35.2919
R14461 vss.n14990 vss.n14989 35.2919
R14462 vss.n14994 vss.n14989 35.2919
R14463 vss.n15000 vss.n14994 35.2919
R14464 vss.n15001 vss.n15000 35.2919
R14465 vss.n15002 vss.n15001 35.2919
R14466 vss.n15005 vss.n15002 35.2919
R14467 vss.n1060 vss.n1051 35.2919
R14468 vss.n1068 vss.n1051 35.2919
R14469 vss.n1069 vss.n1068 35.2919
R14470 vss.n15043 vss.n1069 35.2919
R14471 vss.n15043 vss.n15042 35.2919
R14472 vss.n15042 vss.n15041 35.2919
R14473 vss.n14907 vss.n14898 35.2919
R14474 vss.n14917 vss.n14898 35.2919
R14475 vss.n14918 vss.n14917 35.2919
R14476 vss.n14929 vss.n14918 35.2919
R14477 vss.n14929 vss.n14928 35.2919
R14478 vss.n14928 vss.n14927 35.2919
R14479 vss.n522 vss.n513 35.2919
R14480 vss.n530 vss.n513 35.2919
R14481 vss.n531 vss.n530 35.2919
R14482 vss.n15437 vss.n531 35.2919
R14483 vss.n15437 vss.n15436 35.2919
R14484 vss.n15436 vss.n15435 35.2919
R14485 vss.n7320 vss.n7311 35.2919
R14486 vss.n7328 vss.n7311 35.2919
R14487 vss.n7329 vss.n7328 35.2919
R14488 vss.n7340 vss.n7329 35.2919
R14489 vss.n7340 vss.n7339 35.2919
R14490 vss.n7339 vss.n7338 35.2919
R14491 vss.n7359 vss.n3062 35.2919
R14492 vss.n7383 vss.n7359 35.2919
R14493 vss.n7383 vss.n7382 35.2919
R14494 vss.n7382 vss.n7381 35.2919
R14495 vss.n7381 vss.n7362 35.2919
R14496 vss.n7369 vss.n7362 35.2919
R14497 vss.n3082 vss.n3074 35.2919
R14498 vss.n3092 vss.n3074 35.2919
R14499 vss.n3093 vss.n3092 35.2919
R14500 vss.n3104 vss.n3093 35.2919
R14501 vss.n3104 vss.n3103 35.2919
R14502 vss.n3103 vss.n3102 35.2919
R14503 vss.n727 vss.n718 35.2919
R14504 vss.n735 vss.n718 35.2919
R14505 vss.n736 vss.n735 35.2919
R14506 vss.n15364 vss.n736 35.2919
R14507 vss.n15364 vss.n15363 35.2919
R14508 vss.n15363 vss.n15362 35.2919
R14509 vss.n780 vss.n771 35.2919
R14510 vss.n788 vss.n771 35.2919
R14511 vss.n789 vss.n788 35.2919
R14512 vss.n15287 vss.n789 35.2919
R14513 vss.n15287 vss.n15286 35.2919
R14514 vss.n15286 vss.n15285 35.2919
R14515 vss.n15145 vss.n976 35.2919
R14516 vss.n15153 vss.n976 35.2919
R14517 vss.n15154 vss.n15153 35.2919
R14518 vss.n15166 vss.n15154 35.2919
R14519 vss.n15166 vss.n15165 35.2919
R14520 vss.n15165 vss.n15164 35.2919
R14521 vss.n15194 vss.n15185 35.2919
R14522 vss.n15202 vss.n15185 35.2919
R14523 vss.n15203 vss.n15202 35.2919
R14524 vss.n15214 vss.n15203 35.2919
R14525 vss.n15214 vss.n15213 35.2919
R14526 vss.n15213 vss.n15212 35.2919
R14527 vss.n937 vss.n928 35.2919
R14528 vss.n945 vss.n928 35.2919
R14529 vss.n946 vss.n945 35.2919
R14530 vss.n958 vss.n946 35.2919
R14531 vss.n958 vss.n957 35.2919
R14532 vss.n957 vss.n956 35.2919
R14533 vss.n828 vss.n820 35.2919
R14534 vss.n838 vss.n820 35.2919
R14535 vss.n839 vss.n838 35.2919
R14536 vss.n841 vss.n839 35.2919
R14537 vss.n841 vss.n840 35.2919
R14538 vss.n840 vss.n808 35.2919
R14539 vss.n15110 vss.n15109 35.2919
R14540 vss.n15133 vss.n15110 35.2919
R14541 vss.n15133 vss.n15132 35.2919
R14542 vss.n15132 vss.n15131 35.2919
R14543 vss.n15131 vss.n15113 35.2919
R14544 vss.n15121 vss.n15113 35.2919
R14545 vss.n7454 vss.n7453 35.2919
R14546 vss.n7478 vss.n7454 35.2919
R14547 vss.n7478 vss.n7477 35.2919
R14548 vss.n7477 vss.n7476 35.2919
R14549 vss.n7476 vss.n7457 35.2919
R14550 vss.n7465 vss.n7457 35.2919
R14551 vss.n15314 vss.n15305 35.2919
R14552 vss.n15322 vss.n15305 35.2919
R14553 vss.n15323 vss.n15322 35.2919
R14554 vss.n15335 vss.n15323 35.2919
R14555 vss.n15335 vss.n15334 35.2919
R14556 vss.n15334 vss.n15333 35.2919
R14557 vss.n680 vss.n671 35.2919
R14558 vss.n688 vss.n671 35.2919
R14559 vss.n689 vss.n688 35.2919
R14560 vss.n701 vss.n689 35.2919
R14561 vss.n701 vss.n700 35.2919
R14562 vss.n700 vss.n699 35.2919
R14563 vss.n7408 vss.n7407 35.2919
R14564 vss.n7431 vss.n7408 35.2919
R14565 vss.n7431 vss.n7430 35.2919
R14566 vss.n7430 vss.n7429 35.2919
R14567 vss.n7429 vss.n7411 35.2919
R14568 vss.n7419 vss.n7411 35.2919
R14569 vss.n7273 vss.n3120 35.2919
R14570 vss.n7281 vss.n3120 35.2919
R14571 vss.n7282 vss.n7281 35.2919
R14572 vss.n7294 vss.n7282 35.2919
R14573 vss.n7294 vss.n7293 35.2919
R14574 vss.n7293 vss.n7292 35.2919
R14575 vss.n571 vss.n563 35.2919
R14576 vss.n581 vss.n563 35.2919
R14577 vss.n582 vss.n581 35.2919
R14578 vss.n584 vss.n582 35.2919
R14579 vss.n584 vss.n583 35.2919
R14580 vss.n583 vss.n550 35.2919
R14581 vss.n472 vss.n463 35.2919
R14582 vss.n480 vss.n463 35.2919
R14583 vss.n481 vss.n480 35.2919
R14584 vss.n493 vss.n481 35.2919
R14585 vss.n493 vss.n492 35.2919
R14586 vss.n492 vss.n491 35.2919
R14587 vss.n4722 vss.n4714 35.2919
R14588 vss.n4732 vss.n4714 35.2919
R14589 vss.n4733 vss.n4732 35.2919
R14590 vss.n4735 vss.n4733 35.2919
R14591 vss.n4735 vss.n4734 35.2919
R14592 vss.n4734 vss.n4557 35.2919
R14593 vss.n4673 vss.n4665 35.2919
R14594 vss.n4683 vss.n4665 35.2919
R14595 vss.n4684 vss.n4683 35.2919
R14596 vss.n4695 vss.n4684 35.2919
R14597 vss.n4695 vss.n4694 35.2919
R14598 vss.n4694 vss.n4693 35.2919
R14599 vss.n4626 vss.n4617 35.2919
R14600 vss.n4634 vss.n4617 35.2919
R14601 vss.n4635 vss.n4634 35.2919
R14602 vss.n4647 vss.n4635 35.2919
R14603 vss.n4647 vss.n4646 35.2919
R14604 vss.n4646 vss.n4645 35.2919
R14605 vss.n4579 vss.n4569 35.2919
R14606 vss.n4587 vss.n4569 35.2919
R14607 vss.n4588 vss.n4587 35.2919
R14608 vss.n4600 vss.n4588 35.2919
R14609 vss.n4600 vss.n4599 35.2919
R14610 vss.n4599 vss.n4598 35.2919
R14611 vss.n4337 vss.n4329 35.2919
R14612 vss.n4347 vss.n4329 35.2919
R14613 vss.n4348 vss.n4347 35.2919
R14614 vss.n4350 vss.n4348 35.2919
R14615 vss.n4350 vss.n4349 35.2919
R14616 vss.n4349 vss.n4317 35.2919
R14617 vss.n7238 vss.n7237 35.2919
R14618 vss.n7261 vss.n7238 35.2919
R14619 vss.n7261 vss.n7260 35.2919
R14620 vss.n7260 vss.n7259 35.2919
R14621 vss.n7259 vss.n7241 35.2919
R14622 vss.n7249 vss.n7241 35.2919
R14623 vss.n6850 vss.n6841 35.2919
R14624 vss.n6858 vss.n6841 35.2919
R14625 vss.n6859 vss.n6858 35.2919
R14626 vss.n6870 vss.n6859 35.2919
R14627 vss.n6870 vss.n6869 35.2919
R14628 vss.n6869 vss.n6868 35.2919
R14629 vss.n6821 vss.n6820 35.2919
R14630 vss.n6820 vss.n6819 35.2919
R14631 vss.n6819 vss.n6811 35.2919
R14632 vss.n6811 vss.n3143 35.2919
R14633 vss.n3143 vss.n3139 35.2919
R14634 vss.n7217 vss.n3139 35.2919
R14635 vss.n6887 vss.n6886 35.2919
R14636 vss.n6910 vss.n6887 35.2919
R14637 vss.n6910 vss.n6909 35.2919
R14638 vss.n6909 vss.n6908 35.2919
R14639 vss.n6908 vss.n6890 35.2919
R14640 vss.n6897 vss.n6890 35.2919
R14641 vss.n2624 vss.n2623 35.2919
R14642 vss.n2625 vss.n2624 35.2919
R14643 vss.n2625 vss.n2603 35.2919
R14644 vss.n2637 vss.n2603 35.2919
R14645 vss.n2638 vss.n2637 35.2919
R14646 vss.n2639 vss.n2638 35.2919
R14647 vss.n1941 vss.n1940 35.2919
R14648 vss.n1940 vss.n1939 35.2919
R14649 vss.n1939 vss.n1902 35.2919
R14650 vss.n1928 vss.n1902 35.2919
R14651 vss.n1928 vss.n1927 35.2919
R14652 vss.n1927 vss.n1926 35.2919
R14653 vss.n2857 vss.n2848 35.2919
R14654 vss.n2865 vss.n2848 35.2919
R14655 vss.n2866 vss.n2865 35.2919
R14656 vss.n2877 vss.n2866 35.2919
R14657 vss.n2877 vss.n2876 35.2919
R14658 vss.n2876 vss.n2875 35.2919
R14659 vss.n7738 vss.n7729 35.2919
R14660 vss.n7747 vss.n7729 35.2919
R14661 vss.n7748 vss.n7747 35.2919
R14662 vss.n7759 vss.n7748 35.2919
R14663 vss.n7759 vss.n7758 35.2919
R14664 vss.n7758 vss.n7757 35.2919
R14665 vss.n2907 vss.n2906 35.2919
R14666 vss.n2906 vss.n2905 35.2919
R14667 vss.n2905 vss.n2893 35.2919
R14668 vss.n2918 vss.n2893 35.2919
R14669 vss.n2919 vss.n2918 35.2919
R14670 vss.n2920 vss.n2919 35.2919
R14671 vss.n7689 vss.n7680 35.2919
R14672 vss.n7698 vss.n7680 35.2919
R14673 vss.n7699 vss.n7698 35.2919
R14674 vss.n7711 vss.n7699 35.2919
R14675 vss.n7711 vss.n7710 35.2919
R14676 vss.n7710 vss.n7709 35.2919
R14677 vss.n3037 vss.n3036 35.2919
R14678 vss.n3038 vss.n3037 35.2919
R14679 vss.n3038 vss.n3017 35.2919
R14680 vss.n3053 vss.n3017 35.2919
R14681 vss.n3054 vss.n3053 35.2919
R14682 vss.n3055 vss.n3054 35.2919
R14683 vss.n7641 vss.n7632 35.2919
R14684 vss.n7649 vss.n7632 35.2919
R14685 vss.n7650 vss.n7649 35.2919
R14686 vss.n7661 vss.n7650 35.2919
R14687 vss.n7661 vss.n7660 35.2919
R14688 vss.n7660 vss.n7659 35.2919
R14689 vss.n2811 vss.n2734 35.2919
R14690 vss.n2819 vss.n2734 35.2919
R14691 vss.n2820 vss.n2819 35.2919
R14692 vss.n2831 vss.n2820 35.2919
R14693 vss.n2831 vss.n2830 35.2919
R14694 vss.n2830 vss.n2829 35.2919
R14695 vss.n2949 vss.n2940 35.2919
R14696 vss.n2957 vss.n2940 35.2919
R14697 vss.n2958 vss.n2957 35.2919
R14698 vss.n2970 vss.n2958 35.2919
R14699 vss.n2970 vss.n2969 35.2919
R14700 vss.n2969 vss.n2968 35.2919
R14701 vss.n2995 vss.n2986 35.2919
R14702 vss.n3004 vss.n2986 35.2919
R14703 vss.n3005 vss.n3004 35.2919
R14704 vss.n7495 vss.n3005 35.2919
R14705 vss.n7495 vss.n7494 35.2919
R14706 vss.n7494 vss.n7493 35.2919
R14707 vss.n7968 vss.n7967 35.2919
R14708 vss.n7967 vss.n7966 35.2919
R14709 vss.n7966 vss.n2463 35.2919
R14710 vss.n7979 vss.n2463 35.2919
R14711 vss.n7980 vss.n7979 35.2919
R14712 vss.n7981 vss.n7980 35.2919
R14713 vss.n7090 vss.n7089 35.2919
R14714 vss.n7114 vss.n7090 35.2919
R14715 vss.n7114 vss.n7113 35.2919
R14716 vss.n7113 vss.n7112 35.2919
R14717 vss.n7112 vss.n7093 35.2919
R14718 vss.n7100 vss.n7093 35.2919
R14719 vss.n7073 vss.n7072 35.2919
R14720 vss.n7072 vss.n7071 35.2919
R14721 vss.n7071 vss.n7037 35.2919
R14722 vss.n7053 vss.n7037 35.2919
R14723 vss.n7054 vss.n7053 35.2919
R14724 vss.n7057 vss.n7054 35.2919
R14725 vss.n7013 vss.n7012 35.2919
R14726 vss.n7014 vss.n7013 35.2919
R14727 vss.n7014 vss.n6992 35.2919
R14728 vss.n7026 vss.n6992 35.2919
R14729 vss.n7027 vss.n7026 35.2919
R14730 vss.n7028 vss.n7027 35.2919
R14731 vss.n7152 vss.n7151 35.2919
R14732 vss.n7153 vss.n7152 35.2919
R14733 vss.n7153 vss.n7129 35.2919
R14734 vss.n7164 vss.n7129 35.2919
R14735 vss.n7165 vss.n7164 35.2919
R14736 vss.n7166 vss.n7165 35.2919
R14737 vss.n6968 vss.n6967 35.2919
R14738 vss.n6969 vss.n6968 35.2919
R14739 vss.n6969 vss.n6925 35.2919
R14740 vss.n6981 vss.n6925 35.2919
R14741 vss.n6982 vss.n6981 35.2919
R14742 vss.n6983 vss.n6982 35.2919
R14743 vss.n7593 vss.n7516 35.2919
R14744 vss.n7601 vss.n7516 35.2919
R14745 vss.n7602 vss.n7601 35.2919
R14746 vss.n7613 vss.n7602 35.2919
R14747 vss.n7613 vss.n7612 35.2919
R14748 vss.n7612 vss.n7611 35.2919
R14749 vss.n7788 vss.n7779 35.2919
R14750 vss.n7796 vss.n7779 35.2919
R14751 vss.n7797 vss.n7796 35.2919
R14752 vss.n7808 vss.n7797 35.2919
R14753 vss.n7808 vss.n7807 35.2919
R14754 vss.n7807 vss.n7806 35.2919
R14755 vss.n7836 vss.n7827 35.2919
R14756 vss.n7844 vss.n7827 35.2919
R14757 vss.n7845 vss.n7844 35.2919
R14758 vss.n7856 vss.n7845 35.2919
R14759 vss.n7856 vss.n7855 35.2919
R14760 vss.n7855 vss.n7854 35.2919
R14761 vss.n7884 vss.n7875 35.2919
R14762 vss.n7893 vss.n7875 35.2919
R14763 vss.n7894 vss.n7893 35.2919
R14764 vss.n7906 vss.n7894 35.2919
R14765 vss.n7906 vss.n7905 35.2919
R14766 vss.n7905 vss.n7904 35.2919
R14767 vss.n7922 vss.n7921 35.2919
R14768 vss.n7921 vss.n7920 35.2919
R14769 vss.n7920 vss.n2648 35.2919
R14770 vss.n2668 vss.n2648 35.2919
R14771 vss.n2669 vss.n2668 35.2919
R14772 vss.n2670 vss.n2669 35.2919
R14773 vss.n2698 vss.n2689 35.2919
R14774 vss.n2706 vss.n2689 35.2919
R14775 vss.n2707 vss.n2706 35.2919
R14776 vss.n2717 vss.n2707 35.2919
R14777 vss.n2717 vss.n2716 35.2919
R14778 vss.n2716 vss.n2715 35.2919
R14779 vss.n2580 vss.n2579 35.2919
R14780 vss.n2581 vss.n2580 35.2919
R14781 vss.n2581 vss.n2488 35.2919
R14782 vss.n2592 vss.n2488 35.2919
R14783 vss.n2593 vss.n2592 35.2919
R14784 vss.n2594 vss.n2593 35.2919
R14785 vss.n7932 vss.n7931 35.2919
R14786 vss.n7934 vss.n7931 35.2919
R14787 vss.n7934 vss.n1151 35.2919
R14788 vss.n14876 vss.n1151 35.2919
R14789 vss.n14876 vss.n14875 35.2919
R14790 vss.n14875 vss.n14874 35.2919
R14791 vss.n7180 vss.n3160 35.2919
R14792 vss.n7188 vss.n3160 35.2919
R14793 vss.n7189 vss.n7188 35.2919
R14794 vss.n7200 vss.n7189 35.2919
R14795 vss.n7200 vss.n7199 35.2919
R14796 vss.n7199 vss.n7198 35.2919
R14797 vss.n3206 vss.n3205 35.2919
R14798 vss.n3205 vss.n3204 35.2919
R14799 vss.n3204 vss.n3174 35.2919
R14800 vss.n6798 vss.n3174 35.2919
R14801 vss.n6799 vss.n6798 35.2919
R14802 vss.n6800 vss.n6799 35.2919
R14803 vss.n6764 vss.n6755 35.2919
R14804 vss.n6772 vss.n6755 35.2919
R14805 vss.n6773 vss.n6772 35.2919
R14806 vss.n6784 vss.n6773 35.2919
R14807 vss.n6784 vss.n6783 35.2919
R14808 vss.n6783 vss.n6782 35.2919
R14809 vss.n14824 vss.n14816 35.2919
R14810 vss.n14834 vss.n14816 35.2919
R14811 vss.n14835 vss.n14834 35.2919
R14812 vss.n14837 vss.n14835 35.2919
R14813 vss.n14837 vss.n14836 35.2919
R14814 vss.n14836 vss.n1165 35.2919
R14815 vss.n14160 vss.n14159 35.2919
R14816 vss.n14164 vss.n14160 35.2919
R14817 vss.n14164 vss.n1178 35.2919
R14818 vss.n14798 vss.n1178 35.2919
R14819 vss.n14798 vss.n14797 35.2919
R14820 vss.n14797 vss.n14796 35.2919
R14821 vss.n14295 vss.n14294 35.2919
R14822 vss.n14299 vss.n14294 35.2919
R14823 vss.n14305 vss.n14299 35.2919
R14824 vss.n14306 vss.n14305 35.2919
R14825 vss.n14307 vss.n14306 35.2919
R14826 vss.n14310 vss.n14307 35.2919
R14827 vss.n1839 vss.n1830 35.2919
R14828 vss.n1847 vss.n1830 35.2919
R14829 vss.n1848 vss.n1847 35.2919
R14830 vss.n14348 vss.n1848 35.2919
R14831 vss.n14348 vss.n14347 35.2919
R14832 vss.n14347 vss.n14346 35.2919
R14833 vss.n14212 vss.n14203 35.2919
R14834 vss.n14222 vss.n14203 35.2919
R14835 vss.n14223 vss.n14222 35.2919
R14836 vss.n14234 vss.n14223 35.2919
R14837 vss.n14234 vss.n14233 35.2919
R14838 vss.n14233 vss.n14232 35.2919
R14839 vss.n1301 vss.n1292 35.2919
R14840 vss.n1309 vss.n1292 35.2919
R14841 vss.n1310 vss.n1309 35.2919
R14842 vss.n14742 vss.n1310 35.2919
R14843 vss.n14742 vss.n14741 35.2919
R14844 vss.n14741 vss.n14740 35.2919
R14845 vss.n14000 vss.n13991 35.2919
R14846 vss.n14008 vss.n13991 35.2919
R14847 vss.n14009 vss.n14008 35.2919
R14848 vss.n14020 vss.n14009 35.2919
R14849 vss.n14020 vss.n14019 35.2919
R14850 vss.n14019 vss.n14018 35.2919
R14851 vss.n8188 vss.n8178 35.2919
R14852 vss.n8212 vss.n8188 35.2919
R14853 vss.n8212 vss.n8211 35.2919
R14854 vss.n8211 vss.n8210 35.2919
R14855 vss.n8210 vss.n8191 35.2919
R14856 vss.n8198 vss.n8191 35.2919
R14857 vss.n8171 vss.n8162 35.2919
R14858 vss.n13962 vss.n8162 35.2919
R14859 vss.n13963 vss.n13962 35.2919
R14860 vss.n13974 vss.n13963 35.2919
R14861 vss.n13974 vss.n13973 35.2919
R14862 vss.n13973 vss.n13972 35.2919
R14863 vss.n1506 vss.n1497 35.2919
R14864 vss.n1514 vss.n1497 35.2919
R14865 vss.n1515 vss.n1514 35.2919
R14866 vss.n14669 vss.n1515 35.2919
R14867 vss.n14669 vss.n14668 35.2919
R14868 vss.n14668 vss.n14667 35.2919
R14869 vss.n1559 vss.n1550 35.2919
R14870 vss.n1567 vss.n1550 35.2919
R14871 vss.n1568 vss.n1567 35.2919
R14872 vss.n14592 vss.n1568 35.2919
R14873 vss.n14592 vss.n14591 35.2919
R14874 vss.n14591 vss.n14590 35.2919
R14875 vss.n14450 vss.n1755 35.2919
R14876 vss.n14458 vss.n1755 35.2919
R14877 vss.n14459 vss.n14458 35.2919
R14878 vss.n14471 vss.n14459 35.2919
R14879 vss.n14471 vss.n14470 35.2919
R14880 vss.n14470 vss.n14469 35.2919
R14881 vss.n14499 vss.n14490 35.2919
R14882 vss.n14507 vss.n14490 35.2919
R14883 vss.n14508 vss.n14507 35.2919
R14884 vss.n14519 vss.n14508 35.2919
R14885 vss.n14519 vss.n14518 35.2919
R14886 vss.n14518 vss.n14517 35.2919
R14887 vss.n1716 vss.n1707 35.2919
R14888 vss.n1724 vss.n1707 35.2919
R14889 vss.n1725 vss.n1724 35.2919
R14890 vss.n1737 vss.n1725 35.2919
R14891 vss.n1737 vss.n1736 35.2919
R14892 vss.n1736 vss.n1735 35.2919
R14893 vss.n1607 vss.n1599 35.2919
R14894 vss.n1617 vss.n1599 35.2919
R14895 vss.n1618 vss.n1617 35.2919
R14896 vss.n1620 vss.n1618 35.2919
R14897 vss.n1620 vss.n1619 35.2919
R14898 vss.n1619 vss.n1587 35.2919
R14899 vss.n14415 vss.n14414 35.2919
R14900 vss.n14438 vss.n14415 35.2919
R14901 vss.n14438 vss.n14437 35.2919
R14902 vss.n14437 vss.n14436 35.2919
R14903 vss.n14436 vss.n14418 35.2919
R14904 vss.n14426 vss.n14418 35.2919
R14905 vss.n13919 vss.n13918 35.2919
R14906 vss.n13943 vss.n13919 35.2919
R14907 vss.n13943 vss.n13942 35.2919
R14908 vss.n13942 vss.n13941 35.2919
R14909 vss.n13941 vss.n13922 35.2919
R14910 vss.n13930 vss.n13922 35.2919
R14911 vss.n14619 vss.n14610 35.2919
R14912 vss.n14627 vss.n14610 35.2919
R14913 vss.n14628 vss.n14627 35.2919
R14914 vss.n14640 vss.n14628 35.2919
R14915 vss.n14640 vss.n14639 35.2919
R14916 vss.n14639 vss.n14638 35.2919
R14917 vss.n1459 vss.n1450 35.2919
R14918 vss.n1467 vss.n1450 35.2919
R14919 vss.n1468 vss.n1467 35.2919
R14920 vss.n1480 vss.n1468 35.2919
R14921 vss.n1480 vss.n1479 35.2919
R14922 vss.n1479 vss.n1478 35.2919
R14923 vss.n13873 vss.n13872 35.2919
R14924 vss.n13896 vss.n13873 35.2919
R14925 vss.n13896 vss.n13895 35.2919
R14926 vss.n13895 vss.n13894 35.2919
R14927 vss.n13894 vss.n13876 35.2919
R14928 vss.n13884 vss.n13876 35.2919
R14929 vss.n14036 vss.n14035 35.2919
R14930 vss.n14060 vss.n14036 35.2919
R14931 vss.n14060 vss.n14059 35.2919
R14932 vss.n14059 vss.n14058 35.2919
R14933 vss.n14058 vss.n14039 35.2919
R14934 vss.n14047 vss.n14039 35.2919
R14935 vss.n1350 vss.n1342 35.2919
R14936 vss.n1360 vss.n1342 35.2919
R14937 vss.n1361 vss.n1360 35.2919
R14938 vss.n1363 vss.n1361 35.2919
R14939 vss.n1363 vss.n1362 35.2919
R14940 vss.n1362 vss.n1329 35.2919
R14941 vss.n1251 vss.n1242 35.2919
R14942 vss.n1259 vss.n1242 35.2919
R14943 vss.n1260 vss.n1259 35.2919
R14944 vss.n1272 vss.n1260 35.2919
R14945 vss.n1272 vss.n1271 35.2919
R14946 vss.n1271 vss.n1270 35.2919
R14947 vss.n2344 vss.n2335 35.2919
R14948 vss.n2352 vss.n2335 35.2919
R14949 vss.n2353 vss.n2352 35.2919
R14950 vss.n8041 vss.n2353 35.2919
R14951 vss.n8041 vss.n8040 35.2919
R14952 vss.n8040 vss.n8039 35.2919
R14953 vss.n2249 vss.n2241 35.2919
R14954 vss.n2259 vss.n2241 35.2919
R14955 vss.n2260 vss.n2259 35.2919
R14956 vss.n2271 vss.n2260 35.2919
R14957 vss.n2271 vss.n2270 35.2919
R14958 vss.n2270 vss.n2269 35.2919
R14959 vss.n8060 vss.n2229 35.2919
R14960 vss.n8084 vss.n8060 35.2919
R14961 vss.n8084 vss.n8083 35.2919
R14962 vss.n8083 vss.n8082 35.2919
R14963 vss.n8082 vss.n8063 35.2919
R14964 vss.n8070 vss.n8063 35.2919
R14965 vss.n2297 vss.n2287 35.2919
R14966 vss.n2305 vss.n2287 35.2919
R14967 vss.n2306 vss.n2305 35.2919
R14968 vss.n2318 vss.n2306 35.2919
R14969 vss.n2318 vss.n2317 35.2919
R14970 vss.n2317 vss.n2316 35.2919
R14971 vss.n2392 vss.n2384 35.2919
R14972 vss.n2402 vss.n2384 35.2919
R14973 vss.n2403 vss.n2402 35.2919
R14974 vss.n2405 vss.n2403 35.2919
R14975 vss.n2405 vss.n2404 35.2919
R14976 vss.n2404 vss.n2372 35.2919
R14977 vss.n8112 vss.n8111 35.2919
R14978 vss.n8135 vss.n8112 35.2919
R14979 vss.n8135 vss.n8134 35.2919
R14980 vss.n8134 vss.n8133 35.2919
R14981 vss.n8133 vss.n8115 35.2919
R14982 vss.n8123 vss.n8115 35.2919
R14983 vss.n11959 vss.n11958 35.2919
R14984 vss.n11958 vss.n11957 35.2919
R14985 vss.n11957 vss.n2097 35.2919
R14986 vss.n14132 vss.n2097 35.2919
R14987 vss.n14132 vss.n14131 35.2919
R14988 vss.n14131 vss.n14130 35.2919
R14989 vss.n13486 vss.n13477 35.2919
R14990 vss.n13494 vss.n13477 35.2919
R14991 vss.n13495 vss.n13494 35.2919
R14992 vss.n13506 vss.n13495 35.2919
R14993 vss.n13506 vss.n13505 35.2919
R14994 vss.n13505 vss.n13504 35.2919
R14995 vss.n12057 vss.n12056 35.2919
R14996 vss.n12056 vss.n12055 35.2919
R14997 vss.n12055 vss.n12020 35.2919
R14998 vss.n12045 vss.n12020 35.2919
R14999 vss.n12045 vss.n12044 35.2919
R15000 vss.n12044 vss.n12043 35.2919
R15001 vss.n13718 vss.n8312 35.2919
R15002 vss.n13726 vss.n8312 35.2919
R15003 vss.n13727 vss.n13726 35.2919
R15004 vss.n13738 vss.n13727 35.2919
R15005 vss.n13738 vss.n13737 35.2919
R15006 vss.n13737 vss.n13736 35.2919
R15007 vss.n8483 vss.n8482 35.2919
R15008 vss.n8482 vss.n8481 35.2919
R15009 vss.n8481 vss.n8446 35.2919
R15010 vss.n8471 vss.n8446 35.2919
R15011 vss.n8471 vss.n8470 35.2919
R15012 vss.n8470 vss.n8469 35.2919
R15013 vss.n8560 vss.n8559 35.2919
R15014 vss.n8559 vss.n8558 35.2919
R15015 vss.n8558 vss.n8523 35.2919
R15016 vss.n8548 vss.n8523 35.2919
R15017 vss.n8548 vss.n8547 35.2919
R15018 vss.n8547 vss.n8546 35.2919
R15019 vss.n13006 vss.n9098 35.2919
R15020 vss.n13014 vss.n9098 35.2919
R15021 vss.n13015 vss.n13014 35.2919
R15022 vss.n13026 vss.n13015 35.2919
R15023 vss.n13026 vss.n13025 35.2919
R15024 vss.n13025 vss.n13024 35.2919
R15025 vss.n8971 vss.n8962 35.2919
R15026 vss.n8979 vss.n8962 35.2919
R15027 vss.n8980 vss.n8979 35.2919
R15028 vss.n8991 vss.n8980 35.2919
R15029 vss.n8991 vss.n8990 35.2919
R15030 vss.n8990 vss.n8989 35.2919
R15031 vss.n9155 vss.n9154 35.2919
R15032 vss.n9154 vss.n9153 35.2919
R15033 vss.n9153 vss.n9118 35.2919
R15034 vss.n9143 vss.n9118 35.2919
R15035 vss.n9143 vss.n9142 35.2919
R15036 vss.n9142 vss.n9141 35.2919
R15037 vss.n12635 vss.n12634 35.2919
R15038 vss.n12634 vss.n12633 35.2919
R15039 vss.n12633 vss.n12549 35.2919
R15040 vss.n12574 vss.n12549 35.2919
R15041 vss.n12574 vss.n12573 35.2919
R15042 vss.n12573 vss.n12572 35.2919
R15043 vss.n2165 vss.n2156 35.2919
R15044 vss.n2173 vss.n2156 35.2919
R15045 vss.n2174 vss.n2173 35.2919
R15046 vss.n14081 vss.n2174 35.2919
R15047 vss.n14081 vss.n14080 35.2919
R15048 vss.n14080 vss.n14079 35.2919
R15049 vss.n12598 vss.n12589 35.2919
R15050 vss.n12607 vss.n12589 35.2919
R15051 vss.n12608 vss.n12607 35.2919
R15052 vss.n12619 vss.n12608 35.2919
R15053 vss.n12619 vss.n12618 35.2919
R15054 vss.n12618 vss.n12617 35.2919
R15055 vss.n9016 vss.n9007 35.2919
R15056 vss.n9024 vss.n9007 35.2919
R15057 vss.n9025 vss.n9024 35.2919
R15058 vss.n9035 vss.n9025 35.2919
R15059 vss.n9035 vss.n9034 35.2919
R15060 vss.n9034 vss.n9033 35.2919
R15061 vss.n13101 vss.n13092 35.2919
R15062 vss.n13110 vss.n13092 35.2919
R15063 vss.n13111 vss.n13110 35.2919
R15064 vss.n13123 vss.n13111 35.2919
R15065 vss.n13123 vss.n13122 35.2919
R15066 vss.n13122 vss.n13121 35.2919
R15067 vss.n13053 vss.n13044 35.2919
R15068 vss.n13061 vss.n13044 35.2919
R15069 vss.n13062 vss.n13061 35.2919
R15070 vss.n13075 vss.n13062 35.2919
R15071 vss.n13075 vss.n13074 35.2919
R15072 vss.n13074 vss.n13073 35.2919
R15073 vss.n9060 vss.n9051 35.2919
R15074 vss.n9069 vss.n9051 35.2919
R15075 vss.n9070 vss.n9069 35.2919
R15076 vss.n9081 vss.n9070 35.2919
R15077 vss.n9081 vss.n9080 35.2919
R15078 vss.n9080 vss.n9079 35.2919
R15079 vss.n8248 vss.n8247 35.2919
R15080 vss.n8249 vss.n8248 35.2919
R15081 vss.n8249 vss.n8228 35.2919
R15082 vss.n13854 vss.n8228 35.2919
R15083 vss.n13855 vss.n13854 35.2919
R15084 vss.n13856 vss.n13855 35.2919
R15085 vss.n13813 vss.n13804 35.2919
R15086 vss.n13822 vss.n13804 35.2919
R15087 vss.n13823 vss.n13822 35.2919
R15088 vss.n13835 vss.n13823 35.2919
R15089 vss.n13835 vss.n13834 35.2919
R15090 vss.n13834 vss.n13833 35.2919
R15091 vss.n13765 vss.n13756 35.2919
R15092 vss.n13773 vss.n13756 35.2919
R15093 vss.n13774 vss.n13773 35.2919
R15094 vss.n13787 vss.n13774 35.2919
R15095 vss.n13787 vss.n13786 35.2919
R15096 vss.n13786 vss.n13785 35.2919
R15097 vss.n8274 vss.n8265 35.2919
R15098 vss.n8283 vss.n8265 35.2919
R15099 vss.n8284 vss.n8283 35.2919
R15100 vss.n8295 vss.n8284 35.2919
R15101 vss.n8295 vss.n8294 35.2919
R15102 vss.n8294 vss.n8293 35.2919
R15103 vss.n13531 vss.n13522 35.2919
R15104 vss.n13539 vss.n13522 35.2919
R15105 vss.n13540 vss.n13539 35.2919
R15106 vss.n13550 vss.n13540 35.2919
R15107 vss.n13550 vss.n13549 35.2919
R15108 vss.n13549 vss.n13548 35.2919
R15109 vss.n13624 vss.n13615 35.2919
R15110 vss.n13633 vss.n13615 35.2919
R15111 vss.n13634 vss.n13633 35.2919
R15112 vss.n13646 vss.n13634 35.2919
R15113 vss.n13646 vss.n13645 35.2919
R15114 vss.n13645 vss.n13644 35.2919
R15115 vss.n13576 vss.n13566 35.2919
R15116 vss.n13584 vss.n13566 35.2919
R15117 vss.n13585 vss.n13584 35.2919
R15118 vss.n13598 vss.n13585 35.2919
R15119 vss.n13598 vss.n13597 35.2919
R15120 vss.n13597 vss.n13596 35.2919
R15121 vss.n2081 vss.n2080 35.2919
R15122 vss.n2082 vss.n2081 35.2919
R15123 vss.n2082 vss.n2059 35.2919
R15124 vss.n14150 vss.n2059 35.2919
R15125 vss.n14151 vss.n14150 35.2919
R15126 vss.n14152 vss.n14151 35.2919
R15127 vss.n2206 vss.n2205 35.2919
R15128 vss.n2207 vss.n2206 35.2919
R15129 vss.n2207 vss.n2185 35.2919
R15130 vss.n2219 vss.n2185 35.2919
R15131 vss.n2220 vss.n2219 35.2919
R15132 vss.n2221 vss.n2220 35.2919
R15133 vss.n9298 vss.n9297 35.2919
R15134 vss.n9297 vss.n9296 35.2919
R15135 vss.n9296 vss.n2133 35.2919
R15136 vss.n14098 vss.n2133 35.2919
R15137 vss.n14099 vss.n14098 35.2919
R15138 vss.n14100 vss.n14099 35.2919
R15139 vss.n12843 vss.n9402 35.2919
R15140 vss.n12851 vss.n9402 35.2919
R15141 vss.n12852 vss.n12851 35.2919
R15142 vss.n12863 vss.n12852 35.2919
R15143 vss.n12863 vss.n12862 35.2919
R15144 vss.n12862 vss.n12861 35.2919
R15145 vss.n12771 vss.n12770 35.2919
R15146 vss.n12770 vss.n12769 35.2919
R15147 vss.n12769 vss.n12733 35.2919
R15148 vss.n12758 vss.n12733 35.2919
R15149 vss.n12758 vss.n12757 35.2919
R15150 vss.n12757 vss.n12756 35.2919
R15151 vss.n13320 vss.n8420 35.2919
R15152 vss.n13328 vss.n8420 35.2919
R15153 vss.n13329 vss.n13328 35.2919
R15154 vss.n13340 vss.n13329 35.2919
R15155 vss.n13340 vss.n13339 35.2919
R15156 vss.n13339 vss.n13338 35.2919
R15157 vss.n13439 vss.n13362 35.2919
R15158 vss.n13447 vss.n13362 35.2919
R15159 vss.n13448 vss.n13447 35.2919
R15160 vss.n13459 vss.n13448 35.2919
R15161 vss.n13459 vss.n13458 35.2919
R15162 vss.n13458 vss.n13457 35.2919
R15163 vss.n11862 vss.n11861 35.2919
R15164 vss.n11861 vss.n11860 35.2919
R15165 vss.n11860 vss.n2045 35.2919
R15166 vss.n14184 vss.n2045 35.2919
R15167 vss.n14184 vss.n14183 35.2919
R15168 vss.n14183 vss.n14182 35.2919
R15169 vss.n1782 vss.n1781 35.2919
R15170 vss.n1805 vss.n1782 35.2919
R15171 vss.n1805 vss.n1804 35.2919
R15172 vss.n1804 vss.n1803 35.2919
R15173 vss.n1803 vss.n1785 35.2919
R15174 vss.n1793 vss.n1785 35.2919
R15175 vss.n14364 vss.n14363 35.2919
R15176 vss.n14388 vss.n14364 35.2919
R15177 vss.n14388 vss.n14387 35.2919
R15178 vss.n14387 vss.n14386 35.2919
R15179 vss.n14386 vss.n14367 35.2919
R15180 vss.n14375 vss.n14367 35.2919
R15181 vss.n2006 vss.n1997 35.2919
R15182 vss.n2014 vss.n1997 35.2919
R15183 vss.n2015 vss.n2014 35.2919
R15184 vss.n2027 vss.n2015 35.2919
R15185 vss.n2027 vss.n2026 35.2919
R15186 vss.n2026 vss.n2025 35.2919
R15187 vss.n14266 vss.n14265 35.2919
R15188 vss.n14267 vss.n14266 35.2919
R15189 vss.n14268 vss.n14267 35.2919
R15190 vss.n14269 vss.n14268 35.2919
R15191 vss.n14269 vss.n14248 35.2919
R15192 vss.n14273 vss.n14248 35.2919
R15193 vss.n1003 vss.n1002 35.2919
R15194 vss.n1026 vss.n1003 35.2919
R15195 vss.n1026 vss.n1025 35.2919
R15196 vss.n1025 vss.n1024 35.2919
R15197 vss.n1024 vss.n1006 35.2919
R15198 vss.n1014 vss.n1006 35.2919
R15199 vss.n15059 vss.n15058 35.2919
R15200 vss.n15083 vss.n15059 35.2919
R15201 vss.n15083 vss.n15082 35.2919
R15202 vss.n15082 vss.n15081 35.2919
R15203 vss.n15081 vss.n15062 35.2919
R15204 vss.n15070 vss.n15062 35.2919
R15205 vss.n1111 vss.n1102 35.2919
R15206 vss.n1119 vss.n1102 35.2919
R15207 vss.n1120 vss.n1119 35.2919
R15208 vss.n1132 vss.n1120 35.2919
R15209 vss.n1132 vss.n1131 35.2919
R15210 vss.n1131 vss.n1130 35.2919
R15211 vss.n14961 vss.n14960 35.2919
R15212 vss.n14962 vss.n14961 35.2919
R15213 vss.n14963 vss.n14962 35.2919
R15214 vss.n14964 vss.n14963 35.2919
R15215 vss.n14964 vss.n14943 35.2919
R15216 vss.n14968 vss.n14943 35.2919
R15217 vss.n6218 vss.n6217 35.2919
R15218 vss.n6242 vss.n6218 35.2919
R15219 vss.n6242 vss.n6241 35.2919
R15220 vss.n6241 vss.n6240 35.2919
R15221 vss.n6240 vss.n6221 35.2919
R15222 vss.n6229 vss.n6221 35.2919
R15223 vss.n3954 vss.n3953 35.2919
R15224 vss.n3955 vss.n3954 35.2919
R15225 vss.n3955 vss.n39 35.2919
R15226 vss.n15863 vss.n39 35.2919
R15227 vss.n15863 vss.n15862 35.2919
R15228 vss.n15862 vss.n15861 35.2919
R15229 vss.n3864 vss.n3863 35.2919
R15230 vss.n3888 vss.n3864 35.2919
R15231 vss.n3888 vss.n3887 35.2919
R15232 vss.n3887 vss.n3886 35.2919
R15233 vss.n3886 vss.n3867 35.2919
R15234 vss.n3876 vss.n3867 35.2919
R15235 vss.n3745 vss.n3744 35.2919
R15236 vss.n3769 vss.n3745 35.2919
R15237 vss.n3769 vss.n3768 35.2919
R15238 vss.n3768 vss.n3767 35.2919
R15239 vss.n3767 vss.n3748 35.2919
R15240 vss.n3757 vss.n3748 35.2919
R15241 vss.n3626 vss.n3625 35.2919
R15242 vss.n3650 vss.n3626 35.2919
R15243 vss.n3650 vss.n3649 35.2919
R15244 vss.n3649 vss.n3648 35.2919
R15245 vss.n3648 vss.n3629 35.2919
R15246 vss.n3638 vss.n3629 35.2919
R15247 vss.n6295 vss.n6294 35.2919
R15248 vss.n6299 vss.n6295 35.2919
R15249 vss.n6299 vss.n254 35.2919
R15250 vss.n15695 vss.n254 35.2919
R15251 vss.n15695 vss.n15694 35.2919
R15252 vss.n15694 vss.n15693 35.2919
R15253 vss.n15604 vss.n15603 35.2919
R15254 vss.n15605 vss.n15604 35.2919
R15255 vss.n15606 vss.n15605 35.2919
R15256 vss.n15607 vss.n15606 35.2919
R15257 vss.n15607 vss.n15586 35.2919
R15258 vss.n15611 vss.n15586 35.2919
R15259 vss.n317 vss.n316 35.2919
R15260 vss.n341 vss.n317 35.2919
R15261 vss.n341 vss.n340 35.2919
R15262 vss.n340 vss.n339 35.2919
R15263 vss.n339 vss.n320 35.2919
R15264 vss.n329 vss.n320 35.2919
R15265 vss.n3587 vss.n3579 35.2919
R15266 vss.n3599 vss.n3579 35.2919
R15267 vss.n3600 vss.n3599 35.2919
R15268 vss.n3602 vss.n3600 35.2919
R15269 vss.n3602 vss.n3601 35.2919
R15270 vss.n3601 vss.n3567 35.2919
R15271 vss.n15549 vss.n370 35.2919
R15272 vss.n15557 vss.n370 35.2919
R15273 vss.n15558 vss.n15557 35.2919
R15274 vss.n15569 vss.n15558 35.2919
R15275 vss.n15569 vss.n15568 35.2919
R15276 vss.n15568 vss.n15567 35.2919
R15277 vss.n12148 vss.n12136 35.2919
R15278 vss.n12171 vss.n12148 35.2919
R15279 vss.n12171 vss.n12170 35.2919
R15280 vss.n12170 vss.n12169 35.2919
R15281 vss.n12169 vss.n12151 35.2919
R15282 vss.n12159 vss.n12151 35.2919
R15283 vss.n11790 vss.n11789 35.2919
R15284 vss.n11789 vss.n11788 35.2919
R15285 vss.n11788 vss.n11772 35.2919
R15286 vss.n11780 vss.n11772 35.2919
R15287 vss.n11781 vss.n11780 35.2919
R15288 vss.n11784 vss.n11781 35.2919
R15289 vss.n10443 vss.n10434 35.2919
R15290 vss.n10451 vss.n10434 35.2919
R15291 vss.n10452 vss.n10451 35.2919
R15292 vss.n10464 vss.n10452 35.2919
R15293 vss.n10464 vss.n10463 35.2919
R15294 vss.n10463 vss.n10462 35.2919
R15295 vss.n10589 vss.n10579 35.2919
R15296 vss.n10597 vss.n10579 35.2919
R15297 vss.n10598 vss.n10597 35.2919
R15298 vss.n10609 vss.n10598 35.2919
R15299 vss.n10609 vss.n10608 35.2919
R15300 vss.n10608 vss.n10607 35.2919
R15301 vss.n10983 vss.n10973 35.2919
R15302 vss.n10991 vss.n10973 35.2919
R15303 vss.n10992 vss.n10991 35.2919
R15304 vss.n11003 vss.n10992 35.2919
R15305 vss.n11003 vss.n11002 35.2919
R15306 vss.n11002 vss.n11001 35.2919
R15307 vss.n10035 vss.n10034 35.2919
R15308 vss.n10034 vss.n10033 35.2919
R15309 vss.n10033 vss.n9997 35.2919
R15310 vss.n10022 vss.n9997 35.2919
R15311 vss.n10022 vss.n10021 35.2919
R15312 vss.n10021 vss.n10020 35.2919
R15313 vss.n11645 vss.n11644 35.2919
R15314 vss.n11644 vss.n11643 35.2919
R15315 vss.n11643 vss.n9953 35.2919
R15316 vss.n11627 vss.n9953 35.2919
R15317 vss.n11628 vss.n11627 35.2919
R15318 vss.n11630 vss.n11628 35.2919
R15319 vss.n9943 vss.n9933 27.0634
R15320 vss.n11669 vss.n9943 27.0634
R15321 vss.n11669 vss.n11668 27.0634
R15322 vss.n11668 vss.n11667 27.0634
R15323 vss.n11667 vss.n9946 27.0634
R15324 vss.n11656 vss.n9946 27.0634
R15325 vss.n11361 vss.n11352 27.0634
R15326 vss.n11432 vss.n11361 27.0634
R15327 vss.n11432 vss.n11431 27.0634
R15328 vss.n11431 vss.n11430 27.0634
R15329 vss.n11430 vss.n11364 27.0634
R15330 vss.n11419 vss.n11364 27.0634
R15331 vss.n11032 vss.n10070 27.0634
R15332 vss.n11310 vss.n10070 27.0634
R15333 vss.n11311 vss.n11310 27.0634
R15334 vss.n11313 vss.n11311 27.0634
R15335 vss.n11313 vss.n11312 27.0634
R15336 vss.n11312 vss.n10059 27.0634
R15337 vss.n10649 vss.n10639 27.0634
R15338 vss.n10775 vss.n10649 27.0634
R15339 vss.n10775 vss.n10774 27.0634
R15340 vss.n10774 vss.n10773 27.0634
R15341 vss.n10773 vss.n10652 27.0634
R15342 vss.n10707 vss.n10652 27.0634
R15343 vss.n13681 vss.n13680 27.0634
R15344 vss.n13680 vss.n13679 27.0634
R15345 vss.n13679 vss.n8362 27.0634
R15346 vss.n13668 vss.n8362 27.0634
R15347 vss.n13668 vss.n13667 27.0634
R15348 vss.n13667 vss.n13666 27.0634
R15349 vss.n13711 vss.n13710 27.0634
R15350 vss.n13710 vss.n13709 27.0634
R15351 vss.n13709 vss.n8326 27.0634
R15352 vss.n13409 vss.n8326 27.0634
R15353 vss.n13410 vss.n13409 27.0634
R15354 vss.n13411 vss.n13410 27.0634
R15355 vss.n13300 vss.n13299 27.0634
R15356 vss.n13299 vss.n13298 27.0634
R15357 vss.n13298 vss.n8492 27.0634
R15358 vss.n8612 vss.n8492 27.0634
R15359 vss.n8612 vss.n8611 27.0634
R15360 vss.n8611 vss.n8610 27.0634
R15361 vss.n12999 vss.n12998 27.0634
R15362 vss.n12998 vss.n12997 27.0634
R15363 vss.n12997 vss.n9178 27.0634
R15364 vss.n12986 vss.n9178 27.0634
R15365 vss.n12986 vss.n12985 27.0634
R15366 vss.n12985 vss.n12984 27.0634
R15367 vss.n13158 vss.n13157 27.0634
R15368 vss.n13157 vss.n13156 27.0634
R15369 vss.n13156 vss.n8906 27.0634
R15370 vss.n13145 vss.n8906 27.0634
R15371 vss.n13145 vss.n13144 27.0634
R15372 vss.n13144 vss.n13143 27.0634
R15373 vss.n12900 vss.n12899 27.0634
R15374 vss.n12899 vss.n12898 27.0634
R15375 vss.n12898 vss.n9307 27.0634
R15376 vss.n9380 vss.n9307 27.0634
R15377 vss.n12879 vss.n9380 27.0634
R15378 vss.n12879 vss.n12878 27.0634
R15379 vss.n12823 vss.n12822 27.0634
R15380 vss.n12822 vss.n12821 27.0634
R15381 vss.n12821 vss.n12644 27.0634
R15382 vss.n12716 vss.n12644 27.0634
R15383 vss.n12802 vss.n12716 27.0634
R15384 vss.n12802 vss.n12801 27.0634
R15385 vss.n15683 vss.n15682 27.0634
R15386 vss.n15682 vss.n284 27.0634
R15387 vss.n299 vss.n284 27.0634
R15388 vss.n15669 vss.n299 27.0634
R15389 vss.n15669 vss.n15668 27.0634
R15390 vss.n15668 vss.n15665 27.0634
R15391 vss.n6267 vss.n6266 27.0634
R15392 vss.n6266 vss.n20 27.0634
R15393 vss.n15886 vss.n20 27.0634
R15394 vss.n15886 vss.n15885 27.0634
R15395 vss.n15885 vss.n21 27.0634
R15396 vss.n15876 vss.n21 27.0634
R15397 vss.n15739 vss.n15738 27.0634
R15398 vss.n15738 vss.n15737 27.0634
R15399 vss.n15737 vss.n206 27.0634
R15400 vss.n15726 vss.n206 27.0634
R15401 vss.n15726 vss.n15725 27.0634
R15402 vss.n15725 vss.n15722 27.0634
R15403 vss.n15795 vss.n15794 27.0634
R15404 vss.n15794 vss.n15793 27.0634
R15405 vss.n15793 vss.n128 27.0634
R15406 vss.n15782 vss.n128 27.0634
R15407 vss.n15782 vss.n15781 27.0634
R15408 vss.n15781 vss.n15778 27.0634
R15409 vss.n15851 vss.n15850 27.0634
R15410 vss.n15850 vss.n15849 27.0634
R15411 vss.n15849 vss.n49 27.0634
R15412 vss.n15838 vss.n49 27.0634
R15413 vss.n15838 vss.n15837 27.0634
R15414 vss.n15837 vss.n15834 27.0634
R15415 vss.n15231 vss.n15230 27.0634
R15416 vss.n15230 vss.n15229 27.0634
R15417 vss.n15229 vss.n906 27.0634
R15418 vss.n6412 vss.n906 27.0634
R15419 vss.n6440 vss.n6412 27.0634
R15420 vss.n6441 vss.n6440 27.0634
R15421 vss.n15274 vss.n15273 27.0634
R15422 vss.n15273 vss.n15272 27.0634
R15423 vss.n15272 vss.n801 27.0634
R15424 vss.n15261 vss.n801 27.0634
R15425 vss.n15261 vss.n15260 27.0634
R15426 vss.n15260 vss.n862 27.0634
R15427 vss.n15351 vss.n15350 27.0634
R15428 vss.n15350 vss.n15349 27.0634
R15429 vss.n15349 vss.n748 27.0634
R15430 vss.n5340 vss.n748 27.0634
R15431 vss.n5368 vss.n5340 27.0634
R15432 vss.n5369 vss.n5368 27.0634
R15433 vss.n15381 vss.n15380 27.0634
R15434 vss.n15380 vss.n15379 27.0634
R15435 vss.n15379 vss.n649 27.0634
R15436 vss.n5128 vss.n649 27.0634
R15437 vss.n5156 vss.n5128 27.0634
R15438 vss.n5157 vss.n5156 27.0634
R15439 vss.n15424 vss.n15423 27.0634
R15440 vss.n15423 vss.n15422 27.0634
R15441 vss.n15422 vss.n543 27.0634
R15442 vss.n15411 vss.n543 27.0634
R15443 vss.n15411 vss.n15410 27.0634
R15444 vss.n15410 vss.n605 27.0634
R15445 vss.n15456 vss.n15455 27.0634
R15446 vss.n15455 vss.n15454 27.0634
R15447 vss.n15454 vss.n442 27.0634
R15448 vss.n4810 vss.n442 27.0634
R15449 vss.n4841 vss.n4810 27.0634
R15450 vss.n4842 vss.n4841 27.0634
R15451 vss.n4864 vss.n4311 27.0634
R15452 vss.n4874 vss.n4311 27.0634
R15453 vss.n4875 vss.n4874 27.0634
R15454 vss.n4875 vss.n4295 27.0634
R15455 vss.n4893 vss.n4295 27.0634
R15456 vss.n4894 vss.n4893 27.0634
R15457 vss.n14536 vss.n14535 27.0634
R15458 vss.n14535 vss.n14534 27.0634
R15459 vss.n14534 vss.n1685 27.0634
R15460 vss.n2520 vss.n1685 27.0634
R15461 vss.n2548 vss.n2520 27.0634
R15462 vss.n2549 vss.n2548 27.0634
R15463 vss.n14579 vss.n14578 27.0634
R15464 vss.n14578 vss.n14577 27.0634
R15465 vss.n14577 vss.n1580 27.0634
R15466 vss.n14566 vss.n1580 27.0634
R15467 vss.n14566 vss.n14565 27.0634
R15468 vss.n14565 vss.n1641 27.0634
R15469 vss.n14656 vss.n14655 27.0634
R15470 vss.n14655 vss.n14654 27.0634
R15471 vss.n14654 vss.n1527 27.0634
R15472 vss.n2754 vss.n1527 27.0634
R15473 vss.n2782 vss.n2754 27.0634
R15474 vss.n2783 vss.n2782 27.0634
R15475 vss.n14686 vss.n14685 27.0634
R15476 vss.n14685 vss.n14684 27.0634
R15477 vss.n14684 vss.n1428 27.0634
R15478 vss.n7536 vss.n1428 27.0634
R15479 vss.n7564 vss.n7536 27.0634
R15480 vss.n7565 vss.n7564 27.0634
R15481 vss.n14729 vss.n14728 27.0634
R15482 vss.n14728 vss.n14727 27.0634
R15483 vss.n14727 vss.n1322 27.0634
R15484 vss.n14716 vss.n1322 27.0634
R15485 vss.n14716 vss.n14715 27.0634
R15486 vss.n14715 vss.n1384 27.0634
R15487 vss.n14761 vss.n14760 27.0634
R15488 vss.n14760 vss.n14759 27.0634
R15489 vss.n14759 vss.n1221 27.0634
R15490 vss.n3232 vss.n1221 27.0634
R15491 vss.n3263 vss.n3232 27.0634
R15492 vss.n3264 vss.n3263 27.0634
R15493 vss.n8028 vss.n8027 27.0634
R15494 vss.n8027 vss.n8026 27.0634
R15495 vss.n8026 vss.n2365 27.0634
R15496 vss.n2437 vss.n2365 27.0634
R15497 vss.n8007 vss.n2437 27.0634
R15498 vss.n8007 vss.n8006 27.0634
R15499 vss.n14335 vss.n14334 27.0634
R15500 vss.n14334 vss.n14333 27.0634
R15501 vss.n14333 vss.n1860 27.0634
R15502 vss.n1982 vss.n1860 27.0634
R15503 vss.n1982 vss.n1981 27.0634
R15504 vss.n1981 vss.n1875 27.0634
R15505 vss.n15030 vss.n15029 27.0634
R15506 vss.n15029 vss.n15028 27.0634
R15507 vss.n15028 vss.n1081 27.0634
R15508 vss.n6527 vss.n1081 27.0634
R15509 vss.n6555 vss.n6527 27.0634
R15510 vss.n6556 vss.n6555 27.0634
R15511 vss.n15824 vss.n15823 27.0634
R15512 vss.n15823 vss.n15822 27.0634
R15513 vss.n15822 vss.n73 27.0634
R15514 vss.n106 vss.n73 27.0634
R15515 vss.n118 vss.n106 27.0634
R15516 vss.n119 vss.n118 27.0634
R15517 vss.n15768 vss.n15767 27.0634
R15518 vss.n15767 vss.n15766 27.0634
R15519 vss.n15766 vss.n152 27.0634
R15520 vss.n184 vss.n152 27.0634
R15521 vss.n196 vss.n184 27.0634
R15522 vss.n197 vss.n196 27.0634
R15523 vss.n15712 vss.n15711 27.0634
R15524 vss.n15711 vss.n15710 27.0634
R15525 vss.n15710 vss.n230 27.0634
R15526 vss.n263 vss.n230 27.0634
R15527 vss.n275 vss.n263 27.0634
R15528 vss.n276 vss.n275 27.0634
R15529 vss.n12082 vss.n12081 27.0634
R15530 vss.n12083 vss.n12082 27.0634
R15531 vss.n12083 vss.n11877 27.0634
R15532 vss.n12111 vss.n11877 27.0634
R15533 vss.n12112 vss.n12111 27.0634
R15534 vss.n12113 vss.n12112 27.0634
R15535 vss.n10390 vss.n10245 27.0634
R15536 vss.n10623 vss.n10245 27.0634
R15537 vss.n10624 vss.n10623 27.0634
R15538 vss.n10626 vss.n10624 27.0634
R15539 vss.n10626 vss.n10625 27.0634
R15540 vss.n10625 vss.n10234 27.0634
R15541 vss.n10758 vss.n10158 27.0634
R15542 vss.n11016 vss.n10158 27.0634
R15543 vss.n11017 vss.n11016 27.0634
R15544 vss.n11019 vss.n11017 27.0634
R15545 vss.n11019 vss.n11018 27.0634
R15546 vss.n11018 vss.n10147 27.0634
R15547 vss.n11325 vss.n10045 27.0634
R15548 vss.n11336 vss.n10045 27.0634
R15549 vss.n11337 vss.n11336 27.0634
R15550 vss.n11339 vss.n11337 27.0634
R15551 vss.n11339 vss.n11338 27.0634
R15552 vss.n11338 vss.n9987 27.0634
R15553 vss.n10363 vss.n10333 27.0634
R15554 vss.n10374 vss.n10333 27.0634
R15555 vss.n10375 vss.n10374 27.0634
R15556 vss.n10377 vss.n10375 27.0634
R15557 vss.n10377 vss.n10376 27.0634
R15558 vss.n10376 vss.n10276 27.0634
R15559 vss.n6579 vss.n6564 23.9548
R15560 vss.n6579 vss.n6578 23.9548
R15561 vss.n6578 vss.n6565 23.9548
R15562 vss.n6541 vss.n6535 23.9548
R15563 vss.n6535 vss.n6520 23.9548
R15564 vss.n6564 vss.n6520 23.9548
R15565 vss.n5391 vss.n5377 23.9548
R15566 vss.n5391 vss.n5390 23.9548
R15567 vss.n5390 vss.n5378 23.9548
R15568 vss.n5354 vss.n5348 23.9548
R15569 vss.n5348 vss.n5333 23.9548
R15570 vss.n5377 vss.n5333 23.9548
R15571 vss.n15403 vss.n611 23.9548
R15572 vss.n635 vss.n611 23.9548
R15573 vss.n635 vss.n633 23.9548
R15574 vss.n614 vss.n610 23.9548
R15575 vss.n15404 vss.n610 23.9548
R15576 vss.n15404 vss.n15403 23.9548
R15577 vss.n4916 vss.n4902 23.9548
R15578 vss.n4916 vss.n4915 23.9548
R15579 vss.n4915 vss.n4903 23.9548
R15580 vss.n4879 vss.n4301 23.9548
R15581 vss.n4301 vss.n4288 23.9548
R15582 vss.n4902 vss.n4288 23.9548
R15583 vss.n5179 vss.n5165 23.9548
R15584 vss.n5179 vss.n5178 23.9548
R15585 vss.n5178 vss.n5166 23.9548
R15586 vss.n5142 vss.n5136 23.9548
R15587 vss.n5136 vss.n5121 23.9548
R15588 vss.n5165 vss.n5121 23.9548
R15589 vss.n15253 vss.n868 23.9548
R15590 vss.n892 vss.n868 23.9548
R15591 vss.n892 vss.n890 23.9548
R15592 vss.n871 vss.n867 23.9548
R15593 vss.n15254 vss.n867 23.9548
R15594 vss.n15254 vss.n15253 23.9548
R15595 vss.n6463 vss.n6449 23.9548
R15596 vss.n6463 vss.n6462 23.9548
R15597 vss.n6462 vss.n6450 23.9548
R15598 vss.n6426 vss.n6420 23.9548
R15599 vss.n6420 vss.n6405 23.9548
R15600 vss.n6449 vss.n6405 23.9548
R15601 vss.n4851 vss.n4849 23.9548
R15602 vss.n4851 vss.n4850 23.9548
R15603 vss.n4850 vss.n4748 23.9548
R15604 vss.n4819 vss.n4818 23.9548
R15605 vss.n4818 vss.n4805 23.9548
R15606 vss.n4849 vss.n4805 23.9548
R15607 vss.n1974 vss.n1895 23.9548
R15608 vss.n1951 vss.n1895 23.9548
R15609 vss.n1951 vss.n1949 23.9548
R15610 vss.n1894 vss.n1880 23.9548
R15611 vss.n1975 vss.n1894 23.9548
R15612 vss.n1975 vss.n1974 23.9548
R15613 vss.n2805 vss.n2791 23.9548
R15614 vss.n2805 vss.n2804 23.9548
R15615 vss.n2804 vss.n2792 23.9548
R15616 vss.n2768 vss.n2762 23.9548
R15617 vss.n2762 vss.n2747 23.9548
R15618 vss.n2791 vss.n2747 23.9548
R15619 vss.n14708 vss.n1390 23.9548
R15620 vss.n1414 vss.n1390 23.9548
R15621 vss.n1414 vss.n1412 23.9548
R15622 vss.n1393 vss.n1389 23.9548
R15623 vss.n14709 vss.n1389 23.9548
R15624 vss.n14709 vss.n14708 23.9548
R15625 vss.n6958 vss.n2444 23.9548
R15626 vss.n6958 vss.n6957 23.9548
R15627 vss.n6957 vss.n6946 23.9548
R15628 vss.n8015 vss.n8014 23.9548
R15629 vss.n8014 vss.n2426 23.9548
R15630 vss.n2444 vss.n2426 23.9548
R15631 vss.n7587 vss.n7573 23.9548
R15632 vss.n7587 vss.n7586 23.9548
R15633 vss.n7586 vss.n7574 23.9548
R15634 vss.n7550 vss.n7544 23.9548
R15635 vss.n7544 vss.n7529 23.9548
R15636 vss.n7573 vss.n7529 23.9548
R15637 vss.n14558 vss.n1647 23.9548
R15638 vss.n1671 vss.n1647 23.9548
R15639 vss.n1671 vss.n1669 23.9548
R15640 vss.n1650 vss.n1646 23.9548
R15641 vss.n14559 vss.n1646 23.9548
R15642 vss.n14559 vss.n14558 23.9548
R15643 vss.n2570 vss.n2511 23.9548
R15644 vss.n2570 vss.n2569 23.9548
R15645 vss.n2569 vss.n2512 23.9548
R15646 vss.n2536 vss.n2530 23.9548
R15647 vss.n2530 vss.n2529 23.9548
R15648 vss.n2529 vss.n2511 23.9548
R15649 vss.n3225 vss.n3187 23.9548
R15650 vss.n3225 vss.n3224 23.9548
R15651 vss.n3224 vss.n3213 23.9548
R15652 vss.n3256 vss.n3239 23.9548
R15653 vss.n3257 vss.n3256 23.9548
R15654 vss.n3257 vss.n3187 23.9548
R15655 vss.n12122 vss.n12120 23.9548
R15656 vss.n12122 vss.n12121 23.9548
R15657 vss.n12121 vss.n11843 23.9548
R15658 vss.n11887 vss.n11886 23.9548
R15659 vss.n11886 vss.n11871 23.9548
R15660 vss.n12120 vss.n11871 23.9548
R15661 vss.n12063 vss.n8386 23.9548
R15662 vss.n12063 vss.n12012 23.9548
R15663 vss.n12012 vss.n12011 23.9548
R15664 vss.n8400 vss.n8397 23.9548
R15665 vss.n8400 vss.n8399 23.9548
R15666 vss.n8399 vss.n8386 23.9548
R15667 vss.n8602 vss.n8582 23.9548
R15668 vss.n8582 vss.n8516 23.9548
R15669 vss.n8568 vss.n8516 23.9548
R15670 vss.n8586 vss.n8583 23.9548
R15671 vss.n8601 vss.n8583 23.9548
R15672 vss.n8602 vss.n8601 23.9548
R15673 vss.n9161 vss.n8930 23.9548
R15674 vss.n9161 vss.n9110 23.9548
R15675 vss.n9110 vss.n9109 23.9548
R15676 vss.n8944 vss.n8941 23.9548
R15677 vss.n8944 vss.n8943 23.9548
R15678 vss.n8943 vss.n8930 23.9548
R15679 vss.n12837 vss.n9387 23.9548
R15680 vss.n12837 vss.n12836 23.9548
R15681 vss.n12836 vss.n9413 23.9548
R15682 vss.n12887 vss.n12886 23.9548
R15683 vss.n12886 vss.n9369 23.9548
R15684 vss.n9387 vss.n9369 23.9548
R15685 vss.n12788 vss.n12723 23.9548
R15686 vss.n12788 vss.n12787 23.9548
R15687 vss.n12787 vss.n12784 23.9548
R15688 vss.n12810 vss.n12809 23.9548
R15689 vss.n12809 vss.n12705 23.9548
R15690 vss.n12723 vss.n12705 23.9548
R15691 vss.n13314 vss.n8433 23.9548
R15692 vss.n13314 vss.n13313 23.9548
R15693 vss.n13313 vss.n8434 23.9548
R15694 vss.n12966 vss.n12959 23.9548
R15695 vss.n12968 vss.n12959 23.9548
R15696 vss.n12968 vss.n8433 23.9548
R15697 vss.n13433 vss.n13419 23.9548
R15698 vss.n13433 vss.n13432 23.9548
R15699 vss.n13432 vss.n13420 23.9548
R15700 vss.n13392 vss.n13390 23.9548
R15701 vss.n13390 vss.n13375 23.9548
R15702 vss.n13419 vss.n13375 23.9548
R15703 vss.n10347 vss.n10346 16.2531
R15704 vss.n10347 vss.n8878 16.2531
R15705 vss.n13185 vss.n8878 16.2531
R15706 vss.n13187 vss.n13185 16.2531
R15707 vss.n13187 vss.n13186 16.2531
R15708 vss.n13186 vss.n8869 16.2531
R15709 vss.n10295 vss.n10284 16.2531
R15710 vss.n10296 vss.n10295 16.2531
R15711 vss.n10315 vss.n10296 16.2531
R15712 vss.n10315 vss.n10314 16.2531
R15713 vss.n10314 vss.n10297 16.2531
R15714 vss.n10300 vss.n10297 16.2531
R15715 vss.n9928 vss.n9927 16.2531
R15716 vss.n9927 vss.n9912 16.2531
R15717 vss.n11707 vss.n9912 16.2531
R15718 vss.n11707 vss.n11706 16.2531
R15719 vss.n11706 vss.n9913 16.2531
R15720 vss.n11696 vss.n9913 16.2531
R15721 vss.n9983 vss.n9982 16.2531
R15722 vss.n9982 vss.n9967 16.2531
R15723 vss.n11470 vss.n9967 16.2531
R15724 vss.n11470 vss.n11469 16.2531
R15725 vss.n11469 vss.n9968 16.2531
R15726 vss.n11459 vss.n9968 16.2531
R15727 vss.n11379 vss.n11369 16.2531
R15728 vss.n11402 vss.n11379 16.2531
R15729 vss.n11402 vss.n11401 16.2531
R15730 vss.n11401 vss.n11400 16.2531
R15731 vss.n11400 vss.n11382 16.2531
R15732 vss.n11390 vss.n11382 16.2531
R15733 vss.n11174 vss.n11173 16.2531
R15734 vss.n11173 vss.n11158 16.2531
R15735 vss.n11201 vss.n11158 16.2531
R15736 vss.n11201 vss.n11200 16.2531
R15737 vss.n11200 vss.n11159 16.2531
R15738 vss.n11190 vss.n11159 16.2531
R15739 vss.n10143 vss.n10142 16.2531
R15740 vss.n10142 vss.n10127 16.2531
R15741 vss.n11065 vss.n10127 16.2531
R15742 vss.n11065 vss.n11064 16.2531
R15743 vss.n11064 vss.n10128 16.2531
R15744 vss.n11054 vss.n10128 16.2531
R15745 vss.n10097 vss.n10096 16.2531
R15746 vss.n10096 vss.n10081 16.2531
R15747 vss.n10125 vss.n10081 16.2531
R15748 vss.n10125 vss.n10124 16.2531
R15749 vss.n10124 vss.n10082 16.2531
R15750 vss.n10114 vss.n10082 16.2531
R15751 vss.n10744 vss.n10713 16.2531
R15752 vss.n10745 vss.n10744 16.2531
R15753 vss.n10745 vss.n10168 16.2531
R15754 vss.n10725 vss.n10168 16.2531
R15755 vss.n10732 vss.n10725 16.2531
R15756 vss.n10733 vss.n10732 16.2531
R15757 vss.n10230 vss.n10229 16.2531
R15758 vss.n10229 vss.n10214 16.2531
R15759 vss.n10813 vss.n10214 16.2531
R15760 vss.n10813 vss.n10812 16.2531
R15761 vss.n10812 vss.n10215 16.2531
R15762 vss.n10802 vss.n10215 16.2531
R15763 vss.n10667 vss.n10657 16.2531
R15764 vss.n10690 vss.n10667 16.2531
R15765 vss.n10690 vss.n10689 16.2531
R15766 vss.n10689 vss.n10688 16.2531
R15767 vss.n10688 vss.n10670 16.2531
R15768 vss.n10678 vss.n10670 16.2531
R15769 vss.n10272 vss.n10271 16.2531
R15770 vss.n10271 vss.n10256 16.2531
R15771 vss.n10423 vss.n10256 16.2531
R15772 vss.n10423 vss.n10422 16.2531
R15773 vss.n10422 vss.n10257 16.2531
R15774 vss.n10412 vss.n10257 16.2531
R15775 vss.n10488 vss.n10487 16.2531
R15776 vss.n10487 vss.n10472 16.2531
R15777 vss.n10517 vss.n10472 16.2531
R15778 vss.n10517 vss.n10516 16.2531
R15779 vss.n10516 vss.n10473 16.2531
R15780 vss.n10504 vss.n10473 16.2531
R15781 vss.n10536 vss.n10535 16.2531
R15782 vss.n10535 vss.n10520 16.2531
R15783 vss.n10564 vss.n10520 16.2531
R15784 vss.n10564 vss.n10563 16.2531
R15785 vss.n10563 vss.n10521 16.2531
R15786 vss.n10553 vss.n10521 16.2531
R15787 vss.n10834 vss.n10833 16.2531
R15788 vss.n10833 vss.n10818 16.2531
R15789 vss.n10863 vss.n10818 16.2531
R15790 vss.n10863 vss.n10862 16.2531
R15791 vss.n10862 vss.n10819 16.2531
R15792 vss.n10851 vss.n10819 16.2531
R15793 vss.n10882 vss.n10881 16.2531
R15794 vss.n10881 vss.n10866 16.2531
R15795 vss.n10911 vss.n10866 16.2531
R15796 vss.n10911 vss.n10910 16.2531
R15797 vss.n10910 vss.n10867 16.2531
R15798 vss.n10898 vss.n10867 16.2531
R15799 vss.n10930 vss.n10929 16.2531
R15800 vss.n10929 vss.n10914 16.2531
R15801 vss.n10958 vss.n10914 16.2531
R15802 vss.n10958 vss.n10957 16.2531
R15803 vss.n10957 vss.n10915 16.2531
R15804 vss.n10947 vss.n10915 16.2531
R15805 vss.n11269 vss.n11268 16.2531
R15806 vss.n11268 vss.n11253 16.2531
R15807 vss.n11298 vss.n11253 16.2531
R15808 vss.n11298 vss.n11297 16.2531
R15809 vss.n11297 vss.n11254 16.2531
R15810 vss.n11286 vss.n11254 16.2531
R15811 vss.n11221 vss.n11220 16.2531
R15812 vss.n11220 vss.n11205 16.2531
R15813 vss.n11250 vss.n11205 16.2531
R15814 vss.n11250 vss.n11249 16.2531
R15815 vss.n11249 vss.n11206 16.2531
R15816 vss.n11237 vss.n11206 16.2531
R15817 vss.n11127 vss.n11126 16.2531
R15818 vss.n11126 vss.n11111 16.2531
R15819 vss.n11155 vss.n11111 16.2531
R15820 vss.n11155 vss.n11154 16.2531
R15821 vss.n11154 vss.n11112 16.2531
R15822 vss.n11144 vss.n11112 16.2531
R15823 vss.n11580 vss.n11579 16.2531
R15824 vss.n11579 vss.n11564 16.2531
R15825 vss.n11609 vss.n11564 16.2531
R15826 vss.n11609 vss.n11608 16.2531
R15827 vss.n11608 vss.n11565 16.2531
R15828 vss.n11597 vss.n11565 16.2531
R15829 vss.n11532 vss.n11531 16.2531
R15830 vss.n11531 vss.n11516 16.2531
R15831 vss.n11561 vss.n11516 16.2531
R15832 vss.n11561 vss.n11560 16.2531
R15833 vss.n11560 vss.n11517 16.2531
R15834 vss.n11548 vss.n11517 16.2531
R15835 vss.n9899 vss.n9891 16.2531
R15836 vss.n9910 vss.n9891 16.2531
R15837 vss.n11711 vss.n9910 16.2531
R15838 vss.n11713 vss.n11711 16.2531
R15839 vss.n11713 vss.n11712 16.2531
R15840 vss.n11712 vss.n9882 16.2531
R15841 vss.n11838 vss.n11837 16.2531
R15842 vss.n11837 vss.n11804 16.2531
R15843 vss.n12187 vss.n11804 16.2531
R15844 vss.n12187 vss.n12186 16.2531
R15845 vss.n12186 vss.n11805 16.2531
R15846 vss.n11828 vss.n11805 16.2531
R15847 vss.n11917 vss.n11916 16.2531
R15848 vss.n11918 vss.n11917 16.2531
R15849 vss.n11918 vss.n11894 16.2531
R15850 vss.n11929 vss.n11894 16.2531
R15851 vss.n11930 vss.n11929 16.2531
R15852 vss.n11931 vss.n11930 16.2531
R15853 vss.n9271 vss.n9270 16.2531
R15854 vss.n9270 vss.n8885 16.2531
R15855 vss.n13176 vss.n8885 16.2531
R15856 vss.n13176 vss.n13175 16.2531
R15857 vss.n13175 vss.n8886 16.2531
R15858 vss.n13165 vss.n8886 16.2531
R15859 vss.n12399 vss.n12398 16.2531
R15860 vss.n12398 vss.n12383 16.2531
R15861 vss.n12427 vss.n12383 16.2531
R15862 vss.n12427 vss.n12426 16.2531
R15863 vss.n12426 vss.n12384 16.2531
R15864 vss.n12416 vss.n12384 16.2531
R15865 vss.n9669 vss.n9668 16.2531
R15866 vss.n9668 vss.n9667 16.2531
R15867 vss.n9667 vss.n9630 16.2531
R15868 vss.n9657 vss.n9630 16.2531
R15869 vss.n9657 vss.n9656 16.2531
R15870 vss.n9656 vss.n9655 16.2531
R15871 vss.n9619 vss.n9618 16.2531
R15872 vss.n9618 vss.n9603 16.2531
R15873 vss.n12380 vss.n9603 16.2531
R15874 vss.n12380 vss.n12379 16.2531
R15875 vss.n12379 vss.n9604 16.2531
R15876 vss.n12369 vss.n9604 16.2531
R15877 vss.n8636 vss.n8635 16.2531
R15878 vss.n8635 vss.n8620 16.2531
R15879 vss.n13288 vss.n8620 16.2531
R15880 vss.n13288 vss.n13287 16.2531
R15881 vss.n13287 vss.n8621 16.2531
R15882 vss.n13277 vss.n8621 16.2531
R15883 vss.n12281 vss.n12280 16.2531
R15884 vss.n12280 vss.n12265 16.2531
R15885 vss.n12309 vss.n12265 16.2531
R15886 vss.n12309 vss.n12308 16.2531
R15887 vss.n12308 vss.n12266 16.2531
R15888 vss.n12298 vss.n12266 16.2531
R15889 vss.n9798 vss.n9797 16.2531
R15890 vss.n9797 vss.n9796 16.2531
R15891 vss.n9796 vss.n9760 16.2531
R15892 vss.n9786 vss.n9760 16.2531
R15893 vss.n9786 vss.n9785 16.2531
R15894 vss.n9785 vss.n9784 16.2531
R15895 vss.n9749 vss.n9748 16.2531
R15896 vss.n9748 vss.n9733 16.2531
R15897 vss.n12262 vss.n9733 16.2531
R15898 vss.n12262 vss.n12261 16.2531
R15899 vss.n12261 vss.n9734 16.2531
R15900 vss.n12251 vss.n9734 16.2531
R15901 vss.n8753 vss.n8752 16.2531
R15902 vss.n8752 vss.n8341 16.2531
R15903 vss.n13699 vss.n8341 16.2531
R15904 vss.n13699 vss.n13698 16.2531
R15905 vss.n13698 vss.n8342 16.2531
R15906 vss.n13688 vss.n8342 16.2531
R15907 vss.n11990 vss.n11989 16.2531
R15908 vss.n11991 vss.n11990 16.2531
R15909 vss.n11991 vss.n9858 16.2531
R15910 vss.n12002 vss.n9858 16.2531
R15911 vss.n12003 vss.n12002 16.2531
R15912 vss.n12004 vss.n12003 16.2531
R15913 vss.n9878 vss.n9877 16.2531
R15914 vss.n9877 vss.n9862 16.2531
R15915 vss.n11756 vss.n9862 16.2531
R15916 vss.n11756 vss.n11755 16.2531
R15917 vss.n11755 vss.n9863 16.2531
R15918 vss.n11745 vss.n9863 16.2531
R15919 vss.n12232 vss.n12231 16.2531
R15920 vss.n12231 vss.n12230 16.2531
R15921 vss.n12230 vss.n12195 16.2531
R15922 vss.n12220 vss.n12195 16.2531
R15923 vss.n12220 vss.n12219 16.2531
R15924 vss.n12219 vss.n12218 16.2531
R15925 vss.n8801 vss.n8800 16.2531
R15926 vss.n8800 vss.n8799 16.2531
R15927 vss.n8799 vss.n8764 16.2531
R15928 vss.n8789 vss.n8764 16.2531
R15929 vss.n8789 vss.n8788 16.2531
R15930 vss.n8788 vss.n8787 16.2531
R15931 vss.n8732 vss.n8731 16.2531
R15932 vss.n8731 vss.n8730 16.2531
R15933 vss.n8730 vss.n8695 16.2531
R15934 vss.n8720 vss.n8695 16.2531
R15935 vss.n8720 vss.n8719 16.2531
R15936 vss.n8719 vss.n8718 16.2531
R15937 vss.n9849 vss.n9848 16.2531
R15938 vss.n9848 vss.n9847 16.2531
R15939 vss.n9847 vss.n9811 16.2531
R15940 vss.n9837 vss.n9811 16.2531
R15941 vss.n9837 vss.n9836 16.2531
R15942 vss.n9836 vss.n9835 16.2531
R15943 vss.n12350 vss.n12349 16.2531
R15944 vss.n12349 vss.n12348 16.2531
R15945 vss.n12348 vss.n12313 16.2531
R15946 vss.n12338 vss.n12313 16.2531
R15947 vss.n12338 vss.n12337 16.2531
R15948 vss.n12337 vss.n12336 16.2531
R15949 vss.n8682 vss.n8681 16.2531
R15950 vss.n8681 vss.n8680 16.2531
R15951 vss.n8680 vss.n8645 16.2531
R15952 vss.n8670 vss.n8645 16.2531
R15953 vss.n8670 vss.n8669 16.2531
R15954 vss.n8669 vss.n8668 16.2531
R15955 vss.n12922 vss.n12921 16.2531
R15956 vss.n12923 vss.n12922 16.2531
R15957 vss.n12923 vss.n9187 16.2531
R15958 vss.n12934 vss.n9187 16.2531
R15959 vss.n12935 vss.n12934 16.2531
R15960 vss.n12936 vss.n12935 16.2531
R15961 vss.n9721 vss.n9720 16.2531
R15962 vss.n9720 vss.n9719 16.2531
R15963 vss.n9719 vss.n9682 16.2531
R15964 vss.n9709 vss.n9682 16.2531
R15965 vss.n9709 vss.n9708 16.2531
R15966 vss.n9708 vss.n9707 16.2531
R15967 vss.n12469 vss.n12468 16.2531
R15968 vss.n12468 vss.n12467 16.2531
R15969 vss.n12467 vss.n12432 16.2531
R15970 vss.n12457 vss.n12432 16.2531
R15971 vss.n12457 vss.n12456 16.2531
R15972 vss.n12456 vss.n12455 16.2531
R15973 vss.n9252 vss.n9251 16.2531
R15974 vss.n9251 vss.n9250 16.2531
R15975 vss.n9250 vss.n9215 16.2531
R15976 vss.n9240 vss.n9215 16.2531
R15977 vss.n9240 vss.n9239 16.2531
R15978 vss.n9239 vss.n9238 16.2531
R15979 vss.n9340 vss.n9339 16.2531
R15980 vss.n9341 vss.n9340 16.2531
R15981 vss.n9341 vss.n9317 16.2531
R15982 vss.n9352 vss.n9317 16.2531
R15983 vss.n9353 vss.n9352 16.2531
R15984 vss.n9354 vss.n9353 16.2531
R15985 vss.n12526 vss.n12525 16.2531
R15986 vss.n12527 vss.n12526 16.2531
R15987 vss.n12527 vss.n12503 16.2531
R15988 vss.n12538 vss.n12503 16.2531
R15989 vss.n12539 vss.n12538 16.2531
R15990 vss.n12540 vss.n12539 16.2531
R15991 vss.n9490 vss.n9489 16.2531
R15992 vss.n9489 vss.n9474 16.2531
R15993 vss.n12499 vss.n9474 16.2531
R15994 vss.n12499 vss.n12498 16.2531
R15995 vss.n12498 vss.n9475 16.2531
R15996 vss.n12488 vss.n9475 16.2531
R15997 vss.n9539 vss.n9538 16.2531
R15998 vss.n9538 vss.n9537 16.2531
R15999 vss.n9537 vss.n9501 16.2531
R16000 vss.n9527 vss.n9501 16.2531
R16001 vss.n9527 vss.n9526 16.2531
R16002 vss.n9526 vss.n9525 16.2531
R16003 vss.n9440 vss.n9439 16.2531
R16004 vss.n9439 vss.n9424 16.2531
R16005 vss.n9469 vss.n9424 16.2531
R16006 vss.n9469 vss.n9468 16.2531
R16007 vss.n9468 vss.n9425 16.2531
R16008 vss.n9457 vss.n9425 16.2531
R16009 vss.n12676 vss.n12675 16.2531
R16010 vss.n12677 vss.n12676 16.2531
R16011 vss.n12677 vss.n12653 16.2531
R16012 vss.n12688 vss.n12653 16.2531
R16013 vss.n12689 vss.n12688 16.2531
R16014 vss.n12690 vss.n12689 16.2531
R16015 vss.n9591 vss.n9590 16.2531
R16016 vss.n9590 vss.n9589 16.2531
R16017 vss.n9589 vss.n9553 16.2531
R16018 vss.n9579 vss.n9553 16.2531
R16019 vss.n9579 vss.n9578 16.2531
R16020 vss.n9578 vss.n9577 16.2531
R16021 vss.n10186 vss.n10185 16.2531
R16022 vss.n10185 vss.n10170 16.2531
R16023 vss.n10212 vss.n10170 16.2531
R16024 vss.n10212 vss.n10211 16.2531
R16025 vss.n10211 vss.n10171 16.2531
R16026 vss.n10201 vss.n10171 16.2531
R16027 vss.n11083 vss.n11082 16.2531
R16028 vss.n11082 vss.n11067 16.2531
R16029 vss.n11109 vss.n11067 16.2531
R16030 vss.n11109 vss.n11108 16.2531
R16031 vss.n11108 vss.n11068 16.2531
R16032 vss.n11098 vss.n11068 16.2531
R16033 vss.n11488 vss.n11487 16.2531
R16034 vss.n11487 vss.n11472 16.2531
R16035 vss.n11514 vss.n11472 16.2531
R16036 vss.n11514 vss.n11513 16.2531
R16037 vss.n11513 vss.n11473 16.2531
R16038 vss.n11503 vss.n11473 16.2531
R16039 vss.n13231 vss.n13230 16.2531
R16040 vss.n13232 vss.n13231 16.2531
R16041 vss.n13232 vss.n8816 16.2531
R16042 vss.n13243 vss.n8816 16.2531
R16043 vss.n13244 vss.n13243 16.2531
R16044 vss.n13245 vss.n13244 16.2531
R16045 vss.n15638 vss.n15637 16.2531
R16046 vss.n15637 vss.n15636 16.2531
R16047 vss.n15636 vss.n15622 16.2531
R16048 vss.n15654 vss.n15622 16.2531
R16049 vss.n15654 vss.n15653 16.2531
R16050 vss.n15653 vss.n15652 16.2531
R16051 vss.n3984 vss.n3983 16.2531
R16052 vss.n3983 vss.n1 16.2531
R16053 vss.n15903 vss.n1 16.2531
R16054 vss.n15903 vss.n15902 16.2531
R16055 vss.n15902 vss.n2 16.2531
R16056 vss.n15892 vss.n2 16.2531
R16057 vss.n5649 vss.n5648 16.2531
R16058 vss.n5648 vss.n5633 16.2531
R16059 vss.n5676 vss.n5633 16.2531
R16060 vss.n5676 vss.n5675 16.2531
R16061 vss.n5675 vss.n5634 16.2531
R16062 vss.n5665 vss.n5634 16.2531
R16063 vss.n3725 vss.n3724 16.2531
R16064 vss.n3724 vss.n166 16.2531
R16065 vss.n15756 vss.n166 16.2531
R16066 vss.n15756 vss.n15755 16.2531
R16067 vss.n15755 vss.n167 16.2531
R16068 vss.n15745 vss.n167 16.2531
R16069 vss.n3706 vss.n3705 16.2531
R16070 vss.n3705 vss.n3704 16.2531
R16071 vss.n3704 vss.n3669 16.2531
R16072 vss.n3694 vss.n3669 16.2531
R16073 vss.n3694 vss.n3693 16.2531
R16074 vss.n3693 vss.n3692 16.2531
R16075 vss.n5841 vss.n5840 16.2531
R16076 vss.n5840 vss.n5825 16.2531
R16077 vss.n5868 vss.n5825 16.2531
R16078 vss.n5868 vss.n5867 16.2531
R16079 vss.n5867 vss.n5826 16.2531
R16080 vss.n5857 vss.n5826 16.2531
R16081 vss.n3844 vss.n3843 16.2531
R16082 vss.n3843 vss.n88 16.2531
R16083 vss.n15812 vss.n88 16.2531
R16084 vss.n15812 vss.n15811 16.2531
R16085 vss.n15811 vss.n89 16.2531
R16086 vss.n15801 vss.n89 16.2531
R16087 vss.n3825 vss.n3824 16.2531
R16088 vss.n3824 vss.n3823 16.2531
R16089 vss.n3823 vss.n3788 16.2531
R16090 vss.n3813 vss.n3788 16.2531
R16091 vss.n3813 vss.n3812 16.2531
R16092 vss.n3812 vss.n3811 16.2531
R16093 vss.n3944 vss.n3943 16.2531
R16094 vss.n3943 vss.n3942 16.2531
R16095 vss.n3942 vss.n3907 16.2531
R16096 vss.n3932 vss.n3907 16.2531
R16097 vss.n3932 vss.n3931 16.2531
R16098 vss.n3931 vss.n3930 16.2531
R16099 vss.n6081 vss.n6080 16.2531
R16100 vss.n6080 vss.n6065 16.2531
R16101 vss.n6108 vss.n6065 16.2531
R16102 vss.n6108 vss.n6107 16.2531
R16103 vss.n6107 vss.n6066 16.2531
R16104 vss.n6097 vss.n6066 16.2531
R16105 vss.n6033 vss.n6032 16.2531
R16106 vss.n6032 vss.n6017 16.2531
R16107 vss.n6061 vss.n6017 16.2531
R16108 vss.n6061 vss.n6060 16.2531
R16109 vss.n6060 vss.n6018 16.2531
R16110 vss.n6049 vss.n6018 16.2531
R16111 vss.n6196 vss.n6195 16.2531
R16112 vss.n6195 vss.n6194 16.2531
R16113 vss.n6194 vss.n6158 16.2531
R16114 vss.n6184 vss.n6158 16.2531
R16115 vss.n6184 vss.n6183 16.2531
R16116 vss.n6183 vss.n6182 16.2531
R16117 vss.n5751 vss.n5750 16.2531
R16118 vss.n5750 vss.n5730 16.2531
R16119 vss.n5774 vss.n5730 16.2531
R16120 vss.n5774 vss.n5773 16.2531
R16121 vss.n5773 vss.n5731 16.2531
R16122 vss.n5763 vss.n5731 16.2531
R16123 vss.n5793 vss.n5792 16.2531
R16124 vss.n5792 vss.n5777 16.2531
R16125 vss.n5821 vss.n5777 16.2531
R16126 vss.n5821 vss.n5820 16.2531
R16127 vss.n5820 vss.n5778 16.2531
R16128 vss.n5809 vss.n5778 16.2531
R16129 vss.n5957 vss.n5956 16.2531
R16130 vss.n5956 vss.n5955 16.2531
R16131 vss.n5955 vss.n5919 16.2531
R16132 vss.n5945 vss.n5919 16.2531
R16133 vss.n5945 vss.n5944 16.2531
R16134 vss.n5944 vss.n5943 16.2531
R16135 vss.n5563 vss.n5562 16.2531
R16136 vss.n5562 vss.n5542 16.2531
R16137 vss.n5586 vss.n5542 16.2531
R16138 vss.n5586 vss.n5585 16.2531
R16139 vss.n5585 vss.n5543 16.2531
R16140 vss.n5575 vss.n5543 16.2531
R16141 vss.n5719 vss.n5718 16.2531
R16142 vss.n5718 vss.n5717 16.2531
R16143 vss.n5717 vss.n5681 16.2531
R16144 vss.n5707 vss.n5681 16.2531
R16145 vss.n5707 vss.n5706 16.2531
R16146 vss.n5706 vss.n5705 16.2531
R16147 vss.n6329 vss.n6328 16.2531
R16148 vss.n6328 vss.n6327 16.2531
R16149 vss.n6327 vss.n3542 16.2531
R16150 vss.n6317 vss.n3542 16.2531
R16151 vss.n6317 vss.n6316 16.2531
R16152 vss.n6316 vss.n6315 16.2531
R16153 vss.n5608 vss.n5607 16.2531
R16154 vss.n5607 vss.n5589 16.2531
R16155 vss.n5631 vss.n5589 16.2531
R16156 vss.n5631 vss.n5630 16.2531
R16157 vss.n5630 vss.n5590 16.2531
R16158 vss.n5620 vss.n5590 16.2531
R16159 vss.n5910 vss.n5909 16.2531
R16160 vss.n5909 vss.n5908 16.2531
R16161 vss.n5908 vss.n5872 16.2531
R16162 vss.n5898 vss.n5872 16.2531
R16163 vss.n5898 vss.n5897 16.2531
R16164 vss.n5897 vss.n5896 16.2531
R16165 vss.n6149 vss.n6148 16.2531
R16166 vss.n6148 vss.n6147 16.2531
R16167 vss.n6147 vss.n6111 16.2531
R16168 vss.n6137 vss.n6111 16.2531
R16169 vss.n6137 vss.n6136 16.2531
R16170 vss.n6136 vss.n6135 16.2531
R16171 vss.n5991 vss.n5990 16.2531
R16172 vss.n5990 vss.n5970 16.2531
R16173 vss.n6014 vss.n5970 16.2531
R16174 vss.n6014 vss.n6013 16.2531
R16175 vss.n6013 vss.n5971 16.2531
R16176 vss.n6003 vss.n5971 16.2531
R16177 vss.n4379 vss.n4369 16.2531
R16178 vss.n4544 vss.n4379 16.2531
R16179 vss.n4544 vss.n4543 16.2531
R16180 vss.n4543 vss.n4400 16.2531
R16181 vss.n4400 vss.n4382 16.2531
R16182 vss.n4390 vss.n4382 16.2531
R16183 vss.n4464 vss.n4463 16.2531
R16184 vss.n4463 vss.n4448 16.2531
R16185 vss.n4492 vss.n4448 16.2531
R16186 vss.n4492 vss.n4491 16.2531
R16187 vss.n4491 vss.n4449 16.2531
R16188 vss.n4480 vss.n4449 16.2531
R16189 vss.n4511 vss.n4510 16.2531
R16190 vss.n4510 vss.n4495 16.2531
R16191 vss.n4539 vss.n4495 16.2531
R16192 vss.n4539 vss.n4538 16.2531
R16193 vss.n4538 vss.n4496 16.2531
R16194 vss.n4528 vss.n4496 16.2531
R16195 vss.n6632 vss.n6631 16.2531
R16196 vss.n6631 vss.n6616 16.2531
R16197 vss.n6659 vss.n6616 16.2531
R16198 vss.n6659 vss.n6658 16.2531
R16199 vss.n6658 vss.n6617 16.2531
R16200 vss.n6648 vss.n6617 16.2531
R16201 vss.n6514 vss.n6513 16.2531
R16202 vss.n6513 vss.n6498 16.2531
R16203 vss.n6611 vss.n6498 16.2531
R16204 vss.n6611 vss.n6610 16.2531
R16205 vss.n6610 vss.n6499 16.2531
R16206 vss.n6600 vss.n6499 16.2531
R16207 vss.n5230 vss.n5229 16.2531
R16208 vss.n5229 vss.n5214 16.2531
R16209 vss.n5257 vss.n5214 16.2531
R16210 vss.n5257 vss.n5256 16.2531
R16211 vss.n5256 vss.n5215 16.2531
R16212 vss.n5246 vss.n5215 16.2531
R16213 vss.n5275 vss.n5274 16.2531
R16214 vss.n5274 vss.n5259 16.2531
R16215 vss.n5304 vss.n5259 16.2531
R16216 vss.n5304 vss.n5303 16.2531
R16217 vss.n5303 vss.n5260 16.2531
R16218 vss.n5292 vss.n5260 16.2531
R16219 vss.n4026 vss.n4018 16.2531
R16220 vss.n4037 vss.n4018 16.2531
R16221 vss.n5521 vss.n4037 16.2531
R16222 vss.n5522 vss.n5521 16.2531
R16223 vss.n5522 vss.n4008 16.2531
R16224 vss.n5532 vss.n4008 16.2531
R16225 vss.n5490 vss.n5489 16.2531
R16226 vss.n5489 vss.n5474 16.2531
R16227 vss.n5518 vss.n5474 16.2531
R16228 vss.n5518 vss.n5517 16.2531
R16229 vss.n5517 vss.n5475 16.2531
R16230 vss.n5507 vss.n5475 16.2531
R16231 vss.n4055 vss.n4054 16.2531
R16232 vss.n4054 vss.n4039 16.2531
R16233 vss.n4081 vss.n4039 16.2531
R16234 vss.n4081 vss.n4080 16.2531
R16235 vss.n4080 vss.n4040 16.2531
R16236 vss.n4070 vss.n4040 16.2531
R16237 vss.n5442 vss.n5441 16.2531
R16238 vss.n5441 vss.n5426 16.2531
R16239 vss.n5469 vss.n5426 16.2531
R16240 vss.n5469 vss.n5468 16.2531
R16241 vss.n5468 vss.n5427 16.2531
R16242 vss.n5458 vss.n5427 16.2531
R16243 vss.n5327 vss.n5326 16.2531
R16244 vss.n5326 vss.n5311 16.2531
R16245 vss.n5422 vss.n5311 16.2531
R16246 vss.n5422 vss.n5421 16.2531
R16247 vss.n5421 vss.n5312 16.2531
R16248 vss.n5411 vss.n5312 16.2531
R16249 vss.n4145 vss.n4144 16.2531
R16250 vss.n4144 vss.n4129 16.2531
R16251 vss.n4172 vss.n4129 16.2531
R16252 vss.n4172 vss.n4171 16.2531
R16253 vss.n4171 vss.n4130 16.2531
R16254 vss.n4161 vss.n4130 16.2531
R16255 vss.n5064 vss.n5063 16.2531
R16256 vss.n5063 vss.n5048 16.2531
R16257 vss.n5092 vss.n5048 16.2531
R16258 vss.n5092 vss.n5091 16.2531
R16259 vss.n5091 vss.n5049 16.2531
R16260 vss.n5081 vss.n5049 16.2531
R16261 vss.n4189 vss.n4188 16.2531
R16262 vss.n4188 vss.n4174 16.2531
R16263 vss.n4218 vss.n4174 16.2531
R16264 vss.n4218 vss.n4217 16.2531
R16265 vss.n4217 vss.n4216 16.2531
R16266 vss.n4216 vss.n4215 16.2531
R16267 vss.n5016 vss.n5015 16.2531
R16268 vss.n5015 vss.n5000 16.2531
R16269 vss.n5044 vss.n5000 16.2531
R16270 vss.n5044 vss.n5043 16.2531
R16271 vss.n5043 vss.n5001 16.2531
R16272 vss.n5033 vss.n5001 16.2531
R16273 vss.n4236 vss.n4235 16.2531
R16274 vss.n4235 vss.n4220 16.2531
R16275 vss.n4262 vss.n4220 16.2531
R16276 vss.n4262 vss.n4261 16.2531
R16277 vss.n4261 vss.n4221 16.2531
R16278 vss.n4251 vss.n4221 16.2531
R16279 vss.n4968 vss.n4967 16.2531
R16280 vss.n4967 vss.n4952 16.2531
R16281 vss.n4995 vss.n4952 16.2531
R16282 vss.n4995 vss.n4994 16.2531
R16283 vss.n4994 vss.n4953 16.2531
R16284 vss.n4984 vss.n4953 16.2531
R16285 vss.n4099 vss.n4098 16.2531
R16286 vss.n4098 vss.n4083 16.2531
R16287 vss.n4126 vss.n4083 16.2531
R16288 vss.n4126 vss.n4125 16.2531
R16289 vss.n4125 vss.n4084 16.2531
R16290 vss.n4115 vss.n4084 16.2531
R16291 vss.n4282 vss.n4281 16.2531
R16292 vss.n4281 vss.n4266 16.2531
R16293 vss.n4947 vss.n4266 16.2531
R16294 vss.n4947 vss.n4946 16.2531
R16295 vss.n4946 vss.n4267 16.2531
R16296 vss.n4936 vss.n4267 16.2531
R16297 vss.n5115 vss.n5114 16.2531
R16298 vss.n5114 vss.n5099 16.2531
R16299 vss.n5210 vss.n5099 16.2531
R16300 vss.n5210 vss.n5209 16.2531
R16301 vss.n5209 vss.n5100 16.2531
R16302 vss.n5199 vss.n5100 16.2531
R16303 vss.n3358 vss.n3357 16.2531
R16304 vss.n3357 vss.n3342 16.2531
R16305 vss.n3385 vss.n3342 16.2531
R16306 vss.n3385 vss.n3384 16.2531
R16307 vss.n3384 vss.n3343 16.2531
R16308 vss.n3374 vss.n3343 16.2531
R16309 vss.n3405 vss.n3404 16.2531
R16310 vss.n3404 vss.n3389 16.2531
R16311 vss.n3432 vss.n3389 16.2531
R16312 vss.n3432 vss.n3431 16.2531
R16313 vss.n3431 vss.n3390 16.2531
R16314 vss.n3421 vss.n3390 16.2531
R16315 vss.n3461 vss.n3460 16.2531
R16316 vss.n3460 vss.n3453 16.2531
R16317 vss.n3453 vss.n3433 16.2531
R16318 vss.n3474 vss.n3433 16.2531
R16319 vss.n3474 vss.n3473 16.2531
R16320 vss.n3473 vss.n3444 16.2531
R16321 vss.n6347 vss.n6343 16.2531
R16322 vss.n6347 vss.n3435 16.2531
R16323 vss.n6374 vss.n3435 16.2531
R16324 vss.n6374 vss.n6373 16.2531
R16325 vss.n6373 vss.n6372 16.2531
R16326 vss.n6372 vss.n6371 16.2531
R16327 vss.n3508 vss.n3500 16.2531
R16328 vss.n3518 vss.n3500 16.2531
R16329 vss.n3519 vss.n3518 16.2531
R16330 vss.n3521 vss.n3519 16.2531
R16331 vss.n3521 vss.n3520 16.2531
R16332 vss.n3520 vss.n3491 16.2531
R16333 vss.n6399 vss.n6398 16.2531
R16334 vss.n6398 vss.n6383 16.2531
R16335 vss.n6494 vss.n6383 16.2531
R16336 vss.n6494 vss.n6493 16.2531
R16337 vss.n6493 vss.n6384 16.2531
R16338 vss.n6483 vss.n6384 16.2531
R16339 vss.n6700 vss.n6699 16.2531
R16340 vss.n6699 vss.n6698 16.2531
R16341 vss.n6698 vss.n6663 16.2531
R16342 vss.n6679 vss.n6663 16.2531
R16343 vss.n6686 vss.n6679 16.2531
R16344 vss.n6686 vss.n6685 16.2531
R16345 vss.n4418 vss.n4417 16.2531
R16346 vss.n4417 vss.n4402 16.2531
R16347 vss.n4445 vss.n4402 16.2531
R16348 vss.n4445 vss.n4444 16.2531
R16349 vss.n4444 vss.n4403 16.2531
R16350 vss.n4434 vss.n4403 16.2531
R16351 vss.n4766 vss.n4756 16.2531
R16352 vss.n4790 vss.n4766 16.2531
R16353 vss.n4790 vss.n4789 16.2531
R16354 vss.n4789 vss.n4787 16.2531
R16355 vss.n4787 vss.n4769 16.2531
R16356 vss.n4777 vss.n4769 16.2531
R16357 vss.n3291 vss.n3290 16.2531
R16358 vss.n3290 vss.n3275 16.2531
R16359 vss.n6738 vss.n3275 16.2531
R16360 vss.n6738 vss.n6737 16.2531
R16361 vss.n6737 vss.n3276 16.2531
R16362 vss.n6727 vss.n3276 16.2531
R16363 vss.n15524 vss.n15523 16.2531
R16364 vss.n15525 vss.n15524 16.2531
R16365 vss.n15525 vss.n15501 16.2531
R16366 vss.n15536 vss.n15501 16.2531
R16367 vss.n15537 vss.n15536 16.2531
R16368 vss.n15538 vss.n15537 16.2531
R16369 vss.n14865 vss.n14864 16.2531
R16370 vss.n14864 vss.n390 16.2531
R16371 vss.n15498 vss.n390 16.2531
R16372 vss.n15498 vss.n15497 16.2531
R16373 vss.n15497 vss.n391 16.2531
R16374 vss.n15487 vss.n391 16.2531
R16375 vss.n15013 vss.n15012 16.2531
R16376 vss.n15012 vss.n14979 16.2531
R16377 vss.n15018 vss.n14979 16.2531
R16378 vss.n15018 vss.n15017 16.2531
R16379 vss.n15017 vss.n14980 16.2531
R16380 vss.n15003 vss.n14980 16.2531
R16381 vss.n1058 vss.n1057 16.2531
R16382 vss.n1057 vss.n1042 16.2531
R16383 vss.n15048 vss.n1042 16.2531
R16384 vss.n15048 vss.n15047 16.2531
R16385 vss.n15047 vss.n1043 16.2531
R16386 vss.n15037 vss.n1043 16.2531
R16387 vss.n14905 vss.n14904 16.2531
R16388 vss.n14904 vss.n14889 16.2531
R16389 vss.n14934 vss.n14889 16.2531
R16390 vss.n14934 vss.n14933 16.2531
R16391 vss.n14933 vss.n14890 16.2531
R16392 vss.n14923 vss.n14890 16.2531
R16393 vss.n520 vss.n519 16.2531
R16394 vss.n519 vss.n504 16.2531
R16395 vss.n15442 vss.n504 16.2531
R16396 vss.n15442 vss.n15441 16.2531
R16397 vss.n15441 vss.n505 16.2531
R16398 vss.n15431 vss.n505 16.2531
R16399 vss.n7318 vss.n7317 16.2531
R16400 vss.n7317 vss.n7302 16.2531
R16401 vss.n7345 vss.n7302 16.2531
R16402 vss.n7345 vss.n7344 16.2531
R16403 vss.n7344 vss.n7303 16.2531
R16404 vss.n7334 vss.n7303 16.2531
R16405 vss.n7389 vss.n7388 16.2531
R16406 vss.n7388 vss.n7387 16.2531
R16407 vss.n7387 vss.n7351 16.2531
R16408 vss.n7377 vss.n7351 16.2531
R16409 vss.n7377 vss.n7376 16.2531
R16410 vss.n7376 vss.n7375 16.2531
R16411 vss.n3086 vss.n3085 16.2531
R16412 vss.n3085 vss.n3065 16.2531
R16413 vss.n3109 vss.n3065 16.2531
R16414 vss.n3109 vss.n3108 16.2531
R16415 vss.n3108 vss.n3066 16.2531
R16416 vss.n3098 vss.n3066 16.2531
R16417 vss.n725 vss.n724 16.2531
R16418 vss.n724 vss.n709 16.2531
R16419 vss.n15369 vss.n709 16.2531
R16420 vss.n15369 vss.n15368 16.2531
R16421 vss.n15368 vss.n710 16.2531
R16422 vss.n15358 vss.n710 16.2531
R16423 vss.n778 vss.n777 16.2531
R16424 vss.n777 vss.n762 16.2531
R16425 vss.n15292 vss.n762 16.2531
R16426 vss.n15292 vss.n15291 16.2531
R16427 vss.n15291 vss.n763 16.2531
R16428 vss.n15281 vss.n763 16.2531
R16429 vss.n983 vss.n982 16.2531
R16430 vss.n982 vss.n967 16.2531
R16431 vss.n15171 vss.n967 16.2531
R16432 vss.n15171 vss.n15170 16.2531
R16433 vss.n15170 vss.n968 16.2531
R16434 vss.n15159 vss.n968 16.2531
R16435 vss.n15192 vss.n15191 16.2531
R16436 vss.n15191 vss.n15176 16.2531
R16437 vss.n15219 vss.n15176 16.2531
R16438 vss.n15219 vss.n15218 16.2531
R16439 vss.n15218 vss.n15177 16.2531
R16440 vss.n15208 vss.n15177 16.2531
R16441 vss.n935 vss.n934 16.2531
R16442 vss.n934 vss.n919 16.2531
R16443 vss.n963 vss.n919 16.2531
R16444 vss.n963 vss.n962 16.2531
R16445 vss.n962 vss.n920 16.2531
R16446 vss.n952 vss.n920 16.2531
R16447 vss.n833 vss.n832 16.2531
R16448 vss.n834 vss.n833 16.2531
R16449 vss.n834 vss.n810 16.2531
R16450 vss.n845 vss.n810 16.2531
R16451 vss.n846 vss.n845 16.2531
R16452 vss.n847 vss.n846 16.2531
R16453 vss.n15139 vss.n15138 16.2531
R16454 vss.n15138 vss.n15137 16.2531
R16455 vss.n15137 vss.n15100 16.2531
R16456 vss.n15127 vss.n15100 16.2531
R16457 vss.n15127 vss.n15126 16.2531
R16458 vss.n15126 vss.n15125 16.2531
R16459 vss.n7484 vss.n7483 16.2531
R16460 vss.n7483 vss.n7482 16.2531
R16461 vss.n7482 vss.n7447 16.2531
R16462 vss.n7472 vss.n7447 16.2531
R16463 vss.n7472 vss.n7471 16.2531
R16464 vss.n7471 vss.n7470 16.2531
R16465 vss.n15312 vss.n15311 16.2531
R16466 vss.n15311 vss.n15296 16.2531
R16467 vss.n15340 vss.n15296 16.2531
R16468 vss.n15340 vss.n15339 16.2531
R16469 vss.n15339 vss.n15297 16.2531
R16470 vss.n15329 vss.n15297 16.2531
R16471 vss.n678 vss.n677 16.2531
R16472 vss.n677 vss.n662 16.2531
R16473 vss.n706 vss.n662 16.2531
R16474 vss.n706 vss.n705 16.2531
R16475 vss.n705 vss.n663 16.2531
R16476 vss.n695 vss.n663 16.2531
R16477 vss.n7437 vss.n7436 16.2531
R16478 vss.n7436 vss.n7435 16.2531
R16479 vss.n7435 vss.n7399 16.2531
R16480 vss.n7425 vss.n7399 16.2531
R16481 vss.n7425 vss.n7424 16.2531
R16482 vss.n7424 vss.n7423 16.2531
R16483 vss.n3127 vss.n3126 16.2531
R16484 vss.n3126 vss.n3111 16.2531
R16485 vss.n7299 vss.n3111 16.2531
R16486 vss.n7299 vss.n7298 16.2531
R16487 vss.n7298 vss.n3112 16.2531
R16488 vss.n7287 vss.n3112 16.2531
R16489 vss.n576 vss.n575 16.2531
R16490 vss.n577 vss.n576 16.2531
R16491 vss.n577 vss.n553 16.2531
R16492 vss.n588 vss.n553 16.2531
R16493 vss.n589 vss.n588 16.2531
R16494 vss.n590 vss.n589 16.2531
R16495 vss.n470 vss.n469 16.2531
R16496 vss.n469 vss.n454 16.2531
R16497 vss.n498 vss.n454 16.2531
R16498 vss.n498 vss.n497 16.2531
R16499 vss.n497 vss.n455 16.2531
R16500 vss.n487 vss.n455 16.2531
R16501 vss.n4727 vss.n4726 16.2531
R16502 vss.n4728 vss.n4727 16.2531
R16503 vss.n4728 vss.n4704 16.2531
R16504 vss.n4739 vss.n4704 16.2531
R16505 vss.n4740 vss.n4739 16.2531
R16506 vss.n4741 vss.n4740 16.2531
R16507 vss.n4677 vss.n4676 16.2531
R16508 vss.n4676 vss.n4656 16.2531
R16509 vss.n4700 vss.n4656 16.2531
R16510 vss.n4700 vss.n4699 16.2531
R16511 vss.n4699 vss.n4657 16.2531
R16512 vss.n4689 vss.n4657 16.2531
R16513 vss.n4624 vss.n4623 16.2531
R16514 vss.n4623 vss.n4608 16.2531
R16515 vss.n4652 vss.n4608 16.2531
R16516 vss.n4652 vss.n4651 16.2531
R16517 vss.n4651 vss.n4609 16.2531
R16518 vss.n4640 vss.n4609 16.2531
R16519 vss.n4576 vss.n4575 16.2531
R16520 vss.n4575 vss.n4560 16.2531
R16521 vss.n4605 vss.n4560 16.2531
R16522 vss.n4605 vss.n4604 16.2531
R16523 vss.n4604 vss.n4561 16.2531
R16524 vss.n4593 vss.n4561 16.2531
R16525 vss.n4342 vss.n4341 16.2531
R16526 vss.n4343 vss.n4342 16.2531
R16527 vss.n4343 vss.n4319 16.2531
R16528 vss.n4354 vss.n4319 16.2531
R16529 vss.n4355 vss.n4354 16.2531
R16530 vss.n4356 vss.n4355 16.2531
R16531 vss.n7267 vss.n7266 16.2531
R16532 vss.n7266 vss.n7265 16.2531
R16533 vss.n7265 vss.n7229 16.2531
R16534 vss.n7255 vss.n7229 16.2531
R16535 vss.n7255 vss.n7254 16.2531
R16536 vss.n7254 vss.n7253 16.2531
R16537 vss.n6848 vss.n6847 16.2531
R16538 vss.n6847 vss.n6832 16.2531
R16539 vss.n6875 vss.n6832 16.2531
R16540 vss.n6875 vss.n6874 16.2531
R16541 vss.n6874 vss.n6833 16.2531
R16542 vss.n6864 vss.n6833 16.2531
R16543 vss.n6809 vss.n6808 16.2531
R16544 vss.n6809 vss.n3148 16.2531
R16545 vss.n7208 vss.n3148 16.2531
R16546 vss.n7209 vss.n7208 16.2531
R16547 vss.n7209 vss.n3138 16.2531
R16548 vss.n7219 vss.n3138 16.2531
R16549 vss.n6916 vss.n6915 16.2531
R16550 vss.n6915 vss.n6914 16.2531
R16551 vss.n6914 vss.n6879 16.2531
R16552 vss.n6895 vss.n6879 16.2531
R16553 vss.n6902 vss.n6895 16.2531
R16554 vss.n6902 vss.n6901 16.2531
R16555 vss.n2619 vss.n2618 16.2531
R16556 vss.n2618 vss.n2611 16.2531
R16557 vss.n2611 vss.n1140 16.2531
R16558 vss.n2633 vss.n1140 16.2531
R16559 vss.n2633 vss.n2632 16.2531
R16560 vss.n2632 vss.n2601 16.2531
R16561 vss.n1910 vss.n1900 16.2531
R16562 vss.n1935 vss.n1910 16.2531
R16563 vss.n1935 vss.n1934 16.2531
R16564 vss.n1934 vss.n1932 16.2531
R16565 vss.n1932 vss.n1913 16.2531
R16566 vss.n1922 vss.n1913 16.2531
R16567 vss.n2855 vss.n2854 16.2531
R16568 vss.n2854 vss.n2839 16.2531
R16569 vss.n2882 vss.n2839 16.2531
R16570 vss.n2882 vss.n2881 16.2531
R16571 vss.n2881 vss.n2840 16.2531
R16572 vss.n2871 vss.n2840 16.2531
R16573 vss.n7736 vss.n7735 16.2531
R16574 vss.n7735 vss.n7720 16.2531
R16575 vss.n7764 vss.n7720 16.2531
R16576 vss.n7764 vss.n7763 16.2531
R16577 vss.n7763 vss.n7721 16.2531
R16578 vss.n7753 vss.n7721 16.2531
R16579 vss.n2902 vss.n2898 16.2531
R16580 vss.n2902 vss.n2884 16.2531
R16581 vss.n2929 vss.n2884 16.2531
R16582 vss.n2929 vss.n2928 16.2531
R16583 vss.n2928 vss.n2927 16.2531
R16584 vss.n2927 vss.n2926 16.2531
R16585 vss.n7687 vss.n7686 16.2531
R16586 vss.n7686 vss.n7671 16.2531
R16587 vss.n7716 vss.n7671 16.2531
R16588 vss.n7716 vss.n7715 16.2531
R16589 vss.n7715 vss.n7672 16.2531
R16590 vss.n7704 vss.n7672 16.2531
R16591 vss.n3032 vss.n3024 16.2531
R16592 vss.n3042 vss.n3024 16.2531
R16593 vss.n3043 vss.n3042 16.2531
R16594 vss.n3045 vss.n3043 16.2531
R16595 vss.n3045 vss.n3044 16.2531
R16596 vss.n3044 vss.n3015 16.2531
R16597 vss.n7639 vss.n7638 16.2531
R16598 vss.n7638 vss.n7623 16.2531
R16599 vss.n7666 vss.n7623 16.2531
R16600 vss.n7666 vss.n7665 16.2531
R16601 vss.n7665 vss.n7624 16.2531
R16602 vss.n7655 vss.n7624 16.2531
R16603 vss.n2741 vss.n2740 16.2531
R16604 vss.n2740 vss.n2725 16.2531
R16605 vss.n2836 vss.n2725 16.2531
R16606 vss.n2836 vss.n2835 16.2531
R16607 vss.n2835 vss.n2726 16.2531
R16608 vss.n2825 vss.n2726 16.2531
R16609 vss.n2947 vss.n2946 16.2531
R16610 vss.n2946 vss.n2931 16.2531
R16611 vss.n2975 vss.n2931 16.2531
R16612 vss.n2975 vss.n2974 16.2531
R16613 vss.n2974 vss.n2932 16.2531
R16614 vss.n2964 vss.n2932 16.2531
R16615 vss.n2993 vss.n2992 16.2531
R16616 vss.n2992 vss.n2977 16.2531
R16617 vss.n7500 vss.n2977 16.2531
R16618 vss.n7500 vss.n7499 16.2531
R16619 vss.n7499 vss.n2978 16.2531
R16620 vss.n3010 vss.n2978 16.2531
R16621 vss.n7963 vss.n2468 16.2531
R16622 vss.n7963 vss.n2453 16.2531
R16623 vss.n7990 vss.n2453 16.2531
R16624 vss.n7990 vss.n7989 16.2531
R16625 vss.n7989 vss.n7988 16.2531
R16626 vss.n7988 vss.n7987 16.2531
R16627 vss.n7120 vss.n7119 16.2531
R16628 vss.n7119 vss.n7118 16.2531
R16629 vss.n7118 vss.n2451 16.2531
R16630 vss.n7098 vss.n2451 16.2531
R16631 vss.n7106 vss.n7098 16.2531
R16632 vss.n7106 vss.n7105 16.2531
R16633 vss.n7046 vss.n7035 16.2531
R16634 vss.n7047 vss.n7046 16.2531
R16635 vss.n7065 vss.n7047 16.2531
R16636 vss.n7065 vss.n7064 16.2531
R16637 vss.n7064 vss.n7048 16.2531
R16638 vss.n7055 vss.n7048 16.2531
R16639 vss.n7008 vss.n7007 16.2531
R16640 vss.n7007 vss.n7000 16.2531
R16641 vss.n7000 vss.n2450 16.2531
R16642 vss.n7022 vss.n2450 16.2531
R16643 vss.n7022 vss.n7021 16.2531
R16644 vss.n7021 vss.n6990 16.2531
R16645 vss.n7147 vss.n7139 16.2531
R16646 vss.n7157 vss.n7139 16.2531
R16647 vss.n7158 vss.n7157 16.2531
R16648 vss.n7160 vss.n7158 16.2531
R16649 vss.n7160 vss.n7159 16.2531
R16650 vss.n7159 vss.n7127 16.2531
R16651 vss.n6963 vss.n6935 16.2531
R16652 vss.n6973 vss.n6935 16.2531
R16653 vss.n6975 vss.n6973 16.2531
R16654 vss.n6977 vss.n6975 16.2531
R16655 vss.n6977 vss.n6976 16.2531
R16656 vss.n6976 vss.n6923 16.2531
R16657 vss.n7523 vss.n7522 16.2531
R16658 vss.n7522 vss.n7507 16.2531
R16659 vss.n7618 vss.n7507 16.2531
R16660 vss.n7618 vss.n7617 16.2531
R16661 vss.n7617 vss.n7508 16.2531
R16662 vss.n7607 vss.n7508 16.2531
R16663 vss.n7786 vss.n7785 16.2531
R16664 vss.n7785 vss.n7770 16.2531
R16665 vss.n7813 vss.n7770 16.2531
R16666 vss.n7813 vss.n7812 16.2531
R16667 vss.n7812 vss.n7771 16.2531
R16668 vss.n7802 vss.n7771 16.2531
R16669 vss.n7834 vss.n7833 16.2531
R16670 vss.n7833 vss.n7818 16.2531
R16671 vss.n7861 vss.n7818 16.2531
R16672 vss.n7861 vss.n7860 16.2531
R16673 vss.n7860 vss.n7819 16.2531
R16674 vss.n7850 vss.n7819 16.2531
R16675 vss.n7882 vss.n7881 16.2531
R16676 vss.n7881 vss.n7866 16.2531
R16677 vss.n7911 vss.n7866 16.2531
R16678 vss.n7911 vss.n7910 16.2531
R16679 vss.n7910 vss.n7867 16.2531
R16680 vss.n7899 vss.n7867 16.2531
R16681 vss.n2657 vss.n2646 16.2531
R16682 vss.n2658 vss.n2657 16.2531
R16683 vss.n7914 vss.n2658 16.2531
R16684 vss.n7914 vss.n2678 16.2531
R16685 vss.n2678 vss.n2677 16.2531
R16686 vss.n2677 vss.n2676 16.2531
R16687 vss.n2696 vss.n2695 16.2531
R16688 vss.n2695 vss.n2680 16.2531
R16689 vss.n2722 vss.n2680 16.2531
R16690 vss.n2722 vss.n2721 16.2531
R16691 vss.n2721 vss.n2681 16.2531
R16692 vss.n2711 vss.n2681 16.2531
R16693 vss.n2575 vss.n2498 16.2531
R16694 vss.n2585 vss.n2498 16.2531
R16695 vss.n2586 vss.n2585 16.2531
R16696 vss.n2588 vss.n2586 16.2531
R16697 vss.n2588 vss.n2587 16.2531
R16698 vss.n2587 vss.n2486 16.2531
R16699 vss.n7942 vss.n7941 16.2531
R16700 vss.n7941 vss.n1142 16.2531
R16701 vss.n14881 vss.n1142 16.2531
R16702 vss.n14881 vss.n14880 16.2531
R16703 vss.n14880 vss.n1143 16.2531
R16704 vss.n1156 vss.n1143 16.2531
R16705 vss.n3167 vss.n3166 16.2531
R16706 vss.n3166 vss.n3151 16.2531
R16707 vss.n7205 vss.n3151 16.2531
R16708 vss.n7205 vss.n7204 16.2531
R16709 vss.n7204 vss.n3152 16.2531
R16710 vss.n7194 vss.n3152 16.2531
R16711 vss.n3195 vss.n3194 16.2531
R16712 vss.n3195 vss.n3184 16.2531
R16713 vss.n6792 vss.n3184 16.2531
R16714 vss.n6794 vss.n6792 16.2531
R16715 vss.n6794 vss.n6793 16.2531
R16716 vss.n6793 vss.n3172 16.2531
R16717 vss.n6762 vss.n6761 16.2531
R16718 vss.n6761 vss.n6746 16.2531
R16719 vss.n6789 vss.n6746 16.2531
R16720 vss.n6789 vss.n6788 16.2531
R16721 vss.n6788 vss.n6747 16.2531
R16722 vss.n6778 vss.n6747 16.2531
R16723 vss.n14829 vss.n14828 16.2531
R16724 vss.n14830 vss.n14829 16.2531
R16725 vss.n14830 vss.n14806 16.2531
R16726 vss.n14841 vss.n14806 16.2531
R16727 vss.n14842 vss.n14841 16.2531
R16728 vss.n14843 vss.n14842 16.2531
R16729 vss.n14171 vss.n14170 16.2531
R16730 vss.n14170 vss.n1169 16.2531
R16731 vss.n14803 vss.n1169 16.2531
R16732 vss.n14803 vss.n14802 16.2531
R16733 vss.n14802 vss.n1170 16.2531
R16734 vss.n14792 vss.n1170 16.2531
R16735 vss.n14318 vss.n14317 16.2531
R16736 vss.n14317 vss.n14284 16.2531
R16737 vss.n14323 vss.n14284 16.2531
R16738 vss.n14323 vss.n14322 16.2531
R16739 vss.n14322 vss.n14285 16.2531
R16740 vss.n14308 vss.n14285 16.2531
R16741 vss.n1837 vss.n1836 16.2531
R16742 vss.n1836 vss.n1821 16.2531
R16743 vss.n14353 vss.n1821 16.2531
R16744 vss.n14353 vss.n14352 16.2531
R16745 vss.n14352 vss.n1822 16.2531
R16746 vss.n14342 vss.n1822 16.2531
R16747 vss.n14210 vss.n14209 16.2531
R16748 vss.n14209 vss.n14194 16.2531
R16749 vss.n14239 vss.n14194 16.2531
R16750 vss.n14239 vss.n14238 16.2531
R16751 vss.n14238 vss.n14195 16.2531
R16752 vss.n14228 vss.n14195 16.2531
R16753 vss.n1299 vss.n1298 16.2531
R16754 vss.n1298 vss.n1283 16.2531
R16755 vss.n14747 vss.n1283 16.2531
R16756 vss.n14747 vss.n14746 16.2531
R16757 vss.n14746 vss.n1284 16.2531
R16758 vss.n14736 vss.n1284 16.2531
R16759 vss.n13998 vss.n13997 16.2531
R16760 vss.n13997 vss.n13982 16.2531
R16761 vss.n14025 vss.n13982 16.2531
R16762 vss.n14025 vss.n14024 16.2531
R16763 vss.n14024 vss.n13983 16.2531
R16764 vss.n14014 vss.n13983 16.2531
R16765 vss.n8218 vss.n8217 16.2531
R16766 vss.n8217 vss.n8216 16.2531
R16767 vss.n8216 vss.n8180 16.2531
R16768 vss.n8206 vss.n8180 16.2531
R16769 vss.n8206 vss.n8205 16.2531
R16770 vss.n8205 vss.n8204 16.2531
R16771 vss.n8169 vss.n8168 16.2531
R16772 vss.n8168 vss.n8153 16.2531
R16773 vss.n13979 vss.n8153 16.2531
R16774 vss.n13979 vss.n13978 16.2531
R16775 vss.n13978 vss.n8154 16.2531
R16776 vss.n13968 vss.n8154 16.2531
R16777 vss.n1504 vss.n1503 16.2531
R16778 vss.n1503 vss.n1488 16.2531
R16779 vss.n14674 vss.n1488 16.2531
R16780 vss.n14674 vss.n14673 16.2531
R16781 vss.n14673 vss.n1489 16.2531
R16782 vss.n14663 vss.n1489 16.2531
R16783 vss.n1557 vss.n1556 16.2531
R16784 vss.n1556 vss.n1541 16.2531
R16785 vss.n14597 vss.n1541 16.2531
R16786 vss.n14597 vss.n14596 16.2531
R16787 vss.n14596 vss.n1542 16.2531
R16788 vss.n14586 vss.n1542 16.2531
R16789 vss.n1762 vss.n1761 16.2531
R16790 vss.n1761 vss.n1746 16.2531
R16791 vss.n14476 vss.n1746 16.2531
R16792 vss.n14476 vss.n14475 16.2531
R16793 vss.n14475 vss.n1747 16.2531
R16794 vss.n14464 vss.n1747 16.2531
R16795 vss.n14497 vss.n14496 16.2531
R16796 vss.n14496 vss.n14481 16.2531
R16797 vss.n14524 vss.n14481 16.2531
R16798 vss.n14524 vss.n14523 16.2531
R16799 vss.n14523 vss.n14482 16.2531
R16800 vss.n14513 vss.n14482 16.2531
R16801 vss.n1714 vss.n1713 16.2531
R16802 vss.n1713 vss.n1698 16.2531
R16803 vss.n1742 vss.n1698 16.2531
R16804 vss.n1742 vss.n1741 16.2531
R16805 vss.n1741 vss.n1699 16.2531
R16806 vss.n1731 vss.n1699 16.2531
R16807 vss.n1612 vss.n1611 16.2531
R16808 vss.n1613 vss.n1612 16.2531
R16809 vss.n1613 vss.n1589 16.2531
R16810 vss.n1624 vss.n1589 16.2531
R16811 vss.n1625 vss.n1624 16.2531
R16812 vss.n1626 vss.n1625 16.2531
R16813 vss.n14444 vss.n14443 16.2531
R16814 vss.n14443 vss.n14442 16.2531
R16815 vss.n14442 vss.n14405 16.2531
R16816 vss.n14432 vss.n14405 16.2531
R16817 vss.n14432 vss.n14431 16.2531
R16818 vss.n14431 vss.n14430 16.2531
R16819 vss.n13949 vss.n13948 16.2531
R16820 vss.n13948 vss.n13947 16.2531
R16821 vss.n13947 vss.n13912 16.2531
R16822 vss.n13937 vss.n13912 16.2531
R16823 vss.n13937 vss.n13936 16.2531
R16824 vss.n13936 vss.n13935 16.2531
R16825 vss.n14617 vss.n14616 16.2531
R16826 vss.n14616 vss.n14601 16.2531
R16827 vss.n14645 vss.n14601 16.2531
R16828 vss.n14645 vss.n14644 16.2531
R16829 vss.n14644 vss.n14602 16.2531
R16830 vss.n14634 vss.n14602 16.2531
R16831 vss.n1457 vss.n1456 16.2531
R16832 vss.n1456 vss.n1441 16.2531
R16833 vss.n1485 vss.n1441 16.2531
R16834 vss.n1485 vss.n1484 16.2531
R16835 vss.n1484 vss.n1442 16.2531
R16836 vss.n1474 vss.n1442 16.2531
R16837 vss.n13902 vss.n13901 16.2531
R16838 vss.n13901 vss.n13900 16.2531
R16839 vss.n13900 vss.n13864 16.2531
R16840 vss.n13890 vss.n13864 16.2531
R16841 vss.n13890 vss.n13889 16.2531
R16842 vss.n13889 vss.n13888 16.2531
R16843 vss.n14066 vss.n14065 16.2531
R16844 vss.n14065 vss.n14064 16.2531
R16845 vss.n14064 vss.n14029 16.2531
R16846 vss.n14054 vss.n14029 16.2531
R16847 vss.n14054 vss.n14053 16.2531
R16848 vss.n14053 vss.n14052 16.2531
R16849 vss.n1355 vss.n1354 16.2531
R16850 vss.n1356 vss.n1355 16.2531
R16851 vss.n1356 vss.n1332 16.2531
R16852 vss.n1367 vss.n1332 16.2531
R16853 vss.n1368 vss.n1367 16.2531
R16854 vss.n1369 vss.n1368 16.2531
R16855 vss.n1249 vss.n1248 16.2531
R16856 vss.n1248 vss.n1233 16.2531
R16857 vss.n1277 vss.n1233 16.2531
R16858 vss.n1277 vss.n1276 16.2531
R16859 vss.n1276 vss.n1234 16.2531
R16860 vss.n1266 vss.n1234 16.2531
R16861 vss.n2342 vss.n2341 16.2531
R16862 vss.n2341 vss.n2326 16.2531
R16863 vss.n8046 vss.n2326 16.2531
R16864 vss.n8046 vss.n8045 16.2531
R16865 vss.n8045 vss.n2327 16.2531
R16866 vss.n8035 vss.n2327 16.2531
R16867 vss.n2253 vss.n2252 16.2531
R16868 vss.n2252 vss.n2232 16.2531
R16869 vss.n2276 vss.n2232 16.2531
R16870 vss.n2276 vss.n2275 16.2531
R16871 vss.n2275 vss.n2233 16.2531
R16872 vss.n2265 vss.n2233 16.2531
R16873 vss.n8090 vss.n8089 16.2531
R16874 vss.n8089 vss.n8088 16.2531
R16875 vss.n8088 vss.n8052 16.2531
R16876 vss.n8078 vss.n8052 16.2531
R16877 vss.n8078 vss.n8077 16.2531
R16878 vss.n8077 vss.n8076 16.2531
R16879 vss.n2294 vss.n2293 16.2531
R16880 vss.n2293 vss.n2278 16.2531
R16881 vss.n2323 vss.n2278 16.2531
R16882 vss.n2323 vss.n2322 16.2531
R16883 vss.n2322 vss.n2279 16.2531
R16884 vss.n2311 vss.n2279 16.2531
R16885 vss.n2397 vss.n2396 16.2531
R16886 vss.n2398 vss.n2397 16.2531
R16887 vss.n2398 vss.n2374 16.2531
R16888 vss.n2409 vss.n2374 16.2531
R16889 vss.n2410 vss.n2409 16.2531
R16890 vss.n2411 vss.n2410 16.2531
R16891 vss.n8141 vss.n8140 16.2531
R16892 vss.n8140 vss.n8139 16.2531
R16893 vss.n8139 vss.n8103 16.2531
R16894 vss.n8129 vss.n8103 16.2531
R16895 vss.n8129 vss.n8128 16.2531
R16896 vss.n8128 vss.n8127 16.2531
R16897 vss.n11948 vss.n11947 16.2531
R16898 vss.n11948 vss.n2088 16.2531
R16899 vss.n14137 vss.n2088 16.2531
R16900 vss.n14137 vss.n14136 16.2531
R16901 vss.n14136 vss.n2089 16.2531
R16902 vss.n14126 vss.n2089 16.2531
R16903 vss.n13484 vss.n13483 16.2531
R16904 vss.n13483 vss.n13468 16.2531
R16905 vss.n13511 vss.n13468 16.2531
R16906 vss.n13511 vss.n13510 16.2531
R16907 vss.n13510 vss.n13469 16.2531
R16908 vss.n13500 vss.n13469 16.2531
R16909 vss.n12028 vss.n12018 16.2531
R16910 vss.n12051 vss.n12028 16.2531
R16911 vss.n12051 vss.n12050 16.2531
R16912 vss.n12050 vss.n12049 16.2531
R16913 vss.n12049 vss.n12031 16.2531
R16914 vss.n12039 vss.n12031 16.2531
R16915 vss.n8319 vss.n8318 16.2531
R16916 vss.n8318 vss.n8303 16.2531
R16917 vss.n13743 vss.n8303 16.2531
R16918 vss.n13743 vss.n13742 16.2531
R16919 vss.n13742 vss.n8304 16.2531
R16920 vss.n13732 vss.n8304 16.2531
R16921 vss.n8454 vss.n8444 16.2531
R16922 vss.n8477 vss.n8454 16.2531
R16923 vss.n8477 vss.n8476 16.2531
R16924 vss.n8476 vss.n8475 16.2531
R16925 vss.n8475 vss.n8457 16.2531
R16926 vss.n8465 vss.n8457 16.2531
R16927 vss.n8531 vss.n8521 16.2531
R16928 vss.n8554 vss.n8531 16.2531
R16929 vss.n8554 vss.n8553 16.2531
R16930 vss.n8553 vss.n8552 16.2531
R16931 vss.n8552 vss.n8534 16.2531
R16932 vss.n8542 vss.n8534 16.2531
R16933 vss.n9105 vss.n9104 16.2531
R16934 vss.n9104 vss.n9089 16.2531
R16935 vss.n13031 vss.n9089 16.2531
R16936 vss.n13031 vss.n13030 16.2531
R16937 vss.n13030 vss.n9090 16.2531
R16938 vss.n13020 vss.n9090 16.2531
R16939 vss.n8969 vss.n8968 16.2531
R16940 vss.n8968 vss.n8953 16.2531
R16941 vss.n8996 vss.n8953 16.2531
R16942 vss.n8996 vss.n8995 16.2531
R16943 vss.n8995 vss.n8954 16.2531
R16944 vss.n8985 vss.n8954 16.2531
R16945 vss.n9126 vss.n9116 16.2531
R16946 vss.n9149 vss.n9126 16.2531
R16947 vss.n9149 vss.n9148 16.2531
R16948 vss.n9148 vss.n9147 16.2531
R16949 vss.n9147 vss.n9129 16.2531
R16950 vss.n9137 vss.n9129 16.2531
R16951 vss.n12557 vss.n12547 16.2531
R16952 vss.n12629 vss.n12557 16.2531
R16953 vss.n12629 vss.n12628 16.2531
R16954 vss.n12628 vss.n12578 16.2531
R16955 vss.n12578 vss.n12560 16.2531
R16956 vss.n12568 vss.n12560 16.2531
R16957 vss.n2163 vss.n2162 16.2531
R16958 vss.n2162 vss.n2147 16.2531
R16959 vss.n14086 vss.n2147 16.2531
R16960 vss.n14086 vss.n14085 16.2531
R16961 vss.n14085 vss.n2148 16.2531
R16962 vss.n2179 vss.n2148 16.2531
R16963 vss.n12596 vss.n12595 16.2531
R16964 vss.n12595 vss.n12580 16.2531
R16965 vss.n12624 vss.n12580 16.2531
R16966 vss.n12624 vss.n12623 16.2531
R16967 vss.n12623 vss.n12581 16.2531
R16968 vss.n12613 vss.n12581 16.2531
R16969 vss.n9014 vss.n9013 16.2531
R16970 vss.n9013 vss.n8998 16.2531
R16971 vss.n9040 vss.n8998 16.2531
R16972 vss.n9040 vss.n9039 16.2531
R16973 vss.n9039 vss.n8999 16.2531
R16974 vss.n9029 vss.n8999 16.2531
R16975 vss.n13099 vss.n13098 16.2531
R16976 vss.n13098 vss.n13083 16.2531
R16977 vss.n13128 vss.n13083 16.2531
R16978 vss.n13128 vss.n13127 16.2531
R16979 vss.n13127 vss.n13084 16.2531
R16980 vss.n13116 vss.n13084 16.2531
R16981 vss.n13051 vss.n13050 16.2531
R16982 vss.n13050 vss.n13035 16.2531
R16983 vss.n13080 vss.n13035 16.2531
R16984 vss.n13080 vss.n13079 16.2531
R16985 vss.n13079 vss.n13036 16.2531
R16986 vss.n13067 vss.n13036 16.2531
R16987 vss.n9058 vss.n9057 16.2531
R16988 vss.n9057 vss.n9042 16.2531
R16989 vss.n9086 vss.n9042 16.2531
R16990 vss.n9086 vss.n9085 16.2531
R16991 vss.n9085 vss.n9043 16.2531
R16992 vss.n9075 vss.n9043 16.2531
R16993 vss.n8243 vss.n8235 16.2531
R16994 vss.n8253 vss.n8235 16.2531
R16995 vss.n13844 vss.n8253 16.2531
R16996 vss.n13846 vss.n13844 16.2531
R16997 vss.n13846 vss.n13845 16.2531
R16998 vss.n13845 vss.n8226 16.2531
R16999 vss.n13811 vss.n13810 16.2531
R17000 vss.n13810 vss.n13795 16.2531
R17001 vss.n13840 vss.n13795 16.2531
R17002 vss.n13840 vss.n13839 16.2531
R17003 vss.n13839 vss.n13796 16.2531
R17004 vss.n13828 vss.n13796 16.2531
R17005 vss.n13763 vss.n13762 16.2531
R17006 vss.n13762 vss.n13747 16.2531
R17007 vss.n13792 vss.n13747 16.2531
R17008 vss.n13792 vss.n13791 16.2531
R17009 vss.n13791 vss.n13748 16.2531
R17010 vss.n13779 vss.n13748 16.2531
R17011 vss.n8272 vss.n8271 16.2531
R17012 vss.n8271 vss.n8256 16.2531
R17013 vss.n8300 vss.n8256 16.2531
R17014 vss.n8300 vss.n8299 16.2531
R17015 vss.n8299 vss.n8257 16.2531
R17016 vss.n8289 vss.n8257 16.2531
R17017 vss.n13529 vss.n13528 16.2531
R17018 vss.n13528 vss.n13513 16.2531
R17019 vss.n13555 vss.n13513 16.2531
R17020 vss.n13555 vss.n13554 16.2531
R17021 vss.n13554 vss.n13514 16.2531
R17022 vss.n13544 vss.n13514 16.2531
R17023 vss.n13622 vss.n13621 16.2531
R17024 vss.n13621 vss.n13606 16.2531
R17025 vss.n13651 vss.n13606 16.2531
R17026 vss.n13651 vss.n13650 16.2531
R17027 vss.n13650 vss.n13607 16.2531
R17028 vss.n13639 vss.n13607 16.2531
R17029 vss.n13573 vss.n13572 16.2531
R17030 vss.n13572 vss.n13557 16.2531
R17031 vss.n13603 vss.n13557 16.2531
R17032 vss.n13603 vss.n13602 16.2531
R17033 vss.n13602 vss.n13558 16.2531
R17034 vss.n13590 vss.n13558 16.2531
R17035 vss.n2075 vss.n2066 16.2531
R17036 vss.n2086 vss.n2066 16.2531
R17037 vss.n14141 vss.n2086 16.2531
R17038 vss.n14143 vss.n14141 16.2531
R17039 vss.n14143 vss.n14142 16.2531
R17040 vss.n14142 vss.n2057 16.2531
R17041 vss.n2201 vss.n2200 16.2531
R17042 vss.n2200 vss.n2193 16.2531
R17043 vss.n2193 vss.n2145 16.2531
R17044 vss.n2215 vss.n2145 16.2531
R17045 vss.n2215 vss.n2214 16.2531
R17046 vss.n2214 vss.n2183 16.2531
R17047 vss.n9287 vss.n9286 16.2531
R17048 vss.n9287 vss.n2143 16.2531
R17049 vss.n14092 vss.n2143 16.2531
R17050 vss.n14094 vss.n14092 16.2531
R17051 vss.n14094 vss.n14093 16.2531
R17052 vss.n14093 vss.n2131 16.2531
R17053 vss.n9409 vss.n9408 16.2531
R17054 vss.n9408 vss.n9393 16.2531
R17055 vss.n12868 vss.n9393 16.2531
R17056 vss.n12868 vss.n12867 16.2531
R17057 vss.n12867 vss.n9394 16.2531
R17058 vss.n12857 vss.n9394 16.2531
R17059 vss.n12741 vss.n12731 16.2531
R17060 vss.n12765 vss.n12741 16.2531
R17061 vss.n12765 vss.n12764 16.2531
R17062 vss.n12764 vss.n12762 16.2531
R17063 vss.n12762 vss.n12744 16.2531
R17064 vss.n12752 vss.n12744 16.2531
R17065 vss.n8427 vss.n8426 16.2531
R17066 vss.n8426 vss.n8411 16.2531
R17067 vss.n13345 vss.n8411 16.2531
R17068 vss.n13345 vss.n13344 16.2531
R17069 vss.n13344 vss.n8412 16.2531
R17070 vss.n13334 vss.n8412 16.2531
R17071 vss.n13369 vss.n13368 16.2531
R17072 vss.n13368 vss.n13353 16.2531
R17073 vss.n13464 vss.n13353 16.2531
R17074 vss.n13464 vss.n13463 16.2531
R17075 vss.n13463 vss.n13354 16.2531
R17076 vss.n13453 vss.n13354 16.2531
R17077 vss.n11851 vss.n11850 16.2531
R17078 vss.n11851 vss.n2036 16.2531
R17079 vss.n14189 vss.n2036 16.2531
R17080 vss.n14189 vss.n14188 16.2531
R17081 vss.n14188 vss.n2037 16.2531
R17082 vss.n2050 vss.n2037 16.2531
R17083 vss.n1811 vss.n1810 16.2531
R17084 vss.n1810 vss.n1809 16.2531
R17085 vss.n1809 vss.n1773 16.2531
R17086 vss.n1799 vss.n1773 16.2531
R17087 vss.n1799 vss.n1798 16.2531
R17088 vss.n1798 vss.n1797 16.2531
R17089 vss.n14394 vss.n14393 16.2531
R17090 vss.n14393 vss.n14392 16.2531
R17091 vss.n14392 vss.n14357 16.2531
R17092 vss.n14382 vss.n14357 16.2531
R17093 vss.n14382 vss.n14381 16.2531
R17094 vss.n14381 vss.n14380 16.2531
R17095 vss.n2004 vss.n2003 16.2531
R17096 vss.n2003 vss.n1988 16.2531
R17097 vss.n2032 vss.n1988 16.2531
R17098 vss.n2032 vss.n2031 16.2531
R17099 vss.n2031 vss.n1989 16.2531
R17100 vss.n2021 vss.n1989 16.2531
R17101 vss.n14257 vss.n14256 16.2531
R17102 vss.n14256 vss.n14242 16.2531
R17103 vss.n14280 vss.n14242 16.2531
R17104 vss.n14280 vss.n14279 16.2531
R17105 vss.n14279 vss.n14243 16.2531
R17106 vss.n14275 vss.n14243 16.2531
R17107 vss.n1032 vss.n1031 16.2531
R17108 vss.n1031 vss.n1030 16.2531
R17109 vss.n1030 vss.n994 16.2531
R17110 vss.n1020 vss.n994 16.2531
R17111 vss.n1020 vss.n1019 16.2531
R17112 vss.n1019 vss.n1018 16.2531
R17113 vss.n15089 vss.n15088 16.2531
R17114 vss.n15088 vss.n15087 16.2531
R17115 vss.n15087 vss.n15052 16.2531
R17116 vss.n15077 vss.n15052 16.2531
R17117 vss.n15077 vss.n15076 16.2531
R17118 vss.n15076 vss.n15075 16.2531
R17119 vss.n1109 vss.n1108 16.2531
R17120 vss.n1108 vss.n1093 16.2531
R17121 vss.n1137 vss.n1093 16.2531
R17122 vss.n1137 vss.n1136 16.2531
R17123 vss.n1136 vss.n1094 16.2531
R17124 vss.n1126 vss.n1094 16.2531
R17125 vss.n14952 vss.n14951 16.2531
R17126 vss.n14951 vss.n14937 16.2531
R17127 vss.n14975 vss.n14937 16.2531
R17128 vss.n14975 vss.n14974 16.2531
R17129 vss.n14974 vss.n14938 16.2531
R17130 vss.n14970 vss.n14938 16.2531
R17131 vss.n6248 vss.n6247 16.2531
R17132 vss.n6247 vss.n6246 16.2531
R17133 vss.n6246 vss.n6211 16.2531
R17134 vss.n6236 vss.n6211 16.2531
R17135 vss.n6236 vss.n6235 16.2531
R17136 vss.n6235 vss.n6234 16.2531
R17137 vss.n3963 vss.n3962 16.2531
R17138 vss.n3962 vss.n30 16.2531
R17139 vss.n15868 vss.n30 16.2531
R17140 vss.n15868 vss.n15867 16.2531
R17141 vss.n15867 vss.n31 16.2531
R17142 vss.n15857 vss.n31 16.2531
R17143 vss.n3894 vss.n3893 16.2531
R17144 vss.n3893 vss.n3892 16.2531
R17145 vss.n3892 vss.n3857 16.2531
R17146 vss.n3882 vss.n3857 16.2531
R17147 vss.n3882 vss.n3881 16.2531
R17148 vss.n3881 vss.n3880 16.2531
R17149 vss.n3775 vss.n3774 16.2531
R17150 vss.n3774 vss.n3773 16.2531
R17151 vss.n3773 vss.n3738 16.2531
R17152 vss.n3763 vss.n3738 16.2531
R17153 vss.n3763 vss.n3762 16.2531
R17154 vss.n3762 vss.n3761 16.2531
R17155 vss.n3656 vss.n3655 16.2531
R17156 vss.n3655 vss.n3654 16.2531
R17157 vss.n3654 vss.n3619 16.2531
R17158 vss.n3644 vss.n3619 16.2531
R17159 vss.n3644 vss.n3643 16.2531
R17160 vss.n3643 vss.n3642 16.2531
R17161 vss.n6306 vss.n6305 16.2531
R17162 vss.n6305 vss.n245 16.2531
R17163 vss.n15700 vss.n245 16.2531
R17164 vss.n15700 vss.n15699 16.2531
R17165 vss.n15699 vss.n246 16.2531
R17166 vss.n15689 vss.n246 16.2531
R17167 vss.n15595 vss.n15594 16.2531
R17168 vss.n15594 vss.n15580 16.2531
R17169 vss.n15618 vss.n15580 16.2531
R17170 vss.n15618 vss.n15617 16.2531
R17171 vss.n15617 vss.n15581 16.2531
R17172 vss.n15613 vss.n15581 16.2531
R17173 vss.n347 vss.n346 16.2531
R17174 vss.n346 vss.n345 16.2531
R17175 vss.n345 vss.n310 16.2531
R17176 vss.n335 vss.n310 16.2531
R17177 vss.n335 vss.n334 16.2531
R17178 vss.n334 vss.n333 16.2531
R17179 vss.n3594 vss.n3593 16.2531
R17180 vss.n3595 vss.n3594 16.2531
R17181 vss.n3595 vss.n3569 16.2531
R17182 vss.n3606 vss.n3569 16.2531
R17183 vss.n3607 vss.n3606 16.2531
R17184 vss.n3608 vss.n3607 16.2531
R17185 vss.n377 vss.n376 16.2531
R17186 vss.n376 vss.n361 16.2531
R17187 vss.n15574 vss.n361 16.2531
R17188 vss.n15574 vss.n15573 16.2531
R17189 vss.n15573 vss.n362 16.2531
R17190 vss.n15563 vss.n362 16.2531
R17191 vss.n12177 vss.n12176 16.2531
R17192 vss.n12176 vss.n12175 16.2531
R17193 vss.n12175 vss.n12140 16.2531
R17194 vss.n12165 vss.n12140 16.2531
R17195 vss.n12165 vss.n12164 16.2531
R17196 vss.n12164 vss.n12163 16.2531
R17197 vss.n11770 vss.n11767 16.2531
R17198 vss.n11770 vss.n11759 16.2531
R17199 vss.n11800 vss.n11759 16.2531
R17200 vss.n11800 vss.n11799 16.2531
R17201 vss.n11799 vss.n11760 16.2531
R17202 vss.n11782 vss.n11760 16.2531
R17203 vss.n10441 vss.n10440 16.2531
R17204 vss.n10440 vss.n10425 16.2531
R17205 vss.n10469 vss.n10425 16.2531
R17206 vss.n10469 vss.n10468 16.2531
R17207 vss.n10468 vss.n10426 16.2531
R17208 vss.n10458 vss.n10426 16.2531
R17209 vss.n10586 vss.n10585 16.2531
R17210 vss.n10585 vss.n10570 16.2531
R17211 vss.n10614 vss.n10570 16.2531
R17212 vss.n10614 vss.n10613 16.2531
R17213 vss.n10613 vss.n10571 16.2531
R17214 vss.n10603 vss.n10571 16.2531
R17215 vss.n10980 vss.n10979 16.2531
R17216 vss.n10979 vss.n10964 16.2531
R17217 vss.n11008 vss.n10964 16.2531
R17218 vss.n11008 vss.n11007 16.2531
R17219 vss.n11007 vss.n10965 16.2531
R17220 vss.n10997 vss.n10965 16.2531
R17221 vss.n10005 vss.n9995 16.2531
R17222 vss.n10029 vss.n10005 16.2531
R17223 vss.n10029 vss.n10028 16.2531
R17224 vss.n10028 vss.n10026 16.2531
R17225 vss.n10026 vss.n10008 16.2531
R17226 vss.n10016 vss.n10008 16.2531
R17227 vss.n9962 vss.n9951 16.2531
R17228 vss.n9963 vss.n9962 16.2531
R17229 vss.n11637 vss.n9963 16.2531
R17230 vss.n11637 vss.n11636 16.2531
R17231 vss.n11636 vss.n11619 16.2531
R17232 vss.n11622 vss.n11619 16.2531
R17233 vss.n11675 vss.n11674 15.2779
R17234 vss.n11674 vss.n11673 15.2779
R17235 vss.n11663 vss.n11652 15.2779
R17236 vss.n11663 vss.n11662 15.2779
R17237 vss.n11662 vss.n11661 15.2779
R17238 vss.n11438 vss.n11437 15.2779
R17239 vss.n11437 vss.n11436 15.2779
R17240 vss.n11426 vss.n11415 15.2779
R17241 vss.n11426 vss.n11425 15.2779
R17242 vss.n11425 vss.n11424 15.2779
R17243 vss.n11033 vss.n10078 15.2779
R17244 vss.n11306 vss.n10078 15.2779
R17245 vss.n11317 vss.n10061 15.2779
R17246 vss.n11318 vss.n11317 15.2779
R17247 vss.n11319 vss.n11318 15.2779
R17248 vss.n10781 vss.n10780 15.2779
R17249 vss.n10780 vss.n10779 15.2779
R17250 vss.n10769 vss.n10703 15.2779
R17251 vss.n10769 vss.n10768 15.2779
R17252 vss.n10768 vss.n10767 15.2779
R17253 vss.n8370 vss.n8360 15.2779
R17254 vss.n13675 vss.n8370 15.2779
R17255 vss.n13675 vss.n13674 15.2779
R17256 vss.n13672 vss.n8372 15.2779
R17257 vss.n13662 vss.n8372 15.2779
R17258 vss.n8334 vss.n8324 15.2779
R17259 vss.n13705 vss.n8334 15.2779
R17260 vss.n13705 vss.n13704 15.2779
R17261 vss.n13381 vss.n8336 15.2779
R17262 vss.n13413 vss.n13381 15.2779
R17263 vss.n8500 vss.n8490 15.2779
R17264 vss.n13294 vss.n8500 15.2779
R17265 vss.n13294 vss.n13293 15.2779
R17266 vss.n8616 vss.n8502 15.2779
R17267 vss.n8606 vss.n8502 15.2779
R17268 vss.n12944 vss.n9176 15.2779
R17269 vss.n12993 vss.n12944 15.2779
R17270 vss.n12993 vss.n12992 15.2779
R17271 vss.n12990 vss.n12946 15.2779
R17272 vss.n12980 vss.n12946 15.2779
R17273 vss.n8914 vss.n8904 15.2779
R17274 vss.n13152 vss.n8914 15.2779
R17275 vss.n13152 vss.n13151 15.2779
R17276 vss.n13149 vss.n8916 15.2779
R17277 vss.n13139 vss.n8916 15.2779
R17278 vss.n9362 vss.n9305 15.2779
R17279 vss.n12894 vss.n9362 15.2779
R17280 vss.n12894 vss.n12893 15.2779
R17281 vss.n9378 vss.n9377 15.2779
R17282 vss.n12874 vss.n9378 15.2779
R17283 vss.n12698 vss.n12642 15.2779
R17284 vss.n12817 vss.n12698 15.2779
R17285 vss.n12817 vss.n12816 15.2779
R17286 vss.n12714 vss.n12713 15.2779
R17287 vss.n12797 vss.n12714 15.2779
R17288 vss.n285 vss.n283 15.2779
R17289 vss.n15676 vss.n285 15.2779
R17290 vss.n15676 vss.n15675 15.2779
R17291 vss.n6257 vss.n6256 15.2779
R17292 vss.n6258 vss.n6257 15.2779
R17293 vss.n6258 vss.n19 15.2779
R17294 vss.n214 vss.n204 15.2779
R17295 vss.n15733 vss.n214 15.2779
R17296 vss.n15733 vss.n15732 15.2779
R17297 vss.n136 vss.n126 15.2779
R17298 vss.n15789 vss.n136 15.2779
R17299 vss.n15789 vss.n15788 15.2779
R17300 vss.n57 vss.n47 15.2779
R17301 vss.n15845 vss.n57 15.2779
R17302 vss.n15845 vss.n15844 15.2779
R17303 vss.n914 vss.n904 15.2779
R17304 vss.n15225 vss.n914 15.2779
R17305 vss.n15225 vss.n15224 15.2779
R17306 vss.n855 vss.n799 15.2779
R17307 vss.n15268 vss.n855 15.2779
R17308 vss.n15268 vss.n15267 15.2779
R17309 vss.n756 vss.n746 15.2779
R17310 vss.n15345 vss.n756 15.2779
R17311 vss.n15345 vss.n15344 15.2779
R17312 vss.n657 vss.n647 15.2779
R17313 vss.n15375 vss.n657 15.2779
R17314 vss.n15375 vss.n15374 15.2779
R17315 vss.n598 vss.n541 15.2779
R17316 vss.n15418 vss.n598 15.2779
R17317 vss.n15418 vss.n15417 15.2779
R17318 vss.n450 vss.n440 15.2779
R17319 vss.n15450 vss.n450 15.2779
R17320 vss.n15450 vss.n15449 15.2779
R17321 vss.n4869 vss.n4868 15.2779
R17322 vss.n4870 vss.n4869 15.2779
R17323 vss.n4870 vss.n4310 15.2779
R17324 vss.n1693 vss.n1683 15.2779
R17325 vss.n14530 vss.n1693 15.2779
R17326 vss.n14530 vss.n14529 15.2779
R17327 vss.n1634 vss.n1578 15.2779
R17328 vss.n14573 vss.n1634 15.2779
R17329 vss.n14573 vss.n14572 15.2779
R17330 vss.n1535 vss.n1525 15.2779
R17331 vss.n14650 vss.n1535 15.2779
R17332 vss.n14650 vss.n14649 15.2779
R17333 vss.n1436 vss.n1426 15.2779
R17334 vss.n14680 vss.n1436 15.2779
R17335 vss.n14680 vss.n14679 15.2779
R17336 vss.n1377 vss.n1320 15.2779
R17337 vss.n14723 vss.n1377 15.2779
R17338 vss.n14723 vss.n14722 15.2779
R17339 vss.n1229 vss.n1219 15.2779
R17340 vss.n14755 vss.n1229 15.2779
R17341 vss.n14755 vss.n14754 15.2779
R17342 vss.n2419 vss.n2363 15.2779
R17343 vss.n8022 vss.n2419 15.2779
R17344 vss.n8022 vss.n8021 15.2779
R17345 vss.n1868 vss.n1858 15.2779
R17346 vss.n14329 vss.n1868 15.2779
R17347 vss.n14329 vss.n14328 15.2779
R17348 vss.n1089 vss.n1079 15.2779
R17349 vss.n15024 vss.n1089 15.2779
R17350 vss.n15024 vss.n15023 15.2779
R17351 vss.n81 vss.n71 15.2779
R17352 vss.n15818 vss.n81 15.2779
R17353 vss.n15818 vss.n15817 15.2779
R17354 vss.n160 vss.n150 15.2779
R17355 vss.n15762 vss.n160 15.2779
R17356 vss.n15762 vss.n15761 15.2779
R17357 vss.n238 vss.n228 15.2779
R17358 vss.n15706 vss.n238 15.2779
R17359 vss.n15706 vss.n15705 15.2779
R17360 vss.n12077 vss.n11936 15.2779
R17361 vss.n12087 vss.n11936 15.2779
R17362 vss.n12088 vss.n12087 15.2779
R17363 vss.n12107 vss.n12106 15.2779
R17364 vss.n12106 vss.n11875 15.2779
R17365 vss.n10391 vss.n10253 15.2779
R17366 vss.n10619 vss.n10253 15.2779
R17367 vss.n10630 vss.n10236 15.2779
R17368 vss.n10631 vss.n10630 15.2779
R17369 vss.n10632 vss.n10631 15.2779
R17370 vss.n10759 vss.n10166 15.2779
R17371 vss.n11012 vss.n10166 15.2779
R17372 vss.n11023 vss.n10149 15.2779
R17373 vss.n11024 vss.n11023 15.2779
R17374 vss.n11025 vss.n11024 15.2779
R17375 vss.n11330 vss.n11329 15.2779
R17376 vss.n11332 vss.n11330 15.2779
R17377 vss.n11343 vss.n9989 15.2779
R17378 vss.n11344 vss.n11343 15.2779
R17379 vss.n11345 vss.n11344 15.2779
R17380 vss.n10368 vss.n10367 15.2779
R17381 vss.n10370 vss.n10368 15.2779
R17382 vss.n10381 vss.n10278 15.2779
R17383 vss.n10382 vss.n10381 15.2779
R17384 vss.n10383 vss.n10382 15.2779
R17385 vss.n11673 vss.n9935 14.9682
R17386 vss.n11436 vss.n9964 14.9682
R17387 vss.n11306 vss.n11305 14.9682
R17388 vss.n10779 vss.n10641 14.9682
R17389 vss.n13673 vss.n13672 14.9682
R17390 vss.n13703 vss.n8336 14.9682
R17391 vss.n13292 vss.n8616 14.9682
R17392 vss.n12991 vss.n12990 14.9682
R17393 vss.n13150 vss.n13149 14.9682
R17394 vss.n9377 vss.n8880 14.9682
R17395 vss.n12713 vss.n8881 14.9682
R17396 vss.n15674 vss.n15673 14.9682
R17397 vss.n15874 vss.n15872 14.9682
R17398 vss.n15731 vss.n15730 14.9682
R17399 vss.n15787 vss.n15786 14.9682
R17400 vss.n15843 vss.n15842 14.9682
R17401 vss.n15223 vss.n916 14.9682
R17402 vss.n15266 vss.n15265 14.9682
R17403 vss.n15343 vss.n758 14.9682
R17404 vss.n15373 vss.n659 14.9682
R17405 vss.n15416 vss.n15415 14.9682
R17406 vss.n15448 vss.n452 14.9682
R17407 vss.n4305 vss.n500 14.9682
R17408 vss.n14528 vss.n1695 14.9682
R17409 vss.n14571 vss.n14570 14.9682
R17410 vss.n14648 vss.n1537 14.9682
R17411 vss.n14678 vss.n1438 14.9682
R17412 vss.n14721 vss.n14720 14.9682
R17413 vss.n14753 vss.n1231 14.9682
R17414 vss.n2434 vss.n1279 14.9682
R17415 vss.n14327 vss.n1986 14.9682
R17416 vss.n15022 vss.n1091 14.9682
R17417 vss.n15816 vss.n83 14.9682
R17418 vss.n15760 vss.n162 14.9682
R17419 vss.n15704 vss.n240 14.9682
R17420 vss.n12107 vss.n9859 14.9682
R17421 vss.n10619 vss.n10618 14.9682
R17422 vss.n11012 vss.n11011 14.9682
R17423 vss.n11332 vss.n11331 14.9682
R17424 vss.n10370 vss.n10369 14.9682
R17425 vss.n15661 vss.n292 13.5231
R17426 vss.n15673 vss.n292 13.5231
R17427 vss.n15878 vss.n15875 13.5231
R17428 vss.n15875 vss.n15874 13.5231
R17429 vss.n15718 vss.n216 13.5231
R17430 vss.n15730 vss.n216 13.5231
R17431 vss.n15774 vss.n138 13.5231
R17432 vss.n15786 vss.n138 13.5231
R17433 vss.n15830 vss.n59 13.5231
R17434 vss.n15842 vss.n59 13.5231
R17435 vss.n6570 vss.n6567 13.5231
R17436 vss.n6548 vss.n6545 13.5231
R17437 vss.n6548 vss.n6547 13.5231
R17438 vss.n6547 vss.n6496 13.5231
R17439 vss.n6566 vss.n6496 13.5231
R17440 vss.n6567 vss.n6566 13.5231
R17441 vss.n5383 vss.n5380 13.5231
R17442 vss.n5361 vss.n5358 13.5231
R17443 vss.n5361 vss.n5360 13.5231
R17444 vss.n5360 vss.n5309 13.5231
R17445 vss.n5379 vss.n5309 13.5231
R17446 vss.n5380 vss.n5379 13.5231
R17447 vss.n640 vss.n638 13.5231
R17448 vss.n624 vss.n612 13.5231
R17449 vss.n625 vss.n624 13.5231
R17450 vss.n626 vss.n625 13.5231
R17451 vss.n637 vss.n626 13.5231
R17452 vss.n638 vss.n637 13.5231
R17453 vss.n4908 vss.n4905 13.5231
R17454 vss.n4886 vss.n4883 13.5231
R17455 vss.n4886 vss.n4885 13.5231
R17456 vss.n4885 vss.n4264 13.5231
R17457 vss.n4904 vss.n4264 13.5231
R17458 vss.n4905 vss.n4904 13.5231
R17459 vss.n5171 vss.n5168 13.5231
R17460 vss.n5149 vss.n5146 13.5231
R17461 vss.n5149 vss.n5148 13.5231
R17462 vss.n5148 vss.n5097 13.5231
R17463 vss.n5167 vss.n5097 13.5231
R17464 vss.n5168 vss.n5167 13.5231
R17465 vss.n897 vss.n895 13.5231
R17466 vss.n881 vss.n869 13.5231
R17467 vss.n882 vss.n881 13.5231
R17468 vss.n883 vss.n882 13.5231
R17469 vss.n894 vss.n883 13.5231
R17470 vss.n895 vss.n894 13.5231
R17471 vss.n6455 vss.n6452 13.5231
R17472 vss.n6433 vss.n6430 13.5231
R17473 vss.n6433 vss.n6432 13.5231
R17474 vss.n6432 vss.n6381 13.5231
R17475 vss.n6451 vss.n6381 13.5231
R17476 vss.n6452 vss.n6451 13.5231
R17477 vss.n4857 vss.n4856 13.5231
R17478 vss.n4832 vss.n4830 13.5231
R17479 vss.n4832 vss.n4831 13.5231
R17480 vss.n4831 vss.n4750 13.5231
R17481 vss.n4855 vss.n4750 13.5231
R17482 vss.n4856 vss.n4855 13.5231
R17483 vss.n6443 vss.n6411 13.5231
R17484 vss.n6411 vss.n916 13.5231
R17485 vss.n15246 vss.n857 13.5231
R17486 vss.n15265 vss.n857 13.5231
R17487 vss.n5371 vss.n5339 13.5231
R17488 vss.n5339 vss.n758 13.5231
R17489 vss.n5159 vss.n5127 13.5231
R17490 vss.n5127 vss.n659 13.5231
R17491 vss.n15396 vss.n600 13.5231
R17492 vss.n15415 vss.n600 13.5231
R17493 vss.n4811 vss.n4809 13.5231
R17494 vss.n4811 vss.n452 13.5231
R17495 vss.n4896 vss.n4294 13.5231
R17496 vss.n4305 vss.n4294 13.5231
R17497 vss.n1956 vss.n1954 13.5231
R17498 vss.n1889 vss.n1882 13.5231
R17499 vss.n1882 vss.n1881 13.5231
R17500 vss.n1881 vss.n1138 13.5231
R17501 vss.n1953 vss.n1138 13.5231
R17502 vss.n1954 vss.n1953 13.5231
R17503 vss.n2797 vss.n2794 13.5231
R17504 vss.n2775 vss.n2772 13.5231
R17505 vss.n2775 vss.n2774 13.5231
R17506 vss.n2774 vss.n2723 13.5231
R17507 vss.n2793 vss.n2723 13.5231
R17508 vss.n2794 vss.n2793 13.5231
R17509 vss.n1419 vss.n1417 13.5231
R17510 vss.n1403 vss.n1391 13.5231
R17511 vss.n1404 vss.n1403 13.5231
R17512 vss.n1405 vss.n1404 13.5231
R17513 vss.n1416 vss.n1405 13.5231
R17514 vss.n1417 vss.n1416 13.5231
R17515 vss.n6950 vss.n6947 13.5231
R17516 vss.n2428 vss.n2427 13.5231
R17517 vss.n2446 vss.n2428 13.5231
R17518 vss.n7998 vss.n2446 13.5231
R17519 vss.n7998 vss.n2447 13.5231
R17520 vss.n6947 vss.n2447 13.5231
R17521 vss.n7579 vss.n7576 13.5231
R17522 vss.n7557 vss.n7554 13.5231
R17523 vss.n7557 vss.n7556 13.5231
R17524 vss.n7556 vss.n7505 13.5231
R17525 vss.n7575 vss.n7505 13.5231
R17526 vss.n7576 vss.n7575 13.5231
R17527 vss.n1676 vss.n1674 13.5231
R17528 vss.n1660 vss.n1648 13.5231
R17529 vss.n1661 vss.n1660 13.5231
R17530 vss.n1662 vss.n1661 13.5231
R17531 vss.n1673 vss.n1662 13.5231
R17532 vss.n1674 vss.n1673 13.5231
R17533 vss.n2562 vss.n2559 13.5231
R17534 vss.n2541 vss.n2540 13.5231
R17535 vss.n2541 vss.n2513 13.5231
R17536 vss.n2557 vss.n2513 13.5231
R17537 vss.n2558 vss.n2557 13.5231
R17538 vss.n2559 vss.n2558 13.5231
R17539 vss.n3217 vss.n3214 13.5231
R17540 vss.n3243 vss.n3240 13.5231
R17541 vss.n3240 vss.n3185 13.5231
R17542 vss.n3271 vss.n3185 13.5231
R17543 vss.n3271 vss.n3186 13.5231
R17544 vss.n3214 vss.n3186 13.5231
R17545 vss.n2551 vss.n2519 13.5231
R17546 vss.n2519 vss.n1695 13.5231
R17547 vss.n14551 vss.n1636 13.5231
R17548 vss.n14570 vss.n1636 13.5231
R17549 vss.n2785 vss.n2753 13.5231
R17550 vss.n2753 vss.n1537 13.5231
R17551 vss.n7567 vss.n7535 13.5231
R17552 vss.n7535 vss.n1438 13.5231
R17553 vss.n14701 vss.n1379 13.5231
R17554 vss.n14720 vss.n1379 13.5231
R17555 vss.n3233 vss.n3231 13.5231
R17556 vss.n3233 vss.n1231 13.5231
R17557 vss.n8002 vss.n2435 13.5231
R17558 vss.n2435 vss.n2434 13.5231
R17559 vss.n12128 vss.n12127 13.5231
R17560 vss.n12097 vss.n12095 13.5231
R17561 vss.n12097 vss.n12096 13.5231
R17562 vss.n12096 vss.n2034 13.5231
R17563 vss.n12126 vss.n2034 13.5231
R17564 vss.n12127 vss.n12126 13.5231
R17565 vss.n12070 vss.n12069 13.5231
R17566 vss.n8390 vss.n8387 13.5231
R17567 vss.n8405 vss.n8387 13.5231
R17568 vss.n13658 vss.n8405 13.5231
R17569 vss.n13658 vss.n8406 13.5231
R17570 vss.n12069 vss.n8406 13.5231
R17571 vss.n8577 vss.n8574 13.5231
R17572 vss.n8596 vss.n8593 13.5231
R17573 vss.n8596 vss.n8595 13.5231
R17574 vss.n8595 vss.n8407 13.5231
R17575 vss.n8578 vss.n8407 13.5231
R17576 vss.n8578 vss.n8577 13.5231
R17577 vss.n9168 vss.n9167 13.5231
R17578 vss.n8934 vss.n8931 13.5231
R17579 vss.n8949 vss.n8931 13.5231
R17580 vss.n13135 vss.n8949 13.5231
R17581 vss.n13135 vss.n8950 13.5231
R17582 vss.n9167 vss.n8950 13.5231
R17583 vss.n9417 vss.n9414 13.5231
R17584 vss.n9371 vss.n9370 13.5231
R17585 vss.n9389 vss.n9371 13.5231
R17586 vss.n12870 vss.n9389 13.5231
R17587 vss.n12870 vss.n9390 13.5231
R17588 vss.n9414 vss.n9390 13.5231
R17589 vss.n12780 vss.n12726 13.5231
R17590 vss.n12707 vss.n12706 13.5231
R17591 vss.n12725 vss.n12707 13.5231
R17592 vss.n12793 vss.n12725 13.5231
R17593 vss.n12793 vss.n12792 13.5231
R17594 vss.n12792 vss.n12726 13.5231
R17595 vss.n8439 vss.n8436 13.5231
R17596 vss.n12973 vss.n12958 13.5231
R17597 vss.n12974 vss.n12973 13.5231
R17598 vss.n12974 vss.n8409 13.5231
R17599 vss.n8435 vss.n8409 13.5231
R17600 vss.n8436 vss.n8435 13.5231
R17601 vss.n13425 vss.n13422 13.5231
R17602 vss.n13402 vss.n13399 13.5231
R17603 vss.n13402 vss.n13401 13.5231
R17604 vss.n13401 vss.n13351 13.5231
R17605 vss.n13421 vss.n13351 13.5231
R17606 vss.n13422 vss.n13421 13.5231
R17607 vss.n1967 vss.n1870 13.5231
R17608 vss.n1986 vss.n1870 13.5231
R17609 vss.n6558 vss.n6526 13.5231
R17610 vss.n6526 vss.n1091 13.5231
R17611 vss.n107 vss.n105 13.5231
R17612 vss.n107 vss.n83 13.5231
R17613 vss.n185 vss.n183 13.5231
R17614 vss.n185 vss.n162 13.5231
R17615 vss.n264 vss.n262 13.5231
R17616 vss.n264 vss.n240 13.5231
R17617 vss.n3244 vss.n1225 13.0005
R17618 vss.n3267 vss.n3228 13.0005
R17619 vss.n2420 vss.n2415 13.0005
R17620 vss.n6961 vss.n2440 13.0005
R17621 vss.n1397 vss.n1373 13.0005
R17622 vss.n14704 vss.n14698 13.0005
R17623 vss.n7547 vss.n1432 13.0005
R17624 vss.n7590 vss.n7524 13.0005
R17625 vss.n2765 vss.n1531 13.0005
R17626 vss.n2808 vss.n2742 13.0005
R17627 vss.n1654 vss.n1630 13.0005
R17628 vss.n14554 vss.n14548 13.0005
R17629 vss.n2533 vss.n1689 13.0005
R17630 vss.n2573 vss.n2506 13.0005
R17631 vss.n1886 vss.n1864 13.0005
R17632 vss.n1970 vss.n1964 13.0005
R17633 vss.n4822 vss.n446 13.0005
R17634 vss.n4845 vss.n4800 13.0005
R17635 vss.n4360 vss.n4304 13.0005
R17636 vss.n4919 vss.n4283 13.0005
R17637 vss.n618 vss.n594 13.0005
R17638 vss.n15399 vss.n15393 13.0005
R17639 vss.n5139 vss.n653 13.0005
R17640 vss.n5182 vss.n5116 13.0005
R17641 vss.n5351 vss.n752 13.0005
R17642 vss.n5394 vss.n5328 13.0005
R17643 vss.n875 vss.n851 13.0005
R17644 vss.n15249 vss.n15243 13.0005
R17645 vss.n6423 vss.n910 13.0005
R17646 vss.n6466 vss.n6400 13.0005
R17647 vss.n6538 vss.n1085 13.0005
R17648 vss.n6582 vss.n6515 13.0005
R17649 vss.n9363 vss.n9358 13.0005
R17650 vss.n12840 vss.n9383 13.0005
R17651 vss.n12699 vss.n12694 13.0005
R17652 vss.n12775 vss.n12719 13.0005
R17653 vss.n8938 vss.n8910 13.0005
R17654 vss.n9159 vss.n8927 13.0005
R17655 vss.n12963 vss.n12940 13.0005
R17656 vss.n13317 vss.n8428 13.0005
R17657 vss.n8590 vss.n8496 13.0005
R17658 vss.n8564 vss.n8513 13.0005
R17659 vss.n13396 vss.n8330 13.0005
R17660 vss.n13436 vss.n13370 13.0005
R17661 vss.n8394 vss.n8366 13.0005
R17662 vss.n12061 vss.n8383 13.0005
R17663 vss.n12092 vss.n11935 13.0005
R17664 vss.n12116 vss.n11866 13.0005
R17665 vss.n6741 vss 7.1255
R17666 vss.n13183 vss.n13182 7.05642
R17667 vss.n3272 vss.n2144 6.93142
R17668 vss.n6743 vss.n6742 6.93142
R17669 vss.n12189 vss.n9860 5.17978
R17670 vss.n15578 vss.n15577 5.17978
R17671 vss.n15020 vss.n14887 5.17978
R17672 vss.n14325 vss.n14192 5.17978
R17673 vss.n13182 vss.n2144 5.10905
R17674 vss.n6743 vss.n3272 5.10905
R17675 vss.n6742 vss.n6741 5.10905
R17676 vss.n14805 vss 4.95527
R17677 vss vss.n1167 4.83932
R17678 vss.n15576 vss 4.83932
R17679 vss.n12139 vss 4.7579
R17680 vss.n15500 vss 4.7579
R17681 vss vss.n388 4.64195
R17682 vss vss.n9860 4.35741
R17683 vss.n15577 vss 4.35741
R17684 vss.n14887 vss 4.35741
R17685 vss.n14192 vss 4.35741
R17686 vss.n12138 vss.n9860 3.55067
R17687 vss.n11801 vss.n11757 2.88866
R17688 vss.n12500 vss.n9472 2.88866
R17689 vss.n5046 vss.n5045 2.88866
R17690 vss.n5520 vss.n5519 2.88866
R17691 vss.n4493 vss.n4446 2.88866
R17692 vss.n14976 vss.n14935 2.88866
R17693 vss.n15172 vss.n965 2.88866
R17694 vss.n4701 vss.n4654 2.88866
R17695 vss.n7992 vss.n7991 2.88866
R17696 vss.n7718 vss.n7717 2.88866
R17697 vss.n7207 vss.n7206 2.88866
R17698 vss.n14281 vss.n14240 2.88866
R17699 vss.n14477 vss.n1744 2.88866
R17700 vss.n8051 vss.n8049 2.88866
R17701 vss.n14088 vss.n14087 2.88866
R17702 vss.n13129 vss.n13081 2.88866
R17703 vss.n13841 vss.n13793 2.88866
R17704 vss.n13652 vss.n13604 2.88866
R17705 vss.n15621 vss.n359 2.88866
R17706 vss.n10518 vss.n10470 2.88866
R17707 vss.n10912 vss.n10864 2.88866
R17708 vss.n11299 vss.n11251 2.88866
R17709 vss.n11610 vss.n11562 2.88866
R17710 vss.n12381 vss.n9601 2.88866
R17711 vss.n12263 vss.n9731 2.88866
R17712 vss.n6376 vss.n6375 2.88866
R17713 vss.n7350 vss.n7348 2.88866
R17714 vss.n7913 vss.n7912 2.88866
R17715 vss.n13980 vss.n8151 2.88866
R17716 vss.n6062 vss.n6015 2.88866
R17717 vss.n5822 vss.n5775 2.88866
R17718 vss.n5680 vss.n5587 2.88866
R17719 vss.n15577 vss.n15576 2.43143
R17720 vss.n14887 vss.n388 2.43143
R17721 vss.n14192 vss.n1167 2.43143
R17722 vss.n14324 vss.n14282 1.89112
R17723 vss.n15019 vss.n14977 1.89112
R17724 vss.n15620 vss.n15619 1.89112
R17725 vss.n12188 vss.n11802 1.89112
R17726 vss.n4788 vss 1.87386
R17727 vss.n6791 vss 1.87386
R17728 vss.n12869 vss 1.87386
R17729 vss.n10254 vss 1.87386
R17730 vss.n6613 vss.n6496 1.52776
R17731 vss.n5423 vss.n5309 1.52776
R17732 vss.n4127 vss.n626 1.52776
R17733 vss.n4949 vss.n4264 1.52776
R17734 vss.n5212 vss.n5097 1.52776
R17735 vss.n3387 vss.n883 1.52776
R17736 vss.n6495 vss.n6381 1.52776
R17737 vss.n4788 vss.n4750 1.52776
R17738 vss.n14886 vss.n1138 1.52776
R17739 vss.n2837 vss.n2723 1.52776
R17740 vss.n2449 vss.n1405 1.52776
R17741 vss.n7998 vss.n7997 1.52776
R17742 vss.n7620 vss.n7505 1.52776
R17743 vss.n7815 vss.n1662 1.52776
R17744 vss.n2557 vss.n1139 1.52776
R17745 vss.n6791 vss.n3271 1.52776
R17746 vss.n14191 vss.n2034 1.52776
R17747 vss.n13658 vss.n13657 1.52776
R17748 vss.n13349 vss.n8407 1.52776
R17749 vss.n13135 vss.n13134 1.52776
R17750 vss.n12870 vss.n12869 1.52776
R17751 vss.n12793 vss.n8951 1.52776
R17752 vss.n13347 vss.n8409 1.52776
R17753 vss.n13466 vss.n13351 1.52776
R17754 vss.n11616 vss.n11615 1.44293
R17755 vss.n11304 vss.n10079 1.44293
R17756 vss.n10962 vss.n10167 1.44293
R17757 vss.n10568 vss.n10254 1.44293
R17758 vss.n12191 vss.n12190 1.44293
R17759 vss.n12191 vss.n8338 1.44293
R17760 vss.n13702 vss.n8337 1.44293
R17761 vss.n13702 vss.n13701 1.44293
R17762 vss.n13701 vss.n8338 1.44293
R17763 vss.n13291 vss.n8337 1.44293
R17764 vss.n12428 vss.n8617 1.44293
R17765 vss.n13290 vss.n8617 1.44293
R17766 vss.n12428 vss.n8882 1.44293
R17767 vss.n13181 vss.n13180 1.44293
R17768 vss.n13180 vss.n13179 1.44293
R17769 vss.n13179 vss.n13178 1.44293
R17770 vss.n13178 vss.n8882 1.44293
R17771 vss.n241 vss.n163 1.44293
R17772 vss.n5869 vss.n85 1.44293
R17773 vss.n15870 vss.n27 1.44293
R17774 vss.n84 vss.n27 1.44293
R17775 vss.n5423 vss.n5308 1.44293
R17776 vss.n5096 vss.n4127 1.44293
R17777 vss.n4949 vss.n4263 1.44293
R17778 vss.n4950 vss.n4949 1.44293
R17779 vss.n4950 vss.n4127 1.44293
R17780 vss.n5212 vss.n5096 1.44293
R17781 vss.n5424 vss.n5423 1.44293
R17782 vss.n5308 vss.n3387 1.44293
R17783 vss.n6380 vss.n3387 1.44293
R17784 vss.n6495 vss.n6380 1.44293
R17785 vss.n6614 vss.n6495 1.44293
R17786 vss.n6614 vss.n6613 1.44293
R17787 vss.n4788 vss.n4263 1.44293
R17788 vss.n15222 vss.n917 1.44293
R17789 vss.n15294 vss.n759 1.44293
R17790 vss.n15221 vss.n759 1.44293
R17791 vss.n15222 vss.n15221 1.44293
R17792 vss.n15342 vss.n15294 1.44293
R17793 vss.n15372 vss.n660 1.44293
R17794 vss.n15372 vss.n15371 1.44293
R17795 vss.n660 vss.n501 1.44293
R17796 vss.n15447 vss.n15446 1.44293
R17797 vss.n15446 vss.n15445 1.44293
R17798 vss.n15445 vss.n15444 1.44293
R17799 vss.n15444 vss.n501 1.44293
R17800 vss.n7768 vss.n2837 1.44293
R17801 vss.n7504 vss.n2449 1.44293
R17802 vss.n7997 vss.n2448 1.44293
R17803 vss.n7997 vss.n7996 1.44293
R17804 vss.n7996 vss.n2449 1.44293
R17805 vss.n7620 vss.n7504 1.44293
R17806 vss.n7621 vss.n2837 1.44293
R17807 vss.n7815 vss.n7768 1.44293
R17808 vss.n7816 vss.n7815 1.44293
R17809 vss.n7816 vss.n1139 1.44293
R17810 vss.n14885 vss.n1139 1.44293
R17811 vss.n14886 vss.n14885 1.44293
R17812 vss.n6791 vss.n2448 1.44293
R17813 vss.n14527 vss.n1696 1.44293
R17814 vss.n14599 vss.n1538 1.44293
R17815 vss.n14526 vss.n1538 1.44293
R17816 vss.n14527 vss.n14526 1.44293
R17817 vss.n14647 vss.n14599 1.44293
R17818 vss.n14677 vss.n1439 1.44293
R17819 vss.n14677 vss.n14676 1.44293
R17820 vss.n1439 vss.n1280 1.44293
R17821 vss.n14752 vss.n14751 1.44293
R17822 vss.n14751 vss.n14750 1.44293
R17823 vss.n14750 vss.n14749 1.44293
R17824 vss.n14749 vss.n1280 1.44293
R17825 vss.n13657 vss.n2033 1.44293
R17826 vss.n13350 vss.n13349 1.44293
R17827 vss.n13134 vss.n8408 1.44293
R17828 vss.n12869 vss.n9391 1.44293
R17829 vss.n9391 vss.n8951 1.44293
R17830 vss.n13133 vss.n8951 1.44293
R17831 vss.n13134 vss.n13133 1.44293
R17832 vss.n13347 vss.n8408 1.44293
R17833 vss.n13349 vss.n13348 1.44293
R17834 vss.n13466 vss.n13350 1.44293
R17835 vss.n13656 vss.n13466 1.44293
R17836 vss.n13657 vss.n13656 1.44293
R17837 vss.n14191 vss.n2033 1.44293
R17838 vss.n14326 vss.n1696 1.44293
R17839 vss.n14326 vss.n14325 1.44293
R17840 vss.n15021 vss.n917 1.44293
R17841 vss.n15021 vss.n15020 1.44293
R17842 vss.n15815 vss.n84 1.44293
R17843 vss.n15815 vss.n15814 1.44293
R17844 vss.n15814 vss.n85 1.44293
R17845 vss.n15759 vss.n15758 1.44293
R17846 vss.n15758 vss.n163 1.44293
R17847 vss.n15703 vss.n241 1.44293
R17848 vss.n15703 vss.n15702 1.44293
R17849 vss.n15702 vss.n242 1.44293
R17850 vss.n15578 vss.n242 1.44293
R17851 vss.n12190 vss.n12189 1.44293
R17852 vss.n10617 vss.n10568 1.44293
R17853 vss.n10617 vss.n10616 1.44293
R17854 vss.n10616 vss.n10167 1.44293
R17855 vss.n11010 vss.n10962 1.44293
R17856 vss.n11304 vss.n11303 1.44293
R17857 vss.n10079 vss.n9965 1.44293
R17858 vss.n11614 vss.n9965 1.44293
R17859 vss.n11615 vss.n11614 1.44293
R17860 vss.n11617 vss.n11616 1.44293
R17861 vss.n15871 vss.n15870 1.44293
R17862 vss.n12193 vss.n12192 1.19376
R17863 vss.n13700 vss.n8339 1.19376
R17864 vss.n12311 vss.n12310 1.19376
R17865 vss.n13289 vss.n8618 1.19376
R17866 vss.n12430 vss.n12429 1.19376
R17867 vss.n12502 vss.n12501 1.19376
R17868 vss.n13177 vss.n8883 1.19376
R17869 vss.n4997 vss.n4996 1.19376
R17870 vss.n5095 vss.n5094 1.19376
R17871 vss.n5471 vss.n5470 1.19376
R17872 vss.n5307 vss.n5306 1.19376
R17873 vss.n6379 vss.n6378 1.19376
R17874 vss.n6661 vss.n6660 1.19376
R17875 vss.n4542 vss.n4541 1.19376
R17876 vss.n6740 vss.n6739 1.19376
R17877 vss.n15220 vss.n15174 1.19376
R17878 vss.n15293 vss.n760 1.19376
R17879 vss.n15370 vss.n707 1.19376
R17880 vss.n7347 vss.n7346 1.19376
R17881 vss.n4703 vss.n4702 1.19376
R17882 vss.n15443 vss.n502 1.19376
R17883 vss.n7995 vss.n7994 1.19376
R17884 vss.n7503 vss.n7502 1.19376
R17885 vss.n7668 vss.n7667 1.19376
R17886 vss.n7767 vss.n7766 1.19376
R17887 vss.n7863 vss.n7862 1.19376
R17888 vss.n14884 vss.n14883 1.19376
R17889 vss.n6877 vss.n6876 1.19376
R17890 vss.n6790 vss.n6744 1.19376
R17891 vss.n14525 vss.n14479 1.19376
R17892 vss.n14598 vss.n1539 1.19376
R17893 vss.n14675 vss.n1486 1.19376
R17894 vss.n14027 vss.n14026 1.19376
R17895 vss.n8048 vss.n8047 1.19376
R17896 vss.n14748 vss.n1281 1.19376
R17897 vss.n14091 vss.n14090 1.19376
R17898 vss.n12627 vss.n12626 1.19376
R17899 vss.n13132 vss.n13131 1.19376
R17900 vss.n13033 vss.n13032 1.19376
R17901 vss.n13843 vss.n8254 1.19376
R17902 vss.n13745 vss.n13744 1.19376
R17903 vss.n13655 vss.n13654 1.19376
R17904 vss.n14139 vss.n14138 1.19376
R17905 vss.n14355 vss.n14354 1.19376
R17906 vss.n15050 vss.n15049 1.19376
R17907 vss.n15869 vss.n28 1.19376
R17908 vss.n6110 vss.n6109 1.19376
R17909 vss.n15813 vss.n86 1.19376
R17910 vss.n5871 vss.n5870 1.19376
R17911 vss.n15757 vss.n164 1.19376
R17912 vss.n5678 vss.n5677 1.19376
R17913 vss.n15701 vss.n243 1.19376
R17914 vss.n10567 vss.n10566 1.19376
R17915 vss.n10815 vss.n10814 1.19376
R17916 vss.n10961 vss.n10960 1.19376
R17917 vss.n11302 vss.n11301 1.19376
R17918 vss.n11203 vss.n11202 1.19376
R17919 vss.n11613 vss.n11612 1.19376
R17920 vss.n11709 vss.n11708 1.19376
R17921 vss.n13184 vss.n13183 1.19376
R17922 vss.n14804 vss.n1167 1.11974
R17923 vss.n15499 vss.n388 1.11974
R17924 vss.n15576 vss.n15575 1.11974
R17925 vss.n6613 vss 1.0778
R17926 vss vss.n5212 1.0778
R17927 vss vss.n14886 1.0778
R17928 vss vss.n7620 1.0778
R17929 vss vss.n13347 1.0778
R17930 vss vss.n14191 1.0778
R17931 vss.n11010 vss 1.0778
R17932 vss.n11617 vss 1.0778
R17933 vss.n13291 vss 1.04491
R17934 vss.n15342 vss 1.04491
R17935 vss.n14647 vss 1.04491
R17936 vss.n15759 vss 1.04491
R17937 vss vss.n13181 1.02517
R17938 vss.n15447 vss 1.02517
R17939 vss.n14752 vss 1.02517
R17940 vss.n15871 vss 1.02517
R17941 vss.n5094 vss 0.887013
R17942 vss.n5306 vss 0.887013
R17943 vss.n6661 vss 0.887013
R17944 vss.n4541 vss 0.887013
R17945 vss.n7502 vss 0.887013
R17946 vss.n7766 vss 0.887013
R17947 vss.n14883 vss 0.887013
R17948 vss.n6877 vss 0.887013
R17949 vss.n12626 vss 0.887013
R17950 vss vss.n13033 0.887013
R17951 vss vss.n13745 0.887013
R17952 vss.n14139 vss 0.887013
R17953 vss.n10566 vss 0.887013
R17954 vss.n10960 vss 0.887013
R17955 vss vss.n11203 0.887013
R17956 vss.n11709 vss 0.887013
R17957 vss.n12430 vss 0.854118
R17958 vss.n12311 vss 0.854118
R17959 vss.n12193 vss 0.854118
R17960 vss.n12501 vss 0.854118
R17961 vss.n10815 vss 0.854118
R17962 vss.n11301 vss 0.854118
R17963 vss.n11612 vss 0.854118
R17964 vss vss.n243 0.854118
R17965 vss.n5471 vss 0.854118
R17966 vss.n4997 vss 0.854118
R17967 vss.n6378 vss 0.854118
R17968 vss.n15050 vss 0.854118
R17969 vss vss.n7347 0.854118
R17970 vss vss.n760 0.854118
R17971 vss.n4702 vss 0.854118
R17972 vss.n7668 vss 0.854118
R17973 vss.n7994 vss 0.854118
R17974 vss.n7863 vss 0.854118
R17975 vss.n14355 vss 0.854118
R17976 vss.n14027 vss 0.854118
R17977 vss vss.n1539 0.854118
R17978 vss vss.n8048 0.854118
R17979 vss.n13131 vss 0.854118
R17980 vss vss.n13843 0.854118
R17981 vss.n13654 vss 0.854118
R17982 vss vss.n28 0.854118
R17983 vss vss.n86 0.854118
R17984 vss vss.n164 0.854118
R17985 vss vss.n8339 0.821224
R17986 vss vss.n8618 0.821224
R17987 vss vss.n8883 0.821224
R17988 vss.n5678 vss 0.821224
R17989 vss vss.n5871 0.821224
R17990 vss vss.n6110 0.821224
R17991 vss.n15174 vss 0.821224
R17992 vss vss.n707 0.821224
R17993 vss vss.n502 0.821224
R17994 vss.n14479 vss 0.821224
R17995 vss vss.n1486 0.821224
R17996 vss vss.n1281 0.821224
R17997 vss.n9600 vss.n8618 0.697868
R17998 vss.n9730 vss.n8339 0.697868
R17999 vss.n12194 vss.n12193 0.697868
R18000 vss.n12312 vss.n12311 0.697868
R18001 vss.n12431 vss.n12430 0.697868
R18002 vss.n9471 vss.n8883 0.697868
R18003 vss.n12501 vss.n9470 0.697868
R18004 vss.n6157 vss.n86 0.697868
R18005 vss.n5918 vss.n164 0.697868
R18006 vss.n3541 vss.n243 0.697868
R18007 vss.n4998 vss.n4997 0.697868
R18008 vss.n5094 vss.n5093 0.697868
R18009 vss.n5472 vss.n5471 0.697868
R18010 vss.n5306 vss.n5305 0.697868
R18011 vss.n6378 vss.n6377 0.697868
R18012 vss.n6662 vss.n6661 0.697868
R18013 vss.n6740 vss.n3273 0.697868
R18014 vss.n4541 vss.n4540 0.697868
R18015 vss.n7349 vss.n707 0.697868
R18016 vss.n15174 vss.n15173 0.697868
R18017 vss.n7446 vss.n760 0.697868
R18018 vss.n7347 vss.n7300 0.697868
R18019 vss.n4653 vss.n502 0.697868
R18020 vss.n4702 vss.n4606 0.697868
R18021 vss.n7994 vss.n7993 0.697868
R18022 vss.n7502 vss.n7501 0.697868
R18023 vss.n7669 vss.n7668 0.697868
R18024 vss.n7766 vss.n7765 0.697868
R18025 vss.n7864 vss.n7863 0.697868
R18026 vss.n14883 vss.n14882 0.697868
R18027 vss.n6744 vss.n3149 0.697868
R18028 vss.n6878 vss.n6877 0.697868
R18029 vss.n8150 vss.n1486 0.697868
R18030 vss.n14479 vss.n14478 0.697868
R18031 vss.n13911 vss.n1539 0.697868
R18032 vss.n14028 vss.n14027 0.697868
R18033 vss.n8050 vss.n1281 0.697868
R18034 vss.n8048 vss.n2324 0.697868
R18035 vss.n14090 vss.n14089 0.697868
R18036 vss.n12626 vss.n12625 0.697868
R18037 vss.n13131 vss.n13130 0.697868
R18038 vss.n13033 vss.n9087 0.697868
R18039 vss.n13843 vss.n13842 0.697868
R18040 vss.n13745 vss.n8301 0.697868
R18041 vss.n13654 vss.n13653 0.697868
R18042 vss.n14140 vss.n14139 0.697868
R18043 vss.n14356 vss.n14355 0.697868
R18044 vss.n15051 vss.n15050 0.697868
R18045 vss.n6210 vss.n28 0.697868
R18046 vss.n6110 vss.n6063 0.697868
R18047 vss.n5871 vss.n5823 0.697868
R18048 vss.n5679 vss.n5678 0.697868
R18049 vss.n13183 vss.n8879 0.697868
R18050 vss.n10566 vss.n10565 0.697868
R18051 vss.n10816 vss.n10815 0.697868
R18052 vss.n10960 vss.n10959 0.697868
R18053 vss.n11301 vss.n11300 0.697868
R18054 vss.n11203 vss.n11156 0.697868
R18055 vss.n11612 vss.n11611 0.697868
R18056 vss.n11710 vss.n11709 0.697868
R18057 vss.n6612 vss 0.672375
R18058 vss.n4948 vss 0.672375
R18059 vss.n5211 vss 0.672375
R18060 vss.n3386 vss 0.672375
R18061 vss.n1933 vss 0.672375
R18062 vss.n6974 vss 0.672375
R18063 vss.n7619 vss 0.672375
R18064 vss.n7814 vss 0.672375
R18065 vss.n12763 vss 0.672375
R18066 vss.n13346 vss 0.672375
R18067 vss.n13465 vss 0.672375
R18068 vss.n14190 vss 0.672375
R18069 vss.n10615 vss 0.672375
R18070 vss.n11009 vss 0.672375
R18071 vss.n10027 vss 0.672375
R18072 vss.n11618 vss 0.672375
R18073 vss.n8695 vss 0.662508
R18074 vss.n9811 vss 0.662508
R18075 vss.n9187 vss 0.662508
R18076 vss.n9682 vss 0.662508
R18077 vss.n12653 vss 0.662508
R18078 vss.n9553 vss 0.662508
R18079 vss.n3669 vss 0.662508
R18080 vss.n3788 vss 0.662508
R18081 vss.n3907 vss 0.662508
R18082 vss vss.n5631 0.662508
R18083 vss.n5872 vss 0.662508
R18084 vss.n6111 vss 0.662508
R18085 vss.n994 vss 0.662508
R18086 vss.n810 vss 0.662508
R18087 vss vss.n706 0.662508
R18088 vss.n7399 vss 0.662508
R18089 vss.n4319 vss 0.662508
R18090 vss.n7229 vss 0.662508
R18091 vss.n1773 vss 0.662508
R18092 vss.n1589 vss 0.662508
R18093 vss vss.n1485 0.662508
R18094 vss.n13864 vss 0.662508
R18095 vss.n2374 vss 0.662508
R18096 vss.n8103 vss 0.662508
R18097 vss vss.n2032 0.662508
R18098 vss vss.n1137 0.662508
R18099 vss.n310 vss 0.662508
R18100 vss.n11894 vss 0.662508
R18101 vss vss.n12381 0.662507
R18102 vss vss.n12263 0.662507
R18103 vss.n11757 vss 0.662507
R18104 vss.n12192 vss 0.662507
R18105 vss.n8763 vss 0.662507
R18106 vss vss.n13700 0.662507
R18107 vss.n12310 vss 0.662507
R18108 vss.n8644 vss 0.662507
R18109 vss vss.n13289 0.662507
R18110 vss.n12429 vss 0.662507
R18111 vss.n9214 vss 0.662507
R18112 vss.n9316 vss 0.662507
R18113 vss vss.n12500 0.662507
R18114 vss.n12502 vss 0.662507
R18115 vss vss.n13177 0.662507
R18116 vss.n14935 vss 0.662507
R18117 vss.n7348 vss 0.662507
R18118 vss vss.n964 0.662507
R18119 vss vss.n15220 0.662507
R18120 vss.n965 vss 0.662507
R18121 vss vss.n15293 0.662507
R18122 vss vss.n15341 0.662507
R18123 vss vss.n15370 0.662507
R18124 vss.n7346 vss 0.662507
R18125 vss.n552 vss 0.662507
R18126 vss vss.n499 0.662507
R18127 vss vss.n4701 0.662507
R18128 vss.n4703 vss 0.662507
R18129 vss vss.n15443 0.662507
R18130 vss.n14240 vss 0.662507
R18131 vss vss.n13980 0.662507
R18132 vss vss.n1743 0.662507
R18133 vss vss.n14525 0.662507
R18134 vss.n1744 vss 0.662507
R18135 vss vss.n14598 0.662507
R18136 vss vss.n14646 0.662507
R18137 vss vss.n14675 0.662507
R18138 vss.n14026 vss 0.662507
R18139 vss.n1331 vss 0.662507
R18140 vss vss.n1278 0.662507
R18141 vss.n8049 vss 0.662507
R18142 vss.n8047 vss 0.662507
R18143 vss vss.n14748 0.662507
R18144 vss.n14354 vss 0.662507
R18145 vss vss.n14324 0.662507
R18146 vss.n15049 vss 0.662507
R18147 vss vss.n15019 0.662507
R18148 vss vss.n15869 0.662507
R18149 vss.n6015 vss 0.662507
R18150 vss.n6109 vss 0.662507
R18151 vss.n3856 vss 0.662507
R18152 vss vss.n15813 0.662507
R18153 vss.n5775 vss 0.662507
R18154 vss.n5870 vss 0.662507
R18155 vss.n3737 vss 0.662507
R18156 vss vss.n15757 0.662507
R18157 vss.n5587 vss 0.662507
R18158 vss.n5677 vss 0.662507
R18159 vss.n3618 vss 0.662507
R18160 vss vss.n15701 0.662507
R18161 vss.n15619 vss 0.662507
R18162 vss.n359 vss 0.662507
R18163 vss vss.n12138 0.662507
R18164 vss.n12139 vss 0.662507
R18165 vss vss.n14804 0.662507
R18166 vss.n14805 vss 0.662507
R18167 vss vss.n15499 0.662507
R18168 vss.n15500 vss 0.662507
R18169 vss.n15575 vss 0.662507
R18170 vss vss.n12188 0.662507
R18171 vss.n15904 vss 0.662507
R18172 vss.n11401 vss 0.629613
R18173 vss vss.n10125 0.629613
R18174 vss.n10689 vss 0.629613
R18175 vss vss.n10212 0.629613
R18176 vss vss.n11109 0.629613
R18177 vss vss.n11514 0.629613
R18178 vss vss.n4081 0.629613
R18179 vss vss.n5422 0.629613
R18180 vss vss.n4262 0.629613
R18181 vss vss.n4126 0.629613
R18182 vss.n3519 vss 0.629613
R18183 vss vss.n6494 0.629613
R18184 vss.n4789 vss 0.629613
R18185 vss.n3043 vss 0.629613
R18186 vss vss.n2836 0.629613
R18187 vss.n7065 vss 0.629613
R18188 vss.n7158 vss 0.629613
R18189 vss vss.n2722 0.629613
R18190 vss.n2586 vss 0.629613
R18191 vss.n6792 vss 0.629613
R18192 vss.n12050 vss 0.629613
R18193 vss.n8553 vss 0.629613
R18194 vss.n9148 vss 0.629613
R18195 vss vss.n9040 0.629613
R18196 vss.n13844 vss 0.629613
R18197 vss vss.n13555 0.629613
R18198 vss vss.n12868 0.629613
R18199 vss.n10315 vss 0.629613
R18200 vss vss.n6612 0.629612
R18201 vss vss.n4948 0.629612
R18202 vss.n4996 vss 0.629612
R18203 vss vss.n5046 0.629612
R18204 vss vss.n5095 0.629612
R18205 vss vss.n5211 0.629612
R18206 vss.n5470 vss 0.629612
R18207 vss.n5520 vss 0.629612
R18208 vss vss.n5307 0.629612
R18209 vss vss.n3386 0.629612
R18210 vss.n6375 vss 0.629612
R18211 vss vss.n6379 0.629612
R18212 vss.n6660 vss 0.629612
R18213 vss vss.n4493 0.629612
R18214 vss.n4542 vss 0.629612
R18215 vss.n6739 vss 0.629612
R18216 vss.n1933 vss 0.629612
R18217 vss.n6974 vss 0.629612
R18218 vss vss.n7995 0.629612
R18219 vss.n7991 vss 0.629612
R18220 vss vss.n7503 0.629612
R18221 vss vss.n7619 0.629612
R18222 vss.n7667 vss 0.629612
R18223 vss vss.n7718 0.629612
R18224 vss vss.n7767 0.629612
R18225 vss vss.n7814 0.629612
R18226 vss.n7913 vss 0.629612
R18227 vss.n7862 vss 0.629612
R18228 vss vss.n14884 0.629612
R18229 vss.n7207 vss 0.629612
R18230 vss.n6876 vss 0.629612
R18231 vss vss.n6790 0.629612
R18232 vss.n14091 vss 0.629612
R18233 vss.n14087 vss 0.629612
R18234 vss.n12627 vss 0.629612
R18235 vss.n12763 vss 0.629612
R18236 vss vss.n13132 0.629612
R18237 vss.n13081 vss 0.629612
R18238 vss.n13032 vss 0.629612
R18239 vss vss.n13346 0.629612
R18240 vss vss.n8254 0.629612
R18241 vss.n13793 vss 0.629612
R18242 vss.n13744 vss 0.629612
R18243 vss vss.n13465 0.629612
R18244 vss vss.n13655 0.629612
R18245 vss.n13604 vss 0.629612
R18246 vss.n14138 vss 0.629612
R18247 vss vss.n14190 0.629612
R18248 vss vss.n10518 0.629612
R18249 vss vss.n10567 0.629612
R18250 vss vss.n10615 0.629612
R18251 vss.n10814 vss 0.629612
R18252 vss vss.n10912 0.629612
R18253 vss vss.n10961 0.629612
R18254 vss vss.n11009 0.629612
R18255 vss vss.n11302 0.629612
R18256 vss.n11251 vss 0.629612
R18257 vss.n11202 vss 0.629612
R18258 vss.n10027 vss 0.629612
R18259 vss vss.n11613 0.629612
R18260 vss.n11562 vss 0.629612
R18261 vss.n11708 vss 0.629612
R18262 vss.n11618 vss 0.629612
R18263 vss.n13184 vss 0.629612
R18264 vss.n10565 vss.n10564 0.616455
R18265 vss.n10959 vss.n10958 0.616455
R18266 vss.n11156 vss.n11155 0.616455
R18267 vss.n11711 vss.n11710 0.616455
R18268 vss.n12195 vss.n12194 0.616455
R18269 vss.n12313 vss.n12312 0.616455
R18270 vss.n12432 vss.n12431 0.616455
R18271 vss.n9470 vss.n9469 0.616455
R18272 vss.n6158 vss.n6157 0.616455
R18273 vss.n5919 vss.n5918 0.616455
R18274 vss.n3542 vss.n3541 0.616455
R18275 vss.n4540 vss.n4539 0.616455
R18276 vss.n5305 vss.n5304 0.616455
R18277 vss.n5093 vss.n5092 0.616455
R18278 vss.n6663 vss.n6662 0.616455
R18279 vss.n7447 vss.n7446 0.616455
R18280 vss.n7300 vss.n7299 0.616455
R18281 vss.n4606 vss.n4605 0.616455
R18282 vss.n6879 vss.n6878 0.616455
R18283 vss.n7765 vss.n7764 0.616455
R18284 vss.n7501 vss.n7500 0.616455
R18285 vss.n14882 vss.n14881 0.616455
R18286 vss.n13912 vss.n13911 0.616455
R18287 vss.n14029 vss.n14028 0.616455
R18288 vss.n2324 vss.n2323 0.616455
R18289 vss.n12625 vss.n12624 0.616455
R18290 vss.n9087 vss.n9086 0.616455
R18291 vss.n8301 vss.n8300 0.616455
R18292 vss.n14141 vss.n14140 0.616455
R18293 vss.n14357 vss.n14356 0.616455
R18294 vss.n15052 vss.n15051 0.616455
R18295 vss.n6211 vss.n6210 0.616455
R18296 vss.n9601 vss.n9600 0.616454
R18297 vss.n9731 vss.n9730 0.616454
R18298 vss.n9472 vss.n9471 0.616454
R18299 vss.n5045 vss.n4998 0.616454
R18300 vss.n5519 vss.n5472 0.616454
R18301 vss.n6377 vss.n6376 0.616454
R18302 vss.n4446 vss.n3273 0.616454
R18303 vss.n7350 vss.n7349 0.616454
R18304 vss.n15173 vss.n15172 0.616454
R18305 vss.n4654 vss.n4653 0.616454
R18306 vss.n7993 vss.n7992 0.616454
R18307 vss.n7717 vss.n7669 0.616454
R18308 vss.n7912 vss.n7864 0.616454
R18309 vss.n7206 vss.n3149 0.616454
R18310 vss.n8151 vss.n8150 0.616454
R18311 vss.n14478 vss.n14477 0.616454
R18312 vss.n8051 vss.n8050 0.616454
R18313 vss.n14089 vss.n14088 0.616454
R18314 vss.n13130 vss.n13129 0.616454
R18315 vss.n13842 vss.n13841 0.616454
R18316 vss.n13653 vss.n13652 0.616454
R18317 vss.n14282 vss.n14281 0.616454
R18318 vss.n14977 vss.n14976 0.616454
R18319 vss.n6063 vss.n6062 0.616454
R18320 vss.n5823 vss.n5822 0.616454
R18321 vss.n5680 vss.n5679 0.616454
R18322 vss.n15621 vss.n15620 0.616454
R18323 vss.n11802 vss.n11801 0.616454
R18324 vss.n10470 vss.n8879 0.616454
R18325 vss.n10864 vss.n10816 0.616454
R18326 vss.n11300 vss.n11299 0.616454
R18327 vss.n11611 vss.n11610 0.616454
R18328 vss.n8763 vss 0.606586
R18329 vss.n8644 vss 0.606586
R18330 vss.n9214 vss 0.606586
R18331 vss.n964 vss 0.606586
R18332 vss.n15341 vss 0.606586
R18333 vss.n552 vss 0.606586
R18334 vss.n1743 vss 0.606586
R18335 vss.n14646 vss 0.606586
R18336 vss.n1331 vss 0.606586
R18337 vss.n3856 vss 0.606586
R18338 vss.n3737 vss 0.606586
R18339 vss.n3618 vss 0.606586
R18340 vss.n9316 vss 0.588493
R18341 vss.n499 vss 0.588493
R18342 vss.n1278 vss 0.588493
R18343 vss vss.n15904 0.588493
R18344 vss.n11615 vss 0.431421
R18345 vss.n11304 vss 0.431421
R18346 vss vss.n10167 0.431421
R18347 vss.n6613 vss 0.431421
R18348 vss.n5423 vss 0.431421
R18349 vss.n4127 vss 0.431421
R18350 vss.n4949 vss 0.431421
R18351 vss vss.n4950 0.431421
R18352 vss.n5096 vss 0.431421
R18353 vss.n5212 vss 0.431421
R18354 vss vss.n5424 0.431421
R18355 vss.n5308 vss 0.431421
R18356 vss.n3387 vss 0.431421
R18357 vss.n6380 vss 0.431421
R18358 vss.n6495 vss 0.431421
R18359 vss vss.n6614 0.431421
R18360 vss vss.n4263 0.431421
R18361 vss vss.n4788 0.431421
R18362 vss.n14886 vss 0.431421
R18363 vss.n2837 vss 0.431421
R18364 vss vss.n2449 0.431421
R18365 vss.n7997 vss 0.431421
R18366 vss.n7996 vss 0.431421
R18367 vss.n7504 vss 0.431421
R18368 vss.n7620 vss 0.431421
R18369 vss vss.n7621 0.431421
R18370 vss.n7768 vss 0.431421
R18371 vss.n7815 vss 0.431421
R18372 vss vss.n7816 0.431421
R18373 vss vss.n1139 0.431421
R18374 vss.n14885 vss 0.431421
R18375 vss vss.n2448 0.431421
R18376 vss vss.n6791 0.431421
R18377 vss.n13657 vss 0.431421
R18378 vss.n13349 vss 0.431421
R18379 vss.n13134 vss 0.431421
R18380 vss.n12869 vss 0.431421
R18381 vss vss.n9391 0.431421
R18382 vss vss.n8951 0.431421
R18383 vss.n13133 vss 0.431421
R18384 vss vss.n8408 0.431421
R18385 vss.n13347 vss 0.431421
R18386 vss.n13348 vss 0.431421
R18387 vss.n13350 vss 0.431421
R18388 vss.n13466 vss 0.431421
R18389 vss.n13656 vss 0.431421
R18390 vss vss.n2033 0.431421
R18391 vss.n14191 vss 0.431421
R18392 vss.n10568 vss 0.431421
R18393 vss.n10617 vss 0.431421
R18394 vss.n10616 vss 0.431421
R18395 vss.n10962 vss 0.431421
R18396 vss.n11010 vss 0.431421
R18397 vss.n11303 vss 0.431421
R18398 vss vss.n10079 0.431421
R18399 vss vss.n9965 0.431421
R18400 vss.n11614 vss 0.431421
R18401 vss.n11616 vss 0.431421
R18402 vss vss.n11617 0.431421
R18403 vss vss.n10254 0.431421
R18404 vss vss.n12191 0.398526
R18405 vss vss.n8338 0.398526
R18406 vss.n13702 vss 0.398526
R18407 vss.n13701 vss 0.398526
R18408 vss vss.n8337 0.398526
R18409 vss.n13291 vss 0.398526
R18410 vss vss.n8617 0.398526
R18411 vss vss.n13290 0.398526
R18412 vss.n13290 vss 0.398526
R18413 vss vss.n12428 0.398526
R18414 vss vss.n8882 0.398526
R18415 vss.n13181 vss 0.398526
R18416 vss.n13180 vss 0.398526
R18417 vss.n13179 vss 0.398526
R18418 vss.n13178 vss 0.398526
R18419 vss vss.n163 0.398526
R18420 vss vss.n85 0.398526
R18421 vss vss.n27 0.398526
R18422 vss.n15222 vss 0.398526
R18423 vss vss.n759 0.398526
R18424 vss.n15221 vss 0.398526
R18425 vss.n15294 vss 0.398526
R18426 vss.n15342 vss 0.398526
R18427 vss.n15372 vss 0.398526
R18428 vss.n15371 vss 0.398526
R18429 vss.n15371 vss 0.398526
R18430 vss vss.n660 0.398526
R18431 vss vss.n501 0.398526
R18432 vss.n15447 vss 0.398526
R18433 vss.n15446 vss 0.398526
R18434 vss.n15445 vss 0.398526
R18435 vss.n15444 vss 0.398526
R18436 vss.n14527 vss 0.398526
R18437 vss vss.n1538 0.398526
R18438 vss.n14526 vss 0.398526
R18439 vss.n14599 vss 0.398526
R18440 vss.n14647 vss 0.398526
R18441 vss.n14677 vss 0.398526
R18442 vss.n14676 vss 0.398526
R18443 vss.n14676 vss 0.398526
R18444 vss vss.n1439 0.398526
R18445 vss vss.n1280 0.398526
R18446 vss.n14752 vss 0.398526
R18447 vss.n14751 vss 0.398526
R18448 vss.n14750 vss 0.398526
R18449 vss.n14749 vss 0.398526
R18450 vss vss.n1696 0.398526
R18451 vss.n14326 vss 0.398526
R18452 vss.n14325 vss 0.398526
R18453 vss vss.n917 0.398526
R18454 vss.n15021 vss 0.398526
R18455 vss.n15020 vss 0.398526
R18456 vss.n15870 vss 0.398526
R18457 vss vss.n84 0.398526
R18458 vss.n15815 vss 0.398526
R18459 vss.n15814 vss 0.398526
R18460 vss vss.n5869 0.398526
R18461 vss.n5869 vss 0.398526
R18462 vss.n15759 vss 0.398526
R18463 vss.n15758 vss 0.398526
R18464 vss vss.n241 0.398526
R18465 vss.n15703 vss 0.398526
R18466 vss.n15702 vss 0.398526
R18467 vss vss.n242 0.398526
R18468 vss vss.n15578 0.398526
R18469 vss.n12190 vss 0.398526
R18470 vss.n12189 vss 0.398526
R18471 vss.n15871 vss 0.398526
R18472 vss.n5424 vss 0.365632
R18473 vss.n7621 vss 0.365632
R18474 vss.n13348 vss 0.365632
R18475 vss.n11303 vss 0.365632
R18476 vss.n11652 vss.n9935 0.310177
R18477 vss.n11415 vss.n9964 0.310177
R18478 vss.n11305 vss.n10061 0.310177
R18479 vss.n10703 vss.n10641 0.310177
R18480 vss.n13674 vss.n13673 0.310177
R18481 vss.n13704 vss.n13703 0.310177
R18482 vss.n13293 vss.n13292 0.310177
R18483 vss.n12992 vss.n12991 0.310177
R18484 vss.n13151 vss.n13150 0.310177
R18485 vss.n12893 vss.n8880 0.310177
R18486 vss.n12816 vss.n8881 0.310177
R18487 vss.n15675 vss.n15674 0.310177
R18488 vss.n15872 vss.n19 0.310177
R18489 vss.n15732 vss.n15731 0.310177
R18490 vss.n15788 vss.n15787 0.310177
R18491 vss.n15844 vss.n15843 0.310177
R18492 vss.n15224 vss.n15223 0.310177
R18493 vss.n15267 vss.n15266 0.310177
R18494 vss.n15344 vss.n15343 0.310177
R18495 vss.n15374 vss.n15373 0.310177
R18496 vss.n15417 vss.n15416 0.310177
R18497 vss.n15449 vss.n15448 0.310177
R18498 vss.n4310 vss.n500 0.310177
R18499 vss.n14529 vss.n14528 0.310177
R18500 vss.n14572 vss.n14571 0.310177
R18501 vss.n14649 vss.n14648 0.310177
R18502 vss.n14679 vss.n14678 0.310177
R18503 vss.n14722 vss.n14721 0.310177
R18504 vss.n14754 vss.n14753 0.310177
R18505 vss.n8021 vss.n1279 0.310177
R18506 vss.n14328 vss.n14327 0.310177
R18507 vss.n15023 vss.n15022 0.310177
R18508 vss.n15817 vss.n15816 0.310177
R18509 vss.n15761 vss.n15760 0.310177
R18510 vss.n15705 vss.n15704 0.310177
R18511 vss.n12088 vss.n9859 0.310177
R18512 vss.n10618 vss.n10236 0.310177
R18513 vss.n11011 vss.n10149 0.310177
R18514 vss.n11331 vss.n9989 0.310177
R18515 vss.n10369 vss.n10278 0.310177
R18516 vss.n13182 vss 0.194579
R18517 vss.n6742 vss 0.194579
R18518 vss.n3272 vss 0.194579
R18519 vss.n3220 vss.n3217 0.1305
R18520 vss.n3220 vss.n3219 0.1305
R18521 vss.n3211 vss.n3186 0.1305
R18522 vss.n3227 vss.n3211 0.1305
R18523 vss.n3237 vss.n3185 0.1305
R18524 vss.n3259 vss.n3237 0.1305
R18525 vss.n3252 vss.n3243 0.1305
R18526 vss.n3252 vss.n3251 0.1305
R18527 vss.n3250 vss.n3239 0.1305
R18528 vss.n3251 vss.n3250 0.1305
R18529 vss.n3258 vss.n3257 0.1305
R18530 vss.n3259 vss.n3258 0.1305
R18531 vss.n3226 vss.n3225 0.1305
R18532 vss.n3227 vss.n3226 0.1305
R18533 vss.n3218 vss.n3213 0.1305
R18534 vss.n3219 vss.n3218 0.1305
R18535 vss.n6953 vss.n6950 0.1305
R18536 vss.n6953 vss.n6952 0.1305
R18537 vss.n6944 vss.n2447 0.1305
R18538 vss.n6960 vss.n6944 0.1305
R18539 vss.n2446 vss.n2445 0.1305
R18540 vss.n2445 vss.n2430 0.1305
R18541 vss.n2427 vss.n2422 0.1305
R18542 vss.n8017 vss.n2422 0.1305
R18543 vss.n8016 vss.n8015 0.1305
R18544 vss.n8017 vss.n8016 0.1305
R18545 vss.n2441 vss.n2426 0.1305
R18546 vss.n2441 vss.n2430 0.1305
R18547 vss.n6959 vss.n6958 0.1305
R18548 vss.n6960 vss.n6959 0.1305
R18549 vss.n6951 vss.n6946 0.1305
R18550 vss.n6952 vss.n6951 0.1305
R18551 vss.n1420 vss.n1419 0.1305
R18552 vss.n14693 vss.n1420 0.1305
R18553 vss.n1416 vss.n1409 0.1305
R18554 vss.n14697 vss.n1409 0.1305
R18555 vss.n1404 vss.n1386 0.1305
R18556 vss.n14711 vss.n1386 0.1305
R18557 vss.n1399 vss.n1391 0.1305
R18558 vss.n1399 vss.n1381 0.1305
R18559 vss.n1393 vss.n1392 0.1305
R18560 vss.n1392 vss.n1381 0.1305
R18561 vss.n14710 vss.n14709 0.1305
R18562 vss.n14711 vss.n14710 0.1305
R18563 vss.n14696 vss.n1390 0.1305
R18564 vss.n14697 vss.n14696 0.1305
R18565 vss.n14694 vss.n1412 0.1305
R18566 vss.n14694 vss.n14693 0.1305
R18567 vss.n7582 vss.n7579 0.1305
R18568 vss.n7582 vss.n7581 0.1305
R18569 vss.n7575 vss.n7526 0.1305
R18570 vss.n7589 vss.n7526 0.1305
R18571 vss.n7556 vss.n7555 0.1305
R18572 vss.n7555 vss.n7531 0.1305
R18573 vss.n7554 vss.n7553 0.1305
R18574 vss.n7553 vss.n7552 0.1305
R18575 vss.n7551 vss.n7550 0.1305
R18576 vss.n7552 vss.n7551 0.1305
R18577 vss.n7541 vss.n7529 0.1305
R18578 vss.n7541 vss.n7531 0.1305
R18579 vss.n7588 vss.n7587 0.1305
R18580 vss.n7589 vss.n7588 0.1305
R18581 vss.n7580 vss.n7574 0.1305
R18582 vss.n7581 vss.n7580 0.1305
R18583 vss.n2800 vss.n2797 0.1305
R18584 vss.n2800 vss.n2799 0.1305
R18585 vss.n2793 vss.n2744 0.1305
R18586 vss.n2807 vss.n2744 0.1305
R18587 vss.n2774 vss.n2773 0.1305
R18588 vss.n2773 vss.n2749 0.1305
R18589 vss.n2772 vss.n2771 0.1305
R18590 vss.n2771 vss.n2770 0.1305
R18591 vss.n2769 vss.n2768 0.1305
R18592 vss.n2770 vss.n2769 0.1305
R18593 vss.n2759 vss.n2747 0.1305
R18594 vss.n2759 vss.n2749 0.1305
R18595 vss.n2806 vss.n2805 0.1305
R18596 vss.n2807 vss.n2806 0.1305
R18597 vss.n2798 vss.n2792 0.1305
R18598 vss.n2799 vss.n2798 0.1305
R18599 vss.n1677 vss.n1676 0.1305
R18600 vss.n14543 vss.n1677 0.1305
R18601 vss.n1673 vss.n1666 0.1305
R18602 vss.n14547 vss.n1666 0.1305
R18603 vss.n1661 vss.n1643 0.1305
R18604 vss.n14561 vss.n1643 0.1305
R18605 vss.n1656 vss.n1648 0.1305
R18606 vss.n1656 vss.n1638 0.1305
R18607 vss.n1650 vss.n1649 0.1305
R18608 vss.n1649 vss.n1638 0.1305
R18609 vss.n14560 vss.n14559 0.1305
R18610 vss.n14561 vss.n14560 0.1305
R18611 vss.n14546 vss.n1647 0.1305
R18612 vss.n14547 vss.n14546 0.1305
R18613 vss.n14544 vss.n1669 0.1305
R18614 vss.n14544 vss.n14543 0.1305
R18615 vss.n2565 vss.n2562 0.1305
R18616 vss.n2565 vss.n2564 0.1305
R18617 vss.n2558 vss.n2508 0.1305
R18618 vss.n2572 vss.n2508 0.1305
R18619 vss.n2526 vss.n2513 0.1305
R18620 vss.n2526 vss.n2515 0.1305
R18621 vss.n2540 vss.n2539 0.1305
R18622 vss.n2539 vss.n2538 0.1305
R18623 vss.n2537 vss.n2536 0.1305
R18624 vss.n2538 vss.n2537 0.1305
R18625 vss.n2529 vss.n2528 0.1305
R18626 vss.n2528 vss.n2515 0.1305
R18627 vss.n2571 vss.n2570 0.1305
R18628 vss.n2572 vss.n2571 0.1305
R18629 vss.n2563 vss.n2512 0.1305
R18630 vss.n2564 vss.n2563 0.1305
R18631 vss.n1957 vss.n1956 0.1305
R18632 vss.n1959 vss.n1957 0.1305
R18633 vss.n1953 vss.n1946 0.1305
R18634 vss.n1963 vss.n1946 0.1305
R18635 vss.n1881 vss.n1877 0.1305
R18636 vss.n1977 vss.n1877 0.1305
R18637 vss.n1890 vss.n1889 0.1305
R18638 vss.n1890 vss.n1872 0.1305
R18639 vss.n1883 vss.n1880 0.1305
R18640 vss.n1883 vss.n1872 0.1305
R18641 vss.n1976 vss.n1975 0.1305
R18642 vss.n1977 vss.n1976 0.1305
R18643 vss.n1962 vss.n1895 0.1305
R18644 vss.n1963 vss.n1962 0.1305
R18645 vss.n1960 vss.n1949 0.1305
R18646 vss.n1960 vss.n1959 0.1305
R18647 vss.n1966 vss.n1875 0.1305
R18648 vss.n1966 vss.n1876 0.1305
R18649 vss.n1983 vss.n1982 0.1305
R18650 vss.n1984 vss.n1983 0.1305
R18651 vss.n14333 vss.n14332 0.1305
R18652 vss.n14332 vss.n14331 0.1305
R18653 vss.n14335 vss.n1857 0.1305
R18654 vss.n1857 vss.n1855 0.1305
R18655 vss.n1967 vss.n1965 0.1305
R18656 vss.n1965 vss.n1876 0.1305
R18657 vss.n1986 vss.n1985 0.1305
R18658 vss.n1985 vss.n1984 0.1305
R18659 vss.n14330 vss.n14329 0.1305
R18660 vss.n14331 vss.n14330 0.1305
R18661 vss.n1858 vss.n1856 0.1305
R18662 vss.n1856 vss.n1855 0.1305
R18663 vss.n2549 vss.n2516 0.1305
R18664 vss.n2553 vss.n2516 0.1305
R18665 vss.n2522 vss.n2520 0.1305
R18666 vss.n2524 vss.n2522 0.1305
R18667 vss.n14534 vss.n14533 0.1305
R18668 vss.n14533 vss.n14532 0.1305
R18669 vss.n14536 vss.n1682 0.1305
R18670 vss.n1682 vss.n1680 0.1305
R18671 vss.n2552 vss.n2551 0.1305
R18672 vss.n2553 vss.n2552 0.1305
R18673 vss.n2523 vss.n1695 0.1305
R18674 vss.n2524 vss.n2523 0.1305
R18675 vss.n14531 vss.n14530 0.1305
R18676 vss.n14532 vss.n14531 0.1305
R18677 vss.n1683 vss.n1681 0.1305
R18678 vss.n1681 vss.n1680 0.1305
R18679 vss.n14550 vss.n1641 0.1305
R18680 vss.n14550 vss.n1642 0.1305
R18681 vss.n14567 vss.n14566 0.1305
R18682 vss.n14568 vss.n14567 0.1305
R18683 vss.n14577 vss.n14576 0.1305
R18684 vss.n14576 vss.n14575 0.1305
R18685 vss.n14579 vss.n1577 0.1305
R18686 vss.n1577 vss.n1575 0.1305
R18687 vss.n14551 vss.n14549 0.1305
R18688 vss.n14549 vss.n1642 0.1305
R18689 vss.n14570 vss.n14569 0.1305
R18690 vss.n14569 vss.n14568 0.1305
R18691 vss.n14574 vss.n14573 0.1305
R18692 vss.n14575 vss.n14574 0.1305
R18693 vss.n1578 vss.n1576 0.1305
R18694 vss.n1576 vss.n1575 0.1305
R18695 vss.n2783 vss.n2750 0.1305
R18696 vss.n2787 vss.n2750 0.1305
R18697 vss.n2756 vss.n2754 0.1305
R18698 vss.n2758 vss.n2756 0.1305
R18699 vss.n14654 vss.n14653 0.1305
R18700 vss.n14653 vss.n14652 0.1305
R18701 vss.n14656 vss.n1524 0.1305
R18702 vss.n1524 vss.n1522 0.1305
R18703 vss.n2786 vss.n2785 0.1305
R18704 vss.n2787 vss.n2786 0.1305
R18705 vss.n2757 vss.n1537 0.1305
R18706 vss.n2758 vss.n2757 0.1305
R18707 vss.n14651 vss.n14650 0.1305
R18708 vss.n14652 vss.n14651 0.1305
R18709 vss.n1525 vss.n1523 0.1305
R18710 vss.n1523 vss.n1522 0.1305
R18711 vss.n7565 vss.n7532 0.1305
R18712 vss.n7569 vss.n7532 0.1305
R18713 vss.n7538 vss.n7536 0.1305
R18714 vss.n7540 vss.n7538 0.1305
R18715 vss.n14684 vss.n14683 0.1305
R18716 vss.n14683 vss.n14682 0.1305
R18717 vss.n14686 vss.n1425 0.1305
R18718 vss.n1425 vss.n1423 0.1305
R18719 vss.n7568 vss.n7567 0.1305
R18720 vss.n7569 vss.n7568 0.1305
R18721 vss.n7539 vss.n1438 0.1305
R18722 vss.n7540 vss.n7539 0.1305
R18723 vss.n14681 vss.n14680 0.1305
R18724 vss.n14682 vss.n14681 0.1305
R18725 vss.n1426 vss.n1424 0.1305
R18726 vss.n1424 vss.n1423 0.1305
R18727 vss.n14700 vss.n1384 0.1305
R18728 vss.n14700 vss.n1385 0.1305
R18729 vss.n14717 vss.n14716 0.1305
R18730 vss.n14718 vss.n14717 0.1305
R18731 vss.n14727 vss.n14726 0.1305
R18732 vss.n14726 vss.n14725 0.1305
R18733 vss.n14729 vss.n1319 0.1305
R18734 vss.n1319 vss.n1317 0.1305
R18735 vss.n14701 vss.n14699 0.1305
R18736 vss.n14699 vss.n1385 0.1305
R18737 vss.n14720 vss.n14719 0.1305
R18738 vss.n14719 vss.n14718 0.1305
R18739 vss.n14724 vss.n14723 0.1305
R18740 vss.n14725 vss.n14724 0.1305
R18741 vss.n1320 vss.n1318 0.1305
R18742 vss.n1318 vss.n1317 0.1305
R18743 vss.n8006 vss.n8005 0.1305
R18744 vss.n8005 vss.n8004 0.1305
R18745 vss.n2437 vss.n2436 0.1305
R18746 vss.n2436 vss.n2421 0.1305
R18747 vss.n8026 vss.n8025 0.1305
R18748 vss.n8025 vss.n8024 0.1305
R18749 vss.n8028 vss.n2362 0.1305
R18750 vss.n2362 vss.n2360 0.1305
R18751 vss.n8003 vss.n8002 0.1305
R18752 vss.n8004 vss.n8003 0.1305
R18753 vss.n2434 vss.n2433 0.1305
R18754 vss.n2433 vss.n2421 0.1305
R18755 vss.n8023 vss.n8022 0.1305
R18756 vss.n8024 vss.n8023 0.1305
R18757 vss.n2363 vss.n2361 0.1305
R18758 vss.n2361 vss.n2360 0.1305
R18759 vss.n3264 vss.n3230 0.1305
R18760 vss.n3230 vss.n3190 0.1305
R18761 vss.n3247 vss.n3232 0.1305
R18762 vss.n3249 vss.n3247 0.1305
R18763 vss.n14759 vss.n14758 0.1305
R18764 vss.n14758 vss.n14757 0.1305
R18765 vss.n14761 vss.n1218 0.1305
R18766 vss.n1218 vss.n1216 0.1305
R18767 vss.n3231 vss.n3229 0.1305
R18768 vss.n3229 vss.n3190 0.1305
R18769 vss.n3248 vss.n1231 0.1305
R18770 vss.n3249 vss.n3248 0.1305
R18771 vss.n14756 vss.n14755 0.1305
R18772 vss.n14757 vss.n14756 0.1305
R18773 vss.n1219 vss.n1217 0.1305
R18774 vss.n1217 vss.n1216 0.1305
R18775 vss.n4857 vss.n4747 0.1305
R18776 vss.n4747 vss.n4745 0.1305
R18777 vss.n4855 vss.n4854 0.1305
R18778 vss.n4854 vss.n4853 0.1305
R18779 vss.n4831 vss.n4815 0.1305
R18780 vss.n4837 vss.n4815 0.1305
R18781 vss.n4830 vss.n4829 0.1305
R18782 vss.n4829 vss.n4828 0.1305
R18783 vss.n4819 vss.n4816 0.1305
R18784 vss.n4828 vss.n4816 0.1305
R18785 vss.n4836 vss.n4805 0.1305
R18786 vss.n4837 vss.n4836 0.1305
R18787 vss.n4852 vss.n4851 0.1305
R18788 vss.n4853 vss.n4852 0.1305
R18789 vss.n4748 vss.n4746 0.1305
R18790 vss.n4746 vss.n4745 0.1305
R18791 vss.n4911 vss.n4908 0.1305
R18792 vss.n4911 vss.n4910 0.1305
R18793 vss.n4904 vss.n4285 0.1305
R18794 vss.n4918 vss.n4285 0.1305
R18795 vss.n4885 vss.n4884 0.1305
R18796 vss.n4884 vss.n4290 0.1305
R18797 vss.n4883 vss.n4882 0.1305
R18798 vss.n4882 vss.n4881 0.1305
R18799 vss.n4880 vss.n4879 0.1305
R18800 vss.n4881 vss.n4880 0.1305
R18801 vss.n4298 vss.n4288 0.1305
R18802 vss.n4298 vss.n4290 0.1305
R18803 vss.n4917 vss.n4916 0.1305
R18804 vss.n4918 vss.n4917 0.1305
R18805 vss.n4909 vss.n4903 0.1305
R18806 vss.n4910 vss.n4909 0.1305
R18807 vss.n641 vss.n640 0.1305
R18808 vss.n15388 vss.n641 0.1305
R18809 vss.n637 vss.n630 0.1305
R18810 vss.n15392 vss.n630 0.1305
R18811 vss.n625 vss.n607 0.1305
R18812 vss.n15406 vss.n607 0.1305
R18813 vss.n620 vss.n612 0.1305
R18814 vss.n620 vss.n602 0.1305
R18815 vss.n614 vss.n613 0.1305
R18816 vss.n613 vss.n602 0.1305
R18817 vss.n15405 vss.n15404 0.1305
R18818 vss.n15406 vss.n15405 0.1305
R18819 vss.n15391 vss.n611 0.1305
R18820 vss.n15392 vss.n15391 0.1305
R18821 vss.n15389 vss.n633 0.1305
R18822 vss.n15389 vss.n15388 0.1305
R18823 vss.n5174 vss.n5171 0.1305
R18824 vss.n5174 vss.n5173 0.1305
R18825 vss.n5167 vss.n5118 0.1305
R18826 vss.n5181 vss.n5118 0.1305
R18827 vss.n5148 vss.n5147 0.1305
R18828 vss.n5147 vss.n5123 0.1305
R18829 vss.n5146 vss.n5145 0.1305
R18830 vss.n5145 vss.n5144 0.1305
R18831 vss.n5143 vss.n5142 0.1305
R18832 vss.n5144 vss.n5143 0.1305
R18833 vss.n5133 vss.n5121 0.1305
R18834 vss.n5133 vss.n5123 0.1305
R18835 vss.n5180 vss.n5179 0.1305
R18836 vss.n5181 vss.n5180 0.1305
R18837 vss.n5172 vss.n5166 0.1305
R18838 vss.n5173 vss.n5172 0.1305
R18839 vss.n5386 vss.n5383 0.1305
R18840 vss.n5386 vss.n5385 0.1305
R18841 vss.n5379 vss.n5330 0.1305
R18842 vss.n5393 vss.n5330 0.1305
R18843 vss.n5360 vss.n5359 0.1305
R18844 vss.n5359 vss.n5335 0.1305
R18845 vss.n5358 vss.n5357 0.1305
R18846 vss.n5357 vss.n5356 0.1305
R18847 vss.n5355 vss.n5354 0.1305
R18848 vss.n5356 vss.n5355 0.1305
R18849 vss.n5345 vss.n5333 0.1305
R18850 vss.n5345 vss.n5335 0.1305
R18851 vss.n5392 vss.n5391 0.1305
R18852 vss.n5393 vss.n5392 0.1305
R18853 vss.n5384 vss.n5378 0.1305
R18854 vss.n5385 vss.n5384 0.1305
R18855 vss.n898 vss.n897 0.1305
R18856 vss.n15238 vss.n898 0.1305
R18857 vss.n894 vss.n887 0.1305
R18858 vss.n15242 vss.n887 0.1305
R18859 vss.n882 vss.n864 0.1305
R18860 vss.n15256 vss.n864 0.1305
R18861 vss.n877 vss.n869 0.1305
R18862 vss.n877 vss.n859 0.1305
R18863 vss.n871 vss.n870 0.1305
R18864 vss.n870 vss.n859 0.1305
R18865 vss.n15255 vss.n15254 0.1305
R18866 vss.n15256 vss.n15255 0.1305
R18867 vss.n15241 vss.n868 0.1305
R18868 vss.n15242 vss.n15241 0.1305
R18869 vss.n15239 vss.n890 0.1305
R18870 vss.n15239 vss.n15238 0.1305
R18871 vss.n6458 vss.n6455 0.1305
R18872 vss.n6458 vss.n6457 0.1305
R18873 vss.n6451 vss.n6402 0.1305
R18874 vss.n6465 vss.n6402 0.1305
R18875 vss.n6432 vss.n6431 0.1305
R18876 vss.n6431 vss.n6407 0.1305
R18877 vss.n6430 vss.n6429 0.1305
R18878 vss.n6429 vss.n6428 0.1305
R18879 vss.n6427 vss.n6426 0.1305
R18880 vss.n6428 vss.n6427 0.1305
R18881 vss.n6417 vss.n6405 0.1305
R18882 vss.n6417 vss.n6407 0.1305
R18883 vss.n6464 vss.n6463 0.1305
R18884 vss.n6465 vss.n6464 0.1305
R18885 vss.n6456 vss.n6450 0.1305
R18886 vss.n6457 vss.n6456 0.1305
R18887 vss.n6574 vss.n6570 0.1305
R18888 vss.n6574 vss.n6573 0.1305
R18889 vss.n6566 vss.n6517 0.1305
R18890 vss.n6581 vss.n6517 0.1305
R18891 vss.n6547 vss.n6546 0.1305
R18892 vss.n6546 vss.n6522 0.1305
R18893 vss.n6545 vss.n6544 0.1305
R18894 vss.n6544 vss.n6543 0.1305
R18895 vss.n6542 vss.n6541 0.1305
R18896 vss.n6543 vss.n6542 0.1305
R18897 vss.n6532 vss.n6520 0.1305
R18898 vss.n6532 vss.n6522 0.1305
R18899 vss.n6580 vss.n6579 0.1305
R18900 vss.n6581 vss.n6580 0.1305
R18901 vss.n6572 vss.n6565 0.1305
R18902 vss.n6573 vss.n6572 0.1305
R18903 vss.n6556 vss.n6523 0.1305
R18904 vss.n6560 vss.n6523 0.1305
R18905 vss.n6529 vss.n6527 0.1305
R18906 vss.n6531 vss.n6529 0.1305
R18907 vss.n15028 vss.n15027 0.1305
R18908 vss.n15027 vss.n15026 0.1305
R18909 vss.n15030 vss.n1078 0.1305
R18910 vss.n1078 vss.n1076 0.1305
R18911 vss.n6559 vss.n6558 0.1305
R18912 vss.n6560 vss.n6559 0.1305
R18913 vss.n6530 vss.n1091 0.1305
R18914 vss.n6531 vss.n6530 0.1305
R18915 vss.n15025 vss.n15024 0.1305
R18916 vss.n15026 vss.n15025 0.1305
R18917 vss.n1079 vss.n1077 0.1305
R18918 vss.n1077 vss.n1076 0.1305
R18919 vss.n6441 vss.n6408 0.1305
R18920 vss.n6445 vss.n6408 0.1305
R18921 vss.n6414 vss.n6412 0.1305
R18922 vss.n6416 vss.n6414 0.1305
R18923 vss.n15229 vss.n15228 0.1305
R18924 vss.n15228 vss.n15227 0.1305
R18925 vss.n15231 vss.n903 0.1305
R18926 vss.n903 vss.n901 0.1305
R18927 vss.n6444 vss.n6443 0.1305
R18928 vss.n6445 vss.n6444 0.1305
R18929 vss.n6415 vss.n916 0.1305
R18930 vss.n6416 vss.n6415 0.1305
R18931 vss.n15226 vss.n15225 0.1305
R18932 vss.n15227 vss.n15226 0.1305
R18933 vss.n904 vss.n902 0.1305
R18934 vss.n902 vss.n901 0.1305
R18935 vss.n15245 vss.n862 0.1305
R18936 vss.n15245 vss.n863 0.1305
R18937 vss.n15262 vss.n15261 0.1305
R18938 vss.n15263 vss.n15262 0.1305
R18939 vss.n15272 vss.n15271 0.1305
R18940 vss.n15271 vss.n15270 0.1305
R18941 vss.n15274 vss.n798 0.1305
R18942 vss.n798 vss.n796 0.1305
R18943 vss.n15246 vss.n15244 0.1305
R18944 vss.n15244 vss.n863 0.1305
R18945 vss.n15265 vss.n15264 0.1305
R18946 vss.n15264 vss.n15263 0.1305
R18947 vss.n15269 vss.n15268 0.1305
R18948 vss.n15270 vss.n15269 0.1305
R18949 vss.n799 vss.n797 0.1305
R18950 vss.n797 vss.n796 0.1305
R18951 vss.n5369 vss.n5336 0.1305
R18952 vss.n5373 vss.n5336 0.1305
R18953 vss.n5342 vss.n5340 0.1305
R18954 vss.n5344 vss.n5342 0.1305
R18955 vss.n15349 vss.n15348 0.1305
R18956 vss.n15348 vss.n15347 0.1305
R18957 vss.n15351 vss.n745 0.1305
R18958 vss.n745 vss.n743 0.1305
R18959 vss.n5372 vss.n5371 0.1305
R18960 vss.n5373 vss.n5372 0.1305
R18961 vss.n5343 vss.n758 0.1305
R18962 vss.n5344 vss.n5343 0.1305
R18963 vss.n15346 vss.n15345 0.1305
R18964 vss.n15347 vss.n15346 0.1305
R18965 vss.n746 vss.n744 0.1305
R18966 vss.n744 vss.n743 0.1305
R18967 vss.n5157 vss.n5124 0.1305
R18968 vss.n5161 vss.n5124 0.1305
R18969 vss.n5130 vss.n5128 0.1305
R18970 vss.n5132 vss.n5130 0.1305
R18971 vss.n15379 vss.n15378 0.1305
R18972 vss.n15378 vss.n15377 0.1305
R18973 vss.n15381 vss.n646 0.1305
R18974 vss.n646 vss.n644 0.1305
R18975 vss.n5160 vss.n5159 0.1305
R18976 vss.n5161 vss.n5160 0.1305
R18977 vss.n5131 vss.n659 0.1305
R18978 vss.n5132 vss.n5131 0.1305
R18979 vss.n15376 vss.n15375 0.1305
R18980 vss.n15377 vss.n15376 0.1305
R18981 vss.n647 vss.n645 0.1305
R18982 vss.n645 vss.n644 0.1305
R18983 vss.n15395 vss.n605 0.1305
R18984 vss.n15395 vss.n606 0.1305
R18985 vss.n15412 vss.n15411 0.1305
R18986 vss.n15413 vss.n15412 0.1305
R18987 vss.n15422 vss.n15421 0.1305
R18988 vss.n15421 vss.n15420 0.1305
R18989 vss.n15424 vss.n540 0.1305
R18990 vss.n540 vss.n538 0.1305
R18991 vss.n15396 vss.n15394 0.1305
R18992 vss.n15394 vss.n606 0.1305
R18993 vss.n15415 vss.n15414 0.1305
R18994 vss.n15414 vss.n15413 0.1305
R18995 vss.n15419 vss.n15418 0.1305
R18996 vss.n15420 vss.n15419 0.1305
R18997 vss.n541 vss.n539 0.1305
R18998 vss.n539 vss.n538 0.1305
R18999 vss.n4894 vss.n4291 0.1305
R19000 vss.n4898 vss.n4291 0.1305
R19001 vss.n4308 vss.n4295 0.1305
R19002 vss.n4308 vss.n4297 0.1305
R19003 vss.n4874 vss.n4873 0.1305
R19004 vss.n4873 vss.n4872 0.1305
R19005 vss.n4865 vss.n4864 0.1305
R19006 vss.n4866 vss.n4865 0.1305
R19007 vss.n4897 vss.n4896 0.1305
R19008 vss.n4898 vss.n4897 0.1305
R19009 vss.n4306 vss.n4305 0.1305
R19010 vss.n4306 vss.n4297 0.1305
R19011 vss.n4871 vss.n4870 0.1305
R19012 vss.n4872 vss.n4871 0.1305
R19013 vss.n4868 vss.n4867 0.1305
R19014 vss.n4867 vss.n4866 0.1305
R19015 vss.n4842 vss.n4808 0.1305
R19016 vss.n4808 vss.n4806 0.1305
R19017 vss.n4825 vss.n4810 0.1305
R19018 vss.n4827 vss.n4825 0.1305
R19019 vss.n15454 vss.n15453 0.1305
R19020 vss.n15453 vss.n15452 0.1305
R19021 vss.n15456 vss.n439 0.1305
R19022 vss.n439 vss.n437 0.1305
R19023 vss.n4809 vss.n4807 0.1305
R19024 vss.n4807 vss.n4806 0.1305
R19025 vss.n4826 vss.n452 0.1305
R19026 vss.n4827 vss.n4826 0.1305
R19027 vss.n15451 vss.n15450 0.1305
R19028 vss.n15452 vss.n15451 0.1305
R19029 vss.n440 vss.n438 0.1305
R19030 vss.n438 vss.n437 0.1305
R19031 vss.n15876 vss.n22 0.1305
R19032 vss.n15880 vss.n22 0.1305
R19033 vss.n15885 vss.n15884 0.1305
R19034 vss.n15884 vss.n16 0.1305
R19035 vss.n6261 vss.n20 0.1305
R19036 vss.n6261 vss.n15 0.1305
R19037 vss.n6267 vss.n6255 0.1305
R19038 vss.n6255 vss.n6253 0.1305
R19039 vss.n15879 vss.n15878 0.1305
R19040 vss.n15880 vss.n15879 0.1305
R19041 vss.n15874 vss.n15873 0.1305
R19042 vss.n15873 vss.n16 0.1305
R19043 vss.n6259 vss.n6258 0.1305
R19044 vss.n6259 vss.n15 0.1305
R19045 vss.n6256 vss.n6254 0.1305
R19046 vss.n6254 vss.n6253 0.1305
R19047 vss.n15834 vss.n15833 0.1305
R19048 vss.n15833 vss.n15832 0.1305
R19049 vss.n15839 vss.n15838 0.1305
R19050 vss.n15840 vss.n15839 0.1305
R19051 vss.n15849 vss.n15848 0.1305
R19052 vss.n15848 vss.n15847 0.1305
R19053 vss.n15851 vss.n46 0.1305
R19054 vss.n46 vss.n44 0.1305
R19055 vss.n15831 vss.n15830 0.1305
R19056 vss.n15832 vss.n15831 0.1305
R19057 vss.n15842 vss.n15841 0.1305
R19058 vss.n15841 vss.n15840 0.1305
R19059 vss.n15846 vss.n15845 0.1305
R19060 vss.n15847 vss.n15846 0.1305
R19061 vss.n47 vss.n45 0.1305
R19062 vss.n45 vss.n44 0.1305
R19063 vss.n119 vss.n104 0.1305
R19064 vss.n104 vss.n102 0.1305
R19065 vss.n112 vss.n106 0.1305
R19066 vss.n114 vss.n112 0.1305
R19067 vss.n15822 vss.n15821 0.1305
R19068 vss.n15821 vss.n15820 0.1305
R19069 vss.n15824 vss.n70 0.1305
R19070 vss.n70 vss.n68 0.1305
R19071 vss.n105 vss.n103 0.1305
R19072 vss.n103 vss.n102 0.1305
R19073 vss.n113 vss.n83 0.1305
R19074 vss.n114 vss.n113 0.1305
R19075 vss.n15819 vss.n15818 0.1305
R19076 vss.n15820 vss.n15819 0.1305
R19077 vss.n71 vss.n69 0.1305
R19078 vss.n69 vss.n68 0.1305
R19079 vss.n15778 vss.n15777 0.1305
R19080 vss.n15777 vss.n15776 0.1305
R19081 vss.n15783 vss.n15782 0.1305
R19082 vss.n15784 vss.n15783 0.1305
R19083 vss.n15793 vss.n15792 0.1305
R19084 vss.n15792 vss.n15791 0.1305
R19085 vss.n15795 vss.n125 0.1305
R19086 vss.n125 vss.n123 0.1305
R19087 vss.n15775 vss.n15774 0.1305
R19088 vss.n15776 vss.n15775 0.1305
R19089 vss.n15786 vss.n15785 0.1305
R19090 vss.n15785 vss.n15784 0.1305
R19091 vss.n15790 vss.n15789 0.1305
R19092 vss.n15791 vss.n15790 0.1305
R19093 vss.n126 vss.n124 0.1305
R19094 vss.n124 vss.n123 0.1305
R19095 vss.n197 vss.n182 0.1305
R19096 vss.n182 vss.n180 0.1305
R19097 vss.n190 vss.n184 0.1305
R19098 vss.n192 vss.n190 0.1305
R19099 vss.n15766 vss.n15765 0.1305
R19100 vss.n15765 vss.n15764 0.1305
R19101 vss.n15768 vss.n149 0.1305
R19102 vss.n149 vss.n147 0.1305
R19103 vss.n183 vss.n181 0.1305
R19104 vss.n181 vss.n180 0.1305
R19105 vss.n191 vss.n162 0.1305
R19106 vss.n192 vss.n191 0.1305
R19107 vss.n15763 vss.n15762 0.1305
R19108 vss.n15764 vss.n15763 0.1305
R19109 vss.n150 vss.n148 0.1305
R19110 vss.n148 vss.n147 0.1305
R19111 vss.n15722 vss.n15721 0.1305
R19112 vss.n15721 vss.n15720 0.1305
R19113 vss.n15727 vss.n15726 0.1305
R19114 vss.n15728 vss.n15727 0.1305
R19115 vss.n15737 vss.n15736 0.1305
R19116 vss.n15736 vss.n15735 0.1305
R19117 vss.n15739 vss.n203 0.1305
R19118 vss.n203 vss.n201 0.1305
R19119 vss.n15719 vss.n15718 0.1305
R19120 vss.n15720 vss.n15719 0.1305
R19121 vss.n15730 vss.n15729 0.1305
R19122 vss.n15729 vss.n15728 0.1305
R19123 vss.n15734 vss.n15733 0.1305
R19124 vss.n15735 vss.n15734 0.1305
R19125 vss.n204 vss.n202 0.1305
R19126 vss.n202 vss.n201 0.1305
R19127 vss.n276 vss.n261 0.1305
R19128 vss.n261 vss.n259 0.1305
R19129 vss.n269 vss.n263 0.1305
R19130 vss.n271 vss.n269 0.1305
R19131 vss.n15710 vss.n15709 0.1305
R19132 vss.n15709 vss.n15708 0.1305
R19133 vss.n15712 vss.n227 0.1305
R19134 vss.n227 vss.n225 0.1305
R19135 vss.n262 vss.n260 0.1305
R19136 vss.n260 vss.n259 0.1305
R19137 vss.n270 vss.n240 0.1305
R19138 vss.n271 vss.n270 0.1305
R19139 vss.n15707 vss.n15706 0.1305
R19140 vss.n15708 vss.n15707 0.1305
R19141 vss.n228 vss.n226 0.1305
R19142 vss.n226 vss.n225 0.1305
R19143 vss.n15665 vss.n15664 0.1305
R19144 vss.n15664 vss.n15663 0.1305
R19145 vss.n15670 vss.n15669 0.1305
R19146 vss.n15671 vss.n15670 0.1305
R19147 vss.n289 vss.n284 0.1305
R19148 vss.n15678 vss.n289 0.1305
R19149 vss.n15683 vss.n282 0.1305
R19150 vss.n282 vss.n280 0.1305
R19151 vss.n15662 vss.n15661 0.1305
R19152 vss.n15663 vss.n15662 0.1305
R19153 vss.n15673 vss.n15672 0.1305
R19154 vss.n15672 vss.n15671 0.1305
R19155 vss.n15677 vss.n15676 0.1305
R19156 vss.n15678 vss.n15677 0.1305
R19157 vss.n283 vss.n281 0.1305
R19158 vss.n281 vss.n280 0.1305
R19159 vss.n13666 vss.n13665 0.1305
R19160 vss.n13665 vss.n13664 0.1305
R19161 vss.n13669 vss.n13668 0.1305
R19162 vss.n13670 vss.n13669 0.1305
R19163 vss.n13679 vss.n13678 0.1305
R19164 vss.n13678 vss.n13677 0.1305
R19165 vss.n13681 vss.n8359 0.1305
R19166 vss.n8359 vss.n8357 0.1305
R19167 vss.n13663 vss.n13662 0.1305
R19168 vss.n13664 vss.n13663 0.1305
R19169 vss.n13672 vss.n13671 0.1305
R19170 vss.n13671 vss.n13670 0.1305
R19171 vss.n13676 vss.n13675 0.1305
R19172 vss.n13677 vss.n13676 0.1305
R19173 vss.n8360 vss.n8358 0.1305
R19174 vss.n8358 vss.n8357 0.1305
R19175 vss.n13411 vss.n13378 0.1305
R19176 vss.n13415 vss.n13378 0.1305
R19177 vss.n13409 vss.n13408 0.1305
R19178 vss.n13408 vss.n13407 0.1305
R19179 vss.n13709 vss.n13708 0.1305
R19180 vss.n13708 vss.n13707 0.1305
R19181 vss.n13711 vss.n8323 0.1305
R19182 vss.n8323 vss.n8321 0.1305
R19183 vss.n13414 vss.n13413 0.1305
R19184 vss.n13415 vss.n13414 0.1305
R19185 vss.n13406 vss.n8336 0.1305
R19186 vss.n13407 vss.n13406 0.1305
R19187 vss.n13706 vss.n13705 0.1305
R19188 vss.n13707 vss.n13706 0.1305
R19189 vss.n8324 vss.n8322 0.1305
R19190 vss.n8322 vss.n8321 0.1305
R19191 vss.n8610 vss.n8609 0.1305
R19192 vss.n8609 vss.n8608 0.1305
R19193 vss.n8613 vss.n8612 0.1305
R19194 vss.n8614 vss.n8613 0.1305
R19195 vss.n13298 vss.n13297 0.1305
R19196 vss.n13297 vss.n13296 0.1305
R19197 vss.n13300 vss.n8489 0.1305
R19198 vss.n8489 vss.n8487 0.1305
R19199 vss.n8607 vss.n8606 0.1305
R19200 vss.n8608 vss.n8607 0.1305
R19201 vss.n8616 vss.n8615 0.1305
R19202 vss.n8615 vss.n8614 0.1305
R19203 vss.n13295 vss.n13294 0.1305
R19204 vss.n13296 vss.n13295 0.1305
R19205 vss.n8490 vss.n8488 0.1305
R19206 vss.n8488 vss.n8487 0.1305
R19207 vss.n12984 vss.n12983 0.1305
R19208 vss.n12983 vss.n12982 0.1305
R19209 vss.n12987 vss.n12986 0.1305
R19210 vss.n12988 vss.n12987 0.1305
R19211 vss.n12997 vss.n12996 0.1305
R19212 vss.n12996 vss.n12995 0.1305
R19213 vss.n12999 vss.n9175 0.1305
R19214 vss.n9175 vss.n9173 0.1305
R19215 vss.n12981 vss.n12980 0.1305
R19216 vss.n12982 vss.n12981 0.1305
R19217 vss.n12990 vss.n12989 0.1305
R19218 vss.n12989 vss.n12988 0.1305
R19219 vss.n12994 vss.n12993 0.1305
R19220 vss.n12995 vss.n12994 0.1305
R19221 vss.n9176 vss.n9174 0.1305
R19222 vss.n9174 vss.n9173 0.1305
R19223 vss.n13143 vss.n13142 0.1305
R19224 vss.n13142 vss.n13141 0.1305
R19225 vss.n13146 vss.n13145 0.1305
R19226 vss.n13147 vss.n13146 0.1305
R19227 vss.n13156 vss.n13155 0.1305
R19228 vss.n13155 vss.n13154 0.1305
R19229 vss.n13158 vss.n8903 0.1305
R19230 vss.n8903 vss.n8901 0.1305
R19231 vss.n13140 vss.n13139 0.1305
R19232 vss.n13141 vss.n13140 0.1305
R19233 vss.n13149 vss.n13148 0.1305
R19234 vss.n13148 vss.n13147 0.1305
R19235 vss.n13153 vss.n13152 0.1305
R19236 vss.n13154 vss.n13153 0.1305
R19237 vss.n8904 vss.n8902 0.1305
R19238 vss.n8902 vss.n8901 0.1305
R19239 vss.n12801 vss.n12800 0.1305
R19240 vss.n12800 vss.n12799 0.1305
R19241 vss.n12716 vss.n12715 0.1305
R19242 vss.n12715 vss.n12700 0.1305
R19243 vss.n12821 vss.n12820 0.1305
R19244 vss.n12820 vss.n12819 0.1305
R19245 vss.n12823 vss.n12641 0.1305
R19246 vss.n12641 vss.n12639 0.1305
R19247 vss.n12798 vss.n12797 0.1305
R19248 vss.n12799 vss.n12798 0.1305
R19249 vss.n12713 vss.n12712 0.1305
R19250 vss.n12712 vss.n12700 0.1305
R19251 vss.n12818 vss.n12817 0.1305
R19252 vss.n12819 vss.n12818 0.1305
R19253 vss.n12642 vss.n12640 0.1305
R19254 vss.n12640 vss.n12639 0.1305
R19255 vss.n12878 vss.n12877 0.1305
R19256 vss.n12877 vss.n12876 0.1305
R19257 vss.n9380 vss.n9379 0.1305
R19258 vss.n9379 vss.n9364 0.1305
R19259 vss.n12898 vss.n12897 0.1305
R19260 vss.n12897 vss.n12896 0.1305
R19261 vss.n12900 vss.n9304 0.1305
R19262 vss.n9304 vss.n9302 0.1305
R19263 vss.n12875 vss.n12874 0.1305
R19264 vss.n12876 vss.n12875 0.1305
R19265 vss.n9377 vss.n9376 0.1305
R19266 vss.n9376 vss.n9364 0.1305
R19267 vss.n12895 vss.n12894 0.1305
R19268 vss.n12896 vss.n12895 0.1305
R19269 vss.n9305 vss.n9303 0.1305
R19270 vss.n9303 vss.n9302 0.1305
R19271 vss.n12832 vss.n9417 0.1305
R19272 vss.n12832 vss.n12831 0.1305
R19273 vss.n9411 vss.n9390 0.1305
R19274 vss.n12839 vss.n9411 0.1305
R19275 vss.n9389 vss.n9388 0.1305
R19276 vss.n9388 vss.n9373 0.1305
R19277 vss.n9370 vss.n9365 0.1305
R19278 vss.n12889 vss.n9365 0.1305
R19279 vss.n12888 vss.n12887 0.1305
R19280 vss.n12889 vss.n12888 0.1305
R19281 vss.n9384 vss.n9369 0.1305
R19282 vss.n9384 vss.n9373 0.1305
R19283 vss.n12838 vss.n12837 0.1305
R19284 vss.n12839 vss.n12838 0.1305
R19285 vss.n12830 vss.n9413 0.1305
R19286 vss.n12831 vss.n12830 0.1305
R19287 vss.n12781 vss.n12780 0.1305
R19288 vss.n12782 vss.n12781 0.1305
R19289 vss.n12792 vss.n12791 0.1305
R19290 vss.n12791 vss.n12790 0.1305
R19291 vss.n12725 vss.n12724 0.1305
R19292 vss.n12724 vss.n12709 0.1305
R19293 vss.n12706 vss.n12701 0.1305
R19294 vss.n12812 vss.n12701 0.1305
R19295 vss.n12811 vss.n12810 0.1305
R19296 vss.n12812 vss.n12811 0.1305
R19297 vss.n12720 vss.n12705 0.1305
R19298 vss.n12720 vss.n12709 0.1305
R19299 vss.n12789 vss.n12788 0.1305
R19300 vss.n12790 vss.n12789 0.1305
R19301 vss.n12784 vss.n12783 0.1305
R19302 vss.n12783 vss.n12782 0.1305
R19303 vss.n9168 vss.n9108 0.1305
R19304 vss.n9108 vss.n9106 0.1305
R19305 vss.n9160 vss.n8950 0.1305
R19306 vss.n9163 vss.n9160 0.1305
R19307 vss.n8949 vss.n8948 0.1305
R19308 vss.n8948 vss.n8926 0.1305
R19309 vss.n8934 vss.n8932 0.1305
R19310 vss.n8932 vss.n8918 0.1305
R19311 vss.n8941 vss.n8940 0.1305
R19312 vss.n8940 vss.n8918 0.1305
R19313 vss.n8943 vss.n8942 0.1305
R19314 vss.n8942 vss.n8926 0.1305
R19315 vss.n9162 vss.n9161 0.1305
R19316 vss.n9163 vss.n9162 0.1305
R19317 vss.n9109 vss.n9107 0.1305
R19318 vss.n9107 vss.n9106 0.1305
R19319 vss.n13309 vss.n8439 0.1305
R19320 vss.n13309 vss.n13308 0.1305
R19321 vss.n8435 vss.n8430 0.1305
R19322 vss.n13316 vss.n8430 0.1305
R19323 vss.n12975 vss.n12974 0.1305
R19324 vss.n12975 vss.n12956 0.1305
R19325 vss.n12960 vss.n12958 0.1305
R19326 vss.n12960 vss.n12948 0.1305
R19327 vss.n12967 vss.n12966 0.1305
R19328 vss.n12967 vss.n12948 0.1305
R19329 vss.n12969 vss.n12968 0.1305
R19330 vss.n12969 vss.n12956 0.1305
R19331 vss.n13315 vss.n13314 0.1305
R19332 vss.n13316 vss.n13315 0.1305
R19333 vss.n13307 vss.n8434 0.1305
R19334 vss.n13308 vss.n13307 0.1305
R19335 vss.n8574 vss.n8567 0.1305
R19336 vss.n8570 vss.n8567 0.1305
R19337 vss.n8579 vss.n8578 0.1305
R19338 vss.n8580 vss.n8579 0.1305
R19339 vss.n8595 vss.n8594 0.1305
R19340 vss.n8594 vss.n8512 0.1305
R19341 vss.n8593 vss.n8592 0.1305
R19342 vss.n8592 vss.n8504 0.1305
R19343 vss.n8586 vss.n8584 0.1305
R19344 vss.n8584 vss.n8504 0.1305
R19345 vss.n8601 vss.n8600 0.1305
R19346 vss.n8600 vss.n8512 0.1305
R19347 vss.n8582 vss.n8581 0.1305
R19348 vss.n8581 vss.n8580 0.1305
R19349 vss.n8569 vss.n8568 0.1305
R19350 vss.n8570 vss.n8569 0.1305
R19351 vss.n13428 vss.n13425 0.1305
R19352 vss.n13428 vss.n13427 0.1305
R19353 vss.n13421 vss.n13372 0.1305
R19354 vss.n13435 vss.n13372 0.1305
R19355 vss.n13401 vss.n13400 0.1305
R19356 vss.n13400 vss.n13377 0.1305
R19357 vss.n13399 vss.n13398 0.1305
R19358 vss.n13398 vss.n13384 0.1305
R19359 vss.n13393 vss.n13392 0.1305
R19360 vss.n13393 vss.n13384 0.1305
R19361 vss.n13387 vss.n13375 0.1305
R19362 vss.n13387 vss.n13377 0.1305
R19363 vss.n13434 vss.n13433 0.1305
R19364 vss.n13435 vss.n13434 0.1305
R19365 vss.n13426 vss.n13420 0.1305
R19366 vss.n13427 vss.n13426 0.1305
R19367 vss.n12070 vss.n12010 0.1305
R19368 vss.n12010 vss.n12008 0.1305
R19369 vss.n12062 vss.n8406 0.1305
R19370 vss.n12065 vss.n12062 0.1305
R19371 vss.n8405 vss.n8404 0.1305
R19372 vss.n8404 vss.n8382 0.1305
R19373 vss.n8390 vss.n8388 0.1305
R19374 vss.n8388 vss.n8374 0.1305
R19375 vss.n8397 vss.n8396 0.1305
R19376 vss.n8396 vss.n8374 0.1305
R19377 vss.n8399 vss.n8398 0.1305
R19378 vss.n8398 vss.n8382 0.1305
R19379 vss.n12064 vss.n12063 0.1305
R19380 vss.n12065 vss.n12064 0.1305
R19381 vss.n12011 vss.n12009 0.1305
R19382 vss.n12009 vss.n12008 0.1305
R19383 vss.n12128 vss.n11842 0.1305
R19384 vss.n11842 vss.n11840 0.1305
R19385 vss.n12126 vss.n12125 0.1305
R19386 vss.n12125 vss.n12124 0.1305
R19387 vss.n12096 vss.n11883 0.1305
R19388 vss.n12102 vss.n11883 0.1305
R19389 vss.n12095 vss.n12094 0.1305
R19390 vss.n12094 vss.n11880 0.1305
R19391 vss.n11887 vss.n11884 0.1305
R19392 vss.n11884 vss.n11880 0.1305
R19393 vss.n12101 vss.n11871 0.1305
R19394 vss.n12102 vss.n12101 0.1305
R19395 vss.n12123 vss.n12122 0.1305
R19396 vss.n12124 vss.n12123 0.1305
R19397 vss.n11843 vss.n11841 0.1305
R19398 vss.n11841 vss.n11840 0.1305
R19399 vss.n12113 vss.n11874 0.1305
R19400 vss.n11874 vss.n11872 0.1305
R19401 vss.n12111 vss.n12110 0.1305
R19402 vss.n12110 vss.n12109 0.1305
R19403 vss.n12084 vss.n12083 0.1305
R19404 vss.n12085 vss.n12084 0.1305
R19405 vss.n12081 vss.n12080 0.1305
R19406 vss.n12080 vss.n12079 0.1305
R19407 vss.n11875 vss.n11873 0.1305
R19408 vss.n11873 vss.n11872 0.1305
R19409 vss.n12108 vss.n12107 0.1305
R19410 vss.n12109 vss.n12108 0.1305
R19411 vss.n12087 vss.n12086 0.1305
R19412 vss.n12086 vss.n12085 0.1305
R19413 vss.n12078 vss.n12077 0.1305
R19414 vss.n12079 vss.n12078 0.1305
R19415 vss.n10632 vss.n10233 0.1305
R19416 vss.n10233 vss.n10231 0.1305
R19417 vss.n10630 vss.n10629 0.1305
R19418 vss.n10629 vss.n10628 0.1305
R19419 vss.n10620 vss.n10619 0.1305
R19420 vss.n10621 vss.n10620 0.1305
R19421 vss.n10391 vss.n10389 0.1305
R19422 vss.n10389 vss.n10387 0.1305
R19423 vss.n10390 vss.n10388 0.1305
R19424 vss.n10388 vss.n10387 0.1305
R19425 vss.n10623 vss.n10622 0.1305
R19426 vss.n10622 vss.n10621 0.1305
R19427 vss.n10627 vss.n10626 0.1305
R19428 vss.n10628 vss.n10627 0.1305
R19429 vss.n10234 vss.n10232 0.1305
R19430 vss.n10232 vss.n10231 0.1305
R19431 vss.n10767 vss.n10706 0.1305
R19432 vss.n10709 vss.n10706 0.1305
R19433 vss.n10770 vss.n10769 0.1305
R19434 vss.n10771 vss.n10770 0.1305
R19435 vss.n10779 vss.n10778 0.1305
R19436 vss.n10778 vss.n10777 0.1305
R19437 vss.n10781 vss.n10638 0.1305
R19438 vss.n10638 vss.n10636 0.1305
R19439 vss.n10639 vss.n10637 0.1305
R19440 vss.n10637 vss.n10636 0.1305
R19441 vss.n10776 vss.n10775 0.1305
R19442 vss.n10777 vss.n10776 0.1305
R19443 vss.n10773 vss.n10772 0.1305
R19444 vss.n10772 vss.n10771 0.1305
R19445 vss.n10708 vss.n10707 0.1305
R19446 vss.n10709 vss.n10708 0.1305
R19447 vss.n11025 vss.n10146 0.1305
R19448 vss.n10146 vss.n10144 0.1305
R19449 vss.n11023 vss.n11022 0.1305
R19450 vss.n11022 vss.n11021 0.1305
R19451 vss.n11013 vss.n11012 0.1305
R19452 vss.n11014 vss.n11013 0.1305
R19453 vss.n10759 vss.n10757 0.1305
R19454 vss.n10757 vss.n10755 0.1305
R19455 vss.n10758 vss.n10756 0.1305
R19456 vss.n10756 vss.n10755 0.1305
R19457 vss.n11016 vss.n11015 0.1305
R19458 vss.n11015 vss.n11014 0.1305
R19459 vss.n11020 vss.n11019 0.1305
R19460 vss.n11021 vss.n11020 0.1305
R19461 vss.n10147 vss.n10145 0.1305
R19462 vss.n10145 vss.n10144 0.1305
R19463 vss.n11319 vss.n10058 0.1305
R19464 vss.n10058 vss.n10056 0.1305
R19465 vss.n11317 vss.n11316 0.1305
R19466 vss.n11316 vss.n11315 0.1305
R19467 vss.n11307 vss.n11306 0.1305
R19468 vss.n11308 vss.n11307 0.1305
R19469 vss.n11033 vss.n11031 0.1305
R19470 vss.n11031 vss.n11029 0.1305
R19471 vss.n11032 vss.n11030 0.1305
R19472 vss.n11030 vss.n11029 0.1305
R19473 vss.n11310 vss.n11309 0.1305
R19474 vss.n11309 vss.n11308 0.1305
R19475 vss.n11314 vss.n11313 0.1305
R19476 vss.n11315 vss.n11314 0.1305
R19477 vss.n10059 vss.n10057 0.1305
R19478 vss.n10057 vss.n10056 0.1305
R19479 vss.n11345 vss.n9986 0.1305
R19480 vss.n9986 vss.n9984 0.1305
R19481 vss.n11343 vss.n11342 0.1305
R19482 vss.n11342 vss.n11341 0.1305
R19483 vss.n11333 vss.n11332 0.1305
R19484 vss.n11334 vss.n11333 0.1305
R19485 vss.n11329 vss.n11328 0.1305
R19486 vss.n11328 vss.n11327 0.1305
R19487 vss.n11326 vss.n11325 0.1305
R19488 vss.n11327 vss.n11326 0.1305
R19489 vss.n11336 vss.n11335 0.1305
R19490 vss.n11335 vss.n11334 0.1305
R19491 vss.n11340 vss.n11339 0.1305
R19492 vss.n11341 vss.n11340 0.1305
R19493 vss.n9987 vss.n9985 0.1305
R19494 vss.n9985 vss.n9984 0.1305
R19495 vss.n11424 vss.n11418 0.1305
R19496 vss.n11420 vss.n11418 0.1305
R19497 vss.n11427 vss.n11426 0.1305
R19498 vss.n11428 vss.n11427 0.1305
R19499 vss.n11436 vss.n11435 0.1305
R19500 vss.n11435 vss.n11434 0.1305
R19501 vss.n11438 vss.n11351 0.1305
R19502 vss.n11351 vss.n11349 0.1305
R19503 vss.n11352 vss.n11350 0.1305
R19504 vss.n11350 vss.n11349 0.1305
R19505 vss.n11433 vss.n11432 0.1305
R19506 vss.n11434 vss.n11433 0.1305
R19507 vss.n11430 vss.n11429 0.1305
R19508 vss.n11429 vss.n11428 0.1305
R19509 vss.n11421 vss.n11419 0.1305
R19510 vss.n11421 vss.n11420 0.1305
R19511 vss.n11661 vss.n11655 0.1305
R19512 vss.n11657 vss.n11655 0.1305
R19513 vss.n11664 vss.n11663 0.1305
R19514 vss.n11665 vss.n11664 0.1305
R19515 vss.n11673 vss.n11672 0.1305
R19516 vss.n11672 vss.n11671 0.1305
R19517 vss.n11675 vss.n9932 0.1305
R19518 vss.n9932 vss.n9930 0.1305
R19519 vss.n9933 vss.n9931 0.1305
R19520 vss.n9931 vss.n9930 0.1305
R19521 vss.n11670 vss.n11669 0.1305
R19522 vss.n11671 vss.n11670 0.1305
R19523 vss.n11667 vss.n11666 0.1305
R19524 vss.n11666 vss.n11665 0.1305
R19525 vss.n11658 vss.n11656 0.1305
R19526 vss.n11658 vss.n11657 0.1305
R19527 vss.n10364 vss.n10363 0.1305
R19528 vss.n10365 vss.n10364 0.1305
R19529 vss.n10374 vss.n10373 0.1305
R19530 vss.n10373 vss.n10372 0.1305
R19531 vss.n10378 vss.n10377 0.1305
R19532 vss.n10379 vss.n10378 0.1305
R19533 vss.n10276 vss.n10274 0.1305
R19534 vss.n10274 vss.n10273 0.1305
R19535 vss.n10383 vss.n10275 0.1305
R19536 vss.n10275 vss.n10273 0.1305
R19537 vss.n10381 vss.n10380 0.1305
R19538 vss.n10380 vss.n10379 0.1305
R19539 vss.n10371 vss.n10370 0.1305
R19540 vss.n10372 vss.n10371 0.1305
R19541 vss.n10367 vss.n10366 0.1305
R19542 vss.n10366 vss.n10365 0.1305
R19543 vss.n6741 vss.n6740 0.1255
R19544 vss.n6744 vss.n6743 0.1255
R19545 vss.n14090 vss.n2144 0.1255
R19546 vss.n8869 vss.n8867 0.0702092
R19547 vss.n8867 vss.n8866 0.0702092
R19548 vss.n13188 vss.n13187 0.0702092
R19549 vss.n13192 vss.n13188 0.0702092
R19550 vss.n10353 vss.n8878 0.0702092
R19551 vss.n10354 vss.n10353 0.0702092
R19552 vss.n10346 vss.n10344 0.0702092
R19553 vss.n10344 vss.n10343 0.0702092
R19554 vss.n10358 vss.n10345 0.0702092
R19555 vss.n10345 vss.n10343 0.0702092
R19556 vss.n10356 vss.n10355 0.0702092
R19557 vss.n10355 vss.n10354 0.0702092
R19558 vss.n13194 vss.n13193 0.0702092
R19559 vss.n13193 vss.n13192 0.0702092
R19560 vss.n13196 vss.n8868 0.0702092
R19561 vss.n8868 vss.n8866 0.0702092
R19562 vss.n10311 vss.n10300 0.0702092
R19563 vss.n10311 vss.n10310 0.0702092
R19564 vss.n10314 vss.n10313 0.0702092
R19565 vss.n10313 vss.n10293 0.0702092
R19566 vss.n10296 vss.n10292 0.0702092
R19567 vss.n10319 vss.n10292 0.0702092
R19568 vss.n10284 vss.n10282 0.0702092
R19569 vss.n10282 vss.n10281 0.0702092
R19570 vss.n10323 vss.n10283 0.0702092
R19571 vss.n10283 vss.n10281 0.0702092
R19572 vss.n10321 vss.n10320 0.0702092
R19573 vss.n10320 vss.n10319 0.0702092
R19574 vss.n10305 vss.n10304 0.0702092
R19575 vss.n10304 vss.n10293 0.0702092
R19576 vss.n10309 vss.n10308 0.0702092
R19577 vss.n10310 vss.n10309 0.0702092
R19578 vss.n11683 vss.n11682 0.0702092
R19579 vss.n11684 vss.n11683 0.0702092
R19580 vss.n11690 vss.n11689 0.0702092
R19581 vss.n11689 vss.n11688 0.0702092
R19582 vss.n11703 vss.n11702 0.0702092
R19583 vss.n11704 vss.n11703 0.0702092
R19584 vss.n11700 vss.n11699 0.0702092
R19585 vss.n11699 vss.n11698 0.0702092
R19586 vss.n11697 vss.n11696 0.0702092
R19587 vss.n11698 vss.n11697 0.0702092
R19588 vss.n11706 vss.n11705 0.0702092
R19589 vss.n11705 vss.n11704 0.0702092
R19590 vss.n11687 vss.n9912 0.0702092
R19591 vss.n11688 vss.n11687 0.0702092
R19592 vss.n11685 vss.n9928 0.0702092
R19593 vss.n11685 vss.n11684 0.0702092
R19594 vss.n11446 vss.n11445 0.0702092
R19595 vss.n11447 vss.n11446 0.0702092
R19596 vss.n11453 vss.n11452 0.0702092
R19597 vss.n11452 vss.n11451 0.0702092
R19598 vss.n11466 vss.n11465 0.0702092
R19599 vss.n11467 vss.n11466 0.0702092
R19600 vss.n11463 vss.n11462 0.0702092
R19601 vss.n11462 vss.n11461 0.0702092
R19602 vss.n11460 vss.n11459 0.0702092
R19603 vss.n11461 vss.n11460 0.0702092
R19604 vss.n11469 vss.n11468 0.0702092
R19605 vss.n11468 vss.n11467 0.0702092
R19606 vss.n11450 vss.n9967 0.0702092
R19607 vss.n11451 vss.n11450 0.0702092
R19608 vss.n11448 vss.n9983 0.0702092
R19609 vss.n11448 vss.n11447 0.0702092
R19610 vss.n11408 vss.n11368 0.0702092
R19611 vss.n11368 vss.n11366 0.0702092
R19612 vss.n11406 vss.n11405 0.0702092
R19613 vss.n11405 vss.n11404 0.0702092
R19614 vss.n11397 vss.n11396 0.0702092
R19615 vss.n11398 vss.n11397 0.0702092
R19616 vss.n11394 vss.n11393 0.0702092
R19617 vss.n11393 vss.n11392 0.0702092
R19618 vss.n11391 vss.n11390 0.0702092
R19619 vss.n11392 vss.n11391 0.0702092
R19620 vss.n11400 vss.n11399 0.0702092
R19621 vss.n11399 vss.n11398 0.0702092
R19622 vss.n11403 vss.n11402 0.0702092
R19623 vss.n11404 vss.n11403 0.0702092
R19624 vss.n11369 vss.n11367 0.0702092
R19625 vss.n11367 vss.n11366 0.0702092
R19626 vss.n11177 vss.n11176 0.0702092
R19627 vss.n11178 vss.n11177 0.0702092
R19628 vss.n11184 vss.n11183 0.0702092
R19629 vss.n11183 vss.n11182 0.0702092
R19630 vss.n11197 vss.n11196 0.0702092
R19631 vss.n11198 vss.n11197 0.0702092
R19632 vss.n11194 vss.n11193 0.0702092
R19633 vss.n11193 vss.n11192 0.0702092
R19634 vss.n11191 vss.n11190 0.0702092
R19635 vss.n11192 vss.n11191 0.0702092
R19636 vss.n11200 vss.n11199 0.0702092
R19637 vss.n11199 vss.n11198 0.0702092
R19638 vss.n11181 vss.n11158 0.0702092
R19639 vss.n11182 vss.n11181 0.0702092
R19640 vss.n11179 vss.n11174 0.0702092
R19641 vss.n11179 vss.n11178 0.0702092
R19642 vss.n11041 vss.n11040 0.0702092
R19643 vss.n11042 vss.n11041 0.0702092
R19644 vss.n11048 vss.n11047 0.0702092
R19645 vss.n11047 vss.n11046 0.0702092
R19646 vss.n11061 vss.n11060 0.0702092
R19647 vss.n11062 vss.n11061 0.0702092
R19648 vss.n11058 vss.n11057 0.0702092
R19649 vss.n11057 vss.n11056 0.0702092
R19650 vss.n11055 vss.n11054 0.0702092
R19651 vss.n11056 vss.n11055 0.0702092
R19652 vss.n11064 vss.n11063 0.0702092
R19653 vss.n11063 vss.n11062 0.0702092
R19654 vss.n11045 vss.n10127 0.0702092
R19655 vss.n11046 vss.n11045 0.0702092
R19656 vss.n11043 vss.n10143 0.0702092
R19657 vss.n11043 vss.n11042 0.0702092
R19658 vss.n10101 vss.n10100 0.0702092
R19659 vss.n10102 vss.n10101 0.0702092
R19660 vss.n10108 vss.n10107 0.0702092
R19661 vss.n10107 vss.n10106 0.0702092
R19662 vss.n10121 vss.n10120 0.0702092
R19663 vss.n10122 vss.n10121 0.0702092
R19664 vss.n10118 vss.n10117 0.0702092
R19665 vss.n10117 vss.n10116 0.0702092
R19666 vss.n10115 vss.n10114 0.0702092
R19667 vss.n10116 vss.n10115 0.0702092
R19668 vss.n10124 vss.n10123 0.0702092
R19669 vss.n10123 vss.n10122 0.0702092
R19670 vss.n10105 vss.n10081 0.0702092
R19671 vss.n10106 vss.n10105 0.0702092
R19672 vss.n10103 vss.n10097 0.0702092
R19673 vss.n10103 vss.n10102 0.0702092
R19674 vss.n10751 vss.n10712 0.0702092
R19675 vss.n10712 vss.n10710 0.0702092
R19676 vss.n10749 vss.n10748 0.0702092
R19677 vss.n10748 vss.n10747 0.0702092
R19678 vss.n10740 vss.n10739 0.0702092
R19679 vss.n10741 vss.n10740 0.0702092
R19680 vss.n10737 vss.n10736 0.0702092
R19681 vss.n10736 vss.n10735 0.0702092
R19682 vss.n10734 vss.n10733 0.0702092
R19683 vss.n10735 vss.n10734 0.0702092
R19684 vss.n10742 vss.n10725 0.0702092
R19685 vss.n10742 vss.n10741 0.0702092
R19686 vss.n10746 vss.n10745 0.0702092
R19687 vss.n10747 vss.n10746 0.0702092
R19688 vss.n10713 vss.n10711 0.0702092
R19689 vss.n10711 vss.n10710 0.0702092
R19690 vss.n10789 vss.n10788 0.0702092
R19691 vss.n10790 vss.n10789 0.0702092
R19692 vss.n10796 vss.n10795 0.0702092
R19693 vss.n10795 vss.n10794 0.0702092
R19694 vss.n10809 vss.n10808 0.0702092
R19695 vss.n10810 vss.n10809 0.0702092
R19696 vss.n10806 vss.n10805 0.0702092
R19697 vss.n10805 vss.n10804 0.0702092
R19698 vss.n10803 vss.n10802 0.0702092
R19699 vss.n10804 vss.n10803 0.0702092
R19700 vss.n10812 vss.n10811 0.0702092
R19701 vss.n10811 vss.n10810 0.0702092
R19702 vss.n10793 vss.n10214 0.0702092
R19703 vss.n10794 vss.n10793 0.0702092
R19704 vss.n10791 vss.n10230 0.0702092
R19705 vss.n10791 vss.n10790 0.0702092
R19706 vss.n10696 vss.n10656 0.0702092
R19707 vss.n10656 vss.n10654 0.0702092
R19708 vss.n10694 vss.n10693 0.0702092
R19709 vss.n10693 vss.n10692 0.0702092
R19710 vss.n10685 vss.n10684 0.0702092
R19711 vss.n10686 vss.n10685 0.0702092
R19712 vss.n10682 vss.n10681 0.0702092
R19713 vss.n10681 vss.n10680 0.0702092
R19714 vss.n10679 vss.n10678 0.0702092
R19715 vss.n10680 vss.n10679 0.0702092
R19716 vss.n10688 vss.n10687 0.0702092
R19717 vss.n10687 vss.n10686 0.0702092
R19718 vss.n10691 vss.n10690 0.0702092
R19719 vss.n10692 vss.n10691 0.0702092
R19720 vss.n10657 vss.n10655 0.0702092
R19721 vss.n10655 vss.n10654 0.0702092
R19722 vss.n10399 vss.n10398 0.0702092
R19723 vss.n10400 vss.n10399 0.0702092
R19724 vss.n10406 vss.n10405 0.0702092
R19725 vss.n10405 vss.n10404 0.0702092
R19726 vss.n10419 vss.n10418 0.0702092
R19727 vss.n10420 vss.n10419 0.0702092
R19728 vss.n10416 vss.n10415 0.0702092
R19729 vss.n10415 vss.n10414 0.0702092
R19730 vss.n10413 vss.n10412 0.0702092
R19731 vss.n10414 vss.n10413 0.0702092
R19732 vss.n10422 vss.n10421 0.0702092
R19733 vss.n10421 vss.n10420 0.0702092
R19734 vss.n10403 vss.n10256 0.0702092
R19735 vss.n10404 vss.n10403 0.0702092
R19736 vss.n10401 vss.n10272 0.0702092
R19737 vss.n10401 vss.n10400 0.0702092
R19738 vss.n11916 vss.n11915 0.0702092
R19739 vss.n11915 vss.n11914 0.0702092
R19740 vss.n11931 vss.n11891 0.0702092
R19741 vss.n11891 vss.n11889 0.0702092
R19742 vss.n11929 vss.n11928 0.0702092
R19743 vss.n11928 vss.n11927 0.0702092
R19744 vss.n11919 vss.n11918 0.0702092
R19745 vss.n11920 vss.n11919 0.0702092
R19746 vss.n11913 vss.n11912 0.0702092
R19747 vss.n11914 vss.n11913 0.0702092
R19748 vss.n11922 vss.n11921 0.0702092
R19749 vss.n11921 vss.n11920 0.0702092
R19750 vss.n11926 vss.n11925 0.0702092
R19751 vss.n11927 vss.n11926 0.0702092
R19752 vss.n11892 vss.n11890 0.0702092
R19753 vss.n11890 vss.n11889 0.0702092
R19754 vss.n9261 vss.n9258 0.0702092
R19755 vss.n9273 vss.n9258 0.0702092
R19756 vss.n9266 vss.n9263 0.0702092
R19757 vss.n9266 vss.n9265 0.0702092
R19758 vss.n13172 vss.n13171 0.0702092
R19759 vss.n13173 vss.n13172 0.0702092
R19760 vss.n13169 vss.n13168 0.0702092
R19761 vss.n13168 vss.n13167 0.0702092
R19762 vss.n13166 vss.n13165 0.0702092
R19763 vss.n13167 vss.n13166 0.0702092
R19764 vss.n13175 vss.n13174 0.0702092
R19765 vss.n13174 vss.n13173 0.0702092
R19766 vss.n9264 vss.n8885 0.0702092
R19767 vss.n9265 vss.n9264 0.0702092
R19768 vss.n9272 vss.n9271 0.0702092
R19769 vss.n9273 vss.n9272 0.0702092
R19770 vss.n12402 vss.n12401 0.0702092
R19771 vss.n12403 vss.n12402 0.0702092
R19772 vss.n12409 vss.n12408 0.0702092
R19773 vss.n12408 vss.n12407 0.0702092
R19774 vss.n12423 vss.n12422 0.0702092
R19775 vss.n12424 vss.n12423 0.0702092
R19776 vss.n12420 vss.n12419 0.0702092
R19777 vss.n12419 vss.n12418 0.0702092
R19778 vss.n12417 vss.n12416 0.0702092
R19779 vss.n12418 vss.n12417 0.0702092
R19780 vss.n12426 vss.n12425 0.0702092
R19781 vss.n12425 vss.n12424 0.0702092
R19782 vss.n12406 vss.n12383 0.0702092
R19783 vss.n12407 vss.n12406 0.0702092
R19784 vss.n12404 vss.n12399 0.0702092
R19785 vss.n12404 vss.n12403 0.0702092
R19786 vss.n13264 vss.n13263 0.0702092
R19787 vss.n13265 vss.n13264 0.0702092
R19788 vss.n13271 vss.n13270 0.0702092
R19789 vss.n13270 vss.n13269 0.0702092
R19790 vss.n13284 vss.n13283 0.0702092
R19791 vss.n13285 vss.n13284 0.0702092
R19792 vss.n13281 vss.n13280 0.0702092
R19793 vss.n13280 vss.n13279 0.0702092
R19794 vss.n13278 vss.n13277 0.0702092
R19795 vss.n13279 vss.n13278 0.0702092
R19796 vss.n13287 vss.n13286 0.0702092
R19797 vss.n13286 vss.n13285 0.0702092
R19798 vss.n13268 vss.n8620 0.0702092
R19799 vss.n13269 vss.n13268 0.0702092
R19800 vss.n13266 vss.n8636 0.0702092
R19801 vss.n13266 vss.n13265 0.0702092
R19802 vss.n12284 vss.n12283 0.0702092
R19803 vss.n12285 vss.n12284 0.0702092
R19804 vss.n12291 vss.n12290 0.0702092
R19805 vss.n12290 vss.n12289 0.0702092
R19806 vss.n12305 vss.n12304 0.0702092
R19807 vss.n12306 vss.n12305 0.0702092
R19808 vss.n12302 vss.n12301 0.0702092
R19809 vss.n12301 vss.n12300 0.0702092
R19810 vss.n12299 vss.n12298 0.0702092
R19811 vss.n12300 vss.n12299 0.0702092
R19812 vss.n12308 vss.n12307 0.0702092
R19813 vss.n12307 vss.n12306 0.0702092
R19814 vss.n12288 vss.n12265 0.0702092
R19815 vss.n12289 vss.n12288 0.0702092
R19816 vss.n12286 vss.n12281 0.0702092
R19817 vss.n12286 vss.n12285 0.0702092
R19818 vss.n8743 vss.n8740 0.0702092
R19819 vss.n8755 vss.n8740 0.0702092
R19820 vss.n8748 vss.n8745 0.0702092
R19821 vss.n8748 vss.n8747 0.0702092
R19822 vss.n13695 vss.n13694 0.0702092
R19823 vss.n13696 vss.n13695 0.0702092
R19824 vss.n13692 vss.n13691 0.0702092
R19825 vss.n13691 vss.n13690 0.0702092
R19826 vss.n13689 vss.n13688 0.0702092
R19827 vss.n13690 vss.n13689 0.0702092
R19828 vss.n13698 vss.n13697 0.0702092
R19829 vss.n13697 vss.n13696 0.0702092
R19830 vss.n8746 vss.n8341 0.0702092
R19831 vss.n8747 vss.n8746 0.0702092
R19832 vss.n8754 vss.n8753 0.0702092
R19833 vss.n8755 vss.n8754 0.0702092
R19834 vss.n11986 vss.n11985 0.0702092
R19835 vss.n11987 vss.n11986 0.0702092
R19836 vss.n11995 vss.n11994 0.0702092
R19837 vss.n11994 vss.n11993 0.0702092
R19838 vss.n11999 vss.n11998 0.0702092
R19839 vss.n12000 vss.n11999 0.0702092
R19840 vss.n11966 vss.n11964 0.0702092
R19841 vss.n11964 vss.n11963 0.0702092
R19842 vss.n12004 vss.n11965 0.0702092
R19843 vss.n11965 vss.n11963 0.0702092
R19844 vss.n12002 vss.n12001 0.0702092
R19845 vss.n12001 vss.n12000 0.0702092
R19846 vss.n11992 vss.n11991 0.0702092
R19847 vss.n11993 vss.n11992 0.0702092
R19848 vss.n11989 vss.n11988 0.0702092
R19849 vss.n11988 vss.n11987 0.0702092
R19850 vss.n12201 vss.n9854 0.0702092
R19851 vss.n12234 vss.n9854 0.0702092
R19852 vss.n12227 vss.n12226 0.0702092
R19853 vss.n12228 vss.n12227 0.0702092
R19854 vss.n12224 vss.n12223 0.0702092
R19855 vss.n12223 vss.n12222 0.0702092
R19856 vss.n12221 vss.n12220 0.0702092
R19857 vss.n12222 vss.n12221 0.0702092
R19858 vss.n12230 vss.n12229 0.0702092
R19859 vss.n12229 vss.n12228 0.0702092
R19860 vss.n12233 vss.n12232 0.0702092
R19861 vss.n12234 vss.n12233 0.0702092
R19862 vss.n8770 vss.n8759 0.0702092
R19863 vss.n8803 vss.n8759 0.0702092
R19864 vss.n8796 vss.n8795 0.0702092
R19865 vss.n8797 vss.n8796 0.0702092
R19866 vss.n8793 vss.n8792 0.0702092
R19867 vss.n8792 vss.n8791 0.0702092
R19868 vss.n8784 vss.n8783 0.0702092
R19869 vss.n8785 vss.n8784 0.0702092
R19870 vss.n8787 vss.n8786 0.0702092
R19871 vss.n8786 vss.n8785 0.0702092
R19872 vss.n8790 vss.n8789 0.0702092
R19873 vss.n8791 vss.n8790 0.0702092
R19874 vss.n8799 vss.n8798 0.0702092
R19875 vss.n8798 vss.n8797 0.0702092
R19876 vss.n8802 vss.n8801 0.0702092
R19877 vss.n8803 vss.n8802 0.0702092
R19878 vss.n8701 vss.n8691 0.0702092
R19879 vss.n8734 vss.n8691 0.0702092
R19880 vss.n8727 vss.n8726 0.0702092
R19881 vss.n8728 vss.n8727 0.0702092
R19882 vss.n8724 vss.n8723 0.0702092
R19883 vss.n8723 vss.n8722 0.0702092
R19884 vss.n8715 vss.n8714 0.0702092
R19885 vss.n8716 vss.n8715 0.0702092
R19886 vss.n8718 vss.n8717 0.0702092
R19887 vss.n8717 vss.n8716 0.0702092
R19888 vss.n8721 vss.n8720 0.0702092
R19889 vss.n8722 vss.n8721 0.0702092
R19890 vss.n8730 vss.n8729 0.0702092
R19891 vss.n8729 vss.n8728 0.0702092
R19892 vss.n8733 vss.n8732 0.0702092
R19893 vss.n8734 vss.n8733 0.0702092
R19894 vss.n9850 vss.n9849 0.0702092
R19895 vss.n9851 vss.n9850 0.0702092
R19896 vss.n9819 vss.n9818 0.0702092
R19897 vss.n9835 vss.n9834 0.0702092
R19898 vss.n9834 vss.n9833 0.0702092
R19899 vss.n9838 vss.n9837 0.0702092
R19900 vss.n9839 vss.n9838 0.0702092
R19901 vss.n9847 vss.n9846 0.0702092
R19902 vss.n9846 vss.n9845 0.0702092
R19903 vss.n9844 vss.n9843 0.0702092
R19904 vss.n9845 vss.n9844 0.0702092
R19905 vss.n9841 vss.n9840 0.0702092
R19906 vss.n9840 vss.n9839 0.0702092
R19907 vss.n9832 vss.n9831 0.0702092
R19908 vss.n9833 vss.n9832 0.0702092
R19909 vss.n9784 vss.n9777 0.0702092
R19910 vss.n9780 vss.n9777 0.0702092
R19911 vss.n9779 vss.n9778 0.0702092
R19912 vss.n9787 vss.n9786 0.0702092
R19913 vss.n9788 vss.n9787 0.0702092
R19914 vss.n9796 vss.n9795 0.0702092
R19915 vss.n9795 vss.n9794 0.0702092
R19916 vss.n9798 vss.n9757 0.0702092
R19917 vss.n9757 vss.n9755 0.0702092
R19918 vss.n9758 vss.n9756 0.0702092
R19919 vss.n9756 vss.n9755 0.0702092
R19920 vss.n9793 vss.n9792 0.0702092
R19921 vss.n9794 vss.n9793 0.0702092
R19922 vss.n9790 vss.n9789 0.0702092
R19923 vss.n9789 vss.n9788 0.0702092
R19924 vss.n12240 vss.n9749 0.0702092
R19925 vss.n12240 vss.n12239 0.0702092
R19926 vss.n9752 vss.n9751 0.0702092
R19927 vss.n12252 vss.n12251 0.0702092
R19928 vss.n12253 vss.n12252 0.0702092
R19929 vss.n12261 vss.n12260 0.0702092
R19930 vss.n12260 vss.n12259 0.0702092
R19931 vss.n12242 vss.n9733 0.0702092
R19932 vss.n12243 vss.n12242 0.0702092
R19933 vss.n12245 vss.n12244 0.0702092
R19934 vss.n12244 vss.n12243 0.0702092
R19935 vss.n12258 vss.n12257 0.0702092
R19936 vss.n12259 vss.n12258 0.0702092
R19937 vss.n12255 vss.n12254 0.0702092
R19938 vss.n12254 vss.n12253 0.0702092
R19939 vss.n12319 vss.n9726 0.0702092
R19940 vss.n12352 vss.n9726 0.0702092
R19941 vss.n12345 vss.n12344 0.0702092
R19942 vss.n12346 vss.n12345 0.0702092
R19943 vss.n12342 vss.n12341 0.0702092
R19944 vss.n12341 vss.n12340 0.0702092
R19945 vss.n12332 vss.n12331 0.0702092
R19946 vss.n12336 vss.n12335 0.0702092
R19947 vss.n12335 vss.n12334 0.0702092
R19948 vss.n12339 vss.n12338 0.0702092
R19949 vss.n12340 vss.n12339 0.0702092
R19950 vss.n12348 vss.n12347 0.0702092
R19951 vss.n12347 vss.n12346 0.0702092
R19952 vss.n12351 vss.n12350 0.0702092
R19953 vss.n12352 vss.n12351 0.0702092
R19954 vss.n8651 vss.n8640 0.0702092
R19955 vss.n8684 vss.n8640 0.0702092
R19956 vss.n8677 vss.n8676 0.0702092
R19957 vss.n8678 vss.n8677 0.0702092
R19958 vss.n8674 vss.n8673 0.0702092
R19959 vss.n8673 vss.n8672 0.0702092
R19960 vss.n8665 vss.n8664 0.0702092
R19961 vss.n8666 vss.n8665 0.0702092
R19962 vss.n8668 vss.n8667 0.0702092
R19963 vss.n8667 vss.n8666 0.0702092
R19964 vss.n8671 vss.n8670 0.0702092
R19965 vss.n8672 vss.n8671 0.0702092
R19966 vss.n8680 vss.n8679 0.0702092
R19967 vss.n8679 vss.n8678 0.0702092
R19968 vss.n8683 vss.n8682 0.0702092
R19969 vss.n8684 vss.n8683 0.0702092
R19970 vss.n12918 vss.n12917 0.0702092
R19971 vss.n12919 vss.n12918 0.0702092
R19972 vss.n12927 vss.n12926 0.0702092
R19973 vss.n12926 vss.n12925 0.0702092
R19974 vss.n12931 vss.n12930 0.0702092
R19975 vss.n12932 vss.n12931 0.0702092
R19976 vss.n9185 vss.n9183 0.0702092
R19977 vss.n9183 vss.n9182 0.0702092
R19978 vss.n12936 vss.n9184 0.0702092
R19979 vss.n9184 vss.n9182 0.0702092
R19980 vss.n12934 vss.n12933 0.0702092
R19981 vss.n12933 vss.n12932 0.0702092
R19982 vss.n12924 vss.n12923 0.0702092
R19983 vss.n12925 vss.n12924 0.0702092
R19984 vss.n12921 vss.n12920 0.0702092
R19985 vss.n12920 vss.n12919 0.0702092
R19986 vss.n9722 vss.n9721 0.0702092
R19987 vss.n9723 vss.n9722 0.0702092
R19988 vss.n9690 vss.n9689 0.0702092
R19989 vss.n9707 vss.n9706 0.0702092
R19990 vss.n9706 vss.n9705 0.0702092
R19991 vss.n9710 vss.n9709 0.0702092
R19992 vss.n9711 vss.n9710 0.0702092
R19993 vss.n9719 vss.n9718 0.0702092
R19994 vss.n9718 vss.n9717 0.0702092
R19995 vss.n9716 vss.n9715 0.0702092
R19996 vss.n9717 vss.n9716 0.0702092
R19997 vss.n9713 vss.n9712 0.0702092
R19998 vss.n9712 vss.n9711 0.0702092
R19999 vss.n9704 vss.n9703 0.0702092
R20000 vss.n9705 vss.n9704 0.0702092
R20001 vss.n9655 vss.n9647 0.0702092
R20002 vss.n9651 vss.n9647 0.0702092
R20003 vss.n9649 vss.n9648 0.0702092
R20004 vss.n9658 vss.n9657 0.0702092
R20005 vss.n9659 vss.n9658 0.0702092
R20006 vss.n9667 vss.n9666 0.0702092
R20007 vss.n9666 vss.n9665 0.0702092
R20008 vss.n9669 vss.n9627 0.0702092
R20009 vss.n9627 vss.n9625 0.0702092
R20010 vss.n9628 vss.n9626 0.0702092
R20011 vss.n9626 vss.n9625 0.0702092
R20012 vss.n9664 vss.n9663 0.0702092
R20013 vss.n9665 vss.n9664 0.0702092
R20014 vss.n9661 vss.n9660 0.0702092
R20015 vss.n9660 vss.n9659 0.0702092
R20016 vss.n12358 vss.n9619 0.0702092
R20017 vss.n12358 vss.n12357 0.0702092
R20018 vss.n9622 vss.n9621 0.0702092
R20019 vss.n12370 vss.n12369 0.0702092
R20020 vss.n12371 vss.n12370 0.0702092
R20021 vss.n12379 vss.n12378 0.0702092
R20022 vss.n12378 vss.n12377 0.0702092
R20023 vss.n12360 vss.n9603 0.0702092
R20024 vss.n12361 vss.n12360 0.0702092
R20025 vss.n12363 vss.n12362 0.0702092
R20026 vss.n12362 vss.n12361 0.0702092
R20027 vss.n12376 vss.n12375 0.0702092
R20028 vss.n12377 vss.n12376 0.0702092
R20029 vss.n12373 vss.n12372 0.0702092
R20030 vss.n12372 vss.n12371 0.0702092
R20031 vss.n12438 vss.n9596 0.0702092
R20032 vss.n12471 vss.n9596 0.0702092
R20033 vss.n12464 vss.n12463 0.0702092
R20034 vss.n12465 vss.n12464 0.0702092
R20035 vss.n12461 vss.n12460 0.0702092
R20036 vss.n12460 vss.n12459 0.0702092
R20037 vss.n12451 vss.n12450 0.0702092
R20038 vss.n12455 vss.n12454 0.0702092
R20039 vss.n12454 vss.n12453 0.0702092
R20040 vss.n12458 vss.n12457 0.0702092
R20041 vss.n12459 vss.n12458 0.0702092
R20042 vss.n12467 vss.n12466 0.0702092
R20043 vss.n12466 vss.n12465 0.0702092
R20044 vss.n12470 vss.n12469 0.0702092
R20045 vss.n12471 vss.n12470 0.0702092
R20046 vss.n9221 vss.n9210 0.0702092
R20047 vss.n9254 vss.n9210 0.0702092
R20048 vss.n9247 vss.n9246 0.0702092
R20049 vss.n9248 vss.n9247 0.0702092
R20050 vss.n9244 vss.n9243 0.0702092
R20051 vss.n9243 vss.n9242 0.0702092
R20052 vss.n9235 vss.n9234 0.0702092
R20053 vss.n9236 vss.n9235 0.0702092
R20054 vss.n9238 vss.n9237 0.0702092
R20055 vss.n9237 vss.n9236 0.0702092
R20056 vss.n9241 vss.n9240 0.0702092
R20057 vss.n9242 vss.n9241 0.0702092
R20058 vss.n9250 vss.n9249 0.0702092
R20059 vss.n9249 vss.n9248 0.0702092
R20060 vss.n9253 vss.n9252 0.0702092
R20061 vss.n9254 vss.n9253 0.0702092
R20062 vss.n9336 vss.n9335 0.0702092
R20063 vss.n9337 vss.n9336 0.0702092
R20064 vss.n9345 vss.n9344 0.0702092
R20065 vss.n9344 vss.n9343 0.0702092
R20066 vss.n9349 vss.n9348 0.0702092
R20067 vss.n9350 vss.n9349 0.0702092
R20068 vss.n9314 vss.n9312 0.0702092
R20069 vss.n9312 vss.n9311 0.0702092
R20070 vss.n9354 vss.n9313 0.0702092
R20071 vss.n9313 vss.n9311 0.0702092
R20072 vss.n9352 vss.n9351 0.0702092
R20073 vss.n9351 vss.n9350 0.0702092
R20074 vss.n9342 vss.n9341 0.0702092
R20075 vss.n9343 vss.n9342 0.0702092
R20076 vss.n9339 vss.n9338 0.0702092
R20077 vss.n9338 vss.n9337 0.0702092
R20078 vss.n12522 vss.n12521 0.0702092
R20079 vss.n12523 vss.n12522 0.0702092
R20080 vss.n12531 vss.n12530 0.0702092
R20081 vss.n12530 vss.n12529 0.0702092
R20082 vss.n12535 vss.n12534 0.0702092
R20083 vss.n12536 vss.n12535 0.0702092
R20084 vss.n9421 vss.n9419 0.0702092
R20085 vss.n9419 vss.n9418 0.0702092
R20086 vss.n12540 vss.n9420 0.0702092
R20087 vss.n9420 vss.n9418 0.0702092
R20088 vss.n12538 vss.n12537 0.0702092
R20089 vss.n12537 vss.n12536 0.0702092
R20090 vss.n12528 vss.n12527 0.0702092
R20091 vss.n12529 vss.n12528 0.0702092
R20092 vss.n12525 vss.n12524 0.0702092
R20093 vss.n12524 vss.n12523 0.0702092
R20094 vss.n12672 vss.n12671 0.0702092
R20095 vss.n12673 vss.n12672 0.0702092
R20096 vss.n12681 vss.n12680 0.0702092
R20097 vss.n12680 vss.n12679 0.0702092
R20098 vss.n12685 vss.n12684 0.0702092
R20099 vss.n12686 vss.n12685 0.0702092
R20100 vss.n12651 vss.n12649 0.0702092
R20101 vss.n12649 vss.n12648 0.0702092
R20102 vss.n12690 vss.n12650 0.0702092
R20103 vss.n12650 vss.n12648 0.0702092
R20104 vss.n12688 vss.n12687 0.0702092
R20105 vss.n12687 vss.n12686 0.0702092
R20106 vss.n12678 vss.n12677 0.0702092
R20107 vss.n12679 vss.n12678 0.0702092
R20108 vss.n12675 vss.n12674 0.0702092
R20109 vss.n12674 vss.n12673 0.0702092
R20110 vss.n9592 vss.n9591 0.0702092
R20111 vss.n9593 vss.n9592 0.0702092
R20112 vss.n9561 vss.n9560 0.0702092
R20113 vss.n9577 vss.n9576 0.0702092
R20114 vss.n9576 vss.n9575 0.0702092
R20115 vss.n9580 vss.n9579 0.0702092
R20116 vss.n9581 vss.n9580 0.0702092
R20117 vss.n9589 vss.n9588 0.0702092
R20118 vss.n9588 vss.n9587 0.0702092
R20119 vss.n9586 vss.n9585 0.0702092
R20120 vss.n9587 vss.n9586 0.0702092
R20121 vss.n9583 vss.n9582 0.0702092
R20122 vss.n9582 vss.n9581 0.0702092
R20123 vss.n9574 vss.n9573 0.0702092
R20124 vss.n9575 vss.n9574 0.0702092
R20125 vss.n9525 vss.n9518 0.0702092
R20126 vss.n9521 vss.n9518 0.0702092
R20127 vss.n9520 vss.n9519 0.0702092
R20128 vss.n9528 vss.n9527 0.0702092
R20129 vss.n9529 vss.n9528 0.0702092
R20130 vss.n9537 vss.n9536 0.0702092
R20131 vss.n9536 vss.n9535 0.0702092
R20132 vss.n9539 vss.n9498 0.0702092
R20133 vss.n9498 vss.n9496 0.0702092
R20134 vss.n9499 vss.n9497 0.0702092
R20135 vss.n9497 vss.n9496 0.0702092
R20136 vss.n9534 vss.n9533 0.0702092
R20137 vss.n9535 vss.n9534 0.0702092
R20138 vss.n9531 vss.n9530 0.0702092
R20139 vss.n9530 vss.n9529 0.0702092
R20140 vss.n12477 vss.n9490 0.0702092
R20141 vss.n12477 vss.n12476 0.0702092
R20142 vss.n9493 vss.n9492 0.0702092
R20143 vss.n12489 vss.n12488 0.0702092
R20144 vss.n12490 vss.n12489 0.0702092
R20145 vss.n12498 vss.n12497 0.0702092
R20146 vss.n12497 vss.n12496 0.0702092
R20147 vss.n12479 vss.n9474 0.0702092
R20148 vss.n12480 vss.n12479 0.0702092
R20149 vss.n12482 vss.n12481 0.0702092
R20150 vss.n12481 vss.n12480 0.0702092
R20151 vss.n12495 vss.n12494 0.0702092
R20152 vss.n12496 vss.n12495 0.0702092
R20153 vss.n12492 vss.n12491 0.0702092
R20154 vss.n12491 vss.n12490 0.0702092
R20155 vss.n9458 vss.n9457 0.0702092
R20156 vss.n9459 vss.n9458 0.0702092
R20157 vss.n9462 vss.n9461 0.0702092
R20158 vss.n9468 vss.n9467 0.0702092
R20159 vss.n9467 vss.n9466 0.0702092
R20160 vss.n9448 vss.n9424 0.0702092
R20161 vss.n9449 vss.n9448 0.0702092
R20162 vss.n9446 vss.n9440 0.0702092
R20163 vss.n9446 vss.n9445 0.0702092
R20164 vss.n9444 vss.n9443 0.0702092
R20165 vss.n9445 vss.n9444 0.0702092
R20166 vss.n9451 vss.n9450 0.0702092
R20167 vss.n9450 vss.n9449 0.0702092
R20168 vss.n9465 vss.n9464 0.0702092
R20169 vss.n9466 vss.n9465 0.0702092
R20170 vss.n11734 vss.n9878 0.0702092
R20171 vss.n11734 vss.n11733 0.0702092
R20172 vss.n11729 vss.n11728 0.0702092
R20173 vss.n11746 vss.n11745 0.0702092
R20174 vss.n11747 vss.n11746 0.0702092
R20175 vss.n11755 vss.n11754 0.0702092
R20176 vss.n11754 vss.n11753 0.0702092
R20177 vss.n11736 vss.n9862 0.0702092
R20178 vss.n11737 vss.n11736 0.0702092
R20179 vss.n11739 vss.n11738 0.0702092
R20180 vss.n11738 vss.n11737 0.0702092
R20181 vss.n11752 vss.n11751 0.0702092
R20182 vss.n11753 vss.n11752 0.0702092
R20183 vss.n11749 vss.n11748 0.0702092
R20184 vss.n11748 vss.n11747 0.0702092
R20185 vss.n12218 vss.n12217 0.0702092
R20186 vss.n12217 vss.n12216 0.0702092
R20187 vss.n12214 vss.n12213 0.0702092
R20188 vss.n11839 vss.n11838 0.0702092
R20189 vss.n12184 vss.n11839 0.0702092
R20190 vss.n11828 vss.n11810 0.0702092
R20191 vss.n12184 vss.n11810 0.0702092
R20192 vss.n12186 vss.n12185 0.0702092
R20193 vss.n12185 vss.n12184 0.0702092
R20194 vss.n11809 vss.n11804 0.0702092
R20195 vss.n12184 vss.n11809 0.0702092
R20196 vss.n11816 vss.n11815 0.0702092
R20197 vss.n11832 vss.n11816 0.0702092
R20198 vss.n11833 vss.n11819 0.0702092
R20199 vss.n11833 vss.n11832 0.0702092
R20200 vss.n11826 vss.n11820 0.0702092
R20201 vss.n11832 vss.n11820 0.0702092
R20202 vss.n11831 vss.n11830 0.0702092
R20203 vss.n11832 vss.n11831 0.0702092
R20204 vss.n3984 vss.n3971 0.0702092
R20205 vss.n3971 vss.n3969 0.0702092
R20206 vss.n15893 vss.n15892 0.0702092
R20207 vss.n15894 vss.n15893 0.0702092
R20208 vss.n15902 vss.n15901 0.0702092
R20209 vss.n15901 vss.n15900 0.0702092
R20210 vss.n3976 vss.n1 0.0702092
R20211 vss.n3979 vss.n3976 0.0702092
R20212 vss.n3972 vss.n3970 0.0702092
R20213 vss.n3970 vss.n3969 0.0702092
R20214 vss.n3978 vss.n3977 0.0702092
R20215 vss.n3979 vss.n3978 0.0702092
R20216 vss.n15899 vss.n15898 0.0702092
R20217 vss.n15900 vss.n15899 0.0702092
R20218 vss.n15896 vss.n15895 0.0702092
R20219 vss.n15895 vss.n15894 0.0702092
R20220 vss.n5652 vss.n5651 0.0702092
R20221 vss.n5653 vss.n5652 0.0702092
R20222 vss.n5659 vss.n5658 0.0702092
R20223 vss.n5658 vss.n5657 0.0702092
R20224 vss.n5672 vss.n5671 0.0702092
R20225 vss.n5673 vss.n5672 0.0702092
R20226 vss.n5669 vss.n5668 0.0702092
R20227 vss.n5668 vss.n5667 0.0702092
R20228 vss.n5666 vss.n5665 0.0702092
R20229 vss.n5667 vss.n5666 0.0702092
R20230 vss.n5675 vss.n5674 0.0702092
R20231 vss.n5674 vss.n5673 0.0702092
R20232 vss.n5656 vss.n5633 0.0702092
R20233 vss.n5657 vss.n5656 0.0702092
R20234 vss.n5654 vss.n5649 0.0702092
R20235 vss.n5654 vss.n5653 0.0702092
R20236 vss.n3715 vss.n3712 0.0702092
R20237 vss.n3727 vss.n3712 0.0702092
R20238 vss.n3720 vss.n3717 0.0702092
R20239 vss.n3720 vss.n3719 0.0702092
R20240 vss.n15752 vss.n15751 0.0702092
R20241 vss.n15753 vss.n15752 0.0702092
R20242 vss.n15749 vss.n15748 0.0702092
R20243 vss.n15748 vss.n15747 0.0702092
R20244 vss.n15746 vss.n15745 0.0702092
R20245 vss.n15747 vss.n15746 0.0702092
R20246 vss.n15755 vss.n15754 0.0702092
R20247 vss.n15754 vss.n15753 0.0702092
R20248 vss.n3718 vss.n166 0.0702092
R20249 vss.n3719 vss.n3718 0.0702092
R20250 vss.n3726 vss.n3725 0.0702092
R20251 vss.n3727 vss.n3726 0.0702092
R20252 vss.n3675 vss.n3665 0.0702092
R20253 vss.n3708 vss.n3665 0.0702092
R20254 vss.n3701 vss.n3700 0.0702092
R20255 vss.n3702 vss.n3701 0.0702092
R20256 vss.n3698 vss.n3697 0.0702092
R20257 vss.n3697 vss.n3696 0.0702092
R20258 vss.n3689 vss.n3688 0.0702092
R20259 vss.n3690 vss.n3689 0.0702092
R20260 vss.n3692 vss.n3691 0.0702092
R20261 vss.n3691 vss.n3690 0.0702092
R20262 vss.n3695 vss.n3694 0.0702092
R20263 vss.n3696 vss.n3695 0.0702092
R20264 vss.n3704 vss.n3703 0.0702092
R20265 vss.n3703 vss.n3702 0.0702092
R20266 vss.n3707 vss.n3706 0.0702092
R20267 vss.n3708 vss.n3707 0.0702092
R20268 vss.n5844 vss.n5843 0.0702092
R20269 vss.n5845 vss.n5844 0.0702092
R20270 vss.n5851 vss.n5850 0.0702092
R20271 vss.n5850 vss.n5849 0.0702092
R20272 vss.n5864 vss.n5863 0.0702092
R20273 vss.n5865 vss.n5864 0.0702092
R20274 vss.n5861 vss.n5860 0.0702092
R20275 vss.n5860 vss.n5859 0.0702092
R20276 vss.n5858 vss.n5857 0.0702092
R20277 vss.n5859 vss.n5858 0.0702092
R20278 vss.n5867 vss.n5866 0.0702092
R20279 vss.n5866 vss.n5865 0.0702092
R20280 vss.n5848 vss.n5825 0.0702092
R20281 vss.n5849 vss.n5848 0.0702092
R20282 vss.n5846 vss.n5841 0.0702092
R20283 vss.n5846 vss.n5845 0.0702092
R20284 vss.n3834 vss.n3831 0.0702092
R20285 vss.n3846 vss.n3831 0.0702092
R20286 vss.n3839 vss.n3836 0.0702092
R20287 vss.n3839 vss.n3838 0.0702092
R20288 vss.n15808 vss.n15807 0.0702092
R20289 vss.n15809 vss.n15808 0.0702092
R20290 vss.n15805 vss.n15804 0.0702092
R20291 vss.n15804 vss.n15803 0.0702092
R20292 vss.n15802 vss.n15801 0.0702092
R20293 vss.n15803 vss.n15802 0.0702092
R20294 vss.n15811 vss.n15810 0.0702092
R20295 vss.n15810 vss.n15809 0.0702092
R20296 vss.n3837 vss.n88 0.0702092
R20297 vss.n3838 vss.n3837 0.0702092
R20298 vss.n3845 vss.n3844 0.0702092
R20299 vss.n3846 vss.n3845 0.0702092
R20300 vss.n3794 vss.n3784 0.0702092
R20301 vss.n3827 vss.n3784 0.0702092
R20302 vss.n3820 vss.n3819 0.0702092
R20303 vss.n3821 vss.n3820 0.0702092
R20304 vss.n3817 vss.n3816 0.0702092
R20305 vss.n3816 vss.n3815 0.0702092
R20306 vss.n3808 vss.n3807 0.0702092
R20307 vss.n3809 vss.n3808 0.0702092
R20308 vss.n3811 vss.n3810 0.0702092
R20309 vss.n3810 vss.n3809 0.0702092
R20310 vss.n3814 vss.n3813 0.0702092
R20311 vss.n3815 vss.n3814 0.0702092
R20312 vss.n3823 vss.n3822 0.0702092
R20313 vss.n3822 vss.n3821 0.0702092
R20314 vss.n3826 vss.n3825 0.0702092
R20315 vss.n3827 vss.n3826 0.0702092
R20316 vss.n3913 vss.n3903 0.0702092
R20317 vss.n3946 vss.n3903 0.0702092
R20318 vss.n3939 vss.n3938 0.0702092
R20319 vss.n3940 vss.n3939 0.0702092
R20320 vss.n3936 vss.n3935 0.0702092
R20321 vss.n3935 vss.n3934 0.0702092
R20322 vss.n3927 vss.n3926 0.0702092
R20323 vss.n3928 vss.n3927 0.0702092
R20324 vss.n3930 vss.n3929 0.0702092
R20325 vss.n3929 vss.n3928 0.0702092
R20326 vss.n3933 vss.n3932 0.0702092
R20327 vss.n3934 vss.n3933 0.0702092
R20328 vss.n3942 vss.n3941 0.0702092
R20329 vss.n3941 vss.n3940 0.0702092
R20330 vss.n3945 vss.n3944 0.0702092
R20331 vss.n3946 vss.n3945 0.0702092
R20332 vss.n6084 vss.n6083 0.0702092
R20333 vss.n6085 vss.n6084 0.0702092
R20334 vss.n6091 vss.n6090 0.0702092
R20335 vss.n6090 vss.n6089 0.0702092
R20336 vss.n6104 vss.n6103 0.0702092
R20337 vss.n6105 vss.n6104 0.0702092
R20338 vss.n6101 vss.n6100 0.0702092
R20339 vss.n6100 vss.n6099 0.0702092
R20340 vss.n6098 vss.n6097 0.0702092
R20341 vss.n6099 vss.n6098 0.0702092
R20342 vss.n6107 vss.n6106 0.0702092
R20343 vss.n6106 vss.n6105 0.0702092
R20344 vss.n6088 vss.n6065 0.0702092
R20345 vss.n6089 vss.n6088 0.0702092
R20346 vss.n6086 vss.n6081 0.0702092
R20347 vss.n6086 vss.n6085 0.0702092
R20348 vss.n6329 vss.n3538 0.0702092
R20349 vss.n3538 vss.n3536 0.0702092
R20350 vss.n6318 vss.n6317 0.0702092
R20351 vss.n6319 vss.n6318 0.0702092
R20352 vss.n6327 vss.n6326 0.0702092
R20353 vss.n6326 vss.n6325 0.0702092
R20354 vss.n3539 vss.n3537 0.0702092
R20355 vss.n3537 vss.n3536 0.0702092
R20356 vss.n6324 vss.n6323 0.0702092
R20357 vss.n6325 vss.n6324 0.0702092
R20358 vss.n6321 vss.n6320 0.0702092
R20359 vss.n6320 vss.n6319 0.0702092
R20360 vss.n5609 vss.n5608 0.0702092
R20361 vss.n5609 vss.n3535 0.0702092
R20362 vss.n5604 vss.n5603 0.0702092
R20363 vss.n5621 vss.n5620 0.0702092
R20364 vss.n5622 vss.n5621 0.0702092
R20365 vss.n5630 vss.n5629 0.0702092
R20366 vss.n5629 vss.n5628 0.0702092
R20367 vss.n5611 vss.n5589 0.0702092
R20368 vss.n5612 vss.n5611 0.0702092
R20369 vss.n5614 vss.n5613 0.0702092
R20370 vss.n5613 vss.n5612 0.0702092
R20371 vss.n5627 vss.n5626 0.0702092
R20372 vss.n5628 vss.n5627 0.0702092
R20373 vss.n5624 vss.n5623 0.0702092
R20374 vss.n5623 vss.n5622 0.0702092
R20375 vss.n5705 vss.n5704 0.0702092
R20376 vss.n5704 vss.n5703 0.0702092
R20377 vss.n5701 vss.n5700 0.0702092
R20378 vss.n5708 vss.n5707 0.0702092
R20379 vss.n5709 vss.n5708 0.0702092
R20380 vss.n5717 vss.n5716 0.0702092
R20381 vss.n5716 vss.n5715 0.0702092
R20382 vss.n5719 vss.n5538 0.0702092
R20383 vss.n5538 vss.n5536 0.0702092
R20384 vss.n5539 vss.n5537 0.0702092
R20385 vss.n5537 vss.n5536 0.0702092
R20386 vss.n5714 vss.n5713 0.0702092
R20387 vss.n5715 vss.n5714 0.0702092
R20388 vss.n5711 vss.n5710 0.0702092
R20389 vss.n5710 vss.n5709 0.0702092
R20390 vss.n5564 vss.n5563 0.0702092
R20391 vss.n5564 vss.n5535 0.0702092
R20392 vss.n5559 vss.n5558 0.0702092
R20393 vss.n5576 vss.n5575 0.0702092
R20394 vss.n5577 vss.n5576 0.0702092
R20395 vss.n5585 vss.n5584 0.0702092
R20396 vss.n5584 vss.n5583 0.0702092
R20397 vss.n5566 vss.n5542 0.0702092
R20398 vss.n5567 vss.n5566 0.0702092
R20399 vss.n5569 vss.n5568 0.0702092
R20400 vss.n5568 vss.n5567 0.0702092
R20401 vss.n5582 vss.n5581 0.0702092
R20402 vss.n5583 vss.n5582 0.0702092
R20403 vss.n5579 vss.n5578 0.0702092
R20404 vss.n5578 vss.n5577 0.0702092
R20405 vss.n5943 vss.n5942 0.0702092
R20406 vss.n5942 vss.n5941 0.0702092
R20407 vss.n5939 vss.n5938 0.0702092
R20408 vss.n5946 vss.n5945 0.0702092
R20409 vss.n5947 vss.n5946 0.0702092
R20410 vss.n5955 vss.n5954 0.0702092
R20411 vss.n5954 vss.n5953 0.0702092
R20412 vss.n5957 vss.n5915 0.0702092
R20413 vss.n5915 vss.n5913 0.0702092
R20414 vss.n5916 vss.n5914 0.0702092
R20415 vss.n5914 vss.n5913 0.0702092
R20416 vss.n5952 vss.n5951 0.0702092
R20417 vss.n5953 vss.n5952 0.0702092
R20418 vss.n5949 vss.n5948 0.0702092
R20419 vss.n5948 vss.n5947 0.0702092
R20420 vss.n5911 vss.n5910 0.0702092
R20421 vss.n5912 vss.n5911 0.0702092
R20422 vss.n5880 vss.n5879 0.0702092
R20423 vss.n5896 vss.n5895 0.0702092
R20424 vss.n5895 vss.n5894 0.0702092
R20425 vss.n5899 vss.n5898 0.0702092
R20426 vss.n5900 vss.n5899 0.0702092
R20427 vss.n5908 vss.n5907 0.0702092
R20428 vss.n5907 vss.n5906 0.0702092
R20429 vss.n5905 vss.n5904 0.0702092
R20430 vss.n5906 vss.n5905 0.0702092
R20431 vss.n5902 vss.n5901 0.0702092
R20432 vss.n5901 vss.n5900 0.0702092
R20433 vss.n5893 vss.n5892 0.0702092
R20434 vss.n5894 vss.n5893 0.0702092
R20435 vss.n5810 vss.n5809 0.0702092
R20436 vss.n5811 vss.n5810 0.0702092
R20437 vss.n5814 vss.n5813 0.0702092
R20438 vss.n5820 vss.n5819 0.0702092
R20439 vss.n5819 vss.n5818 0.0702092
R20440 vss.n5800 vss.n5777 0.0702092
R20441 vss.n5801 vss.n5800 0.0702092
R20442 vss.n5798 vss.n5793 0.0702092
R20443 vss.n5798 vss.n5797 0.0702092
R20444 vss.n5796 vss.n5795 0.0702092
R20445 vss.n5797 vss.n5796 0.0702092
R20446 vss.n5803 vss.n5802 0.0702092
R20447 vss.n5802 vss.n5801 0.0702092
R20448 vss.n5817 vss.n5816 0.0702092
R20449 vss.n5818 vss.n5817 0.0702092
R20450 vss.n5752 vss.n5751 0.0702092
R20451 vss.n5752 vss.n3998 0.0702092
R20452 vss.n5747 vss.n5746 0.0702092
R20453 vss.n5764 vss.n5763 0.0702092
R20454 vss.n5765 vss.n5764 0.0702092
R20455 vss.n5773 vss.n5772 0.0702092
R20456 vss.n5772 vss.n5771 0.0702092
R20457 vss.n5754 vss.n5730 0.0702092
R20458 vss.n5755 vss.n5754 0.0702092
R20459 vss.n5757 vss.n5756 0.0702092
R20460 vss.n5756 vss.n5755 0.0702092
R20461 vss.n5770 vss.n5769 0.0702092
R20462 vss.n5771 vss.n5770 0.0702092
R20463 vss.n5767 vss.n5766 0.0702092
R20464 vss.n5766 vss.n5765 0.0702092
R20465 vss.n6182 vss.n6181 0.0702092
R20466 vss.n6181 vss.n6180 0.0702092
R20467 vss.n6178 vss.n6177 0.0702092
R20468 vss.n6185 vss.n6184 0.0702092
R20469 vss.n6186 vss.n6185 0.0702092
R20470 vss.n6194 vss.n6193 0.0702092
R20471 vss.n6193 vss.n6192 0.0702092
R20472 vss.n6196 vss.n6154 0.0702092
R20473 vss.n6154 vss.n6152 0.0702092
R20474 vss.n6155 vss.n6153 0.0702092
R20475 vss.n6153 vss.n6152 0.0702092
R20476 vss.n6191 vss.n6190 0.0702092
R20477 vss.n6192 vss.n6191 0.0702092
R20478 vss.n6188 vss.n6187 0.0702092
R20479 vss.n6187 vss.n6186 0.0702092
R20480 vss.n6150 vss.n6149 0.0702092
R20481 vss.n6151 vss.n6150 0.0702092
R20482 vss.n6119 vss.n6118 0.0702092
R20483 vss.n6135 vss.n6134 0.0702092
R20484 vss.n6134 vss.n6133 0.0702092
R20485 vss.n6138 vss.n6137 0.0702092
R20486 vss.n6139 vss.n6138 0.0702092
R20487 vss.n6147 vss.n6146 0.0702092
R20488 vss.n6146 vss.n6145 0.0702092
R20489 vss.n6144 vss.n6143 0.0702092
R20490 vss.n6145 vss.n6144 0.0702092
R20491 vss.n6141 vss.n6140 0.0702092
R20492 vss.n6140 vss.n6139 0.0702092
R20493 vss.n6132 vss.n6131 0.0702092
R20494 vss.n6133 vss.n6132 0.0702092
R20495 vss.n6050 vss.n6049 0.0702092
R20496 vss.n6051 vss.n6050 0.0702092
R20497 vss.n6054 vss.n6053 0.0702092
R20498 vss.n6060 vss.n6059 0.0702092
R20499 vss.n6059 vss.n6058 0.0702092
R20500 vss.n6040 vss.n6017 0.0702092
R20501 vss.n6041 vss.n6040 0.0702092
R20502 vss.n6038 vss.n6033 0.0702092
R20503 vss.n6038 vss.n6037 0.0702092
R20504 vss.n6036 vss.n6035 0.0702092
R20505 vss.n6037 vss.n6036 0.0702092
R20506 vss.n6043 vss.n6042 0.0702092
R20507 vss.n6042 vss.n6041 0.0702092
R20508 vss.n6057 vss.n6056 0.0702092
R20509 vss.n6058 vss.n6057 0.0702092
R20510 vss.n5994 vss.n5970 0.0702092
R20511 vss.n5995 vss.n5994 0.0702092
R20512 vss.n6004 vss.n6003 0.0702092
R20513 vss.n6005 vss.n6004 0.0702092
R20514 vss.n6013 vss.n6012 0.0702092
R20515 vss.n6012 vss.n6011 0.0702092
R20516 vss.n5997 vss.n5996 0.0702092
R20517 vss.n5996 vss.n5995 0.0702092
R20518 vss.n6010 vss.n6009 0.0702092
R20519 vss.n6011 vss.n6010 0.0702092
R20520 vss.n6007 vss.n6006 0.0702092
R20521 vss.n6006 vss.n6005 0.0702092
R20522 vss.n5992 vss.n5991 0.0702092
R20523 vss.n5992 vss.n3990 0.0702092
R20524 vss.n5987 vss.n5986 0.0702092
R20525 vss.n4550 vss.n4368 0.0702092
R20526 vss.n4368 vss.n4366 0.0702092
R20527 vss.n4548 vss.n4547 0.0702092
R20528 vss.n4547 vss.n4546 0.0702092
R20529 vss.n4397 vss.n4396 0.0702092
R20530 vss.n4398 vss.n4397 0.0702092
R20531 vss.n4394 vss.n4393 0.0702092
R20532 vss.n4393 vss.n4392 0.0702092
R20533 vss.n4391 vss.n4390 0.0702092
R20534 vss.n4392 vss.n4391 0.0702092
R20535 vss.n4400 vss.n4399 0.0702092
R20536 vss.n4399 vss.n4398 0.0702092
R20537 vss.n4545 vss.n4544 0.0702092
R20538 vss.n4546 vss.n4545 0.0702092
R20539 vss.n4369 vss.n4367 0.0702092
R20540 vss.n4367 vss.n4366 0.0702092
R20541 vss.n6635 vss.n6634 0.0702092
R20542 vss.n6636 vss.n6635 0.0702092
R20543 vss.n6642 vss.n6641 0.0702092
R20544 vss.n6641 vss.n6640 0.0702092
R20545 vss.n6655 vss.n6654 0.0702092
R20546 vss.n6656 vss.n6655 0.0702092
R20547 vss.n6652 vss.n6651 0.0702092
R20548 vss.n6651 vss.n6650 0.0702092
R20549 vss.n6649 vss.n6648 0.0702092
R20550 vss.n6650 vss.n6649 0.0702092
R20551 vss.n6658 vss.n6657 0.0702092
R20552 vss.n6657 vss.n6656 0.0702092
R20553 vss.n6639 vss.n6616 0.0702092
R20554 vss.n6640 vss.n6639 0.0702092
R20555 vss.n6637 vss.n6632 0.0702092
R20556 vss.n6637 vss.n6636 0.0702092
R20557 vss.n6586 vss.n6585 0.0702092
R20558 vss.n6587 vss.n6586 0.0702092
R20559 vss.n6593 vss.n6592 0.0702092
R20560 vss.n6592 vss.n6591 0.0702092
R20561 vss.n6607 vss.n6606 0.0702092
R20562 vss.n6608 vss.n6607 0.0702092
R20563 vss.n6604 vss.n6603 0.0702092
R20564 vss.n6603 vss.n6602 0.0702092
R20565 vss.n6601 vss.n6600 0.0702092
R20566 vss.n6602 vss.n6601 0.0702092
R20567 vss.n6610 vss.n6609 0.0702092
R20568 vss.n6609 vss.n6608 0.0702092
R20569 vss.n6590 vss.n6498 0.0702092
R20570 vss.n6591 vss.n6590 0.0702092
R20571 vss.n6588 vss.n6514 0.0702092
R20572 vss.n6588 vss.n6587 0.0702092
R20573 vss.n5233 vss.n5232 0.0702092
R20574 vss.n5234 vss.n5233 0.0702092
R20575 vss.n5240 vss.n5239 0.0702092
R20576 vss.n5239 vss.n5238 0.0702092
R20577 vss.n5253 vss.n5252 0.0702092
R20578 vss.n5254 vss.n5253 0.0702092
R20579 vss.n5250 vss.n5249 0.0702092
R20580 vss.n5249 vss.n5248 0.0702092
R20581 vss.n5247 vss.n5246 0.0702092
R20582 vss.n5248 vss.n5247 0.0702092
R20583 vss.n5256 vss.n5255 0.0702092
R20584 vss.n5255 vss.n5254 0.0702092
R20585 vss.n5237 vss.n5214 0.0702092
R20586 vss.n5238 vss.n5237 0.0702092
R20587 vss.n5235 vss.n5230 0.0702092
R20588 vss.n5235 vss.n5234 0.0702092
R20589 vss.n5445 vss.n5444 0.0702092
R20590 vss.n5446 vss.n5445 0.0702092
R20591 vss.n5452 vss.n5451 0.0702092
R20592 vss.n5451 vss.n5450 0.0702092
R20593 vss.n5465 vss.n5464 0.0702092
R20594 vss.n5466 vss.n5465 0.0702092
R20595 vss.n5462 vss.n5461 0.0702092
R20596 vss.n5461 vss.n5460 0.0702092
R20597 vss.n5459 vss.n5458 0.0702092
R20598 vss.n5460 vss.n5459 0.0702092
R20599 vss.n5468 vss.n5467 0.0702092
R20600 vss.n5467 vss.n5466 0.0702092
R20601 vss.n5449 vss.n5426 0.0702092
R20602 vss.n5450 vss.n5449 0.0702092
R20603 vss.n5447 vss.n5442 0.0702092
R20604 vss.n5447 vss.n5446 0.0702092
R20605 vss.n5398 vss.n5397 0.0702092
R20606 vss.n5399 vss.n5398 0.0702092
R20607 vss.n5405 vss.n5404 0.0702092
R20608 vss.n5404 vss.n5403 0.0702092
R20609 vss.n5418 vss.n5417 0.0702092
R20610 vss.n5419 vss.n5418 0.0702092
R20611 vss.n5415 vss.n5414 0.0702092
R20612 vss.n5414 vss.n5413 0.0702092
R20613 vss.n5412 vss.n5411 0.0702092
R20614 vss.n5413 vss.n5412 0.0702092
R20615 vss.n5421 vss.n5420 0.0702092
R20616 vss.n5420 vss.n5419 0.0702092
R20617 vss.n5402 vss.n5311 0.0702092
R20618 vss.n5403 vss.n5402 0.0702092
R20619 vss.n5400 vss.n5327 0.0702092
R20620 vss.n5400 vss.n5399 0.0702092
R20621 vss.n4148 vss.n4147 0.0702092
R20622 vss.n4149 vss.n4148 0.0702092
R20623 vss.n4155 vss.n4154 0.0702092
R20624 vss.n4154 vss.n4153 0.0702092
R20625 vss.n4168 vss.n4167 0.0702092
R20626 vss.n4169 vss.n4168 0.0702092
R20627 vss.n4165 vss.n4164 0.0702092
R20628 vss.n4164 vss.n4163 0.0702092
R20629 vss.n4162 vss.n4161 0.0702092
R20630 vss.n4163 vss.n4162 0.0702092
R20631 vss.n4171 vss.n4170 0.0702092
R20632 vss.n4170 vss.n4169 0.0702092
R20633 vss.n4152 vss.n4129 0.0702092
R20634 vss.n4153 vss.n4152 0.0702092
R20635 vss.n4150 vss.n4145 0.0702092
R20636 vss.n4150 vss.n4149 0.0702092
R20637 vss.n4971 vss.n4970 0.0702092
R20638 vss.n4972 vss.n4971 0.0702092
R20639 vss.n4978 vss.n4977 0.0702092
R20640 vss.n4977 vss.n4976 0.0702092
R20641 vss.n4991 vss.n4990 0.0702092
R20642 vss.n4992 vss.n4991 0.0702092
R20643 vss.n4988 vss.n4987 0.0702092
R20644 vss.n4987 vss.n4986 0.0702092
R20645 vss.n4985 vss.n4984 0.0702092
R20646 vss.n4986 vss.n4985 0.0702092
R20647 vss.n4994 vss.n4993 0.0702092
R20648 vss.n4993 vss.n4992 0.0702092
R20649 vss.n4975 vss.n4952 0.0702092
R20650 vss.n4976 vss.n4975 0.0702092
R20651 vss.n4973 vss.n4968 0.0702092
R20652 vss.n4973 vss.n4972 0.0702092
R20653 vss.n4102 vss.n4101 0.0702092
R20654 vss.n4103 vss.n4102 0.0702092
R20655 vss.n4109 vss.n4108 0.0702092
R20656 vss.n4108 vss.n4107 0.0702092
R20657 vss.n4122 vss.n4121 0.0702092
R20658 vss.n4123 vss.n4122 0.0702092
R20659 vss.n4119 vss.n4118 0.0702092
R20660 vss.n4118 vss.n4117 0.0702092
R20661 vss.n4116 vss.n4115 0.0702092
R20662 vss.n4117 vss.n4116 0.0702092
R20663 vss.n4125 vss.n4124 0.0702092
R20664 vss.n4124 vss.n4123 0.0702092
R20665 vss.n4106 vss.n4083 0.0702092
R20666 vss.n4107 vss.n4106 0.0702092
R20667 vss.n4104 vss.n4099 0.0702092
R20668 vss.n4104 vss.n4103 0.0702092
R20669 vss.n4923 vss.n4922 0.0702092
R20670 vss.n4924 vss.n4923 0.0702092
R20671 vss.n4930 vss.n4929 0.0702092
R20672 vss.n4929 vss.n4928 0.0702092
R20673 vss.n4943 vss.n4942 0.0702092
R20674 vss.n4944 vss.n4943 0.0702092
R20675 vss.n4940 vss.n4939 0.0702092
R20676 vss.n4939 vss.n4938 0.0702092
R20677 vss.n4937 vss.n4936 0.0702092
R20678 vss.n4938 vss.n4937 0.0702092
R20679 vss.n4946 vss.n4945 0.0702092
R20680 vss.n4945 vss.n4944 0.0702092
R20681 vss.n4927 vss.n4266 0.0702092
R20682 vss.n4928 vss.n4927 0.0702092
R20683 vss.n4925 vss.n4282 0.0702092
R20684 vss.n4925 vss.n4924 0.0702092
R20685 vss.n5186 vss.n5185 0.0702092
R20686 vss.n5187 vss.n5186 0.0702092
R20687 vss.n5193 vss.n5192 0.0702092
R20688 vss.n5192 vss.n5191 0.0702092
R20689 vss.n5206 vss.n5205 0.0702092
R20690 vss.n5207 vss.n5206 0.0702092
R20691 vss.n5203 vss.n5202 0.0702092
R20692 vss.n5202 vss.n5201 0.0702092
R20693 vss.n5200 vss.n5199 0.0702092
R20694 vss.n5201 vss.n5200 0.0702092
R20695 vss.n5209 vss.n5208 0.0702092
R20696 vss.n5208 vss.n5207 0.0702092
R20697 vss.n5190 vss.n5099 0.0702092
R20698 vss.n5191 vss.n5190 0.0702092
R20699 vss.n5188 vss.n5115 0.0702092
R20700 vss.n5188 vss.n5187 0.0702092
R20701 vss.n3361 vss.n3360 0.0702092
R20702 vss.n3362 vss.n3361 0.0702092
R20703 vss.n3368 vss.n3367 0.0702092
R20704 vss.n3367 vss.n3366 0.0702092
R20705 vss.n3381 vss.n3380 0.0702092
R20706 vss.n3382 vss.n3381 0.0702092
R20707 vss.n3378 vss.n3377 0.0702092
R20708 vss.n3377 vss.n3376 0.0702092
R20709 vss.n3375 vss.n3374 0.0702092
R20710 vss.n3376 vss.n3375 0.0702092
R20711 vss.n3384 vss.n3383 0.0702092
R20712 vss.n3383 vss.n3382 0.0702092
R20713 vss.n3365 vss.n3342 0.0702092
R20714 vss.n3366 vss.n3365 0.0702092
R20715 vss.n3363 vss.n3358 0.0702092
R20716 vss.n3363 vss.n3362 0.0702092
R20717 vss.n3408 vss.n3407 0.0702092
R20718 vss.n3409 vss.n3408 0.0702092
R20719 vss.n3415 vss.n3414 0.0702092
R20720 vss.n3414 vss.n3413 0.0702092
R20721 vss.n3428 vss.n3427 0.0702092
R20722 vss.n3429 vss.n3428 0.0702092
R20723 vss.n3425 vss.n3424 0.0702092
R20724 vss.n3424 vss.n3423 0.0702092
R20725 vss.n3422 vss.n3421 0.0702092
R20726 vss.n3423 vss.n3422 0.0702092
R20727 vss.n3431 vss.n3430 0.0702092
R20728 vss.n3430 vss.n3429 0.0702092
R20729 vss.n3412 vss.n3389 0.0702092
R20730 vss.n3413 vss.n3412 0.0702092
R20731 vss.n3410 vss.n3405 0.0702092
R20732 vss.n3410 vss.n3409 0.0702092
R20733 vss.n6470 vss.n6469 0.0702092
R20734 vss.n6471 vss.n6470 0.0702092
R20735 vss.n6477 vss.n6476 0.0702092
R20736 vss.n6476 vss.n6475 0.0702092
R20737 vss.n6490 vss.n6489 0.0702092
R20738 vss.n6491 vss.n6490 0.0702092
R20739 vss.n6487 vss.n6486 0.0702092
R20740 vss.n6486 vss.n6485 0.0702092
R20741 vss.n6484 vss.n6483 0.0702092
R20742 vss.n6485 vss.n6484 0.0702092
R20743 vss.n6493 vss.n6492 0.0702092
R20744 vss.n6492 vss.n6491 0.0702092
R20745 vss.n6474 vss.n6383 0.0702092
R20746 vss.n6475 vss.n6474 0.0702092
R20747 vss.n6472 vss.n6399 0.0702092
R20748 vss.n6472 vss.n6471 0.0702092
R20749 vss.n6685 vss.n6684 0.0702092
R20750 vss.n6684 vss.n6677 0.0702092
R20751 vss.n6679 vss.n6676 0.0702092
R20752 vss.n6690 vss.n6676 0.0702092
R20753 vss.n6698 vss.n6697 0.0702092
R20754 vss.n6697 vss.n6696 0.0702092
R20755 vss.n6695 vss.n6694 0.0702092
R20756 vss.n6696 vss.n6695 0.0702092
R20757 vss.n6692 vss.n6691 0.0702092
R20758 vss.n6691 vss.n6690 0.0702092
R20759 vss.n6682 vss.n6681 0.0702092
R20760 vss.n6682 vss.n6677 0.0702092
R20761 vss.n6701 vss.n6700 0.0702092
R20762 vss.n6702 vss.n6701 0.0702092
R20763 vss.n6670 vss.n6669 0.0702092
R20764 vss.n6373 vss.n3436 0.0702092
R20765 vss.n6361 vss.n3436 0.0702092
R20766 vss.n6357 vss.n3435 0.0702092
R20767 vss.n6357 vss.n6340 0.0702092
R20768 vss.n6355 vss.n6343 0.0702092
R20769 vss.n6355 vss.n6354 0.0702092
R20770 vss.n6353 vss.n6352 0.0702092
R20771 vss.n6354 vss.n6353 0.0702092
R20772 vss.n6350 vss.n6349 0.0702092
R20773 vss.n6349 vss.n6340 0.0702092
R20774 vss.n6363 vss.n6362 0.0702092
R20775 vss.n6362 vss.n6361 0.0702092
R20776 vss.n6371 vss.n6370 0.0702092
R20777 vss.n6370 vss.n6369 0.0702092
R20778 vss.n6366 vss.n6365 0.0702092
R20779 vss.n3444 vss.n3442 0.0702092
R20780 vss.n3442 vss.n3441 0.0702092
R20781 vss.n3475 vss.n3474 0.0702092
R20782 vss.n3479 vss.n3475 0.0702092
R20783 vss.n3471 vss.n3453 0.0702092
R20784 vss.n3471 vss.n3470 0.0702092
R20785 vss.n3469 vss.n3468 0.0702092
R20786 vss.n3470 vss.n3469 0.0702092
R20787 vss.n3481 vss.n3480 0.0702092
R20788 vss.n3480 vss.n3479 0.0702092
R20789 vss.n3483 vss.n3443 0.0702092
R20790 vss.n3443 vss.n3441 0.0702092
R20791 vss.n3462 vss.n3461 0.0702092
R20792 vss.n3463 vss.n3462 0.0702092
R20793 vss.n3466 vss.n3465 0.0702092
R20794 vss.n3522 vss.n3521 0.0702092
R20795 vss.n3527 vss.n3522 0.0702092
R20796 vss.n3518 vss.n3517 0.0702092
R20797 vss.n3517 vss.n3516 0.0702092
R20798 vss.n3509 vss.n3508 0.0702092
R20799 vss.n3510 vss.n3509 0.0702092
R20800 vss.n3512 vss.n3511 0.0702092
R20801 vss.n3511 vss.n3510 0.0702092
R20802 vss.n3515 vss.n3514 0.0702092
R20803 vss.n3516 vss.n3515 0.0702092
R20804 vss.n3529 vss.n3528 0.0702092
R20805 vss.n3528 vss.n3527 0.0702092
R20806 vss.n3491 vss.n3489 0.0702092
R20807 vss.n3489 vss.n3488 0.0702092
R20808 vss.n3531 vss.n3490 0.0702092
R20809 vss.n5293 vss.n5292 0.0702092
R20810 vss.n5295 vss.n5293 0.0702092
R20811 vss.n5303 vss.n5302 0.0702092
R20812 vss.n5302 vss.n5301 0.0702092
R20813 vss.n5283 vss.n5259 0.0702092
R20814 vss.n5284 vss.n5283 0.0702092
R20815 vss.n5286 vss.n5285 0.0702092
R20816 vss.n5285 vss.n5284 0.0702092
R20817 vss.n5300 vss.n5299 0.0702092
R20818 vss.n5301 vss.n5300 0.0702092
R20819 vss.n5297 vss.n5296 0.0702092
R20820 vss.n5296 vss.n5295 0.0702092
R20821 vss.n5281 vss.n5275 0.0702092
R20822 vss.n5281 vss.n5280 0.0702092
R20823 vss.n5278 vss.n5277 0.0702092
R20824 vss.n5523 vss.n5522 0.0702092
R20825 vss.n5525 vss.n5523 0.0702092
R20826 vss.n4037 vss.n4036 0.0702092
R20827 vss.n4036 vss.n4035 0.0702092
R20828 vss.n4027 vss.n4026 0.0702092
R20829 vss.n4028 vss.n4027 0.0702092
R20830 vss.n4030 vss.n4029 0.0702092
R20831 vss.n4029 vss.n4028 0.0702092
R20832 vss.n4034 vss.n4033 0.0702092
R20833 vss.n4035 vss.n4034 0.0702092
R20834 vss.n5526 vss.n4013 0.0702092
R20835 vss.n5526 vss.n5525 0.0702092
R20836 vss.n5533 vss.n5532 0.0702092
R20837 vss.n5534 vss.n5533 0.0702092
R20838 vss.n5530 vss.n5529 0.0702092
R20839 vss.n5508 vss.n5507 0.0702092
R20840 vss.n5509 vss.n5508 0.0702092
R20841 vss.n5517 vss.n5516 0.0702092
R20842 vss.n5516 vss.n5515 0.0702092
R20843 vss.n5498 vss.n5474 0.0702092
R20844 vss.n5499 vss.n5498 0.0702092
R20845 vss.n5501 vss.n5500 0.0702092
R20846 vss.n5500 vss.n5499 0.0702092
R20847 vss.n5514 vss.n5513 0.0702092
R20848 vss.n5515 vss.n5514 0.0702092
R20849 vss.n5511 vss.n5510 0.0702092
R20850 vss.n5510 vss.n5509 0.0702092
R20851 vss.n5496 vss.n5490 0.0702092
R20852 vss.n5496 vss.n5495 0.0702092
R20853 vss.n5493 vss.n5492 0.0702092
R20854 vss.n4080 vss.n4079 0.0702092
R20855 vss.n4079 vss.n4078 0.0702092
R20856 vss.n4062 vss.n4039 0.0702092
R20857 vss.n4063 vss.n4062 0.0702092
R20858 vss.n4060 vss.n4055 0.0702092
R20859 vss.n4060 vss.n4059 0.0702092
R20860 vss.n4058 vss.n4057 0.0702092
R20861 vss.n4059 vss.n4058 0.0702092
R20862 vss.n4065 vss.n4064 0.0702092
R20863 vss.n4064 vss.n4063 0.0702092
R20864 vss.n4077 vss.n4076 0.0702092
R20865 vss.n4078 vss.n4077 0.0702092
R20866 vss.n4070 vss.n4069 0.0702092
R20867 vss.n4069 vss.n4000 0.0702092
R20868 vss.n4074 vss.n4073 0.0702092
R20869 vss.n5082 vss.n5081 0.0702092
R20870 vss.n5083 vss.n5082 0.0702092
R20871 vss.n5091 vss.n5090 0.0702092
R20872 vss.n5090 vss.n5089 0.0702092
R20873 vss.n5072 vss.n5048 0.0702092
R20874 vss.n5073 vss.n5072 0.0702092
R20875 vss.n5075 vss.n5074 0.0702092
R20876 vss.n5074 vss.n5073 0.0702092
R20877 vss.n5088 vss.n5087 0.0702092
R20878 vss.n5089 vss.n5088 0.0702092
R20879 vss.n5085 vss.n5084 0.0702092
R20880 vss.n5084 vss.n5083 0.0702092
R20881 vss.n5070 vss.n5064 0.0702092
R20882 vss.n5070 vss.n5069 0.0702092
R20883 vss.n5067 vss.n5066 0.0702092
R20884 vss.n4217 vss.n4175 0.0702092
R20885 vss.n4180 vss.n4175 0.0702092
R20886 vss.n4196 vss.n4174 0.0702092
R20887 vss.n4200 vss.n4196 0.0702092
R20888 vss.n4194 vss.n4189 0.0702092
R20889 vss.n4194 vss.n4193 0.0702092
R20890 vss.n4192 vss.n4191 0.0702092
R20891 vss.n4193 vss.n4192 0.0702092
R20892 vss.n4202 vss.n4201 0.0702092
R20893 vss.n4201 vss.n4200 0.0702092
R20894 vss.n4207 vss.n4206 0.0702092
R20895 vss.n4207 vss.n4180 0.0702092
R20896 vss.n4215 vss.n4214 0.0702092
R20897 vss.n4214 vss.n3997 0.0702092
R20898 vss.n4204 vss.n4179 0.0702092
R20899 vss.n5034 vss.n5033 0.0702092
R20900 vss.n5035 vss.n5034 0.0702092
R20901 vss.n5043 vss.n5042 0.0702092
R20902 vss.n5042 vss.n5041 0.0702092
R20903 vss.n5024 vss.n5000 0.0702092
R20904 vss.n5025 vss.n5024 0.0702092
R20905 vss.n5027 vss.n5026 0.0702092
R20906 vss.n5026 vss.n5025 0.0702092
R20907 vss.n5040 vss.n5039 0.0702092
R20908 vss.n5041 vss.n5040 0.0702092
R20909 vss.n5037 vss.n5036 0.0702092
R20910 vss.n5036 vss.n5035 0.0702092
R20911 vss.n5022 vss.n5016 0.0702092
R20912 vss.n5022 vss.n5021 0.0702092
R20913 vss.n5019 vss.n5018 0.0702092
R20914 vss.n4261 vss.n4260 0.0702092
R20915 vss.n4260 vss.n4259 0.0702092
R20916 vss.n4243 vss.n4220 0.0702092
R20917 vss.n4244 vss.n4243 0.0702092
R20918 vss.n4241 vss.n4236 0.0702092
R20919 vss.n4241 vss.n4240 0.0702092
R20920 vss.n4239 vss.n4238 0.0702092
R20921 vss.n4240 vss.n4239 0.0702092
R20922 vss.n4246 vss.n4245 0.0702092
R20923 vss.n4245 vss.n4244 0.0702092
R20924 vss.n4258 vss.n4257 0.0702092
R20925 vss.n4259 vss.n4258 0.0702092
R20926 vss.n4251 vss.n4250 0.0702092
R20927 vss.n4250 vss.n3992 0.0702092
R20928 vss.n4255 vss.n4254 0.0702092
R20929 vss.n4529 vss.n4528 0.0702092
R20930 vss.n4530 vss.n4529 0.0702092
R20931 vss.n4538 vss.n4537 0.0702092
R20932 vss.n4537 vss.n4536 0.0702092
R20933 vss.n4519 vss.n4495 0.0702092
R20934 vss.n4520 vss.n4519 0.0702092
R20935 vss.n4522 vss.n4521 0.0702092
R20936 vss.n4521 vss.n4520 0.0702092
R20937 vss.n4535 vss.n4534 0.0702092
R20938 vss.n4536 vss.n4535 0.0702092
R20939 vss.n4532 vss.n4531 0.0702092
R20940 vss.n4531 vss.n4530 0.0702092
R20941 vss.n4517 vss.n4511 0.0702092
R20942 vss.n4517 vss.n4516 0.0702092
R20943 vss.n4514 vss.n4513 0.0702092
R20944 vss.n4491 vss.n4490 0.0702092
R20945 vss.n4490 vss.n4489 0.0702092
R20946 vss.n4471 vss.n4448 0.0702092
R20947 vss.n4472 vss.n4471 0.0702092
R20948 vss.n4469 vss.n4464 0.0702092
R20949 vss.n4469 vss.n4468 0.0702092
R20950 vss.n4467 vss.n4466 0.0702092
R20951 vss.n4468 vss.n4467 0.0702092
R20952 vss.n4474 vss.n4473 0.0702092
R20953 vss.n4473 vss.n4472 0.0702092
R20954 vss.n4488 vss.n4487 0.0702092
R20955 vss.n4489 vss.n4488 0.0702092
R20956 vss.n4481 vss.n4480 0.0702092
R20957 vss.n4481 vss.n3989 0.0702092
R20958 vss.n4485 vss.n4484 0.0702092
R20959 vss.n4421 vss.n4420 0.0702092
R20960 vss.n4422 vss.n4421 0.0702092
R20961 vss.n4428 vss.n4427 0.0702092
R20962 vss.n4427 vss.n4426 0.0702092
R20963 vss.n4441 vss.n4440 0.0702092
R20964 vss.n4442 vss.n4441 0.0702092
R20965 vss.n4438 vss.n4437 0.0702092
R20966 vss.n4437 vss.n4436 0.0702092
R20967 vss.n4435 vss.n4434 0.0702092
R20968 vss.n4436 vss.n4435 0.0702092
R20969 vss.n4444 vss.n4443 0.0702092
R20970 vss.n4443 vss.n4442 0.0702092
R20971 vss.n4425 vss.n4402 0.0702092
R20972 vss.n4426 vss.n4425 0.0702092
R20973 vss.n4423 vss.n4418 0.0702092
R20974 vss.n4423 vss.n4422 0.0702092
R20975 vss.n4796 vss.n4755 0.0702092
R20976 vss.n4755 vss.n4753 0.0702092
R20977 vss.n4794 vss.n4793 0.0702092
R20978 vss.n4793 vss.n4792 0.0702092
R20979 vss.n4784 vss.n4783 0.0702092
R20980 vss.n4785 vss.n4784 0.0702092
R20981 vss.n4781 vss.n4780 0.0702092
R20982 vss.n4780 vss.n4779 0.0702092
R20983 vss.n4778 vss.n4777 0.0702092
R20984 vss.n4779 vss.n4778 0.0702092
R20985 vss.n4787 vss.n4786 0.0702092
R20986 vss.n4786 vss.n4785 0.0702092
R20987 vss.n4791 vss.n4790 0.0702092
R20988 vss.n4792 vss.n4791 0.0702092
R20989 vss.n4756 vss.n4754 0.0702092
R20990 vss.n4754 vss.n4753 0.0702092
R20991 vss.n3294 vss.n3293 0.0702092
R20992 vss.n3295 vss.n3294 0.0702092
R20993 vss.n3301 vss.n3300 0.0702092
R20994 vss.n3300 vss.n3299 0.0702092
R20995 vss.n6734 vss.n6733 0.0702092
R20996 vss.n6735 vss.n6734 0.0702092
R20997 vss.n6731 vss.n6730 0.0702092
R20998 vss.n6730 vss.n6729 0.0702092
R20999 vss.n3296 vss.n3291 0.0702092
R21000 vss.n3296 vss.n3295 0.0702092
R21001 vss.n3298 vss.n3275 0.0702092
R21002 vss.n3299 vss.n3298 0.0702092
R21003 vss.n6737 vss.n6736 0.0702092
R21004 vss.n6736 vss.n6735 0.0702092
R21005 vss.n6728 vss.n6727 0.0702092
R21006 vss.n6729 vss.n6728 0.0702092
R21007 vss.n15526 vss.n15525 0.0702092
R21008 vss.n15527 vss.n15526 0.0702092
R21009 vss.n15529 vss.n15528 0.0702092
R21010 vss.n15528 vss.n15527 0.0702092
R21011 vss.n15523 vss.n15522 0.0702092
R21012 vss.n15522 vss.n15521 0.0702092
R21013 vss.n15520 vss.n15519 0.0702092
R21014 vss.n15521 vss.n15520 0.0702092
R21015 vss.n1061 vss.n1060 0.0702092
R21016 vss.n1062 vss.n1061 0.0702092
R21017 vss.n1068 vss.n1067 0.0702092
R21018 vss.n1067 vss.n1066 0.0702092
R21019 vss.n15044 vss.n15043 0.0702092
R21020 vss.n15045 vss.n15044 0.0702092
R21021 vss.n15041 vss.n15040 0.0702092
R21022 vss.n15040 vss.n15039 0.0702092
R21023 vss.n15038 vss.n15037 0.0702092
R21024 vss.n15039 vss.n15038 0.0702092
R21025 vss.n15047 vss.n15046 0.0702092
R21026 vss.n15046 vss.n15045 0.0702092
R21027 vss.n1065 vss.n1042 0.0702092
R21028 vss.n1066 vss.n1065 0.0702092
R21029 vss.n1063 vss.n1058 0.0702092
R21030 vss.n1063 vss.n1062 0.0702092
R21031 vss.n14914 vss.n14889 0.0702092
R21032 vss.n14915 vss.n14914 0.0702092
R21033 vss.n14924 vss.n14923 0.0702092
R21034 vss.n14925 vss.n14924 0.0702092
R21035 vss.n14933 vss.n14932 0.0702092
R21036 vss.n14932 vss.n14931 0.0702092
R21037 vss.n14917 vss.n14916 0.0702092
R21038 vss.n14916 vss.n14915 0.0702092
R21039 vss.n14930 vss.n14929 0.0702092
R21040 vss.n14931 vss.n14930 0.0702092
R21041 vss.n14927 vss.n14926 0.0702092
R21042 vss.n14926 vss.n14925 0.0702092
R21043 vss.n14912 vss.n14905 0.0702092
R21044 vss.n14912 vss.n14911 0.0702092
R21045 vss.n14908 vss.n14907 0.0702092
R21046 vss.n523 vss.n522 0.0702092
R21047 vss.n524 vss.n523 0.0702092
R21048 vss.n530 vss.n529 0.0702092
R21049 vss.n529 vss.n528 0.0702092
R21050 vss.n15438 vss.n15437 0.0702092
R21051 vss.n15439 vss.n15438 0.0702092
R21052 vss.n15435 vss.n15434 0.0702092
R21053 vss.n15434 vss.n15433 0.0702092
R21054 vss.n15432 vss.n15431 0.0702092
R21055 vss.n15433 vss.n15432 0.0702092
R21056 vss.n15441 vss.n15440 0.0702092
R21057 vss.n15440 vss.n15439 0.0702092
R21058 vss.n527 vss.n504 0.0702092
R21059 vss.n528 vss.n527 0.0702092
R21060 vss.n525 vss.n520 0.0702092
R21061 vss.n525 vss.n524 0.0702092
R21062 vss.n7321 vss.n7320 0.0702092
R21063 vss.n7322 vss.n7321 0.0702092
R21064 vss.n7328 vss.n7327 0.0702092
R21065 vss.n7327 vss.n7326 0.0702092
R21066 vss.n7341 vss.n7340 0.0702092
R21067 vss.n7342 vss.n7341 0.0702092
R21068 vss.n7338 vss.n7337 0.0702092
R21069 vss.n7337 vss.n7336 0.0702092
R21070 vss.n7335 vss.n7334 0.0702092
R21071 vss.n7336 vss.n7335 0.0702092
R21072 vss.n7344 vss.n7343 0.0702092
R21073 vss.n7343 vss.n7342 0.0702092
R21074 vss.n7325 vss.n7302 0.0702092
R21075 vss.n7326 vss.n7325 0.0702092
R21076 vss.n7323 vss.n7318 0.0702092
R21077 vss.n7323 vss.n7322 0.0702092
R21078 vss.n728 vss.n727 0.0702092
R21079 vss.n729 vss.n728 0.0702092
R21080 vss.n735 vss.n734 0.0702092
R21081 vss.n734 vss.n733 0.0702092
R21082 vss.n15365 vss.n15364 0.0702092
R21083 vss.n15366 vss.n15365 0.0702092
R21084 vss.n15362 vss.n15361 0.0702092
R21085 vss.n15361 vss.n15360 0.0702092
R21086 vss.n15359 vss.n15358 0.0702092
R21087 vss.n15360 vss.n15359 0.0702092
R21088 vss.n15368 vss.n15367 0.0702092
R21089 vss.n15367 vss.n15366 0.0702092
R21090 vss.n732 vss.n709 0.0702092
R21091 vss.n733 vss.n732 0.0702092
R21092 vss.n730 vss.n725 0.0702092
R21093 vss.n730 vss.n729 0.0702092
R21094 vss.n781 vss.n780 0.0702092
R21095 vss.n782 vss.n781 0.0702092
R21096 vss.n788 vss.n787 0.0702092
R21097 vss.n787 vss.n786 0.0702092
R21098 vss.n15288 vss.n15287 0.0702092
R21099 vss.n15289 vss.n15288 0.0702092
R21100 vss.n15285 vss.n15284 0.0702092
R21101 vss.n15284 vss.n15283 0.0702092
R21102 vss.n15282 vss.n15281 0.0702092
R21103 vss.n15283 vss.n15282 0.0702092
R21104 vss.n15291 vss.n15290 0.0702092
R21105 vss.n15290 vss.n15289 0.0702092
R21106 vss.n785 vss.n762 0.0702092
R21107 vss.n786 vss.n785 0.0702092
R21108 vss.n783 vss.n778 0.0702092
R21109 vss.n783 vss.n782 0.0702092
R21110 vss.n15195 vss.n15194 0.0702092
R21111 vss.n15196 vss.n15195 0.0702092
R21112 vss.n15202 vss.n15201 0.0702092
R21113 vss.n15201 vss.n15200 0.0702092
R21114 vss.n15215 vss.n15214 0.0702092
R21115 vss.n15216 vss.n15215 0.0702092
R21116 vss.n15212 vss.n15211 0.0702092
R21117 vss.n15211 vss.n15210 0.0702092
R21118 vss.n15209 vss.n15208 0.0702092
R21119 vss.n15210 vss.n15209 0.0702092
R21120 vss.n15218 vss.n15217 0.0702092
R21121 vss.n15217 vss.n15216 0.0702092
R21122 vss.n15199 vss.n15176 0.0702092
R21123 vss.n15200 vss.n15199 0.0702092
R21124 vss.n15197 vss.n15192 0.0702092
R21125 vss.n15197 vss.n15196 0.0702092
R21126 vss.n938 vss.n937 0.0702092
R21127 vss.n939 vss.n938 0.0702092
R21128 vss.n945 vss.n944 0.0702092
R21129 vss.n944 vss.n943 0.0702092
R21130 vss.n959 vss.n958 0.0702092
R21131 vss.n960 vss.n959 0.0702092
R21132 vss.n956 vss.n955 0.0702092
R21133 vss.n955 vss.n954 0.0702092
R21134 vss.n953 vss.n952 0.0702092
R21135 vss.n954 vss.n953 0.0702092
R21136 vss.n962 vss.n961 0.0702092
R21137 vss.n961 vss.n960 0.0702092
R21138 vss.n942 vss.n919 0.0702092
R21139 vss.n943 vss.n942 0.0702092
R21140 vss.n940 vss.n935 0.0702092
R21141 vss.n940 vss.n939 0.0702092
R21142 vss.n829 vss.n828 0.0702092
R21143 vss.n830 vss.n829 0.0702092
R21144 vss.n838 vss.n837 0.0702092
R21145 vss.n837 vss.n836 0.0702092
R21146 vss.n842 vss.n841 0.0702092
R21147 vss.n843 vss.n842 0.0702092
R21148 vss.n808 vss.n806 0.0702092
R21149 vss.n806 vss.n805 0.0702092
R21150 vss.n847 vss.n807 0.0702092
R21151 vss.n807 vss.n805 0.0702092
R21152 vss.n845 vss.n844 0.0702092
R21153 vss.n844 vss.n843 0.0702092
R21154 vss.n835 vss.n834 0.0702092
R21155 vss.n836 vss.n835 0.0702092
R21156 vss.n832 vss.n831 0.0702092
R21157 vss.n831 vss.n830 0.0702092
R21158 vss.n15137 vss.n15136 0.0702092
R21159 vss.n15136 vss.n15135 0.0702092
R21160 vss.n15125 vss.n15124 0.0702092
R21161 vss.n15124 vss.n15123 0.0702092
R21162 vss.n15128 vss.n15127 0.0702092
R21163 vss.n15129 vss.n15128 0.0702092
R21164 vss.n15134 vss.n15133 0.0702092
R21165 vss.n15135 vss.n15134 0.0702092
R21166 vss.n15131 vss.n15130 0.0702092
R21167 vss.n15130 vss.n15129 0.0702092
R21168 vss.n15122 vss.n15121 0.0702092
R21169 vss.n15123 vss.n15122 0.0702092
R21170 vss.n7453 vss.n7442 0.0702092
R21171 vss.n7486 vss.n7442 0.0702092
R21172 vss.n7479 vss.n7478 0.0702092
R21173 vss.n7480 vss.n7479 0.0702092
R21174 vss.n7476 vss.n7475 0.0702092
R21175 vss.n7475 vss.n7474 0.0702092
R21176 vss.n7466 vss.n7465 0.0702092
R21177 vss.n7470 vss.n7469 0.0702092
R21178 vss.n7469 vss.n7468 0.0702092
R21179 vss.n7473 vss.n7472 0.0702092
R21180 vss.n7474 vss.n7473 0.0702092
R21181 vss.n7482 vss.n7481 0.0702092
R21182 vss.n7481 vss.n7480 0.0702092
R21183 vss.n7485 vss.n7484 0.0702092
R21184 vss.n7486 vss.n7485 0.0702092
R21185 vss.n15315 vss.n15314 0.0702092
R21186 vss.n15316 vss.n15315 0.0702092
R21187 vss.n15322 vss.n15321 0.0702092
R21188 vss.n15321 vss.n15320 0.0702092
R21189 vss.n15336 vss.n15335 0.0702092
R21190 vss.n15337 vss.n15336 0.0702092
R21191 vss.n15333 vss.n15332 0.0702092
R21192 vss.n15332 vss.n15331 0.0702092
R21193 vss.n15330 vss.n15329 0.0702092
R21194 vss.n15331 vss.n15330 0.0702092
R21195 vss.n15339 vss.n15338 0.0702092
R21196 vss.n15338 vss.n15337 0.0702092
R21197 vss.n15319 vss.n15296 0.0702092
R21198 vss.n15320 vss.n15319 0.0702092
R21199 vss.n15317 vss.n15312 0.0702092
R21200 vss.n15317 vss.n15316 0.0702092
R21201 vss.n681 vss.n680 0.0702092
R21202 vss.n682 vss.n681 0.0702092
R21203 vss.n688 vss.n687 0.0702092
R21204 vss.n687 vss.n686 0.0702092
R21205 vss.n702 vss.n701 0.0702092
R21206 vss.n703 vss.n702 0.0702092
R21207 vss.n699 vss.n698 0.0702092
R21208 vss.n698 vss.n697 0.0702092
R21209 vss.n696 vss.n695 0.0702092
R21210 vss.n697 vss.n696 0.0702092
R21211 vss.n705 vss.n704 0.0702092
R21212 vss.n704 vss.n703 0.0702092
R21213 vss.n685 vss.n662 0.0702092
R21214 vss.n686 vss.n685 0.0702092
R21215 vss.n683 vss.n678 0.0702092
R21216 vss.n683 vss.n682 0.0702092
R21217 vss.n7438 vss.n7437 0.0702092
R21218 vss.n7439 vss.n7438 0.0702092
R21219 vss.n7407 vss.n7406 0.0702092
R21220 vss.n7423 vss.n7422 0.0702092
R21221 vss.n7422 vss.n7421 0.0702092
R21222 vss.n7426 vss.n7425 0.0702092
R21223 vss.n7427 vss.n7426 0.0702092
R21224 vss.n7435 vss.n7434 0.0702092
R21225 vss.n7434 vss.n7433 0.0702092
R21226 vss.n7432 vss.n7431 0.0702092
R21227 vss.n7433 vss.n7432 0.0702092
R21228 vss.n7429 vss.n7428 0.0702092
R21229 vss.n7428 vss.n7427 0.0702092
R21230 vss.n7420 vss.n7419 0.0702092
R21231 vss.n7421 vss.n7420 0.0702092
R21232 vss.n7375 vss.n7368 0.0702092
R21233 vss.n7371 vss.n7368 0.0702092
R21234 vss.n7370 vss.n7369 0.0702092
R21235 vss.n7378 vss.n7377 0.0702092
R21236 vss.n7379 vss.n7378 0.0702092
R21237 vss.n7387 vss.n7386 0.0702092
R21238 vss.n7386 vss.n7385 0.0702092
R21239 vss.n7389 vss.n3061 0.0702092
R21240 vss.n3061 vss.n3059 0.0702092
R21241 vss.n3062 vss.n3060 0.0702092
R21242 vss.n3060 vss.n3059 0.0702092
R21243 vss.n7384 vss.n7383 0.0702092
R21244 vss.n7385 vss.n7384 0.0702092
R21245 vss.n7381 vss.n7380 0.0702092
R21246 vss.n7380 vss.n7379 0.0702092
R21247 vss.n3087 vss.n3086 0.0702092
R21248 vss.n3087 vss.n3058 0.0702092
R21249 vss.n3082 vss.n3081 0.0702092
R21250 vss.n3099 vss.n3098 0.0702092
R21251 vss.n3100 vss.n3099 0.0702092
R21252 vss.n3108 vss.n3107 0.0702092
R21253 vss.n3107 vss.n3106 0.0702092
R21254 vss.n3089 vss.n3065 0.0702092
R21255 vss.n3090 vss.n3089 0.0702092
R21256 vss.n3092 vss.n3091 0.0702092
R21257 vss.n3091 vss.n3090 0.0702092
R21258 vss.n3105 vss.n3104 0.0702092
R21259 vss.n3106 vss.n3105 0.0702092
R21260 vss.n3102 vss.n3101 0.0702092
R21261 vss.n3101 vss.n3100 0.0702092
R21262 vss.n7274 vss.n7273 0.0702092
R21263 vss.n7275 vss.n7274 0.0702092
R21264 vss.n7281 vss.n7280 0.0702092
R21265 vss.n7280 vss.n7279 0.0702092
R21266 vss.n7295 vss.n7294 0.0702092
R21267 vss.n7296 vss.n7295 0.0702092
R21268 vss.n7292 vss.n7291 0.0702092
R21269 vss.n7288 vss.n7287 0.0702092
R21270 vss.n7288 vss.n7286 0.0702092
R21271 vss.n7298 vss.n7297 0.0702092
R21272 vss.n7297 vss.n7296 0.0702092
R21273 vss.n7278 vss.n3111 0.0702092
R21274 vss.n7279 vss.n7278 0.0702092
R21275 vss.n7276 vss.n3127 0.0702092
R21276 vss.n7276 vss.n7275 0.0702092
R21277 vss.n572 vss.n571 0.0702092
R21278 vss.n573 vss.n572 0.0702092
R21279 vss.n581 vss.n580 0.0702092
R21280 vss.n580 vss.n579 0.0702092
R21281 vss.n585 vss.n584 0.0702092
R21282 vss.n586 vss.n585 0.0702092
R21283 vss.n550 vss.n548 0.0702092
R21284 vss.n548 vss.n547 0.0702092
R21285 vss.n590 vss.n549 0.0702092
R21286 vss.n549 vss.n547 0.0702092
R21287 vss.n588 vss.n587 0.0702092
R21288 vss.n587 vss.n586 0.0702092
R21289 vss.n578 vss.n577 0.0702092
R21290 vss.n579 vss.n578 0.0702092
R21291 vss.n575 vss.n574 0.0702092
R21292 vss.n574 vss.n573 0.0702092
R21293 vss.n473 vss.n472 0.0702092
R21294 vss.n474 vss.n473 0.0702092
R21295 vss.n480 vss.n479 0.0702092
R21296 vss.n479 vss.n478 0.0702092
R21297 vss.n494 vss.n493 0.0702092
R21298 vss.n495 vss.n494 0.0702092
R21299 vss.n491 vss.n490 0.0702092
R21300 vss.n490 vss.n489 0.0702092
R21301 vss.n488 vss.n487 0.0702092
R21302 vss.n489 vss.n488 0.0702092
R21303 vss.n497 vss.n496 0.0702092
R21304 vss.n496 vss.n495 0.0702092
R21305 vss.n477 vss.n454 0.0702092
R21306 vss.n478 vss.n477 0.0702092
R21307 vss.n475 vss.n470 0.0702092
R21308 vss.n475 vss.n474 0.0702092
R21309 vss.n4723 vss.n4722 0.0702092
R21310 vss.n4724 vss.n4723 0.0702092
R21311 vss.n4732 vss.n4731 0.0702092
R21312 vss.n4731 vss.n4730 0.0702092
R21313 vss.n4736 vss.n4735 0.0702092
R21314 vss.n4737 vss.n4736 0.0702092
R21315 vss.n4557 vss.n4555 0.0702092
R21316 vss.n4555 vss.n4554 0.0702092
R21317 vss.n4741 vss.n4556 0.0702092
R21318 vss.n4556 vss.n4554 0.0702092
R21319 vss.n4739 vss.n4738 0.0702092
R21320 vss.n4738 vss.n4737 0.0702092
R21321 vss.n4729 vss.n4728 0.0702092
R21322 vss.n4730 vss.n4729 0.0702092
R21323 vss.n4726 vss.n4725 0.0702092
R21324 vss.n4725 vss.n4724 0.0702092
R21325 vss.n4338 vss.n4337 0.0702092
R21326 vss.n4339 vss.n4338 0.0702092
R21327 vss.n4347 vss.n4346 0.0702092
R21328 vss.n4346 vss.n4345 0.0702092
R21329 vss.n4351 vss.n4350 0.0702092
R21330 vss.n4352 vss.n4351 0.0702092
R21331 vss.n4317 vss.n4315 0.0702092
R21332 vss.n4315 vss.n4314 0.0702092
R21333 vss.n4356 vss.n4316 0.0702092
R21334 vss.n4316 vss.n4314 0.0702092
R21335 vss.n4354 vss.n4353 0.0702092
R21336 vss.n4353 vss.n4352 0.0702092
R21337 vss.n4344 vss.n4343 0.0702092
R21338 vss.n4345 vss.n4344 0.0702092
R21339 vss.n4341 vss.n4340 0.0702092
R21340 vss.n4340 vss.n4339 0.0702092
R21341 vss.n7268 vss.n7267 0.0702092
R21342 vss.n7269 vss.n7268 0.0702092
R21343 vss.n7237 vss.n7236 0.0702092
R21344 vss.n7253 vss.n7252 0.0702092
R21345 vss.n7252 vss.n7251 0.0702092
R21346 vss.n7256 vss.n7255 0.0702092
R21347 vss.n7257 vss.n7256 0.0702092
R21348 vss.n7265 vss.n7264 0.0702092
R21349 vss.n7264 vss.n7263 0.0702092
R21350 vss.n7262 vss.n7261 0.0702092
R21351 vss.n7263 vss.n7262 0.0702092
R21352 vss.n7259 vss.n7258 0.0702092
R21353 vss.n7258 vss.n7257 0.0702092
R21354 vss.n7250 vss.n7249 0.0702092
R21355 vss.n7251 vss.n7250 0.0702092
R21356 vss.n4641 vss.n4640 0.0702092
R21357 vss.n4642 vss.n4641 0.0702092
R21358 vss.n4645 vss.n4644 0.0702092
R21359 vss.n4651 vss.n4650 0.0702092
R21360 vss.n4650 vss.n4649 0.0702092
R21361 vss.n4631 vss.n4608 0.0702092
R21362 vss.n4632 vss.n4631 0.0702092
R21363 vss.n4629 vss.n4624 0.0702092
R21364 vss.n4629 vss.n4628 0.0702092
R21365 vss.n4627 vss.n4626 0.0702092
R21366 vss.n4628 vss.n4627 0.0702092
R21367 vss.n4634 vss.n4633 0.0702092
R21368 vss.n4633 vss.n4632 0.0702092
R21369 vss.n4648 vss.n4647 0.0702092
R21370 vss.n4649 vss.n4648 0.0702092
R21371 vss.n4678 vss.n4677 0.0702092
R21372 vss.n4678 vss.n3132 0.0702092
R21373 vss.n4673 vss.n4672 0.0702092
R21374 vss.n4690 vss.n4689 0.0702092
R21375 vss.n4691 vss.n4690 0.0702092
R21376 vss.n4699 vss.n4698 0.0702092
R21377 vss.n4698 vss.n4697 0.0702092
R21378 vss.n4680 vss.n4656 0.0702092
R21379 vss.n4681 vss.n4680 0.0702092
R21380 vss.n4683 vss.n4682 0.0702092
R21381 vss.n4682 vss.n4681 0.0702092
R21382 vss.n4696 vss.n4695 0.0702092
R21383 vss.n4697 vss.n4696 0.0702092
R21384 vss.n4693 vss.n4692 0.0702092
R21385 vss.n4692 vss.n4691 0.0702092
R21386 vss.n4594 vss.n4593 0.0702092
R21387 vss.n4595 vss.n4594 0.0702092
R21388 vss.n4598 vss.n4597 0.0702092
R21389 vss.n4604 vss.n4603 0.0702092
R21390 vss.n4603 vss.n4602 0.0702092
R21391 vss.n4584 vss.n4560 0.0702092
R21392 vss.n4585 vss.n4584 0.0702092
R21393 vss.n4582 vss.n4576 0.0702092
R21394 vss.n4582 vss.n4581 0.0702092
R21395 vss.n4580 vss.n4579 0.0702092
R21396 vss.n4581 vss.n4580 0.0702092
R21397 vss.n4587 vss.n4586 0.0702092
R21398 vss.n4586 vss.n4585 0.0702092
R21399 vss.n4601 vss.n4600 0.0702092
R21400 vss.n4602 vss.n4601 0.0702092
R21401 vss.n6851 vss.n6850 0.0702092
R21402 vss.n6852 vss.n6851 0.0702092
R21403 vss.n6858 vss.n6857 0.0702092
R21404 vss.n6857 vss.n6856 0.0702092
R21405 vss.n6871 vss.n6870 0.0702092
R21406 vss.n6872 vss.n6871 0.0702092
R21407 vss.n6868 vss.n6867 0.0702092
R21408 vss.n6867 vss.n6866 0.0702092
R21409 vss.n6865 vss.n6864 0.0702092
R21410 vss.n6866 vss.n6865 0.0702092
R21411 vss.n6874 vss.n6873 0.0702092
R21412 vss.n6873 vss.n6872 0.0702092
R21413 vss.n6855 vss.n6832 0.0702092
R21414 vss.n6856 vss.n6855 0.0702092
R21415 vss.n6853 vss.n6848 0.0702092
R21416 vss.n6853 vss.n6852 0.0702092
R21417 vss.n2623 vss.n2622 0.0702092
R21418 vss.n2622 vss.n2621 0.0702092
R21419 vss.n2626 vss.n2625 0.0702092
R21420 vss.n2627 vss.n2626 0.0702092
R21421 vss.n2637 vss.n2636 0.0702092
R21422 vss.n2636 vss.n2635 0.0702092
R21423 vss.n2639 vss.n2600 0.0702092
R21424 vss.n2600 vss.n2598 0.0702092
R21425 vss.n2601 vss.n2599 0.0702092
R21426 vss.n2599 vss.n2598 0.0702092
R21427 vss.n2634 vss.n2633 0.0702092
R21428 vss.n2635 vss.n2634 0.0702092
R21429 vss.n2628 vss.n2611 0.0702092
R21430 vss.n2628 vss.n2627 0.0702092
R21431 vss.n2620 vss.n2619 0.0702092
R21432 vss.n2621 vss.n2620 0.0702092
R21433 vss.n1941 vss.n1899 0.0702092
R21434 vss.n1899 vss.n1897 0.0702092
R21435 vss.n1939 vss.n1938 0.0702092
R21436 vss.n1938 vss.n1937 0.0702092
R21437 vss.n1929 vss.n1928 0.0702092
R21438 vss.n1930 vss.n1929 0.0702092
R21439 vss.n1926 vss.n1925 0.0702092
R21440 vss.n1925 vss.n1924 0.0702092
R21441 vss.n1923 vss.n1922 0.0702092
R21442 vss.n1924 vss.n1923 0.0702092
R21443 vss.n1932 vss.n1931 0.0702092
R21444 vss.n1931 vss.n1930 0.0702092
R21445 vss.n1936 vss.n1935 0.0702092
R21446 vss.n1937 vss.n1936 0.0702092
R21447 vss.n1900 vss.n1898 0.0702092
R21448 vss.n1898 vss.n1897 0.0702092
R21449 vss.n2858 vss.n2857 0.0702092
R21450 vss.n2859 vss.n2858 0.0702092
R21451 vss.n2865 vss.n2864 0.0702092
R21452 vss.n2864 vss.n2863 0.0702092
R21453 vss.n2878 vss.n2877 0.0702092
R21454 vss.n2879 vss.n2878 0.0702092
R21455 vss.n2875 vss.n2874 0.0702092
R21456 vss.n2874 vss.n2873 0.0702092
R21457 vss.n2872 vss.n2871 0.0702092
R21458 vss.n2873 vss.n2872 0.0702092
R21459 vss.n2881 vss.n2880 0.0702092
R21460 vss.n2880 vss.n2879 0.0702092
R21461 vss.n2862 vss.n2839 0.0702092
R21462 vss.n2863 vss.n2862 0.0702092
R21463 vss.n2860 vss.n2855 0.0702092
R21464 vss.n2860 vss.n2859 0.0702092
R21465 vss.n7642 vss.n7641 0.0702092
R21466 vss.n7643 vss.n7642 0.0702092
R21467 vss.n7649 vss.n7648 0.0702092
R21468 vss.n7648 vss.n7647 0.0702092
R21469 vss.n7662 vss.n7661 0.0702092
R21470 vss.n7663 vss.n7662 0.0702092
R21471 vss.n7659 vss.n7658 0.0702092
R21472 vss.n7658 vss.n7657 0.0702092
R21473 vss.n7656 vss.n7655 0.0702092
R21474 vss.n7657 vss.n7656 0.0702092
R21475 vss.n7665 vss.n7664 0.0702092
R21476 vss.n7664 vss.n7663 0.0702092
R21477 vss.n7646 vss.n7623 0.0702092
R21478 vss.n7647 vss.n7646 0.0702092
R21479 vss.n7644 vss.n7639 0.0702092
R21480 vss.n7644 vss.n7643 0.0702092
R21481 vss.n2812 vss.n2811 0.0702092
R21482 vss.n2813 vss.n2812 0.0702092
R21483 vss.n2819 vss.n2818 0.0702092
R21484 vss.n2818 vss.n2817 0.0702092
R21485 vss.n2832 vss.n2831 0.0702092
R21486 vss.n2833 vss.n2832 0.0702092
R21487 vss.n2829 vss.n2828 0.0702092
R21488 vss.n2828 vss.n2827 0.0702092
R21489 vss.n2826 vss.n2825 0.0702092
R21490 vss.n2827 vss.n2826 0.0702092
R21491 vss.n2835 vss.n2834 0.0702092
R21492 vss.n2834 vss.n2833 0.0702092
R21493 vss.n2816 vss.n2725 0.0702092
R21494 vss.n2817 vss.n2816 0.0702092
R21495 vss.n2814 vss.n2741 0.0702092
R21496 vss.n2814 vss.n2813 0.0702092
R21497 vss.n2950 vss.n2949 0.0702092
R21498 vss.n2951 vss.n2950 0.0702092
R21499 vss.n2957 vss.n2956 0.0702092
R21500 vss.n2956 vss.n2955 0.0702092
R21501 vss.n2971 vss.n2970 0.0702092
R21502 vss.n2972 vss.n2971 0.0702092
R21503 vss.n2968 vss.n2967 0.0702092
R21504 vss.n2967 vss.n2966 0.0702092
R21505 vss.n2965 vss.n2964 0.0702092
R21506 vss.n2966 vss.n2965 0.0702092
R21507 vss.n2974 vss.n2973 0.0702092
R21508 vss.n2973 vss.n2972 0.0702092
R21509 vss.n2954 vss.n2931 0.0702092
R21510 vss.n2955 vss.n2954 0.0702092
R21511 vss.n2952 vss.n2947 0.0702092
R21512 vss.n2952 vss.n2951 0.0702092
R21513 vss.n7012 vss.n7011 0.0702092
R21514 vss.n7011 vss.n7010 0.0702092
R21515 vss.n7015 vss.n7014 0.0702092
R21516 vss.n7016 vss.n7015 0.0702092
R21517 vss.n7026 vss.n7025 0.0702092
R21518 vss.n7025 vss.n7024 0.0702092
R21519 vss.n7028 vss.n6989 0.0702092
R21520 vss.n6989 vss.n6987 0.0702092
R21521 vss.n6990 vss.n6988 0.0702092
R21522 vss.n6988 vss.n6987 0.0702092
R21523 vss.n7023 vss.n7022 0.0702092
R21524 vss.n7024 vss.n7023 0.0702092
R21525 vss.n7017 vss.n7000 0.0702092
R21526 vss.n7017 vss.n7016 0.0702092
R21527 vss.n7009 vss.n7008 0.0702092
R21528 vss.n7010 vss.n7009 0.0702092
R21529 vss.n7151 vss.n7150 0.0702092
R21530 vss.n7150 vss.n7149 0.0702092
R21531 vss.n7154 vss.n7153 0.0702092
R21532 vss.n7155 vss.n7154 0.0702092
R21533 vss.n7164 vss.n7163 0.0702092
R21534 vss.n7163 vss.n7162 0.0702092
R21535 vss.n7166 vss.n7126 0.0702092
R21536 vss.n7126 vss.n7124 0.0702092
R21537 vss.n7127 vss.n7125 0.0702092
R21538 vss.n7125 vss.n7124 0.0702092
R21539 vss.n7161 vss.n7160 0.0702092
R21540 vss.n7162 vss.n7161 0.0702092
R21541 vss.n7157 vss.n7156 0.0702092
R21542 vss.n7156 vss.n7155 0.0702092
R21543 vss.n7148 vss.n7147 0.0702092
R21544 vss.n7149 vss.n7148 0.0702092
R21545 vss.n6967 vss.n6966 0.0702092
R21546 vss.n6966 vss.n6965 0.0702092
R21547 vss.n6970 vss.n6969 0.0702092
R21548 vss.n6971 vss.n6970 0.0702092
R21549 vss.n6981 vss.n6980 0.0702092
R21550 vss.n6980 vss.n6979 0.0702092
R21551 vss.n6983 vss.n6922 0.0702092
R21552 vss.n6922 vss.n6920 0.0702092
R21553 vss.n6923 vss.n6921 0.0702092
R21554 vss.n6921 vss.n6920 0.0702092
R21555 vss.n6978 vss.n6977 0.0702092
R21556 vss.n6979 vss.n6978 0.0702092
R21557 vss.n6973 vss.n6972 0.0702092
R21558 vss.n6972 vss.n6971 0.0702092
R21559 vss.n6964 vss.n6963 0.0702092
R21560 vss.n6965 vss.n6964 0.0702092
R21561 vss.n7594 vss.n7593 0.0702092
R21562 vss.n7595 vss.n7594 0.0702092
R21563 vss.n7601 vss.n7600 0.0702092
R21564 vss.n7600 vss.n7599 0.0702092
R21565 vss.n7614 vss.n7613 0.0702092
R21566 vss.n7615 vss.n7614 0.0702092
R21567 vss.n7611 vss.n7610 0.0702092
R21568 vss.n7610 vss.n7609 0.0702092
R21569 vss.n7608 vss.n7607 0.0702092
R21570 vss.n7609 vss.n7608 0.0702092
R21571 vss.n7617 vss.n7616 0.0702092
R21572 vss.n7616 vss.n7615 0.0702092
R21573 vss.n7598 vss.n7507 0.0702092
R21574 vss.n7599 vss.n7598 0.0702092
R21575 vss.n7596 vss.n7523 0.0702092
R21576 vss.n7596 vss.n7595 0.0702092
R21577 vss.n7789 vss.n7788 0.0702092
R21578 vss.n7790 vss.n7789 0.0702092
R21579 vss.n7796 vss.n7795 0.0702092
R21580 vss.n7795 vss.n7794 0.0702092
R21581 vss.n7809 vss.n7808 0.0702092
R21582 vss.n7810 vss.n7809 0.0702092
R21583 vss.n7806 vss.n7805 0.0702092
R21584 vss.n7805 vss.n7804 0.0702092
R21585 vss.n7803 vss.n7802 0.0702092
R21586 vss.n7804 vss.n7803 0.0702092
R21587 vss.n7812 vss.n7811 0.0702092
R21588 vss.n7811 vss.n7810 0.0702092
R21589 vss.n7793 vss.n7770 0.0702092
R21590 vss.n7794 vss.n7793 0.0702092
R21591 vss.n7791 vss.n7786 0.0702092
R21592 vss.n7791 vss.n7790 0.0702092
R21593 vss.n7837 vss.n7836 0.0702092
R21594 vss.n7838 vss.n7837 0.0702092
R21595 vss.n7844 vss.n7843 0.0702092
R21596 vss.n7843 vss.n7842 0.0702092
R21597 vss.n7857 vss.n7856 0.0702092
R21598 vss.n7858 vss.n7857 0.0702092
R21599 vss.n7854 vss.n7853 0.0702092
R21600 vss.n7853 vss.n7852 0.0702092
R21601 vss.n7851 vss.n7850 0.0702092
R21602 vss.n7852 vss.n7851 0.0702092
R21603 vss.n7860 vss.n7859 0.0702092
R21604 vss.n7859 vss.n7858 0.0702092
R21605 vss.n7841 vss.n7818 0.0702092
R21606 vss.n7842 vss.n7841 0.0702092
R21607 vss.n7839 vss.n7834 0.0702092
R21608 vss.n7839 vss.n7838 0.0702092
R21609 vss.n2579 vss.n2578 0.0702092
R21610 vss.n2578 vss.n2577 0.0702092
R21611 vss.n2582 vss.n2581 0.0702092
R21612 vss.n2583 vss.n2582 0.0702092
R21613 vss.n2592 vss.n2591 0.0702092
R21614 vss.n2591 vss.n2590 0.0702092
R21615 vss.n2594 vss.n2485 0.0702092
R21616 vss.n2485 vss.n2483 0.0702092
R21617 vss.n2486 vss.n2484 0.0702092
R21618 vss.n2484 vss.n2483 0.0702092
R21619 vss.n2589 vss.n2588 0.0702092
R21620 vss.n2590 vss.n2589 0.0702092
R21621 vss.n2585 vss.n2584 0.0702092
R21622 vss.n2584 vss.n2583 0.0702092
R21623 vss.n2576 vss.n2575 0.0702092
R21624 vss.n2577 vss.n2576 0.0702092
R21625 vss.n1157 vss.n1156 0.0702092
R21626 vss.n14872 vss.n1157 0.0702092
R21627 vss.n14880 vss.n14879 0.0702092
R21628 vss.n14879 vss.n14878 0.0702092
R21629 vss.n7935 vss.n1142 0.0702092
R21630 vss.n7936 vss.n7935 0.0702092
R21631 vss.n7937 vss.n7934 0.0702092
R21632 vss.n7937 vss.n7936 0.0702092
R21633 vss.n14877 vss.n14876 0.0702092
R21634 vss.n14878 vss.n14877 0.0702092
R21635 vss.n14874 vss.n14873 0.0702092
R21636 vss.n14873 vss.n14872 0.0702092
R21637 vss.n7943 vss.n7942 0.0702092
R21638 vss.n7944 vss.n7943 0.0702092
R21639 vss.n7933 vss.n7932 0.0702092
R21640 vss.n2678 vss.n2659 0.0702092
R21641 vss.n2659 vss.n2655 0.0702092
R21642 vss.n2658 vss.n2654 0.0702092
R21643 vss.n7918 vss.n2654 0.0702092
R21644 vss.n2646 vss.n2644 0.0702092
R21645 vss.n2644 vss.n2643 0.0702092
R21646 vss.n7922 vss.n2645 0.0702092
R21647 vss.n2645 vss.n2643 0.0702092
R21648 vss.n7920 vss.n7919 0.0702092
R21649 vss.n7919 vss.n7918 0.0702092
R21650 vss.n2668 vss.n2667 0.0702092
R21651 vss.n2667 vss.n2655 0.0702092
R21652 vss.n2676 vss.n2675 0.0702092
R21653 vss.n2675 vss.n2674 0.0702092
R21654 vss.n2671 vss.n2670 0.0702092
R21655 vss.n7900 vss.n7899 0.0702092
R21656 vss.n7902 vss.n7900 0.0702092
R21657 vss.n7910 vss.n7909 0.0702092
R21658 vss.n7909 vss.n7908 0.0702092
R21659 vss.n7890 vss.n7866 0.0702092
R21660 vss.n7891 vss.n7890 0.0702092
R21661 vss.n7893 vss.n7892 0.0702092
R21662 vss.n7892 vss.n7891 0.0702092
R21663 vss.n7907 vss.n7906 0.0702092
R21664 vss.n7908 vss.n7907 0.0702092
R21665 vss.n7904 vss.n7903 0.0702092
R21666 vss.n7903 vss.n7902 0.0702092
R21667 vss.n7888 vss.n7882 0.0702092
R21668 vss.n7888 vss.n7887 0.0702092
R21669 vss.n7885 vss.n7884 0.0702092
R21670 vss.n2721 vss.n2720 0.0702092
R21671 vss.n2720 vss.n2719 0.0702092
R21672 vss.n2703 vss.n2680 0.0702092
R21673 vss.n2704 vss.n2703 0.0702092
R21674 vss.n2701 vss.n2696 0.0702092
R21675 vss.n2701 vss.n2700 0.0702092
R21676 vss.n2699 vss.n2698 0.0702092
R21677 vss.n2700 vss.n2699 0.0702092
R21678 vss.n2706 vss.n2705 0.0702092
R21679 vss.n2705 vss.n2704 0.0702092
R21680 vss.n2718 vss.n2717 0.0702092
R21681 vss.n2719 vss.n2718 0.0702092
R21682 vss.n2711 vss.n2710 0.0702092
R21683 vss.n2710 vss.n985 0.0702092
R21684 vss.n2715 vss.n2714 0.0702092
R21685 vss.n7754 vss.n7753 0.0702092
R21686 vss.n7755 vss.n7754 0.0702092
R21687 vss.n7763 vss.n7762 0.0702092
R21688 vss.n7762 vss.n7761 0.0702092
R21689 vss.n7744 vss.n7720 0.0702092
R21690 vss.n7745 vss.n7744 0.0702092
R21691 vss.n7747 vss.n7746 0.0702092
R21692 vss.n7746 vss.n7745 0.0702092
R21693 vss.n7760 vss.n7759 0.0702092
R21694 vss.n7761 vss.n7760 0.0702092
R21695 vss.n7757 vss.n7756 0.0702092
R21696 vss.n7756 vss.n7755 0.0702092
R21697 vss.n7742 vss.n7736 0.0702092
R21698 vss.n7742 vss.n7741 0.0702092
R21699 vss.n7739 vss.n7738 0.0702092
R21700 vss.n2928 vss.n2885 0.0702092
R21701 vss.n2916 vss.n2885 0.0702092
R21702 vss.n2912 vss.n2884 0.0702092
R21703 vss.n2912 vss.n2895 0.0702092
R21704 vss.n2910 vss.n2898 0.0702092
R21705 vss.n2910 vss.n2909 0.0702092
R21706 vss.n2908 vss.n2907 0.0702092
R21707 vss.n2909 vss.n2908 0.0702092
R21708 vss.n2905 vss.n2904 0.0702092
R21709 vss.n2904 vss.n2895 0.0702092
R21710 vss.n2918 vss.n2917 0.0702092
R21711 vss.n2917 vss.n2916 0.0702092
R21712 vss.n2926 vss.n2925 0.0702092
R21713 vss.n2925 vss.n2924 0.0702092
R21714 vss.n2921 vss.n2920 0.0702092
R21715 vss.n7705 vss.n7704 0.0702092
R21716 vss.n7707 vss.n7705 0.0702092
R21717 vss.n7715 vss.n7714 0.0702092
R21718 vss.n7714 vss.n7713 0.0702092
R21719 vss.n7695 vss.n7671 0.0702092
R21720 vss.n7696 vss.n7695 0.0702092
R21721 vss.n7698 vss.n7697 0.0702092
R21722 vss.n7697 vss.n7696 0.0702092
R21723 vss.n7712 vss.n7711 0.0702092
R21724 vss.n7713 vss.n7712 0.0702092
R21725 vss.n7709 vss.n7708 0.0702092
R21726 vss.n7708 vss.n7707 0.0702092
R21727 vss.n7693 vss.n7687 0.0702092
R21728 vss.n7693 vss.n7692 0.0702092
R21729 vss.n7690 vss.n7689 0.0702092
R21730 vss.n3046 vss.n3045 0.0702092
R21731 vss.n3051 vss.n3046 0.0702092
R21732 vss.n3042 vss.n3041 0.0702092
R21733 vss.n3041 vss.n3040 0.0702092
R21734 vss.n3033 vss.n3032 0.0702092
R21735 vss.n3034 vss.n3033 0.0702092
R21736 vss.n3036 vss.n3035 0.0702092
R21737 vss.n3035 vss.n3034 0.0702092
R21738 vss.n3039 vss.n3038 0.0702092
R21739 vss.n3040 vss.n3039 0.0702092
R21740 vss.n3053 vss.n3052 0.0702092
R21741 vss.n3052 vss.n3051 0.0702092
R21742 vss.n3015 vss.n3013 0.0702092
R21743 vss.n3013 vss.n3012 0.0702092
R21744 vss.n3055 vss.n3014 0.0702092
R21745 vss.n3011 vss.n3010 0.0702092
R21746 vss.n7491 vss.n3011 0.0702092
R21747 vss.n7499 vss.n7498 0.0702092
R21748 vss.n7498 vss.n7497 0.0702092
R21749 vss.n3001 vss.n2977 0.0702092
R21750 vss.n3002 vss.n3001 0.0702092
R21751 vss.n3004 vss.n3003 0.0702092
R21752 vss.n3003 vss.n3002 0.0702092
R21753 vss.n7496 vss.n7495 0.0702092
R21754 vss.n7497 vss.n7496 0.0702092
R21755 vss.n7493 vss.n7492 0.0702092
R21756 vss.n7492 vss.n7491 0.0702092
R21757 vss.n2999 vss.n2993 0.0702092
R21758 vss.n2999 vss.n2998 0.0702092
R21759 vss.n2996 vss.n2995 0.0702092
R21760 vss.n7989 vss.n2454 0.0702092
R21761 vss.n7977 vss.n2454 0.0702092
R21762 vss.n7973 vss.n2453 0.0702092
R21763 vss.n7973 vss.n2465 0.0702092
R21764 vss.n7971 vss.n2468 0.0702092
R21765 vss.n7971 vss.n7970 0.0702092
R21766 vss.n7969 vss.n7968 0.0702092
R21767 vss.n7970 vss.n7969 0.0702092
R21768 vss.n7966 vss.n7965 0.0702092
R21769 vss.n7965 vss.n2465 0.0702092
R21770 vss.n7979 vss.n7978 0.0702092
R21771 vss.n7978 vss.n7977 0.0702092
R21772 vss.n7987 vss.n7986 0.0702092
R21773 vss.n7986 vss.n7985 0.0702092
R21774 vss.n7982 vss.n7981 0.0702092
R21775 vss.n7105 vss.n7099 0.0702092
R21776 vss.n7099 vss.n7096 0.0702092
R21777 vss.n7098 vss.n7095 0.0702092
R21778 vss.n7110 vss.n7095 0.0702092
R21779 vss.n7118 vss.n7117 0.0702092
R21780 vss.n7117 vss.n7116 0.0702092
R21781 vss.n7115 vss.n7114 0.0702092
R21782 vss.n7116 vss.n7115 0.0702092
R21783 vss.n7112 vss.n7111 0.0702092
R21784 vss.n7111 vss.n7110 0.0702092
R21785 vss.n7101 vss.n7100 0.0702092
R21786 vss.n7101 vss.n7096 0.0702092
R21787 vss.n7121 vss.n7120 0.0702092
R21788 vss.n7122 vss.n7121 0.0702092
R21789 vss.n7089 vss.n7088 0.0702092
R21790 vss.n7064 vss.n7063 0.0702092
R21791 vss.n7063 vss.n7044 0.0702092
R21792 vss.n7047 vss.n7043 0.0702092
R21793 vss.n7069 vss.n7043 0.0702092
R21794 vss.n7035 vss.n7033 0.0702092
R21795 vss.n7033 vss.n7032 0.0702092
R21796 vss.n7073 vss.n7034 0.0702092
R21797 vss.n7034 vss.n7032 0.0702092
R21798 vss.n7071 vss.n7070 0.0702092
R21799 vss.n7070 vss.n7069 0.0702092
R21800 vss.n7053 vss.n7052 0.0702092
R21801 vss.n7052 vss.n7044 0.0702092
R21802 vss.n7055 vss.n7049 0.0702092
R21803 vss.n7049 vss.n3129 0.0702092
R21804 vss.n7058 vss.n7057 0.0702092
R21805 vss.n6901 vss.n6900 0.0702092
R21806 vss.n6900 vss.n6893 0.0702092
R21807 vss.n6895 vss.n6892 0.0702092
R21808 vss.n6906 vss.n6892 0.0702092
R21809 vss.n6914 vss.n6913 0.0702092
R21810 vss.n6913 vss.n6912 0.0702092
R21811 vss.n6911 vss.n6910 0.0702092
R21812 vss.n6912 vss.n6911 0.0702092
R21813 vss.n6908 vss.n6907 0.0702092
R21814 vss.n6907 vss.n6906 0.0702092
R21815 vss.n6898 vss.n6897 0.0702092
R21816 vss.n6898 vss.n6893 0.0702092
R21817 vss.n6917 vss.n6916 0.0702092
R21818 vss.n6918 vss.n6917 0.0702092
R21819 vss.n6886 vss.n6885 0.0702092
R21820 vss.n7210 vss.n7209 0.0702092
R21821 vss.n7212 vss.n7210 0.0702092
R21822 vss.n6816 vss.n3148 0.0702092
R21823 vss.n6817 vss.n6816 0.0702092
R21824 vss.n6808 vss.n6806 0.0702092
R21825 vss.n6806 vss.n6805 0.0702092
R21826 vss.n6821 vss.n6807 0.0702092
R21827 vss.n6807 vss.n6805 0.0702092
R21828 vss.n6819 vss.n6818 0.0702092
R21829 vss.n6818 vss.n6817 0.0702092
R21830 vss.n7213 vss.n3143 0.0702092
R21831 vss.n7213 vss.n7212 0.0702092
R21832 vss.n7220 vss.n7219 0.0702092
R21833 vss.n7221 vss.n7220 0.0702092
R21834 vss.n7217 vss.n7216 0.0702092
R21835 vss.n7181 vss.n7180 0.0702092
R21836 vss.n7182 vss.n7181 0.0702092
R21837 vss.n7188 vss.n7187 0.0702092
R21838 vss.n7187 vss.n7186 0.0702092
R21839 vss.n7201 vss.n7200 0.0702092
R21840 vss.n7202 vss.n7201 0.0702092
R21841 vss.n7198 vss.n7197 0.0702092
R21842 vss.n7197 vss.n7196 0.0702092
R21843 vss.n7195 vss.n7194 0.0702092
R21844 vss.n7196 vss.n7195 0.0702092
R21845 vss.n7204 vss.n7203 0.0702092
R21846 vss.n7203 vss.n7202 0.0702092
R21847 vss.n7185 vss.n3151 0.0702092
R21848 vss.n7186 vss.n7185 0.0702092
R21849 vss.n7183 vss.n3167 0.0702092
R21850 vss.n7183 vss.n7182 0.0702092
R21851 vss.n3206 vss.n3193 0.0702092
R21852 vss.n3193 vss.n3191 0.0702092
R21853 vss.n3204 vss.n3203 0.0702092
R21854 vss.n3203 vss.n3202 0.0702092
R21855 vss.n6798 vss.n6797 0.0702092
R21856 vss.n6797 vss.n6796 0.0702092
R21857 vss.n6800 vss.n3171 0.0702092
R21858 vss.n3171 vss.n3169 0.0702092
R21859 vss.n3172 vss.n3170 0.0702092
R21860 vss.n3170 vss.n3169 0.0702092
R21861 vss.n6795 vss.n6794 0.0702092
R21862 vss.n6796 vss.n6795 0.0702092
R21863 vss.n3201 vss.n3184 0.0702092
R21864 vss.n3202 vss.n3201 0.0702092
R21865 vss.n3194 vss.n3192 0.0702092
R21866 vss.n3192 vss.n3191 0.0702092
R21867 vss.n6779 vss.n6778 0.0702092
R21868 vss.n6780 vss.n6779 0.0702092
R21869 vss.n6788 vss.n6787 0.0702092
R21870 vss.n6787 vss.n6786 0.0702092
R21871 vss.n6769 vss.n6746 0.0702092
R21872 vss.n6770 vss.n6769 0.0702092
R21873 vss.n6767 vss.n6762 0.0702092
R21874 vss.n6767 vss.n6766 0.0702092
R21875 vss.n6765 vss.n6764 0.0702092
R21876 vss.n6766 vss.n6765 0.0702092
R21877 vss.n6772 vss.n6771 0.0702092
R21878 vss.n6771 vss.n6770 0.0702092
R21879 vss.n6785 vss.n6784 0.0702092
R21880 vss.n6786 vss.n6785 0.0702092
R21881 vss.n6782 vss.n6781 0.0702092
R21882 vss.n6781 vss.n6780 0.0702092
R21883 vss.n14828 vss.n14827 0.0702092
R21884 vss.n14827 vss.n14826 0.0702092
R21885 vss.n14831 vss.n14830 0.0702092
R21886 vss.n14832 vss.n14831 0.0702092
R21887 vss.n14825 vss.n14824 0.0702092
R21888 vss.n14826 vss.n14825 0.0702092
R21889 vss.n14834 vss.n14833 0.0702092
R21890 vss.n14833 vss.n14832 0.0702092
R21891 vss.n1840 vss.n1839 0.0702092
R21892 vss.n1841 vss.n1840 0.0702092
R21893 vss.n1847 vss.n1846 0.0702092
R21894 vss.n1846 vss.n1845 0.0702092
R21895 vss.n14349 vss.n14348 0.0702092
R21896 vss.n14350 vss.n14349 0.0702092
R21897 vss.n14346 vss.n14345 0.0702092
R21898 vss.n14345 vss.n14344 0.0702092
R21899 vss.n14343 vss.n14342 0.0702092
R21900 vss.n14344 vss.n14343 0.0702092
R21901 vss.n14352 vss.n14351 0.0702092
R21902 vss.n14351 vss.n14350 0.0702092
R21903 vss.n1844 vss.n1821 0.0702092
R21904 vss.n1845 vss.n1844 0.0702092
R21905 vss.n1842 vss.n1837 0.0702092
R21906 vss.n1842 vss.n1841 0.0702092
R21907 vss.n14219 vss.n14194 0.0702092
R21908 vss.n14220 vss.n14219 0.0702092
R21909 vss.n14229 vss.n14228 0.0702092
R21910 vss.n14230 vss.n14229 0.0702092
R21911 vss.n14238 vss.n14237 0.0702092
R21912 vss.n14237 vss.n14236 0.0702092
R21913 vss.n14222 vss.n14221 0.0702092
R21914 vss.n14221 vss.n14220 0.0702092
R21915 vss.n14235 vss.n14234 0.0702092
R21916 vss.n14236 vss.n14235 0.0702092
R21917 vss.n14232 vss.n14231 0.0702092
R21918 vss.n14231 vss.n14230 0.0702092
R21919 vss.n14217 vss.n14210 0.0702092
R21920 vss.n14217 vss.n14216 0.0702092
R21921 vss.n14213 vss.n14212 0.0702092
R21922 vss.n1302 vss.n1301 0.0702092
R21923 vss.n1303 vss.n1302 0.0702092
R21924 vss.n1309 vss.n1308 0.0702092
R21925 vss.n1308 vss.n1307 0.0702092
R21926 vss.n14743 vss.n14742 0.0702092
R21927 vss.n14744 vss.n14743 0.0702092
R21928 vss.n14740 vss.n14739 0.0702092
R21929 vss.n14739 vss.n14738 0.0702092
R21930 vss.n14737 vss.n14736 0.0702092
R21931 vss.n14738 vss.n14737 0.0702092
R21932 vss.n14746 vss.n14745 0.0702092
R21933 vss.n14745 vss.n14744 0.0702092
R21934 vss.n1306 vss.n1283 0.0702092
R21935 vss.n1307 vss.n1306 0.0702092
R21936 vss.n1304 vss.n1299 0.0702092
R21937 vss.n1304 vss.n1303 0.0702092
R21938 vss.n14001 vss.n14000 0.0702092
R21939 vss.n14002 vss.n14001 0.0702092
R21940 vss.n14008 vss.n14007 0.0702092
R21941 vss.n14007 vss.n14006 0.0702092
R21942 vss.n14021 vss.n14020 0.0702092
R21943 vss.n14022 vss.n14021 0.0702092
R21944 vss.n14018 vss.n14017 0.0702092
R21945 vss.n14017 vss.n14016 0.0702092
R21946 vss.n14015 vss.n14014 0.0702092
R21947 vss.n14016 vss.n14015 0.0702092
R21948 vss.n14024 vss.n14023 0.0702092
R21949 vss.n14023 vss.n14022 0.0702092
R21950 vss.n14005 vss.n13982 0.0702092
R21951 vss.n14006 vss.n14005 0.0702092
R21952 vss.n14003 vss.n13998 0.0702092
R21953 vss.n14003 vss.n14002 0.0702092
R21954 vss.n1507 vss.n1506 0.0702092
R21955 vss.n1508 vss.n1507 0.0702092
R21956 vss.n1514 vss.n1513 0.0702092
R21957 vss.n1513 vss.n1512 0.0702092
R21958 vss.n14670 vss.n14669 0.0702092
R21959 vss.n14671 vss.n14670 0.0702092
R21960 vss.n14667 vss.n14666 0.0702092
R21961 vss.n14666 vss.n14665 0.0702092
R21962 vss.n14664 vss.n14663 0.0702092
R21963 vss.n14665 vss.n14664 0.0702092
R21964 vss.n14673 vss.n14672 0.0702092
R21965 vss.n14672 vss.n14671 0.0702092
R21966 vss.n1511 vss.n1488 0.0702092
R21967 vss.n1512 vss.n1511 0.0702092
R21968 vss.n1509 vss.n1504 0.0702092
R21969 vss.n1509 vss.n1508 0.0702092
R21970 vss.n1560 vss.n1559 0.0702092
R21971 vss.n1561 vss.n1560 0.0702092
R21972 vss.n1567 vss.n1566 0.0702092
R21973 vss.n1566 vss.n1565 0.0702092
R21974 vss.n14593 vss.n14592 0.0702092
R21975 vss.n14594 vss.n14593 0.0702092
R21976 vss.n14590 vss.n14589 0.0702092
R21977 vss.n14589 vss.n14588 0.0702092
R21978 vss.n14587 vss.n14586 0.0702092
R21979 vss.n14588 vss.n14587 0.0702092
R21980 vss.n14596 vss.n14595 0.0702092
R21981 vss.n14595 vss.n14594 0.0702092
R21982 vss.n1564 vss.n1541 0.0702092
R21983 vss.n1565 vss.n1564 0.0702092
R21984 vss.n1562 vss.n1557 0.0702092
R21985 vss.n1562 vss.n1561 0.0702092
R21986 vss.n14500 vss.n14499 0.0702092
R21987 vss.n14501 vss.n14500 0.0702092
R21988 vss.n14507 vss.n14506 0.0702092
R21989 vss.n14506 vss.n14505 0.0702092
R21990 vss.n14520 vss.n14519 0.0702092
R21991 vss.n14521 vss.n14520 0.0702092
R21992 vss.n14517 vss.n14516 0.0702092
R21993 vss.n14516 vss.n14515 0.0702092
R21994 vss.n14514 vss.n14513 0.0702092
R21995 vss.n14515 vss.n14514 0.0702092
R21996 vss.n14523 vss.n14522 0.0702092
R21997 vss.n14522 vss.n14521 0.0702092
R21998 vss.n14504 vss.n14481 0.0702092
R21999 vss.n14505 vss.n14504 0.0702092
R22000 vss.n14502 vss.n14497 0.0702092
R22001 vss.n14502 vss.n14501 0.0702092
R22002 vss.n1717 vss.n1716 0.0702092
R22003 vss.n1718 vss.n1717 0.0702092
R22004 vss.n1724 vss.n1723 0.0702092
R22005 vss.n1723 vss.n1722 0.0702092
R22006 vss.n1738 vss.n1737 0.0702092
R22007 vss.n1739 vss.n1738 0.0702092
R22008 vss.n1735 vss.n1734 0.0702092
R22009 vss.n1734 vss.n1733 0.0702092
R22010 vss.n1732 vss.n1731 0.0702092
R22011 vss.n1733 vss.n1732 0.0702092
R22012 vss.n1741 vss.n1740 0.0702092
R22013 vss.n1740 vss.n1739 0.0702092
R22014 vss.n1721 vss.n1698 0.0702092
R22015 vss.n1722 vss.n1721 0.0702092
R22016 vss.n1719 vss.n1714 0.0702092
R22017 vss.n1719 vss.n1718 0.0702092
R22018 vss.n1608 vss.n1607 0.0702092
R22019 vss.n1609 vss.n1608 0.0702092
R22020 vss.n1617 vss.n1616 0.0702092
R22021 vss.n1616 vss.n1615 0.0702092
R22022 vss.n1621 vss.n1620 0.0702092
R22023 vss.n1622 vss.n1621 0.0702092
R22024 vss.n1587 vss.n1585 0.0702092
R22025 vss.n1585 vss.n1584 0.0702092
R22026 vss.n1626 vss.n1586 0.0702092
R22027 vss.n1586 vss.n1584 0.0702092
R22028 vss.n1624 vss.n1623 0.0702092
R22029 vss.n1623 vss.n1622 0.0702092
R22030 vss.n1614 vss.n1613 0.0702092
R22031 vss.n1615 vss.n1614 0.0702092
R22032 vss.n1611 vss.n1610 0.0702092
R22033 vss.n1610 vss.n1609 0.0702092
R22034 vss.n14442 vss.n14441 0.0702092
R22035 vss.n14441 vss.n14440 0.0702092
R22036 vss.n14430 vss.n14429 0.0702092
R22037 vss.n14429 vss.n14428 0.0702092
R22038 vss.n14433 vss.n14432 0.0702092
R22039 vss.n14434 vss.n14433 0.0702092
R22040 vss.n14439 vss.n14438 0.0702092
R22041 vss.n14440 vss.n14439 0.0702092
R22042 vss.n14436 vss.n14435 0.0702092
R22043 vss.n14435 vss.n14434 0.0702092
R22044 vss.n14427 vss.n14426 0.0702092
R22045 vss.n14428 vss.n14427 0.0702092
R22046 vss.n13918 vss.n13907 0.0702092
R22047 vss.n13951 vss.n13907 0.0702092
R22048 vss.n13944 vss.n13943 0.0702092
R22049 vss.n13945 vss.n13944 0.0702092
R22050 vss.n13941 vss.n13940 0.0702092
R22051 vss.n13940 vss.n13939 0.0702092
R22052 vss.n13931 vss.n13930 0.0702092
R22053 vss.n13935 vss.n13934 0.0702092
R22054 vss.n13934 vss.n13933 0.0702092
R22055 vss.n13938 vss.n13937 0.0702092
R22056 vss.n13939 vss.n13938 0.0702092
R22057 vss.n13947 vss.n13946 0.0702092
R22058 vss.n13946 vss.n13945 0.0702092
R22059 vss.n13950 vss.n13949 0.0702092
R22060 vss.n13951 vss.n13950 0.0702092
R22061 vss.n14620 vss.n14619 0.0702092
R22062 vss.n14621 vss.n14620 0.0702092
R22063 vss.n14627 vss.n14626 0.0702092
R22064 vss.n14626 vss.n14625 0.0702092
R22065 vss.n14641 vss.n14640 0.0702092
R22066 vss.n14642 vss.n14641 0.0702092
R22067 vss.n14638 vss.n14637 0.0702092
R22068 vss.n14637 vss.n14636 0.0702092
R22069 vss.n14635 vss.n14634 0.0702092
R22070 vss.n14636 vss.n14635 0.0702092
R22071 vss.n14644 vss.n14643 0.0702092
R22072 vss.n14643 vss.n14642 0.0702092
R22073 vss.n14624 vss.n14601 0.0702092
R22074 vss.n14625 vss.n14624 0.0702092
R22075 vss.n14622 vss.n14617 0.0702092
R22076 vss.n14622 vss.n14621 0.0702092
R22077 vss.n1460 vss.n1459 0.0702092
R22078 vss.n1461 vss.n1460 0.0702092
R22079 vss.n1467 vss.n1466 0.0702092
R22080 vss.n1466 vss.n1465 0.0702092
R22081 vss.n1481 vss.n1480 0.0702092
R22082 vss.n1482 vss.n1481 0.0702092
R22083 vss.n1478 vss.n1477 0.0702092
R22084 vss.n1477 vss.n1476 0.0702092
R22085 vss.n1475 vss.n1474 0.0702092
R22086 vss.n1476 vss.n1475 0.0702092
R22087 vss.n1484 vss.n1483 0.0702092
R22088 vss.n1483 vss.n1482 0.0702092
R22089 vss.n1464 vss.n1441 0.0702092
R22090 vss.n1465 vss.n1464 0.0702092
R22091 vss.n1462 vss.n1457 0.0702092
R22092 vss.n1462 vss.n1461 0.0702092
R22093 vss.n13903 vss.n13902 0.0702092
R22094 vss.n13904 vss.n13903 0.0702092
R22095 vss.n13872 vss.n13871 0.0702092
R22096 vss.n13888 vss.n13887 0.0702092
R22097 vss.n13887 vss.n13886 0.0702092
R22098 vss.n13891 vss.n13890 0.0702092
R22099 vss.n13892 vss.n13891 0.0702092
R22100 vss.n13900 vss.n13899 0.0702092
R22101 vss.n13899 vss.n13898 0.0702092
R22102 vss.n13897 vss.n13896 0.0702092
R22103 vss.n13898 vss.n13897 0.0702092
R22104 vss.n13894 vss.n13893 0.0702092
R22105 vss.n13893 vss.n13892 0.0702092
R22106 vss.n13885 vss.n13884 0.0702092
R22107 vss.n13886 vss.n13885 0.0702092
R22108 vss.n8204 vss.n8197 0.0702092
R22109 vss.n8200 vss.n8197 0.0702092
R22110 vss.n8199 vss.n8198 0.0702092
R22111 vss.n8207 vss.n8206 0.0702092
R22112 vss.n8208 vss.n8207 0.0702092
R22113 vss.n8216 vss.n8215 0.0702092
R22114 vss.n8215 vss.n8214 0.0702092
R22115 vss.n8218 vss.n8177 0.0702092
R22116 vss.n8177 vss.n8175 0.0702092
R22117 vss.n8178 vss.n8176 0.0702092
R22118 vss.n8176 vss.n8175 0.0702092
R22119 vss.n8213 vss.n8212 0.0702092
R22120 vss.n8214 vss.n8213 0.0702092
R22121 vss.n8210 vss.n8209 0.0702092
R22122 vss.n8209 vss.n8208 0.0702092
R22123 vss.n13957 vss.n8169 0.0702092
R22124 vss.n13957 vss.n13956 0.0702092
R22125 vss.n8172 vss.n8171 0.0702092
R22126 vss.n13969 vss.n13968 0.0702092
R22127 vss.n13970 vss.n13969 0.0702092
R22128 vss.n13978 vss.n13977 0.0702092
R22129 vss.n13977 vss.n13976 0.0702092
R22130 vss.n13959 vss.n8153 0.0702092
R22131 vss.n13960 vss.n13959 0.0702092
R22132 vss.n13962 vss.n13961 0.0702092
R22133 vss.n13961 vss.n13960 0.0702092
R22134 vss.n13975 vss.n13974 0.0702092
R22135 vss.n13976 vss.n13975 0.0702092
R22136 vss.n13972 vss.n13971 0.0702092
R22137 vss.n13971 vss.n13970 0.0702092
R22138 vss.n14035 vss.n8146 0.0702092
R22139 vss.n14068 vss.n8146 0.0702092
R22140 vss.n14061 vss.n14060 0.0702092
R22141 vss.n14062 vss.n14061 0.0702092
R22142 vss.n14058 vss.n14057 0.0702092
R22143 vss.n14057 vss.n14056 0.0702092
R22144 vss.n14048 vss.n14047 0.0702092
R22145 vss.n14052 vss.n14051 0.0702092
R22146 vss.n14051 vss.n14050 0.0702092
R22147 vss.n14055 vss.n14054 0.0702092
R22148 vss.n14056 vss.n14055 0.0702092
R22149 vss.n14064 vss.n14063 0.0702092
R22150 vss.n14063 vss.n14062 0.0702092
R22151 vss.n14067 vss.n14066 0.0702092
R22152 vss.n14068 vss.n14067 0.0702092
R22153 vss.n1351 vss.n1350 0.0702092
R22154 vss.n1352 vss.n1351 0.0702092
R22155 vss.n1360 vss.n1359 0.0702092
R22156 vss.n1359 vss.n1358 0.0702092
R22157 vss.n1364 vss.n1363 0.0702092
R22158 vss.n1365 vss.n1364 0.0702092
R22159 vss.n1329 vss.n1327 0.0702092
R22160 vss.n1327 vss.n1326 0.0702092
R22161 vss.n1369 vss.n1328 0.0702092
R22162 vss.n1328 vss.n1326 0.0702092
R22163 vss.n1367 vss.n1366 0.0702092
R22164 vss.n1366 vss.n1365 0.0702092
R22165 vss.n1357 vss.n1356 0.0702092
R22166 vss.n1358 vss.n1357 0.0702092
R22167 vss.n1354 vss.n1353 0.0702092
R22168 vss.n1353 vss.n1352 0.0702092
R22169 vss.n1252 vss.n1251 0.0702092
R22170 vss.n1253 vss.n1252 0.0702092
R22171 vss.n1259 vss.n1258 0.0702092
R22172 vss.n1258 vss.n1257 0.0702092
R22173 vss.n1273 vss.n1272 0.0702092
R22174 vss.n1274 vss.n1273 0.0702092
R22175 vss.n1270 vss.n1269 0.0702092
R22176 vss.n1269 vss.n1268 0.0702092
R22177 vss.n1267 vss.n1266 0.0702092
R22178 vss.n1268 vss.n1267 0.0702092
R22179 vss.n1276 vss.n1275 0.0702092
R22180 vss.n1275 vss.n1274 0.0702092
R22181 vss.n1256 vss.n1233 0.0702092
R22182 vss.n1257 vss.n1256 0.0702092
R22183 vss.n1254 vss.n1249 0.0702092
R22184 vss.n1254 vss.n1253 0.0702092
R22185 vss.n2345 vss.n2344 0.0702092
R22186 vss.n2346 vss.n2345 0.0702092
R22187 vss.n2352 vss.n2351 0.0702092
R22188 vss.n2351 vss.n2350 0.0702092
R22189 vss.n8042 vss.n8041 0.0702092
R22190 vss.n8043 vss.n8042 0.0702092
R22191 vss.n8039 vss.n8038 0.0702092
R22192 vss.n8038 vss.n8037 0.0702092
R22193 vss.n8036 vss.n8035 0.0702092
R22194 vss.n8037 vss.n8036 0.0702092
R22195 vss.n8045 vss.n8044 0.0702092
R22196 vss.n8044 vss.n8043 0.0702092
R22197 vss.n2349 vss.n2326 0.0702092
R22198 vss.n2350 vss.n2349 0.0702092
R22199 vss.n2347 vss.n2342 0.0702092
R22200 vss.n2347 vss.n2346 0.0702092
R22201 vss.n2393 vss.n2392 0.0702092
R22202 vss.n2394 vss.n2393 0.0702092
R22203 vss.n2402 vss.n2401 0.0702092
R22204 vss.n2401 vss.n2400 0.0702092
R22205 vss.n2406 vss.n2405 0.0702092
R22206 vss.n2407 vss.n2406 0.0702092
R22207 vss.n2372 vss.n2370 0.0702092
R22208 vss.n2370 vss.n2369 0.0702092
R22209 vss.n2411 vss.n2371 0.0702092
R22210 vss.n2371 vss.n2369 0.0702092
R22211 vss.n2409 vss.n2408 0.0702092
R22212 vss.n2408 vss.n2407 0.0702092
R22213 vss.n2399 vss.n2398 0.0702092
R22214 vss.n2400 vss.n2399 0.0702092
R22215 vss.n2396 vss.n2395 0.0702092
R22216 vss.n2395 vss.n2394 0.0702092
R22217 vss.n8142 vss.n8141 0.0702092
R22218 vss.n8143 vss.n8142 0.0702092
R22219 vss.n8111 vss.n8110 0.0702092
R22220 vss.n8127 vss.n8126 0.0702092
R22221 vss.n8126 vss.n8125 0.0702092
R22222 vss.n8130 vss.n8129 0.0702092
R22223 vss.n8131 vss.n8130 0.0702092
R22224 vss.n8139 vss.n8138 0.0702092
R22225 vss.n8138 vss.n8137 0.0702092
R22226 vss.n8136 vss.n8135 0.0702092
R22227 vss.n8137 vss.n8136 0.0702092
R22228 vss.n8133 vss.n8132 0.0702092
R22229 vss.n8132 vss.n8131 0.0702092
R22230 vss.n8124 vss.n8123 0.0702092
R22231 vss.n8125 vss.n8124 0.0702092
R22232 vss.n8076 vss.n8069 0.0702092
R22233 vss.n8072 vss.n8069 0.0702092
R22234 vss.n8071 vss.n8070 0.0702092
R22235 vss.n8079 vss.n8078 0.0702092
R22236 vss.n8080 vss.n8079 0.0702092
R22237 vss.n8088 vss.n8087 0.0702092
R22238 vss.n8087 vss.n8086 0.0702092
R22239 vss.n8090 vss.n2228 0.0702092
R22240 vss.n2228 vss.n2226 0.0702092
R22241 vss.n2229 vss.n2227 0.0702092
R22242 vss.n2227 vss.n2226 0.0702092
R22243 vss.n8085 vss.n8084 0.0702092
R22244 vss.n8086 vss.n8085 0.0702092
R22245 vss.n8082 vss.n8081 0.0702092
R22246 vss.n8081 vss.n8080 0.0702092
R22247 vss.n2254 vss.n2253 0.0702092
R22248 vss.n2254 vss.n2225 0.0702092
R22249 vss.n2249 vss.n2248 0.0702092
R22250 vss.n2266 vss.n2265 0.0702092
R22251 vss.n2267 vss.n2266 0.0702092
R22252 vss.n2275 vss.n2274 0.0702092
R22253 vss.n2274 vss.n2273 0.0702092
R22254 vss.n2256 vss.n2232 0.0702092
R22255 vss.n2257 vss.n2256 0.0702092
R22256 vss.n2259 vss.n2258 0.0702092
R22257 vss.n2258 vss.n2257 0.0702092
R22258 vss.n2272 vss.n2271 0.0702092
R22259 vss.n2273 vss.n2272 0.0702092
R22260 vss.n2269 vss.n2268 0.0702092
R22261 vss.n2268 vss.n2267 0.0702092
R22262 vss.n2312 vss.n2311 0.0702092
R22263 vss.n2313 vss.n2312 0.0702092
R22264 vss.n2316 vss.n2315 0.0702092
R22265 vss.n2322 vss.n2321 0.0702092
R22266 vss.n2321 vss.n2320 0.0702092
R22267 vss.n2302 vss.n2278 0.0702092
R22268 vss.n2303 vss.n2302 0.0702092
R22269 vss.n2300 vss.n2294 0.0702092
R22270 vss.n2300 vss.n2299 0.0702092
R22271 vss.n2298 vss.n2297 0.0702092
R22272 vss.n2299 vss.n2298 0.0702092
R22273 vss.n2305 vss.n2304 0.0702092
R22274 vss.n2304 vss.n2303 0.0702092
R22275 vss.n2319 vss.n2318 0.0702092
R22276 vss.n2320 vss.n2319 0.0702092
R22277 vss.n11959 vss.n11946 0.0702092
R22278 vss.n11946 vss.n11944 0.0702092
R22279 vss.n11957 vss.n11956 0.0702092
R22280 vss.n11956 vss.n11955 0.0702092
R22281 vss.n14133 vss.n14132 0.0702092
R22282 vss.n14134 vss.n14133 0.0702092
R22283 vss.n14130 vss.n14129 0.0702092
R22284 vss.n14129 vss.n14128 0.0702092
R22285 vss.n14127 vss.n14126 0.0702092
R22286 vss.n14128 vss.n14127 0.0702092
R22287 vss.n14136 vss.n14135 0.0702092
R22288 vss.n14135 vss.n14134 0.0702092
R22289 vss.n11954 vss.n2088 0.0702092
R22290 vss.n11955 vss.n11954 0.0702092
R22291 vss.n11947 vss.n11945 0.0702092
R22292 vss.n11945 vss.n11944 0.0702092
R22293 vss.n13487 vss.n13486 0.0702092
R22294 vss.n13488 vss.n13487 0.0702092
R22295 vss.n13494 vss.n13493 0.0702092
R22296 vss.n13493 vss.n13492 0.0702092
R22297 vss.n13507 vss.n13506 0.0702092
R22298 vss.n13508 vss.n13507 0.0702092
R22299 vss.n13504 vss.n13503 0.0702092
R22300 vss.n13503 vss.n13502 0.0702092
R22301 vss.n13501 vss.n13500 0.0702092
R22302 vss.n13502 vss.n13501 0.0702092
R22303 vss.n13510 vss.n13509 0.0702092
R22304 vss.n13509 vss.n13508 0.0702092
R22305 vss.n13491 vss.n13468 0.0702092
R22306 vss.n13492 vss.n13491 0.0702092
R22307 vss.n13489 vss.n13484 0.0702092
R22308 vss.n13489 vss.n13488 0.0702092
R22309 vss.n12057 vss.n12017 0.0702092
R22310 vss.n12017 vss.n12015 0.0702092
R22311 vss.n12055 vss.n12054 0.0702092
R22312 vss.n12054 vss.n12053 0.0702092
R22313 vss.n12046 vss.n12045 0.0702092
R22314 vss.n12047 vss.n12046 0.0702092
R22315 vss.n12043 vss.n12042 0.0702092
R22316 vss.n12042 vss.n12041 0.0702092
R22317 vss.n12040 vss.n12039 0.0702092
R22318 vss.n12041 vss.n12040 0.0702092
R22319 vss.n12049 vss.n12048 0.0702092
R22320 vss.n12048 vss.n12047 0.0702092
R22321 vss.n12052 vss.n12051 0.0702092
R22322 vss.n12053 vss.n12052 0.0702092
R22323 vss.n12018 vss.n12016 0.0702092
R22324 vss.n12016 vss.n12015 0.0702092
R22325 vss.n13719 vss.n13718 0.0702092
R22326 vss.n13720 vss.n13719 0.0702092
R22327 vss.n13726 vss.n13725 0.0702092
R22328 vss.n13725 vss.n13724 0.0702092
R22329 vss.n13739 vss.n13738 0.0702092
R22330 vss.n13740 vss.n13739 0.0702092
R22331 vss.n13736 vss.n13735 0.0702092
R22332 vss.n13735 vss.n13734 0.0702092
R22333 vss.n13733 vss.n13732 0.0702092
R22334 vss.n13734 vss.n13733 0.0702092
R22335 vss.n13742 vss.n13741 0.0702092
R22336 vss.n13741 vss.n13740 0.0702092
R22337 vss.n13723 vss.n8303 0.0702092
R22338 vss.n13724 vss.n13723 0.0702092
R22339 vss.n13721 vss.n8319 0.0702092
R22340 vss.n13721 vss.n13720 0.0702092
R22341 vss.n8483 vss.n8443 0.0702092
R22342 vss.n8443 vss.n8441 0.0702092
R22343 vss.n8481 vss.n8480 0.0702092
R22344 vss.n8480 vss.n8479 0.0702092
R22345 vss.n8472 vss.n8471 0.0702092
R22346 vss.n8473 vss.n8472 0.0702092
R22347 vss.n8469 vss.n8468 0.0702092
R22348 vss.n8468 vss.n8467 0.0702092
R22349 vss.n8466 vss.n8465 0.0702092
R22350 vss.n8467 vss.n8466 0.0702092
R22351 vss.n8475 vss.n8474 0.0702092
R22352 vss.n8474 vss.n8473 0.0702092
R22353 vss.n8478 vss.n8477 0.0702092
R22354 vss.n8479 vss.n8478 0.0702092
R22355 vss.n8444 vss.n8442 0.0702092
R22356 vss.n8442 vss.n8441 0.0702092
R22357 vss.n8560 vss.n8520 0.0702092
R22358 vss.n8520 vss.n8518 0.0702092
R22359 vss.n8558 vss.n8557 0.0702092
R22360 vss.n8557 vss.n8556 0.0702092
R22361 vss.n8549 vss.n8548 0.0702092
R22362 vss.n8550 vss.n8549 0.0702092
R22363 vss.n8546 vss.n8545 0.0702092
R22364 vss.n8545 vss.n8544 0.0702092
R22365 vss.n8543 vss.n8542 0.0702092
R22366 vss.n8544 vss.n8543 0.0702092
R22367 vss.n8552 vss.n8551 0.0702092
R22368 vss.n8551 vss.n8550 0.0702092
R22369 vss.n8555 vss.n8554 0.0702092
R22370 vss.n8556 vss.n8555 0.0702092
R22371 vss.n8521 vss.n8519 0.0702092
R22372 vss.n8519 vss.n8518 0.0702092
R22373 vss.n13007 vss.n13006 0.0702092
R22374 vss.n13008 vss.n13007 0.0702092
R22375 vss.n13014 vss.n13013 0.0702092
R22376 vss.n13013 vss.n13012 0.0702092
R22377 vss.n13027 vss.n13026 0.0702092
R22378 vss.n13028 vss.n13027 0.0702092
R22379 vss.n13024 vss.n13023 0.0702092
R22380 vss.n13023 vss.n13022 0.0702092
R22381 vss.n13021 vss.n13020 0.0702092
R22382 vss.n13022 vss.n13021 0.0702092
R22383 vss.n13030 vss.n13029 0.0702092
R22384 vss.n13029 vss.n13028 0.0702092
R22385 vss.n13011 vss.n9089 0.0702092
R22386 vss.n13012 vss.n13011 0.0702092
R22387 vss.n13009 vss.n9105 0.0702092
R22388 vss.n13009 vss.n13008 0.0702092
R22389 vss.n8972 vss.n8971 0.0702092
R22390 vss.n8973 vss.n8972 0.0702092
R22391 vss.n8979 vss.n8978 0.0702092
R22392 vss.n8978 vss.n8977 0.0702092
R22393 vss.n8992 vss.n8991 0.0702092
R22394 vss.n8993 vss.n8992 0.0702092
R22395 vss.n8989 vss.n8988 0.0702092
R22396 vss.n8988 vss.n8987 0.0702092
R22397 vss.n8986 vss.n8985 0.0702092
R22398 vss.n8987 vss.n8986 0.0702092
R22399 vss.n8995 vss.n8994 0.0702092
R22400 vss.n8994 vss.n8993 0.0702092
R22401 vss.n8976 vss.n8953 0.0702092
R22402 vss.n8977 vss.n8976 0.0702092
R22403 vss.n8974 vss.n8969 0.0702092
R22404 vss.n8974 vss.n8973 0.0702092
R22405 vss.n9155 vss.n9115 0.0702092
R22406 vss.n9115 vss.n9113 0.0702092
R22407 vss.n9153 vss.n9152 0.0702092
R22408 vss.n9152 vss.n9151 0.0702092
R22409 vss.n9144 vss.n9143 0.0702092
R22410 vss.n9145 vss.n9144 0.0702092
R22411 vss.n9141 vss.n9140 0.0702092
R22412 vss.n9140 vss.n9139 0.0702092
R22413 vss.n9138 vss.n9137 0.0702092
R22414 vss.n9139 vss.n9138 0.0702092
R22415 vss.n9147 vss.n9146 0.0702092
R22416 vss.n9146 vss.n9145 0.0702092
R22417 vss.n9150 vss.n9149 0.0702092
R22418 vss.n9151 vss.n9150 0.0702092
R22419 vss.n9116 vss.n9114 0.0702092
R22420 vss.n9114 vss.n9113 0.0702092
R22421 vss.n12635 vss.n12546 0.0702092
R22422 vss.n12546 vss.n12544 0.0702092
R22423 vss.n12633 vss.n12632 0.0702092
R22424 vss.n12632 vss.n12631 0.0702092
R22425 vss.n12575 vss.n12574 0.0702092
R22426 vss.n12576 vss.n12575 0.0702092
R22427 vss.n12572 vss.n12571 0.0702092
R22428 vss.n12571 vss.n12570 0.0702092
R22429 vss.n12569 vss.n12568 0.0702092
R22430 vss.n12570 vss.n12569 0.0702092
R22431 vss.n12578 vss.n12577 0.0702092
R22432 vss.n12577 vss.n12576 0.0702092
R22433 vss.n12630 vss.n12629 0.0702092
R22434 vss.n12631 vss.n12630 0.0702092
R22435 vss.n12547 vss.n12545 0.0702092
R22436 vss.n12545 vss.n12544 0.0702092
R22437 vss.n2057 vss.n2055 0.0702092
R22438 vss.n2055 vss.n2054 0.0702092
R22439 vss.n14144 vss.n14143 0.0702092
R22440 vss.n14148 vss.n14144 0.0702092
R22441 vss.n2086 vss.n2085 0.0702092
R22442 vss.n2085 vss.n2084 0.0702092
R22443 vss.n2083 vss.n2082 0.0702092
R22444 vss.n2084 vss.n2083 0.0702092
R22445 vss.n14150 vss.n14149 0.0702092
R22446 vss.n14149 vss.n14148 0.0702092
R22447 vss.n14152 vss.n2056 0.0702092
R22448 vss.n2056 vss.n2054 0.0702092
R22449 vss.n2076 vss.n2075 0.0702092
R22450 vss.n2077 vss.n2076 0.0702092
R22451 vss.n2080 vss.n2079 0.0702092
R22452 vss.n13602 vss.n13601 0.0702092
R22453 vss.n13601 vss.n13600 0.0702092
R22454 vss.n13581 vss.n13557 0.0702092
R22455 vss.n13582 vss.n13581 0.0702092
R22456 vss.n13579 vss.n13573 0.0702092
R22457 vss.n13579 vss.n13578 0.0702092
R22458 vss.n13577 vss.n13576 0.0702092
R22459 vss.n13578 vss.n13577 0.0702092
R22460 vss.n13584 vss.n13583 0.0702092
R22461 vss.n13583 vss.n13582 0.0702092
R22462 vss.n13599 vss.n13598 0.0702092
R22463 vss.n13600 vss.n13599 0.0702092
R22464 vss.n13592 vss.n13590 0.0702092
R22465 vss.n13592 vss.n13591 0.0702092
R22466 vss.n13596 vss.n13595 0.0702092
R22467 vss.n13640 vss.n13639 0.0702092
R22468 vss.n13642 vss.n13640 0.0702092
R22469 vss.n13650 vss.n13649 0.0702092
R22470 vss.n13649 vss.n13648 0.0702092
R22471 vss.n13630 vss.n13606 0.0702092
R22472 vss.n13631 vss.n13630 0.0702092
R22473 vss.n13633 vss.n13632 0.0702092
R22474 vss.n13632 vss.n13631 0.0702092
R22475 vss.n13647 vss.n13646 0.0702092
R22476 vss.n13648 vss.n13647 0.0702092
R22477 vss.n13644 vss.n13643 0.0702092
R22478 vss.n13643 vss.n13642 0.0702092
R22479 vss.n13628 vss.n13622 0.0702092
R22480 vss.n13628 vss.n13627 0.0702092
R22481 vss.n13625 vss.n13624 0.0702092
R22482 vss.n13554 vss.n13553 0.0702092
R22483 vss.n13553 vss.n13552 0.0702092
R22484 vss.n13536 vss.n13513 0.0702092
R22485 vss.n13537 vss.n13536 0.0702092
R22486 vss.n13534 vss.n13529 0.0702092
R22487 vss.n13534 vss.n13533 0.0702092
R22488 vss.n13532 vss.n13531 0.0702092
R22489 vss.n13533 vss.n13532 0.0702092
R22490 vss.n13539 vss.n13538 0.0702092
R22491 vss.n13538 vss.n13537 0.0702092
R22492 vss.n13551 vss.n13550 0.0702092
R22493 vss.n13552 vss.n13551 0.0702092
R22494 vss.n13544 vss.n13543 0.0702092
R22495 vss.n13543 vss.n1764 0.0702092
R22496 vss.n13548 vss.n13547 0.0702092
R22497 vss.n8290 vss.n8289 0.0702092
R22498 vss.n8291 vss.n8290 0.0702092
R22499 vss.n8299 vss.n8298 0.0702092
R22500 vss.n8298 vss.n8297 0.0702092
R22501 vss.n8280 vss.n8256 0.0702092
R22502 vss.n8281 vss.n8280 0.0702092
R22503 vss.n8283 vss.n8282 0.0702092
R22504 vss.n8282 vss.n8281 0.0702092
R22505 vss.n8296 vss.n8295 0.0702092
R22506 vss.n8297 vss.n8296 0.0702092
R22507 vss.n8293 vss.n8292 0.0702092
R22508 vss.n8292 vss.n8291 0.0702092
R22509 vss.n8278 vss.n8272 0.0702092
R22510 vss.n8278 vss.n8277 0.0702092
R22511 vss.n8275 vss.n8274 0.0702092
R22512 vss.n13791 vss.n13790 0.0702092
R22513 vss.n13790 vss.n13789 0.0702092
R22514 vss.n13770 vss.n13747 0.0702092
R22515 vss.n13771 vss.n13770 0.0702092
R22516 vss.n13768 vss.n13763 0.0702092
R22517 vss.n13768 vss.n13767 0.0702092
R22518 vss.n13766 vss.n13765 0.0702092
R22519 vss.n13767 vss.n13766 0.0702092
R22520 vss.n13773 vss.n13772 0.0702092
R22521 vss.n13772 vss.n13771 0.0702092
R22522 vss.n13788 vss.n13787 0.0702092
R22523 vss.n13789 vss.n13788 0.0702092
R22524 vss.n13781 vss.n13779 0.0702092
R22525 vss.n13781 vss.n13780 0.0702092
R22526 vss.n13785 vss.n13784 0.0702092
R22527 vss.n13829 vss.n13828 0.0702092
R22528 vss.n13831 vss.n13829 0.0702092
R22529 vss.n13839 vss.n13838 0.0702092
R22530 vss.n13838 vss.n13837 0.0702092
R22531 vss.n13819 vss.n13795 0.0702092
R22532 vss.n13820 vss.n13819 0.0702092
R22533 vss.n13822 vss.n13821 0.0702092
R22534 vss.n13821 vss.n13820 0.0702092
R22535 vss.n13836 vss.n13835 0.0702092
R22536 vss.n13837 vss.n13836 0.0702092
R22537 vss.n13833 vss.n13832 0.0702092
R22538 vss.n13832 vss.n13831 0.0702092
R22539 vss.n13817 vss.n13811 0.0702092
R22540 vss.n13817 vss.n13816 0.0702092
R22541 vss.n13814 vss.n13813 0.0702092
R22542 vss.n13847 vss.n13846 0.0702092
R22543 vss.n13852 vss.n13847 0.0702092
R22544 vss.n8253 vss.n8252 0.0702092
R22545 vss.n8252 vss.n8251 0.0702092
R22546 vss.n8244 vss.n8243 0.0702092
R22547 vss.n8245 vss.n8244 0.0702092
R22548 vss.n8247 vss.n8246 0.0702092
R22549 vss.n8246 vss.n8245 0.0702092
R22550 vss.n8250 vss.n8249 0.0702092
R22551 vss.n8251 vss.n8250 0.0702092
R22552 vss.n13854 vss.n13853 0.0702092
R22553 vss.n13853 vss.n13852 0.0702092
R22554 vss.n8226 vss.n8224 0.0702092
R22555 vss.n8224 vss.n8222 0.0702092
R22556 vss.n13856 vss.n8225 0.0702092
R22557 vss.n9076 vss.n9075 0.0702092
R22558 vss.n9077 vss.n9076 0.0702092
R22559 vss.n9085 vss.n9084 0.0702092
R22560 vss.n9084 vss.n9083 0.0702092
R22561 vss.n9066 vss.n9042 0.0702092
R22562 vss.n9067 vss.n9066 0.0702092
R22563 vss.n9069 vss.n9068 0.0702092
R22564 vss.n9068 vss.n9067 0.0702092
R22565 vss.n9082 vss.n9081 0.0702092
R22566 vss.n9083 vss.n9082 0.0702092
R22567 vss.n9079 vss.n9078 0.0702092
R22568 vss.n9078 vss.n9077 0.0702092
R22569 vss.n9064 vss.n9058 0.0702092
R22570 vss.n9064 vss.n9063 0.0702092
R22571 vss.n9061 vss.n9060 0.0702092
R22572 vss.n13079 vss.n13078 0.0702092
R22573 vss.n13078 vss.n13077 0.0702092
R22574 vss.n13058 vss.n13035 0.0702092
R22575 vss.n13059 vss.n13058 0.0702092
R22576 vss.n13056 vss.n13051 0.0702092
R22577 vss.n13056 vss.n13055 0.0702092
R22578 vss.n13054 vss.n13053 0.0702092
R22579 vss.n13055 vss.n13054 0.0702092
R22580 vss.n13061 vss.n13060 0.0702092
R22581 vss.n13060 vss.n13059 0.0702092
R22582 vss.n13076 vss.n13075 0.0702092
R22583 vss.n13077 vss.n13076 0.0702092
R22584 vss.n13069 vss.n13067 0.0702092
R22585 vss.n13069 vss.n13068 0.0702092
R22586 vss.n13073 vss.n13072 0.0702092
R22587 vss.n13117 vss.n13116 0.0702092
R22588 vss.n13119 vss.n13117 0.0702092
R22589 vss.n13127 vss.n13126 0.0702092
R22590 vss.n13126 vss.n13125 0.0702092
R22591 vss.n13107 vss.n13083 0.0702092
R22592 vss.n13108 vss.n13107 0.0702092
R22593 vss.n13110 vss.n13109 0.0702092
R22594 vss.n13109 vss.n13108 0.0702092
R22595 vss.n13124 vss.n13123 0.0702092
R22596 vss.n13125 vss.n13124 0.0702092
R22597 vss.n13121 vss.n13120 0.0702092
R22598 vss.n13120 vss.n13119 0.0702092
R22599 vss.n13105 vss.n13099 0.0702092
R22600 vss.n13105 vss.n13104 0.0702092
R22601 vss.n13102 vss.n13101 0.0702092
R22602 vss.n9039 vss.n9038 0.0702092
R22603 vss.n9038 vss.n9037 0.0702092
R22604 vss.n9021 vss.n8998 0.0702092
R22605 vss.n9022 vss.n9021 0.0702092
R22606 vss.n9019 vss.n9014 0.0702092
R22607 vss.n9019 vss.n9018 0.0702092
R22608 vss.n9017 vss.n9016 0.0702092
R22609 vss.n9018 vss.n9017 0.0702092
R22610 vss.n9024 vss.n9023 0.0702092
R22611 vss.n9023 vss.n9022 0.0702092
R22612 vss.n9036 vss.n9035 0.0702092
R22613 vss.n9037 vss.n9036 0.0702092
R22614 vss.n9029 vss.n9028 0.0702092
R22615 vss.n9028 vss.n8094 0.0702092
R22616 vss.n9033 vss.n9032 0.0702092
R22617 vss.n12614 vss.n12613 0.0702092
R22618 vss.n12615 vss.n12614 0.0702092
R22619 vss.n12623 vss.n12622 0.0702092
R22620 vss.n12622 vss.n12621 0.0702092
R22621 vss.n12604 vss.n12580 0.0702092
R22622 vss.n12605 vss.n12604 0.0702092
R22623 vss.n12607 vss.n12606 0.0702092
R22624 vss.n12606 vss.n12605 0.0702092
R22625 vss.n12620 vss.n12619 0.0702092
R22626 vss.n12621 vss.n12620 0.0702092
R22627 vss.n12617 vss.n12616 0.0702092
R22628 vss.n12616 vss.n12615 0.0702092
R22629 vss.n12602 vss.n12596 0.0702092
R22630 vss.n12602 vss.n12601 0.0702092
R22631 vss.n12599 vss.n12598 0.0702092
R22632 vss.n14085 vss.n14084 0.0702092
R22633 vss.n14084 vss.n14083 0.0702092
R22634 vss.n2170 vss.n2147 0.0702092
R22635 vss.n2171 vss.n2170 0.0702092
R22636 vss.n2168 vss.n2163 0.0702092
R22637 vss.n2168 vss.n2167 0.0702092
R22638 vss.n2166 vss.n2165 0.0702092
R22639 vss.n2167 vss.n2166 0.0702092
R22640 vss.n2173 vss.n2172 0.0702092
R22641 vss.n2172 vss.n2171 0.0702092
R22642 vss.n14082 vss.n14081 0.0702092
R22643 vss.n14083 vss.n14082 0.0702092
R22644 vss.n14075 vss.n2179 0.0702092
R22645 vss.n14075 vss.n14074 0.0702092
R22646 vss.n14079 vss.n14078 0.0702092
R22647 vss.n2205 vss.n2204 0.0702092
R22648 vss.n2204 vss.n2203 0.0702092
R22649 vss.n2208 vss.n2207 0.0702092
R22650 vss.n2209 vss.n2208 0.0702092
R22651 vss.n2219 vss.n2218 0.0702092
R22652 vss.n2218 vss.n2217 0.0702092
R22653 vss.n2221 vss.n2182 0.0702092
R22654 vss.n2182 vss.n2180 0.0702092
R22655 vss.n2183 vss.n2181 0.0702092
R22656 vss.n2181 vss.n2180 0.0702092
R22657 vss.n2216 vss.n2215 0.0702092
R22658 vss.n2217 vss.n2216 0.0702092
R22659 vss.n2210 vss.n2193 0.0702092
R22660 vss.n2210 vss.n2209 0.0702092
R22661 vss.n2202 vss.n2201 0.0702092
R22662 vss.n2203 vss.n2202 0.0702092
R22663 vss.n9298 vss.n9285 0.0702092
R22664 vss.n9285 vss.n9283 0.0702092
R22665 vss.n9296 vss.n9295 0.0702092
R22666 vss.n9295 vss.n9294 0.0702092
R22667 vss.n14098 vss.n14097 0.0702092
R22668 vss.n14097 vss.n14096 0.0702092
R22669 vss.n14100 vss.n2130 0.0702092
R22670 vss.n2130 vss.n2128 0.0702092
R22671 vss.n2131 vss.n2129 0.0702092
R22672 vss.n2129 vss.n2128 0.0702092
R22673 vss.n14095 vss.n14094 0.0702092
R22674 vss.n14096 vss.n14095 0.0702092
R22675 vss.n9293 vss.n2143 0.0702092
R22676 vss.n9294 vss.n9293 0.0702092
R22677 vss.n9286 vss.n9284 0.0702092
R22678 vss.n9284 vss.n9283 0.0702092
R22679 vss.n12844 vss.n12843 0.0702092
R22680 vss.n12845 vss.n12844 0.0702092
R22681 vss.n12851 vss.n12850 0.0702092
R22682 vss.n12850 vss.n12849 0.0702092
R22683 vss.n12864 vss.n12863 0.0702092
R22684 vss.n12865 vss.n12864 0.0702092
R22685 vss.n12861 vss.n12860 0.0702092
R22686 vss.n12860 vss.n12859 0.0702092
R22687 vss.n12858 vss.n12857 0.0702092
R22688 vss.n12859 vss.n12858 0.0702092
R22689 vss.n12867 vss.n12866 0.0702092
R22690 vss.n12866 vss.n12865 0.0702092
R22691 vss.n12848 vss.n9393 0.0702092
R22692 vss.n12849 vss.n12848 0.0702092
R22693 vss.n12846 vss.n9409 0.0702092
R22694 vss.n12846 vss.n12845 0.0702092
R22695 vss.n12771 vss.n12730 0.0702092
R22696 vss.n12730 vss.n12728 0.0702092
R22697 vss.n12769 vss.n12768 0.0702092
R22698 vss.n12768 vss.n12767 0.0702092
R22699 vss.n12759 vss.n12758 0.0702092
R22700 vss.n12760 vss.n12759 0.0702092
R22701 vss.n12756 vss.n12755 0.0702092
R22702 vss.n12755 vss.n12754 0.0702092
R22703 vss.n12753 vss.n12752 0.0702092
R22704 vss.n12754 vss.n12753 0.0702092
R22705 vss.n12762 vss.n12761 0.0702092
R22706 vss.n12761 vss.n12760 0.0702092
R22707 vss.n12766 vss.n12765 0.0702092
R22708 vss.n12767 vss.n12766 0.0702092
R22709 vss.n12731 vss.n12729 0.0702092
R22710 vss.n12729 vss.n12728 0.0702092
R22711 vss.n13321 vss.n13320 0.0702092
R22712 vss.n13322 vss.n13321 0.0702092
R22713 vss.n13328 vss.n13327 0.0702092
R22714 vss.n13327 vss.n13326 0.0702092
R22715 vss.n13341 vss.n13340 0.0702092
R22716 vss.n13342 vss.n13341 0.0702092
R22717 vss.n13338 vss.n13337 0.0702092
R22718 vss.n13337 vss.n13336 0.0702092
R22719 vss.n13335 vss.n13334 0.0702092
R22720 vss.n13336 vss.n13335 0.0702092
R22721 vss.n13344 vss.n13343 0.0702092
R22722 vss.n13343 vss.n13342 0.0702092
R22723 vss.n13325 vss.n8411 0.0702092
R22724 vss.n13326 vss.n13325 0.0702092
R22725 vss.n13323 vss.n8427 0.0702092
R22726 vss.n13323 vss.n13322 0.0702092
R22727 vss.n13440 vss.n13439 0.0702092
R22728 vss.n13441 vss.n13440 0.0702092
R22729 vss.n13447 vss.n13446 0.0702092
R22730 vss.n13446 vss.n13445 0.0702092
R22731 vss.n13460 vss.n13459 0.0702092
R22732 vss.n13461 vss.n13460 0.0702092
R22733 vss.n13457 vss.n13456 0.0702092
R22734 vss.n13456 vss.n13455 0.0702092
R22735 vss.n13454 vss.n13453 0.0702092
R22736 vss.n13455 vss.n13454 0.0702092
R22737 vss.n13463 vss.n13462 0.0702092
R22738 vss.n13462 vss.n13461 0.0702092
R22739 vss.n13444 vss.n13353 0.0702092
R22740 vss.n13445 vss.n13444 0.0702092
R22741 vss.n13442 vss.n13369 0.0702092
R22742 vss.n13442 vss.n13441 0.0702092
R22743 vss.n2051 vss.n2050 0.0702092
R22744 vss.n14180 vss.n2051 0.0702092
R22745 vss.n14188 vss.n14187 0.0702092
R22746 vss.n14187 vss.n14186 0.0702092
R22747 vss.n11857 vss.n2036 0.0702092
R22748 vss.n11858 vss.n11857 0.0702092
R22749 vss.n11850 vss.n11848 0.0702092
R22750 vss.n11848 vss.n11847 0.0702092
R22751 vss.n11862 vss.n11849 0.0702092
R22752 vss.n11849 vss.n11847 0.0702092
R22753 vss.n11860 vss.n11859 0.0702092
R22754 vss.n11859 vss.n11858 0.0702092
R22755 vss.n14185 vss.n14184 0.0702092
R22756 vss.n14186 vss.n14185 0.0702092
R22757 vss.n14182 vss.n14181 0.0702092
R22758 vss.n14181 vss.n14180 0.0702092
R22759 vss.n14445 vss.n14444 0.0702092
R22760 vss.n14446 vss.n14445 0.0702092
R22761 vss.n14414 vss.n14413 0.0702092
R22762 vss.n14453 vss.n1762 0.0702092
R22763 vss.n14453 vss.n14452 0.0702092
R22764 vss.n14475 vss.n14474 0.0702092
R22765 vss.n14474 vss.n14473 0.0702092
R22766 vss.n14455 vss.n1746 0.0702092
R22767 vss.n14456 vss.n14455 0.0702092
R22768 vss.n14451 vss.n14450 0.0702092
R22769 vss.n14452 vss.n14451 0.0702092
R22770 vss.n14458 vss.n14457 0.0702092
R22771 vss.n14457 vss.n14456 0.0702092
R22772 vss.n14472 vss.n14471 0.0702092
R22773 vss.n14473 vss.n14472 0.0702092
R22774 vss.n14465 vss.n14464 0.0702092
R22775 vss.n14466 vss.n14465 0.0702092
R22776 vss.n14469 vss.n14468 0.0702092
R22777 vss.n1806 vss.n1805 0.0702092
R22778 vss.n1807 vss.n1806 0.0702092
R22779 vss.n1803 vss.n1802 0.0702092
R22780 vss.n1802 vss.n1801 0.0702092
R22781 vss.n1794 vss.n1793 0.0702092
R22782 vss.n1795 vss.n1794 0.0702092
R22783 vss.n1797 vss.n1796 0.0702092
R22784 vss.n1796 vss.n1795 0.0702092
R22785 vss.n1800 vss.n1799 0.0702092
R22786 vss.n1801 vss.n1800 0.0702092
R22787 vss.n1809 vss.n1808 0.0702092
R22788 vss.n1808 vss.n1807 0.0702092
R22789 vss.n1812 vss.n1811 0.0702092
R22790 vss.n1813 vss.n1812 0.0702092
R22791 vss.n1781 vss.n1780 0.0702092
R22792 vss.n14363 vss.n1816 0.0702092
R22793 vss.n14396 vss.n1816 0.0702092
R22794 vss.n14389 vss.n14388 0.0702092
R22795 vss.n14390 vss.n14389 0.0702092
R22796 vss.n14386 vss.n14385 0.0702092
R22797 vss.n14385 vss.n14384 0.0702092
R22798 vss.n14376 vss.n14375 0.0702092
R22799 vss.n14380 vss.n14379 0.0702092
R22800 vss.n14379 vss.n14378 0.0702092
R22801 vss.n14383 vss.n14382 0.0702092
R22802 vss.n14384 vss.n14383 0.0702092
R22803 vss.n14392 vss.n14391 0.0702092
R22804 vss.n14391 vss.n14390 0.0702092
R22805 vss.n14395 vss.n14394 0.0702092
R22806 vss.n14396 vss.n14395 0.0702092
R22807 vss.n2007 vss.n2006 0.0702092
R22808 vss.n2008 vss.n2007 0.0702092
R22809 vss.n2014 vss.n2013 0.0702092
R22810 vss.n2013 vss.n2012 0.0702092
R22811 vss.n2028 vss.n2027 0.0702092
R22812 vss.n2029 vss.n2028 0.0702092
R22813 vss.n2025 vss.n2024 0.0702092
R22814 vss.n2024 vss.n2023 0.0702092
R22815 vss.n2022 vss.n2021 0.0702092
R22816 vss.n2023 vss.n2022 0.0702092
R22817 vss.n2031 vss.n2030 0.0702092
R22818 vss.n2030 vss.n2029 0.0702092
R22819 vss.n2011 vss.n1988 0.0702092
R22820 vss.n2012 vss.n2011 0.0702092
R22821 vss.n2009 vss.n2004 0.0702092
R22822 vss.n2009 vss.n2008 0.0702092
R22823 vss.n14262 vss.n14257 0.0702092
R22824 vss.n14262 vss.n1184 0.0702092
R22825 vss.n14276 vss.n14275 0.0702092
R22826 vss.n14276 vss.n1184 0.0702092
R22827 vss.n14279 vss.n14278 0.0702092
R22828 vss.n14278 vss.n1184 0.0702092
R22829 vss.n14260 vss.n14242 0.0702092
R22830 vss.n14260 vss.n1184 0.0702092
R22831 vss.n14265 vss.n14251 0.0702092
R22832 vss.n14271 vss.n14251 0.0702092
R22833 vss.n14267 vss.n14252 0.0702092
R22834 vss.n14271 vss.n14252 0.0702092
R22835 vss.n14270 vss.n14269 0.0702092
R22836 vss.n14271 vss.n14270 0.0702092
R22837 vss.n14273 vss.n14272 0.0702092
R22838 vss.n14272 vss.n14271 0.0702092
R22839 vss.n14171 vss.n14158 0.0702092
R22840 vss.n14158 vss.n14156 0.0702092
R22841 vss.n14793 vss.n14792 0.0702092
R22842 vss.n14794 vss.n14793 0.0702092
R22843 vss.n14802 vss.n14801 0.0702092
R22844 vss.n14801 vss.n14800 0.0702092
R22845 vss.n14163 vss.n1169 0.0702092
R22846 vss.n14166 vss.n14163 0.0702092
R22847 vss.n14159 vss.n14157 0.0702092
R22848 vss.n14157 vss.n14156 0.0702092
R22849 vss.n14165 vss.n14164 0.0702092
R22850 vss.n14166 vss.n14165 0.0702092
R22851 vss.n14799 vss.n14798 0.0702092
R22852 vss.n14800 vss.n14799 0.0702092
R22853 vss.n14796 vss.n14795 0.0702092
R22854 vss.n14795 vss.n14794 0.0702092
R22855 vss.n14319 vss.n14318 0.0702092
R22856 vss.n14320 vss.n14319 0.0702092
R22857 vss.n14308 vss.n14290 0.0702092
R22858 vss.n14320 vss.n14290 0.0702092
R22859 vss.n14322 vss.n14321 0.0702092
R22860 vss.n14321 vss.n14320 0.0702092
R22861 vss.n14289 vss.n14284 0.0702092
R22862 vss.n14320 vss.n14289 0.0702092
R22863 vss.n14296 vss.n14295 0.0702092
R22864 vss.n14312 vss.n14296 0.0702092
R22865 vss.n14313 vss.n14299 0.0702092
R22866 vss.n14313 vss.n14312 0.0702092
R22867 vss.n14306 vss.n14300 0.0702092
R22868 vss.n14312 vss.n14300 0.0702092
R22869 vss.n14311 vss.n14310 0.0702092
R22870 vss.n14312 vss.n14311 0.0702092
R22871 vss.n14843 vss.n1164 0.0702092
R22872 vss.n1164 vss.n1162 0.0702092
R22873 vss.n14841 vss.n14840 0.0702092
R22874 vss.n14840 vss.n14839 0.0702092
R22875 vss.n14838 vss.n14837 0.0702092
R22876 vss.n14839 vss.n14838 0.0702092
R22877 vss.n1165 vss.n1163 0.0702092
R22878 vss.n1163 vss.n1162 0.0702092
R22879 vss.n15140 vss.n15139 0.0702092
R22880 vss.n15141 vss.n15140 0.0702092
R22881 vss.n15109 vss.n15108 0.0702092
R22882 vss.n15148 vss.n983 0.0702092
R22883 vss.n15148 vss.n15147 0.0702092
R22884 vss.n15170 vss.n15169 0.0702092
R22885 vss.n15169 vss.n15168 0.0702092
R22886 vss.n15150 vss.n967 0.0702092
R22887 vss.n15151 vss.n15150 0.0702092
R22888 vss.n15146 vss.n15145 0.0702092
R22889 vss.n15147 vss.n15146 0.0702092
R22890 vss.n15153 vss.n15152 0.0702092
R22891 vss.n15152 vss.n15151 0.0702092
R22892 vss.n15167 vss.n15166 0.0702092
R22893 vss.n15168 vss.n15167 0.0702092
R22894 vss.n15160 vss.n15159 0.0702092
R22895 vss.n15161 vss.n15160 0.0702092
R22896 vss.n15164 vss.n15163 0.0702092
R22897 vss.n1027 vss.n1026 0.0702092
R22898 vss.n1028 vss.n1027 0.0702092
R22899 vss.n1024 vss.n1023 0.0702092
R22900 vss.n1023 vss.n1022 0.0702092
R22901 vss.n1015 vss.n1014 0.0702092
R22902 vss.n1016 vss.n1015 0.0702092
R22903 vss.n1018 vss.n1017 0.0702092
R22904 vss.n1017 vss.n1016 0.0702092
R22905 vss.n1021 vss.n1020 0.0702092
R22906 vss.n1022 vss.n1021 0.0702092
R22907 vss.n1030 vss.n1029 0.0702092
R22908 vss.n1029 vss.n1028 0.0702092
R22909 vss.n1033 vss.n1032 0.0702092
R22910 vss.n1034 vss.n1033 0.0702092
R22911 vss.n1002 vss.n1001 0.0702092
R22912 vss.n15058 vss.n1037 0.0702092
R22913 vss.n15091 vss.n1037 0.0702092
R22914 vss.n15084 vss.n15083 0.0702092
R22915 vss.n15085 vss.n15084 0.0702092
R22916 vss.n15081 vss.n15080 0.0702092
R22917 vss.n15080 vss.n15079 0.0702092
R22918 vss.n15071 vss.n15070 0.0702092
R22919 vss.n15075 vss.n15074 0.0702092
R22920 vss.n15074 vss.n15073 0.0702092
R22921 vss.n15078 vss.n15077 0.0702092
R22922 vss.n15079 vss.n15078 0.0702092
R22923 vss.n15087 vss.n15086 0.0702092
R22924 vss.n15086 vss.n15085 0.0702092
R22925 vss.n15090 vss.n15089 0.0702092
R22926 vss.n15091 vss.n15090 0.0702092
R22927 vss.n1112 vss.n1111 0.0702092
R22928 vss.n1113 vss.n1112 0.0702092
R22929 vss.n1119 vss.n1118 0.0702092
R22930 vss.n1118 vss.n1117 0.0702092
R22931 vss.n1133 vss.n1132 0.0702092
R22932 vss.n1134 vss.n1133 0.0702092
R22933 vss.n1130 vss.n1129 0.0702092
R22934 vss.n1129 vss.n1128 0.0702092
R22935 vss.n1127 vss.n1126 0.0702092
R22936 vss.n1128 vss.n1127 0.0702092
R22937 vss.n1136 vss.n1135 0.0702092
R22938 vss.n1135 vss.n1134 0.0702092
R22939 vss.n1116 vss.n1093 0.0702092
R22940 vss.n1117 vss.n1116 0.0702092
R22941 vss.n1114 vss.n1109 0.0702092
R22942 vss.n1114 vss.n1113 0.0702092
R22943 vss.n14957 vss.n14952 0.0702092
R22944 vss.n14957 vss.n405 0.0702092
R22945 vss.n14971 vss.n14970 0.0702092
R22946 vss.n14971 vss.n405 0.0702092
R22947 vss.n14974 vss.n14973 0.0702092
R22948 vss.n14973 vss.n405 0.0702092
R22949 vss.n14955 vss.n14937 0.0702092
R22950 vss.n14955 vss.n405 0.0702092
R22951 vss.n14960 vss.n14946 0.0702092
R22952 vss.n14966 vss.n14946 0.0702092
R22953 vss.n14962 vss.n14947 0.0702092
R22954 vss.n14966 vss.n14947 0.0702092
R22955 vss.n14965 vss.n14964 0.0702092
R22956 vss.n14966 vss.n14965 0.0702092
R22957 vss.n14968 vss.n14967 0.0702092
R22958 vss.n14967 vss.n14966 0.0702092
R22959 vss.n14865 vss.n14852 0.0702092
R22960 vss.n14852 vss.n14850 0.0702092
R22961 vss.n15488 vss.n15487 0.0702092
R22962 vss.n15489 vss.n15488 0.0702092
R22963 vss.n15497 vss.n15496 0.0702092
R22964 vss.n15496 vss.n15495 0.0702092
R22965 vss.n14857 vss.n390 0.0702092
R22966 vss.n14860 vss.n14857 0.0702092
R22967 vss.n14853 vss.n14851 0.0702092
R22968 vss.n14851 vss.n14850 0.0702092
R22969 vss.n14859 vss.n14858 0.0702092
R22970 vss.n14860 vss.n14859 0.0702092
R22971 vss.n15494 vss.n15493 0.0702092
R22972 vss.n15495 vss.n15494 0.0702092
R22973 vss.n15491 vss.n15490 0.0702092
R22974 vss.n15490 vss.n15489 0.0702092
R22975 vss.n15014 vss.n15013 0.0702092
R22976 vss.n15015 vss.n15014 0.0702092
R22977 vss.n15003 vss.n14985 0.0702092
R22978 vss.n15015 vss.n14985 0.0702092
R22979 vss.n15017 vss.n15016 0.0702092
R22980 vss.n15016 vss.n15015 0.0702092
R22981 vss.n14984 vss.n14979 0.0702092
R22982 vss.n15015 vss.n14984 0.0702092
R22983 vss.n14991 vss.n14990 0.0702092
R22984 vss.n15007 vss.n14991 0.0702092
R22985 vss.n15008 vss.n14994 0.0702092
R22986 vss.n15008 vss.n15007 0.0702092
R22987 vss.n15001 vss.n14995 0.0702092
R22988 vss.n15007 vss.n14995 0.0702092
R22989 vss.n15006 vss.n15005 0.0702092
R22990 vss.n15007 vss.n15006 0.0702092
R22991 vss.n15538 vss.n385 0.0702092
R22992 vss.n385 vss.n383 0.0702092
R22993 vss.n15536 vss.n15535 0.0702092
R22994 vss.n15535 vss.n15534 0.0702092
R22995 vss.n15533 vss.n15532 0.0702092
R22996 vss.n15534 vss.n15533 0.0702092
R22997 vss.n386 vss.n384 0.0702092
R22998 vss.n384 vss.n383 0.0702092
R22999 vss.n6217 vss.n6206 0.0702092
R23000 vss.n6250 vss.n6206 0.0702092
R23001 vss.n6243 vss.n6242 0.0702092
R23002 vss.n6244 vss.n6243 0.0702092
R23003 vss.n6240 vss.n6239 0.0702092
R23004 vss.n6239 vss.n6238 0.0702092
R23005 vss.n6230 vss.n6229 0.0702092
R23006 vss.n6234 vss.n6233 0.0702092
R23007 vss.n6233 vss.n6232 0.0702092
R23008 vss.n6237 vss.n6236 0.0702092
R23009 vss.n6238 vss.n6237 0.0702092
R23010 vss.n6246 vss.n6245 0.0702092
R23011 vss.n6245 vss.n6244 0.0702092
R23012 vss.n6249 vss.n6248 0.0702092
R23013 vss.n6250 vss.n6249 0.0702092
R23014 vss.n3953 vss.n3950 0.0702092
R23015 vss.n3965 vss.n3950 0.0702092
R23016 vss.n3958 vss.n3955 0.0702092
R23017 vss.n3958 vss.n3957 0.0702092
R23018 vss.n15864 vss.n15863 0.0702092
R23019 vss.n15865 vss.n15864 0.0702092
R23020 vss.n15861 vss.n15860 0.0702092
R23021 vss.n15860 vss.n15859 0.0702092
R23022 vss.n15858 vss.n15857 0.0702092
R23023 vss.n15859 vss.n15858 0.0702092
R23024 vss.n15867 vss.n15866 0.0702092
R23025 vss.n15866 vss.n15865 0.0702092
R23026 vss.n3956 vss.n30 0.0702092
R23027 vss.n3957 vss.n3956 0.0702092
R23028 vss.n3964 vss.n3963 0.0702092
R23029 vss.n3965 vss.n3964 0.0702092
R23030 vss.n3863 vss.n3852 0.0702092
R23031 vss.n3896 vss.n3852 0.0702092
R23032 vss.n3889 vss.n3888 0.0702092
R23033 vss.n3890 vss.n3889 0.0702092
R23034 vss.n3886 vss.n3885 0.0702092
R23035 vss.n3885 vss.n3884 0.0702092
R23036 vss.n3877 vss.n3876 0.0702092
R23037 vss.n3878 vss.n3877 0.0702092
R23038 vss.n3880 vss.n3879 0.0702092
R23039 vss.n3879 vss.n3878 0.0702092
R23040 vss.n3883 vss.n3882 0.0702092
R23041 vss.n3884 vss.n3883 0.0702092
R23042 vss.n3892 vss.n3891 0.0702092
R23043 vss.n3891 vss.n3890 0.0702092
R23044 vss.n3895 vss.n3894 0.0702092
R23045 vss.n3896 vss.n3895 0.0702092
R23046 vss.n3744 vss.n3733 0.0702092
R23047 vss.n3777 vss.n3733 0.0702092
R23048 vss.n3770 vss.n3769 0.0702092
R23049 vss.n3771 vss.n3770 0.0702092
R23050 vss.n3767 vss.n3766 0.0702092
R23051 vss.n3766 vss.n3765 0.0702092
R23052 vss.n3758 vss.n3757 0.0702092
R23053 vss.n3759 vss.n3758 0.0702092
R23054 vss.n3761 vss.n3760 0.0702092
R23055 vss.n3760 vss.n3759 0.0702092
R23056 vss.n3764 vss.n3763 0.0702092
R23057 vss.n3765 vss.n3764 0.0702092
R23058 vss.n3773 vss.n3772 0.0702092
R23059 vss.n3772 vss.n3771 0.0702092
R23060 vss.n3776 vss.n3775 0.0702092
R23061 vss.n3777 vss.n3776 0.0702092
R23062 vss.n3625 vss.n3614 0.0702092
R23063 vss.n3658 vss.n3614 0.0702092
R23064 vss.n3651 vss.n3650 0.0702092
R23065 vss.n3652 vss.n3651 0.0702092
R23066 vss.n3648 vss.n3647 0.0702092
R23067 vss.n3647 vss.n3646 0.0702092
R23068 vss.n3639 vss.n3638 0.0702092
R23069 vss.n3640 vss.n3639 0.0702092
R23070 vss.n3642 vss.n3641 0.0702092
R23071 vss.n3641 vss.n3640 0.0702092
R23072 vss.n3645 vss.n3644 0.0702092
R23073 vss.n3646 vss.n3645 0.0702092
R23074 vss.n3654 vss.n3653 0.0702092
R23075 vss.n3653 vss.n3652 0.0702092
R23076 vss.n3657 vss.n3656 0.0702092
R23077 vss.n3658 vss.n3657 0.0702092
R23078 vss.n6306 vss.n6293 0.0702092
R23079 vss.n6293 vss.n6291 0.0702092
R23080 vss.n15690 vss.n15689 0.0702092
R23081 vss.n15691 vss.n15690 0.0702092
R23082 vss.n15699 vss.n15698 0.0702092
R23083 vss.n15698 vss.n15697 0.0702092
R23084 vss.n6298 vss.n245 0.0702092
R23085 vss.n6301 vss.n6298 0.0702092
R23086 vss.n6294 vss.n6292 0.0702092
R23087 vss.n6292 vss.n6291 0.0702092
R23088 vss.n6300 vss.n6299 0.0702092
R23089 vss.n6301 vss.n6300 0.0702092
R23090 vss.n15696 vss.n15695 0.0702092
R23091 vss.n15697 vss.n15696 0.0702092
R23092 vss.n15693 vss.n15692 0.0702092
R23093 vss.n15692 vss.n15691 0.0702092
R23094 vss.n15600 vss.n15595 0.0702092
R23095 vss.n15600 vss.n302 0.0702092
R23096 vss.n15614 vss.n15613 0.0702092
R23097 vss.n15614 vss.n302 0.0702092
R23098 vss.n15617 vss.n15616 0.0702092
R23099 vss.n15616 vss.n302 0.0702092
R23100 vss.n15598 vss.n15580 0.0702092
R23101 vss.n15598 vss.n302 0.0702092
R23102 vss.n15603 vss.n15589 0.0702092
R23103 vss.n15609 vss.n15589 0.0702092
R23104 vss.n15605 vss.n15590 0.0702092
R23105 vss.n15609 vss.n15590 0.0702092
R23106 vss.n15608 vss.n15607 0.0702092
R23107 vss.n15609 vss.n15608 0.0702092
R23108 vss.n15611 vss.n15610 0.0702092
R23109 vss.n15610 vss.n15609 0.0702092
R23110 vss.n316 vss.n306 0.0702092
R23111 vss.n349 vss.n306 0.0702092
R23112 vss.n342 vss.n341 0.0702092
R23113 vss.n343 vss.n342 0.0702092
R23114 vss.n339 vss.n338 0.0702092
R23115 vss.n338 vss.n337 0.0702092
R23116 vss.n330 vss.n329 0.0702092
R23117 vss.n331 vss.n330 0.0702092
R23118 vss.n333 vss.n332 0.0702092
R23119 vss.n332 vss.n331 0.0702092
R23120 vss.n336 vss.n335 0.0702092
R23121 vss.n337 vss.n336 0.0702092
R23122 vss.n345 vss.n344 0.0702092
R23123 vss.n344 vss.n343 0.0702092
R23124 vss.n348 vss.n347 0.0702092
R23125 vss.n349 vss.n348 0.0702092
R23126 vss.n3596 vss.n3595 0.0702092
R23127 vss.n3597 vss.n3596 0.0702092
R23128 vss.n3608 vss.n3566 0.0702092
R23129 vss.n3566 vss.n3564 0.0702092
R23130 vss.n3606 vss.n3605 0.0702092
R23131 vss.n3605 vss.n3604 0.0702092
R23132 vss.n3599 vss.n3598 0.0702092
R23133 vss.n3598 vss.n3597 0.0702092
R23134 vss.n3603 vss.n3602 0.0702092
R23135 vss.n3604 vss.n3603 0.0702092
R23136 vss.n3567 vss.n3565 0.0702092
R23137 vss.n3565 vss.n3564 0.0702092
R23138 vss.n6315 vss.n6314 0.0702092
R23139 vss.n6314 vss.n6313 0.0702092
R23140 vss.n3562 vss.n3561 0.0702092
R23141 vss.n3593 vss.n3592 0.0702092
R23142 vss.n3592 vss.n3591 0.0702092
R23143 vss.n3588 vss.n3587 0.0702092
R23144 vss.n15638 vss.n356 0.0702092
R23145 vss.n15656 vss.n356 0.0702092
R23146 vss.n15652 vss.n355 0.0702092
R23147 vss.n15656 vss.n355 0.0702092
R23148 vss.n15655 vss.n15654 0.0702092
R23149 vss.n15656 vss.n15655 0.0702092
R23150 vss.n15636 vss.n354 0.0702092
R23151 vss.n15656 vss.n354 0.0702092
R23152 vss.n15641 vss.n15627 0.0702092
R23153 vss.n15648 vss.n15627 0.0702092
R23154 vss.n15643 vss.n15628 0.0702092
R23155 vss.n15648 vss.n15628 0.0702092
R23156 vss.n15647 vss.n15646 0.0702092
R23157 vss.n15648 vss.n15647 0.0702092
R23158 vss.n15649 vss.n15624 0.0702092
R23159 vss.n15649 vss.n15648 0.0702092
R23160 vss.n15550 vss.n15549 0.0702092
R23161 vss.n15551 vss.n15550 0.0702092
R23162 vss.n15557 vss.n15556 0.0702092
R23163 vss.n15556 vss.n15555 0.0702092
R23164 vss.n15570 vss.n15569 0.0702092
R23165 vss.n15571 vss.n15570 0.0702092
R23166 vss.n15567 vss.n15566 0.0702092
R23167 vss.n15566 vss.n15565 0.0702092
R23168 vss.n15564 vss.n15563 0.0702092
R23169 vss.n15565 vss.n15564 0.0702092
R23170 vss.n15573 vss.n15572 0.0702092
R23171 vss.n15572 vss.n15571 0.0702092
R23172 vss.n15554 vss.n361 0.0702092
R23173 vss.n15555 vss.n15554 0.0702092
R23174 vss.n15552 vss.n377 0.0702092
R23175 vss.n15552 vss.n15551 0.0702092
R23176 vss.n12175 vss.n12174 0.0702092
R23177 vss.n12174 vss.n12173 0.0702092
R23178 vss.n12172 vss.n12171 0.0702092
R23179 vss.n12173 vss.n12172 0.0702092
R23180 vss.n12163 vss.n12162 0.0702092
R23181 vss.n12162 vss.n12161 0.0702092
R23182 vss.n12166 vss.n12165 0.0702092
R23183 vss.n12167 vss.n12166 0.0702092
R23184 vss.n12169 vss.n12168 0.0702092
R23185 vss.n12168 vss.n12167 0.0702092
R23186 vss.n12160 vss.n12159 0.0702092
R23187 vss.n12161 vss.n12160 0.0702092
R23188 vss.n12177 vss.n12135 0.0702092
R23189 vss.n12135 vss.n12133 0.0702092
R23190 vss.n12136 vss.n12134 0.0702092
R23191 vss.n12134 vss.n12133 0.0702092
R23192 vss.n11794 vss.n11767 0.0702092
R23193 vss.n11794 vss.n11793 0.0702092
R23194 vss.n11791 vss.n11790 0.0702092
R23195 vss.n11782 vss.n11764 0.0702092
R23196 vss.n11797 vss.n11764 0.0702092
R23197 vss.n11799 vss.n11798 0.0702092
R23198 vss.n11798 vss.n11797 0.0702092
R23199 vss.n11796 vss.n11759 0.0702092
R23200 vss.n11797 vss.n11796 0.0702092
R23201 vss.n11788 vss.n11787 0.0702092
R23202 vss.n11787 vss.n11786 0.0702092
R23203 vss.n11780 vss.n11775 0.0702092
R23204 vss.n11786 vss.n11775 0.0702092
R23205 vss.n11785 vss.n11784 0.0702092
R23206 vss.n11786 vss.n11785 0.0702092
R23207 vss.n13230 vss.n13229 0.0702092
R23208 vss.n13229 vss.n13228 0.0702092
R23209 vss.n13245 vss.n8813 0.0702092
R23210 vss.n8813 vss.n8811 0.0702092
R23211 vss.n13243 vss.n13242 0.0702092
R23212 vss.n13242 vss.n13241 0.0702092
R23213 vss.n13233 vss.n13232 0.0702092
R23214 vss.n13234 vss.n13233 0.0702092
R23215 vss.n13227 vss.n13226 0.0702092
R23216 vss.n13228 vss.n13227 0.0702092
R23217 vss.n13236 vss.n13235 0.0702092
R23218 vss.n13235 vss.n13234 0.0702092
R23219 vss.n13240 vss.n13239 0.0702092
R23220 vss.n13241 vss.n13240 0.0702092
R23221 vss.n8814 vss.n8812 0.0702092
R23222 vss.n8812 vss.n8811 0.0702092
R23223 vss.n9882 vss.n9880 0.0702092
R23224 vss.n9880 vss.n9879 0.0702092
R23225 vss.n11714 vss.n11713 0.0702092
R23226 vss.n11718 vss.n11714 0.0702092
R23227 vss.n9910 vss.n9909 0.0702092
R23228 vss.n9909 vss.n9908 0.0702092
R23229 vss.n9907 vss.n9906 0.0702092
R23230 vss.n9908 vss.n9907 0.0702092
R23231 vss.n11720 vss.n11719 0.0702092
R23232 vss.n11719 vss.n11718 0.0702092
R23233 vss.n11722 vss.n9881 0.0702092
R23234 vss.n9881 vss.n9879 0.0702092
R23235 vss.n9900 vss.n9899 0.0702092
R23236 vss.n9901 vss.n9900 0.0702092
R23237 vss.n9904 vss.n9903 0.0702092
R23238 vss.n11560 vss.n11559 0.0702092
R23239 vss.n11559 vss.n11558 0.0702092
R23240 vss.n11539 vss.n11516 0.0702092
R23241 vss.n11540 vss.n11539 0.0702092
R23242 vss.n11537 vss.n11532 0.0702092
R23243 vss.n11537 vss.n11536 0.0702092
R23244 vss.n11535 vss.n11534 0.0702092
R23245 vss.n11536 vss.n11535 0.0702092
R23246 vss.n11542 vss.n11541 0.0702092
R23247 vss.n11541 vss.n11540 0.0702092
R23248 vss.n11557 vss.n11556 0.0702092
R23249 vss.n11558 vss.n11557 0.0702092
R23250 vss.n11550 vss.n11548 0.0702092
R23251 vss.n11550 vss.n11549 0.0702092
R23252 vss.n11554 vss.n11553 0.0702092
R23253 vss.n11598 vss.n11597 0.0702092
R23254 vss.n11600 vss.n11598 0.0702092
R23255 vss.n11608 vss.n11607 0.0702092
R23256 vss.n11607 vss.n11606 0.0702092
R23257 vss.n11588 vss.n11564 0.0702092
R23258 vss.n11589 vss.n11588 0.0702092
R23259 vss.n11591 vss.n11590 0.0702092
R23260 vss.n11590 vss.n11589 0.0702092
R23261 vss.n11605 vss.n11604 0.0702092
R23262 vss.n11606 vss.n11605 0.0702092
R23263 vss.n11602 vss.n11601 0.0702092
R23264 vss.n11601 vss.n11600 0.0702092
R23265 vss.n11586 vss.n11580 0.0702092
R23266 vss.n11586 vss.n11585 0.0702092
R23267 vss.n11583 vss.n11582 0.0702092
R23268 vss.n11513 vss.n11512 0.0702092
R23269 vss.n11512 vss.n11511 0.0702092
R23270 vss.n11495 vss.n11472 0.0702092
R23271 vss.n11496 vss.n11495 0.0702092
R23272 vss.n11493 vss.n11488 0.0702092
R23273 vss.n11493 vss.n11492 0.0702092
R23274 vss.n11491 vss.n11490 0.0702092
R23275 vss.n11492 vss.n11491 0.0702092
R23276 vss.n11498 vss.n11497 0.0702092
R23277 vss.n11497 vss.n11496 0.0702092
R23278 vss.n11510 vss.n11509 0.0702092
R23279 vss.n11511 vss.n11510 0.0702092
R23280 vss.n11503 vss.n11502 0.0702092
R23281 vss.n11502 vss.n9802 0.0702092
R23282 vss.n11507 vss.n11506 0.0702092
R23283 vss.n11145 vss.n11144 0.0702092
R23284 vss.n11146 vss.n11145 0.0702092
R23285 vss.n11154 vss.n11153 0.0702092
R23286 vss.n11153 vss.n11152 0.0702092
R23287 vss.n11135 vss.n11111 0.0702092
R23288 vss.n11136 vss.n11135 0.0702092
R23289 vss.n11138 vss.n11137 0.0702092
R23290 vss.n11137 vss.n11136 0.0702092
R23291 vss.n11151 vss.n11150 0.0702092
R23292 vss.n11152 vss.n11151 0.0702092
R23293 vss.n11148 vss.n11147 0.0702092
R23294 vss.n11147 vss.n11146 0.0702092
R23295 vss.n11133 vss.n11127 0.0702092
R23296 vss.n11133 vss.n11132 0.0702092
R23297 vss.n11130 vss.n11129 0.0702092
R23298 vss.n11249 vss.n11248 0.0702092
R23299 vss.n11248 vss.n11247 0.0702092
R23300 vss.n11228 vss.n11205 0.0702092
R23301 vss.n11229 vss.n11228 0.0702092
R23302 vss.n11226 vss.n11221 0.0702092
R23303 vss.n11226 vss.n11225 0.0702092
R23304 vss.n11224 vss.n11223 0.0702092
R23305 vss.n11225 vss.n11224 0.0702092
R23306 vss.n11231 vss.n11230 0.0702092
R23307 vss.n11230 vss.n11229 0.0702092
R23308 vss.n11246 vss.n11245 0.0702092
R23309 vss.n11247 vss.n11246 0.0702092
R23310 vss.n11239 vss.n11237 0.0702092
R23311 vss.n11239 vss.n11238 0.0702092
R23312 vss.n11243 vss.n11242 0.0702092
R23313 vss.n11287 vss.n11286 0.0702092
R23314 vss.n11289 vss.n11287 0.0702092
R23315 vss.n11297 vss.n11296 0.0702092
R23316 vss.n11296 vss.n11295 0.0702092
R23317 vss.n11277 vss.n11253 0.0702092
R23318 vss.n11278 vss.n11277 0.0702092
R23319 vss.n11280 vss.n11279 0.0702092
R23320 vss.n11279 vss.n11278 0.0702092
R23321 vss.n11294 vss.n11293 0.0702092
R23322 vss.n11295 vss.n11294 0.0702092
R23323 vss.n11291 vss.n11290 0.0702092
R23324 vss.n11290 vss.n11289 0.0702092
R23325 vss.n11275 vss.n11269 0.0702092
R23326 vss.n11275 vss.n11274 0.0702092
R23327 vss.n11272 vss.n11271 0.0702092
R23328 vss.n11108 vss.n11107 0.0702092
R23329 vss.n11107 vss.n11106 0.0702092
R23330 vss.n11090 vss.n11067 0.0702092
R23331 vss.n11091 vss.n11090 0.0702092
R23332 vss.n11088 vss.n11083 0.0702092
R23333 vss.n11088 vss.n11087 0.0702092
R23334 vss.n11086 vss.n11085 0.0702092
R23335 vss.n11087 vss.n11086 0.0702092
R23336 vss.n11093 vss.n11092 0.0702092
R23337 vss.n11092 vss.n11091 0.0702092
R23338 vss.n11105 vss.n11104 0.0702092
R23339 vss.n11106 vss.n11105 0.0702092
R23340 vss.n11098 vss.n11097 0.0702092
R23341 vss.n11097 vss.n9673 0.0702092
R23342 vss.n11102 vss.n11101 0.0702092
R23343 vss.n10948 vss.n10947 0.0702092
R23344 vss.n10949 vss.n10948 0.0702092
R23345 vss.n10957 vss.n10956 0.0702092
R23346 vss.n10956 vss.n10955 0.0702092
R23347 vss.n10938 vss.n10914 0.0702092
R23348 vss.n10939 vss.n10938 0.0702092
R23349 vss.n10941 vss.n10940 0.0702092
R23350 vss.n10940 vss.n10939 0.0702092
R23351 vss.n10954 vss.n10953 0.0702092
R23352 vss.n10955 vss.n10954 0.0702092
R23353 vss.n10951 vss.n10950 0.0702092
R23354 vss.n10950 vss.n10949 0.0702092
R23355 vss.n10936 vss.n10930 0.0702092
R23356 vss.n10936 vss.n10935 0.0702092
R23357 vss.n10933 vss.n10932 0.0702092
R23358 vss.n10910 vss.n10909 0.0702092
R23359 vss.n10909 vss.n10908 0.0702092
R23360 vss.n10889 vss.n10866 0.0702092
R23361 vss.n10890 vss.n10889 0.0702092
R23362 vss.n10887 vss.n10882 0.0702092
R23363 vss.n10887 vss.n10886 0.0702092
R23364 vss.n10885 vss.n10884 0.0702092
R23365 vss.n10886 vss.n10885 0.0702092
R23366 vss.n10892 vss.n10891 0.0702092
R23367 vss.n10891 vss.n10890 0.0702092
R23368 vss.n10907 vss.n10906 0.0702092
R23369 vss.n10908 vss.n10907 0.0702092
R23370 vss.n10900 vss.n10898 0.0702092
R23371 vss.n10900 vss.n10899 0.0702092
R23372 vss.n10904 vss.n10903 0.0702092
R23373 vss.n10852 vss.n10851 0.0702092
R23374 vss.n10854 vss.n10852 0.0702092
R23375 vss.n10862 vss.n10861 0.0702092
R23376 vss.n10861 vss.n10860 0.0702092
R23377 vss.n10842 vss.n10818 0.0702092
R23378 vss.n10843 vss.n10842 0.0702092
R23379 vss.n10845 vss.n10844 0.0702092
R23380 vss.n10844 vss.n10843 0.0702092
R23381 vss.n10859 vss.n10858 0.0702092
R23382 vss.n10860 vss.n10859 0.0702092
R23383 vss.n10856 vss.n10855 0.0702092
R23384 vss.n10855 vss.n10854 0.0702092
R23385 vss.n10840 vss.n10834 0.0702092
R23386 vss.n10840 vss.n10839 0.0702092
R23387 vss.n10837 vss.n10836 0.0702092
R23388 vss.n10211 vss.n10210 0.0702092
R23389 vss.n10210 vss.n10209 0.0702092
R23390 vss.n10193 vss.n10170 0.0702092
R23391 vss.n10194 vss.n10193 0.0702092
R23392 vss.n10191 vss.n10186 0.0702092
R23393 vss.n10191 vss.n10190 0.0702092
R23394 vss.n10189 vss.n10188 0.0702092
R23395 vss.n10190 vss.n10189 0.0702092
R23396 vss.n10196 vss.n10195 0.0702092
R23397 vss.n10195 vss.n10194 0.0702092
R23398 vss.n10208 vss.n10207 0.0702092
R23399 vss.n10209 vss.n10208 0.0702092
R23400 vss.n10201 vss.n10200 0.0702092
R23401 vss.n10200 vss.n9544 0.0702092
R23402 vss.n10205 vss.n10204 0.0702092
R23403 vss.n10554 vss.n10553 0.0702092
R23404 vss.n10555 vss.n10554 0.0702092
R23405 vss.n10563 vss.n10562 0.0702092
R23406 vss.n10562 vss.n10561 0.0702092
R23407 vss.n10544 vss.n10520 0.0702092
R23408 vss.n10545 vss.n10544 0.0702092
R23409 vss.n10547 vss.n10546 0.0702092
R23410 vss.n10546 vss.n10545 0.0702092
R23411 vss.n10560 vss.n10559 0.0702092
R23412 vss.n10561 vss.n10560 0.0702092
R23413 vss.n10557 vss.n10556 0.0702092
R23414 vss.n10556 vss.n10555 0.0702092
R23415 vss.n10542 vss.n10536 0.0702092
R23416 vss.n10542 vss.n10541 0.0702092
R23417 vss.n10539 vss.n10538 0.0702092
R23418 vss.n10516 vss.n10515 0.0702092
R23419 vss.n10515 vss.n10514 0.0702092
R23420 vss.n10495 vss.n10472 0.0702092
R23421 vss.n10496 vss.n10495 0.0702092
R23422 vss.n10493 vss.n10488 0.0702092
R23423 vss.n10493 vss.n10492 0.0702092
R23424 vss.n10491 vss.n10490 0.0702092
R23425 vss.n10492 vss.n10491 0.0702092
R23426 vss.n10498 vss.n10497 0.0702092
R23427 vss.n10497 vss.n10496 0.0702092
R23428 vss.n10513 vss.n10512 0.0702092
R23429 vss.n10514 vss.n10513 0.0702092
R23430 vss.n10506 vss.n10504 0.0702092
R23431 vss.n10506 vss.n10505 0.0702092
R23432 vss.n10510 vss.n10509 0.0702092
R23433 vss.n10444 vss.n10443 0.0702092
R23434 vss.n10445 vss.n10444 0.0702092
R23435 vss.n10451 vss.n10450 0.0702092
R23436 vss.n10450 vss.n10449 0.0702092
R23437 vss.n10465 vss.n10464 0.0702092
R23438 vss.n10466 vss.n10465 0.0702092
R23439 vss.n10462 vss.n10461 0.0702092
R23440 vss.n10461 vss.n10460 0.0702092
R23441 vss.n10459 vss.n10458 0.0702092
R23442 vss.n10460 vss.n10459 0.0702092
R23443 vss.n10468 vss.n10467 0.0702092
R23444 vss.n10467 vss.n10466 0.0702092
R23445 vss.n10448 vss.n10425 0.0702092
R23446 vss.n10449 vss.n10448 0.0702092
R23447 vss.n10446 vss.n10441 0.0702092
R23448 vss.n10446 vss.n10445 0.0702092
R23449 vss.n10590 vss.n10589 0.0702092
R23450 vss.n10591 vss.n10590 0.0702092
R23451 vss.n10597 vss.n10596 0.0702092
R23452 vss.n10596 vss.n10595 0.0702092
R23453 vss.n10610 vss.n10609 0.0702092
R23454 vss.n10611 vss.n10610 0.0702092
R23455 vss.n10607 vss.n10606 0.0702092
R23456 vss.n10606 vss.n10605 0.0702092
R23457 vss.n10604 vss.n10603 0.0702092
R23458 vss.n10605 vss.n10604 0.0702092
R23459 vss.n10613 vss.n10612 0.0702092
R23460 vss.n10612 vss.n10611 0.0702092
R23461 vss.n10594 vss.n10570 0.0702092
R23462 vss.n10595 vss.n10594 0.0702092
R23463 vss.n10592 vss.n10586 0.0702092
R23464 vss.n10592 vss.n10591 0.0702092
R23465 vss.n10984 vss.n10983 0.0702092
R23466 vss.n10985 vss.n10984 0.0702092
R23467 vss.n10991 vss.n10990 0.0702092
R23468 vss.n10990 vss.n10989 0.0702092
R23469 vss.n11004 vss.n11003 0.0702092
R23470 vss.n11005 vss.n11004 0.0702092
R23471 vss.n11001 vss.n11000 0.0702092
R23472 vss.n11000 vss.n10999 0.0702092
R23473 vss.n10998 vss.n10997 0.0702092
R23474 vss.n10999 vss.n10998 0.0702092
R23475 vss.n11007 vss.n11006 0.0702092
R23476 vss.n11006 vss.n11005 0.0702092
R23477 vss.n10988 vss.n10964 0.0702092
R23478 vss.n10989 vss.n10988 0.0702092
R23479 vss.n10986 vss.n10980 0.0702092
R23480 vss.n10986 vss.n10985 0.0702092
R23481 vss.n10035 vss.n9994 0.0702092
R23482 vss.n9994 vss.n9992 0.0702092
R23483 vss.n10033 vss.n10032 0.0702092
R23484 vss.n10032 vss.n10031 0.0702092
R23485 vss.n10023 vss.n10022 0.0702092
R23486 vss.n10024 vss.n10023 0.0702092
R23487 vss.n10020 vss.n10019 0.0702092
R23488 vss.n10019 vss.n10018 0.0702092
R23489 vss.n10017 vss.n10016 0.0702092
R23490 vss.n10018 vss.n10017 0.0702092
R23491 vss.n10026 vss.n10025 0.0702092
R23492 vss.n10025 vss.n10024 0.0702092
R23493 vss.n10030 vss.n10029 0.0702092
R23494 vss.n10031 vss.n10030 0.0702092
R23495 vss.n9995 vss.n9993 0.0702092
R23496 vss.n9993 vss.n9992 0.0702092
R23497 vss.n11633 vss.n11622 0.0702092
R23498 vss.n11633 vss.n11632 0.0702092
R23499 vss.n11636 vss.n11635 0.0702092
R23500 vss.n11635 vss.n9960 0.0702092
R23501 vss.n9963 vss.n9959 0.0702092
R23502 vss.n11641 vss.n9959 0.0702092
R23503 vss.n9951 vss.n9949 0.0702092
R23504 vss.n9949 vss.n9948 0.0702092
R23505 vss.n11645 vss.n9950 0.0702092
R23506 vss.n9950 vss.n9948 0.0702092
R23507 vss.n11643 vss.n11642 0.0702092
R23508 vss.n11642 vss.n11641 0.0702092
R23509 vss.n11627 vss.n11626 0.0702092
R23510 vss.n11626 vss.n9960 0.0702092
R23511 vss.n11631 vss.n11630 0.0702092
R23512 vss.n11632 vss.n11631 0.0702092
R23513 vss.n13190 vss.n8870 0.0661418
R23514 vss.n13191 vss.n13190 0.0661418
R23515 vss.n8877 vss.n8876 0.0661418
R23516 vss.n8876 vss.n8874 0.0661418
R23517 vss.n10351 vss.n10348 0.0661418
R23518 vss.n10351 vss.n10350 0.0661418
R23519 vss.n10360 vss.n10359 0.0661418
R23520 vss.n10361 vss.n10360 0.0661418
R23521 vss.n13198 vss.n13197 0.0661418
R23522 vss.n13199 vss.n13198 0.0661418
R23523 vss.n10303 vss.n10298 0.0661418
R23524 vss.n10301 vss.n10298 0.0661418
R23525 vss.n10317 vss.n10316 0.0661418
R23526 vss.n10318 vss.n10317 0.0661418
R23527 vss.n10290 vss.n10285 0.0661418
R23528 vss.n10290 vss.n10289 0.0661418
R23529 vss.n10325 vss.n10324 0.0661418
R23530 vss.n10326 vss.n10325 0.0661418
R23531 vss.n10307 vss.n10299 0.0661418
R23532 vss.n10299 vss.n8864 0.0661418
R23533 vss.n9918 vss.n9911 0.0661418
R23534 vss.n9918 vss.n9916 0.0661418
R23535 vss.n9926 vss.n9924 0.0661418
R23536 vss.n9924 vss.n9923 0.0661418
R23537 vss.n11693 vss.n11692 0.0661418
R23538 vss.n11692 vss.n9917 0.0661418
R23539 vss.n11695 vss.n11694 0.0661418
R23540 vss.n11695 vss.n8839 0.0661418
R23541 vss.n11681 vss.n9925 0.0661418
R23542 vss.n11680 vss.n9925 0.0661418
R23543 vss.n9973 vss.n9966 0.0661418
R23544 vss.n9973 vss.n9971 0.0661418
R23545 vss.n9981 vss.n9979 0.0661418
R23546 vss.n9979 vss.n9978 0.0661418
R23547 vss.n11456 vss.n11455 0.0661418
R23548 vss.n11455 vss.n9972 0.0661418
R23549 vss.n11458 vss.n11457 0.0661418
R23550 vss.n11458 vss.n8843 0.0661418
R23551 vss.n11444 vss.n9980 0.0661418
R23552 vss.n11443 vss.n9980 0.0661418
R23553 vss.n11381 vss.n11380 0.0661418
R23554 vss.n11380 vss.n11375 0.0661418
R23555 vss.n11376 vss.n11370 0.0661418
R23556 vss.n11376 vss.n11374 0.0661418
R23557 vss.n11387 vss.n11386 0.0661418
R23558 vss.n11386 vss.n11384 0.0661418
R23559 vss.n11389 vss.n11388 0.0661418
R23560 vss.n11389 vss.n8840 0.0661418
R23561 vss.n11410 vss.n11409 0.0661418
R23562 vss.n11411 vss.n11410 0.0661418
R23563 vss.n11164 vss.n11157 0.0661418
R23564 vss.n11164 vss.n11162 0.0661418
R23565 vss.n11172 vss.n11170 0.0661418
R23566 vss.n11170 vss.n11169 0.0661418
R23567 vss.n11187 vss.n11186 0.0661418
R23568 vss.n11186 vss.n11163 0.0661418
R23569 vss.n11189 vss.n11188 0.0661418
R23570 vss.n11189 vss.n8847 0.0661418
R23571 vss.n11175 vss.n11171 0.0661418
R23572 vss.n11171 vss.n10055 0.0661418
R23573 vss.n10133 vss.n10126 0.0661418
R23574 vss.n10133 vss.n10131 0.0661418
R23575 vss.n10141 vss.n10139 0.0661418
R23576 vss.n10139 vss.n10138 0.0661418
R23577 vss.n11051 vss.n11050 0.0661418
R23578 vss.n11050 vss.n10132 0.0661418
R23579 vss.n11053 vss.n11052 0.0661418
R23580 vss.n11053 vss.n8851 0.0661418
R23581 vss.n11039 vss.n10140 0.0661418
R23582 vss.n11038 vss.n10140 0.0661418
R23583 vss.n10087 vss.n10080 0.0661418
R23584 vss.n10087 vss.n10085 0.0661418
R23585 vss.n10095 vss.n10093 0.0661418
R23586 vss.n10093 vss.n10092 0.0661418
R23587 vss.n10111 vss.n10110 0.0661418
R23588 vss.n10110 vss.n10086 0.0661418
R23589 vss.n10113 vss.n10112 0.0661418
R23590 vss.n10113 vss.n8848 0.0661418
R23591 vss.n10099 vss.n10094 0.0661418
R23592 vss.n10098 vss.n10094 0.0661418
R23593 vss.n10723 vss.n10722 0.0661418
R23594 vss.n10723 vss.n10719 0.0661418
R23595 vss.n10720 vss.n10714 0.0661418
R23596 vss.n10720 vss.n10718 0.0661418
R23597 vss.n10729 vss.n10728 0.0661418
R23598 vss.n10728 vss.n10726 0.0661418
R23599 vss.n10731 vss.n10730 0.0661418
R23600 vss.n10731 vss.n8855 0.0661418
R23601 vss.n10753 vss.n10752 0.0661418
R23602 vss.n10754 vss.n10753 0.0661418
R23603 vss.n10220 vss.n10213 0.0661418
R23604 vss.n10220 vss.n10218 0.0661418
R23605 vss.n10228 vss.n10226 0.0661418
R23606 vss.n10226 vss.n10225 0.0661418
R23607 vss.n10799 vss.n10798 0.0661418
R23608 vss.n10798 vss.n10219 0.0661418
R23609 vss.n10801 vss.n10800 0.0661418
R23610 vss.n10801 vss.n8859 0.0661418
R23611 vss.n10787 vss.n10227 0.0661418
R23612 vss.n10786 vss.n10227 0.0661418
R23613 vss.n10669 vss.n10668 0.0661418
R23614 vss.n10668 vss.n10663 0.0661418
R23615 vss.n10664 vss.n10658 0.0661418
R23616 vss.n10664 vss.n10662 0.0661418
R23617 vss.n10675 vss.n10674 0.0661418
R23618 vss.n10674 vss.n10672 0.0661418
R23619 vss.n10677 vss.n10676 0.0661418
R23620 vss.n10677 vss.n8856 0.0661418
R23621 vss.n10698 vss.n10697 0.0661418
R23622 vss.n10699 vss.n10698 0.0661418
R23623 vss.n10262 vss.n10255 0.0661418
R23624 vss.n10262 vss.n10260 0.0661418
R23625 vss.n10270 vss.n10268 0.0661418
R23626 vss.n10268 vss.n10267 0.0661418
R23627 vss.n10409 vss.n10408 0.0661418
R23628 vss.n10408 vss.n10261 0.0661418
R23629 vss.n10411 vss.n10410 0.0661418
R23630 vss.n10411 vss.n8863 0.0661418
R23631 vss.n10397 vss.n10269 0.0661418
R23632 vss.n10396 vss.n10269 0.0661418
R23633 vss.n11909 vss.n11908 0.0661418
R23634 vss.n11908 vss.n11906 0.0661418
R23635 vss.n11903 vss.n11902 0.0661418
R23636 vss.n11902 vss.n11897 0.0661418
R23637 vss.n11900 vss.n11893 0.0661418
R23638 vss.n11900 vss.n11898 0.0661418
R23639 vss.n11933 vss.n11932 0.0661418
R23640 vss.n11934 vss.n11933 0.0661418
R23641 vss.n11911 vss.n11910 0.0661418
R23642 vss.n11911 vss.n8808 0.0661418
R23643 vss.n8891 vss.n8884 0.0661418
R23644 vss.n8891 vss.n8889 0.0661418
R23645 vss.n8896 vss.n8895 0.0661418
R23646 vss.n8895 vss.n8890 0.0661418
R23647 vss.n9269 vss.n9268 0.0661418
R23648 vss.n9268 vss.n9257 0.0661418
R23649 vss.n9260 vss.n9256 0.0661418
R23650 vss.n9274 vss.n9256 0.0661418
R23651 vss.n8898 vss.n8897 0.0661418
R23652 vss.n13164 vss.n8898 0.0661418
R23653 vss.n12389 vss.n12382 0.0661418
R23654 vss.n12389 vss.n12387 0.0661418
R23655 vss.n12412 vss.n12411 0.0661418
R23656 vss.n12411 vss.n12388 0.0661418
R23657 vss.n12397 vss.n12395 0.0661418
R23658 vss.n12395 vss.n12394 0.0661418
R23659 vss.n12400 vss.n12396 0.0661418
R23660 vss.n12396 vss.n9205 0.0661418
R23661 vss.n12414 vss.n12413 0.0661418
R23662 vss.n12415 vss.n12414 0.0661418
R23663 vss.n8626 vss.n8619 0.0661418
R23664 vss.n8626 vss.n8624 0.0661418
R23665 vss.n13274 vss.n13273 0.0661418
R23666 vss.n13273 vss.n8625 0.0661418
R23667 vss.n8634 vss.n8632 0.0661418
R23668 vss.n8632 vss.n8631 0.0661418
R23669 vss.n13262 vss.n8633 0.0661418
R23670 vss.n13261 vss.n8633 0.0661418
R23671 vss.n13276 vss.n13275 0.0661418
R23672 vss.n13276 vss.n8440 0.0661418
R23673 vss.n12271 vss.n12264 0.0661418
R23674 vss.n12271 vss.n12269 0.0661418
R23675 vss.n12294 vss.n12293 0.0661418
R23676 vss.n12293 vss.n12270 0.0661418
R23677 vss.n12279 vss.n12277 0.0661418
R23678 vss.n12277 vss.n12276 0.0661418
R23679 vss.n12282 vss.n12278 0.0661418
R23680 vss.n12278 vss.n8688 0.0661418
R23681 vss.n12296 vss.n12295 0.0661418
R23682 vss.n12297 vss.n12296 0.0661418
R23683 vss.n8347 vss.n8340 0.0661418
R23684 vss.n8347 vss.n8345 0.0661418
R23685 vss.n8352 vss.n8351 0.0661418
R23686 vss.n8351 vss.n8346 0.0661418
R23687 vss.n8751 vss.n8750 0.0661418
R23688 vss.n8750 vss.n8739 0.0661418
R23689 vss.n8742 vss.n8738 0.0661418
R23690 vss.n8756 vss.n8738 0.0661418
R23691 vss.n8354 vss.n8353 0.0661418
R23692 vss.n13687 vss.n8354 0.0661418
R23693 vss.n11976 vss.n11975 0.0661418
R23694 vss.n11975 vss.n11970 0.0661418
R23695 vss.n11973 vss.n11967 0.0661418
R23696 vss.n11973 vss.n11971 0.0661418
R23697 vss.n11982 vss.n11981 0.0661418
R23698 vss.n11981 vss.n11979 0.0661418
R23699 vss.n11984 vss.n11983 0.0661418
R23700 vss.n11984 vss.n8807 0.0661418
R23701 vss.n12006 vss.n12005 0.0661418
R23702 vss.n12007 vss.n12006 0.0661418
R23703 vss.n12204 vss.n12203 0.0661418
R23704 vss.n12203 vss.n12197 0.0661418
R23705 vss.n12210 vss.n12209 0.0661418
R23706 vss.n12209 vss.n12207 0.0661418
R23707 vss.n12198 vss.n9857 0.0661418
R23708 vss.n12198 vss.n9853 0.0661418
R23709 vss.n9856 vss.n9852 0.0661418
R23710 vss.n12235 vss.n9852 0.0661418
R23711 vss.n8773 vss.n8772 0.0661418
R23712 vss.n8772 vss.n8766 0.0661418
R23713 vss.n8779 vss.n8778 0.0661418
R23714 vss.n8778 vss.n8776 0.0661418
R23715 vss.n8767 vss.n8762 0.0661418
R23716 vss.n8767 vss.n8758 0.0661418
R23717 vss.n8761 vss.n8757 0.0661418
R23718 vss.n8804 vss.n8757 0.0661418
R23719 vss.n8781 vss.n8780 0.0661418
R23720 vss.n8782 vss.n8781 0.0661418
R23721 vss.n8704 vss.n8703 0.0661418
R23722 vss.n8703 vss.n8697 0.0661418
R23723 vss.n8710 vss.n8709 0.0661418
R23724 vss.n8709 vss.n8707 0.0661418
R23725 vss.n8698 vss.n8694 0.0661418
R23726 vss.n8698 vss.n8690 0.0661418
R23727 vss.n8693 vss.n8689 0.0661418
R23728 vss.n8735 vss.n8689 0.0661418
R23729 vss.n8712 vss.n8711 0.0661418
R23730 vss.n8713 vss.n8712 0.0661418
R23731 vss.n9809 vss.n9805 0.0661418
R23732 vss.n9815 vss.n9810 0.0661418
R23733 vss.n9815 vss.n9813 0.0661418
R23734 vss.n9822 vss.n9821 0.0661418
R23735 vss.n9821 vss.n9814 0.0661418
R23736 vss.n9828 vss.n9827 0.0661418
R23737 vss.n9827 vss.n9825 0.0661418
R23738 vss.n9830 vss.n9829 0.0661418
R23739 vss.n9830 vss.n8737 0.0661418
R23740 vss.n9783 vss.n9782 0.0661418
R23741 vss.n9765 vss.n9759 0.0661418
R23742 vss.n9765 vss.n9763 0.0661418
R23743 vss.n9770 vss.n9769 0.0661418
R23744 vss.n9769 vss.n9764 0.0661418
R23745 vss.n9776 vss.n9775 0.0661418
R23746 vss.n9775 vss.n9773 0.0661418
R23747 vss.n9800 vss.n9799 0.0661418
R23748 vss.n9801 vss.n9800 0.0661418
R23749 vss.n9750 vss.n9746 0.0661418
R23750 vss.n9747 vss.n9745 0.0661418
R23751 vss.n9745 vss.n9744 0.0661418
R23752 vss.n9739 vss.n9732 0.0661418
R23753 vss.n9739 vss.n9737 0.0661418
R23754 vss.n12248 vss.n12247 0.0661418
R23755 vss.n12247 vss.n9738 0.0661418
R23756 vss.n12250 vss.n12249 0.0661418
R23757 vss.n12250 vss.n8687 0.0661418
R23758 vss.n12322 vss.n12321 0.0661418
R23759 vss.n12321 vss.n12315 0.0661418
R23760 vss.n12328 vss.n12327 0.0661418
R23761 vss.n12327 vss.n12325 0.0661418
R23762 vss.n12316 vss.n9729 0.0661418
R23763 vss.n12316 vss.n9725 0.0661418
R23764 vss.n9728 vss.n9724 0.0661418
R23765 vss.n12353 vss.n9724 0.0661418
R23766 vss.n12330 vss.n12329 0.0661418
R23767 vss.n8654 vss.n8653 0.0661418
R23768 vss.n8653 vss.n8647 0.0661418
R23769 vss.n8660 vss.n8659 0.0661418
R23770 vss.n8659 vss.n8657 0.0661418
R23771 vss.n8648 vss.n8643 0.0661418
R23772 vss.n8648 vss.n8639 0.0661418
R23773 vss.n8642 vss.n8638 0.0661418
R23774 vss.n8685 vss.n8638 0.0661418
R23775 vss.n8662 vss.n8661 0.0661418
R23776 vss.n8663 vss.n8662 0.0661418
R23777 vss.n9196 vss.n9195 0.0661418
R23778 vss.n9195 vss.n9190 0.0661418
R23779 vss.n9193 vss.n9186 0.0661418
R23780 vss.n9193 vss.n9191 0.0661418
R23781 vss.n9202 vss.n9201 0.0661418
R23782 vss.n9201 vss.n9199 0.0661418
R23783 vss.n9204 vss.n9203 0.0661418
R23784 vss.n12916 vss.n9204 0.0661418
R23785 vss.n12938 vss.n12937 0.0661418
R23786 vss.n12939 vss.n12938 0.0661418
R23787 vss.n9680 vss.n9676 0.0661418
R23788 vss.n9686 vss.n9681 0.0661418
R23789 vss.n9686 vss.n9684 0.0661418
R23790 vss.n9693 vss.n9692 0.0661418
R23791 vss.n9692 vss.n9685 0.0661418
R23792 vss.n9699 vss.n9698 0.0661418
R23793 vss.n9698 vss.n9696 0.0661418
R23794 vss.n9701 vss.n9700 0.0661418
R23795 vss.n9702 vss.n9701 0.0661418
R23796 vss.n9654 vss.n9653 0.0661418
R23797 vss.n9635 vss.n9629 0.0661418
R23798 vss.n9635 vss.n9633 0.0661418
R23799 vss.n9640 vss.n9639 0.0661418
R23800 vss.n9639 vss.n9634 0.0661418
R23801 vss.n9646 vss.n9645 0.0661418
R23802 vss.n9645 vss.n9643 0.0661418
R23803 vss.n9671 vss.n9670 0.0661418
R23804 vss.n9672 vss.n9671 0.0661418
R23805 vss.n9620 vss.n9616 0.0661418
R23806 vss.n9617 vss.n9615 0.0661418
R23807 vss.n9615 vss.n9614 0.0661418
R23808 vss.n9609 vss.n9602 0.0661418
R23809 vss.n9609 vss.n9607 0.0661418
R23810 vss.n12366 vss.n12365 0.0661418
R23811 vss.n12365 vss.n9608 0.0661418
R23812 vss.n12368 vss.n12367 0.0661418
R23813 vss.n12368 vss.n9207 0.0661418
R23814 vss.n12441 vss.n12440 0.0661418
R23815 vss.n12440 vss.n12434 0.0661418
R23816 vss.n12447 vss.n12446 0.0661418
R23817 vss.n12446 vss.n12444 0.0661418
R23818 vss.n12435 vss.n9599 0.0661418
R23819 vss.n12435 vss.n9595 0.0661418
R23820 vss.n9598 vss.n9594 0.0661418
R23821 vss.n12472 vss.n9594 0.0661418
R23822 vss.n12449 vss.n12448 0.0661418
R23823 vss.n9224 vss.n9223 0.0661418
R23824 vss.n9223 vss.n9217 0.0661418
R23825 vss.n9230 vss.n9229 0.0661418
R23826 vss.n9229 vss.n9227 0.0661418
R23827 vss.n9218 vss.n9213 0.0661418
R23828 vss.n9218 vss.n9209 0.0661418
R23829 vss.n9212 vss.n9208 0.0661418
R23830 vss.n9255 vss.n9208 0.0661418
R23831 vss.n9232 vss.n9231 0.0661418
R23832 vss.n9233 vss.n9232 0.0661418
R23833 vss.n9326 vss.n9325 0.0661418
R23834 vss.n9325 vss.n9320 0.0661418
R23835 vss.n9323 vss.n9315 0.0661418
R23836 vss.n9323 vss.n9321 0.0661418
R23837 vss.n9332 vss.n9331 0.0661418
R23838 vss.n9331 vss.n9329 0.0661418
R23839 vss.n9334 vss.n9333 0.0661418
R23840 vss.n9334 vss.n9281 0.0661418
R23841 vss.n9356 vss.n9355 0.0661418
R23842 vss.n9357 vss.n9356 0.0661418
R23843 vss.n12512 vss.n12511 0.0661418
R23844 vss.n12511 vss.n12506 0.0661418
R23845 vss.n12509 vss.n9422 0.0661418
R23846 vss.n12509 vss.n12507 0.0661418
R23847 vss.n12518 vss.n12517 0.0661418
R23848 vss.n12517 vss.n12515 0.0661418
R23849 vss.n12520 vss.n12519 0.0661418
R23850 vss.n12520 vss.n9278 0.0661418
R23851 vss.n12542 vss.n12541 0.0661418
R23852 vss.n12543 vss.n12542 0.0661418
R23853 vss.n12662 vss.n12661 0.0661418
R23854 vss.n12661 vss.n12656 0.0661418
R23855 vss.n12659 vss.n12652 0.0661418
R23856 vss.n12659 vss.n12657 0.0661418
R23857 vss.n12668 vss.n12667 0.0661418
R23858 vss.n12667 vss.n12665 0.0661418
R23859 vss.n12670 vss.n12669 0.0661418
R23860 vss.n12670 vss.n9277 0.0661418
R23861 vss.n12692 vss.n12691 0.0661418
R23862 vss.n12693 vss.n12692 0.0661418
R23863 vss.n9551 vss.n9547 0.0661418
R23864 vss.n9557 vss.n9552 0.0661418
R23865 vss.n9557 vss.n9555 0.0661418
R23866 vss.n9564 vss.n9563 0.0661418
R23867 vss.n9563 vss.n9556 0.0661418
R23868 vss.n9570 vss.n9569 0.0661418
R23869 vss.n9569 vss.n9567 0.0661418
R23870 vss.n9572 vss.n9571 0.0661418
R23871 vss.n9572 vss.n9276 0.0661418
R23872 vss.n9524 vss.n9523 0.0661418
R23873 vss.n9506 vss.n9500 0.0661418
R23874 vss.n9506 vss.n9504 0.0661418
R23875 vss.n9511 vss.n9510 0.0661418
R23876 vss.n9510 vss.n9505 0.0661418
R23877 vss.n9517 vss.n9516 0.0661418
R23878 vss.n9516 vss.n9514 0.0661418
R23879 vss.n9541 vss.n9540 0.0661418
R23880 vss.n9542 vss.n9541 0.0661418
R23881 vss.n9491 vss.n9487 0.0661418
R23882 vss.n9488 vss.n9486 0.0661418
R23883 vss.n9486 vss.n9485 0.0661418
R23884 vss.n9480 vss.n9473 0.0661418
R23885 vss.n9480 vss.n9478 0.0661418
R23886 vss.n12485 vss.n12484 0.0661418
R23887 vss.n12484 vss.n9479 0.0661418
R23888 vss.n12487 vss.n12486 0.0661418
R23889 vss.n12487 vss.n9280 0.0661418
R23890 vss.n9456 vss.n9455 0.0661418
R23891 vss.n9438 vss.n9436 0.0661418
R23892 vss.n9436 vss.n9435 0.0661418
R23893 vss.n9430 vss.n9423 0.0661418
R23894 vss.n9430 vss.n9428 0.0661418
R23895 vss.n9454 vss.n9453 0.0661418
R23896 vss.n9453 vss.n9429 0.0661418
R23897 vss.n9442 vss.n9437 0.0661418
R23898 vss.n9441 vss.n9437 0.0661418
R23899 vss.n10202 vss.n9546 0.0661418
R23900 vss.n11099 vss.n9675 0.0661418
R23901 vss.n11504 vss.n9804 0.0661418
R23902 vss.n11727 vss.n9875 0.0661418
R23903 vss.n11731 vss.n9875 0.0661418
R23904 vss.n9876 vss.n9874 0.0661418
R23905 vss.n9874 vss.n9873 0.0661418
R23906 vss.n9868 vss.n9861 0.0661418
R23907 vss.n9868 vss.n9866 0.0661418
R23908 vss.n11742 vss.n11741 0.0661418
R23909 vss.n11741 vss.n9867 0.0661418
R23910 vss.n11744 vss.n11743 0.0661418
R23911 vss.n11744 vss.n8806 0.0661418
R23912 vss.n12212 vss.n12211 0.0661418
R23913 vss.n11836 vss.n11835 0.0661418
R23914 vss.n11835 vss.n11808 0.0661418
R23915 vss.n11817 vss.n11803 0.0661418
R23916 vss.n11817 vss.n11808 0.0661418
R23917 vss.n11824 vss.n11823 0.0661418
R23918 vss.n11823 vss.n11808 0.0661418
R23919 vss.n11829 vss.n11822 0.0661418
R23920 vss.n11822 vss.n11808 0.0661418
R23921 vss.n11813 vss.n11811 0.0661418
R23922 vss.n11811 vss.n11808 0.0661418
R23923 vss.n3982 vss.n3981 0.0661418
R23924 vss.n3981 vss.n3980 0.0661418
R23925 vss.n7 vss.n0 0.0661418
R23926 vss.n7 vss.n5 0.0661418
R23927 vss.n12 vss.n11 0.0661418
R23928 vss.n11 vss.n6 0.0661418
R23929 vss.n14 vss.n13 0.0661418
R23930 vss.n15891 vss.n14 0.0661418
R23931 vss.n3986 vss.n3985 0.0661418
R23932 vss.n3987 vss.n3986 0.0661418
R23933 vss.n5639 vss.n5632 0.0661418
R23934 vss.n5639 vss.n5637 0.0661418
R23935 vss.n5662 vss.n5661 0.0661418
R23936 vss.n5661 vss.n5638 0.0661418
R23937 vss.n5647 vss.n5645 0.0661418
R23938 vss.n5645 vss.n5644 0.0661418
R23939 vss.n5650 vss.n5646 0.0661418
R23940 vss.n5646 vss.n3660 0.0661418
R23941 vss.n5664 vss.n5663 0.0661418
R23942 vss.n5664 vss.n224 0.0661418
R23943 vss.n172 vss.n165 0.0661418
R23944 vss.n172 vss.n170 0.0661418
R23945 vss.n177 vss.n176 0.0661418
R23946 vss.n176 vss.n171 0.0661418
R23947 vss.n3723 vss.n3722 0.0661418
R23948 vss.n3722 vss.n3711 0.0661418
R23949 vss.n3714 vss.n3710 0.0661418
R23950 vss.n3728 vss.n3710 0.0661418
R23951 vss.n179 vss.n178 0.0661418
R23952 vss.n15744 vss.n179 0.0661418
R23953 vss.n3678 vss.n3677 0.0661418
R23954 vss.n3677 vss.n3671 0.0661418
R23955 vss.n3684 vss.n3683 0.0661418
R23956 vss.n3683 vss.n3681 0.0661418
R23957 vss.n3672 vss.n3668 0.0661418
R23958 vss.n3672 vss.n3664 0.0661418
R23959 vss.n3667 vss.n3663 0.0661418
R23960 vss.n3709 vss.n3663 0.0661418
R23961 vss.n3686 vss.n3685 0.0661418
R23962 vss.n3687 vss.n3686 0.0661418
R23963 vss.n5831 vss.n5824 0.0661418
R23964 vss.n5831 vss.n5829 0.0661418
R23965 vss.n5854 vss.n5853 0.0661418
R23966 vss.n5853 vss.n5830 0.0661418
R23967 vss.n5839 vss.n5837 0.0661418
R23968 vss.n5837 vss.n5836 0.0661418
R23969 vss.n5842 vss.n5838 0.0661418
R23970 vss.n5838 vss.n3779 0.0661418
R23971 vss.n5856 vss.n5855 0.0661418
R23972 vss.n5856 vss.n146 0.0661418
R23973 vss.n94 vss.n87 0.0661418
R23974 vss.n94 vss.n92 0.0661418
R23975 vss.n99 vss.n98 0.0661418
R23976 vss.n98 vss.n93 0.0661418
R23977 vss.n3842 vss.n3841 0.0661418
R23978 vss.n3841 vss.n3830 0.0661418
R23979 vss.n3833 vss.n3829 0.0661418
R23980 vss.n3847 vss.n3829 0.0661418
R23981 vss.n101 vss.n100 0.0661418
R23982 vss.n15800 vss.n101 0.0661418
R23983 vss.n3797 vss.n3796 0.0661418
R23984 vss.n3796 vss.n3790 0.0661418
R23985 vss.n3803 vss.n3802 0.0661418
R23986 vss.n3802 vss.n3800 0.0661418
R23987 vss.n3791 vss.n3787 0.0661418
R23988 vss.n3791 vss.n3783 0.0661418
R23989 vss.n3786 vss.n3782 0.0661418
R23990 vss.n3828 vss.n3782 0.0661418
R23991 vss.n3805 vss.n3804 0.0661418
R23992 vss.n3806 vss.n3805 0.0661418
R23993 vss.n3916 vss.n3915 0.0661418
R23994 vss.n3915 vss.n3909 0.0661418
R23995 vss.n3922 vss.n3921 0.0661418
R23996 vss.n3921 vss.n3919 0.0661418
R23997 vss.n3910 vss.n3906 0.0661418
R23998 vss.n3910 vss.n3902 0.0661418
R23999 vss.n3905 vss.n3901 0.0661418
R24000 vss.n3947 vss.n3901 0.0661418
R24001 vss.n3924 vss.n3923 0.0661418
R24002 vss.n3925 vss.n3924 0.0661418
R24003 vss.n6071 vss.n6064 0.0661418
R24004 vss.n6071 vss.n6069 0.0661418
R24005 vss.n6094 vss.n6093 0.0661418
R24006 vss.n6093 vss.n6070 0.0661418
R24007 vss.n6079 vss.n6077 0.0661418
R24008 vss.n6077 vss.n6076 0.0661418
R24009 vss.n6082 vss.n6078 0.0661418
R24010 vss.n6078 vss.n3898 0.0661418
R24011 vss.n6096 vss.n6095 0.0661418
R24012 vss.n6096 vss.n67 0.0661418
R24013 vss.n3547 vss.n3540 0.0661418
R24014 vss.n3547 vss.n3545 0.0661418
R24015 vss.n3552 vss.n3551 0.0661418
R24016 vss.n3551 vss.n3546 0.0661418
R24017 vss.n3558 vss.n3557 0.0661418
R24018 vss.n3557 vss.n3555 0.0661418
R24019 vss.n6331 vss.n6330 0.0661418
R24020 vss.n6332 vss.n6331 0.0661418
R24021 vss.n5605 vss.n3487 0.0661418
R24022 vss.n5606 vss.n5601 0.0661418
R24023 vss.n5601 vss.n5600 0.0661418
R24024 vss.n5595 vss.n5588 0.0661418
R24025 vss.n5595 vss.n5593 0.0661418
R24026 vss.n5617 vss.n5616 0.0661418
R24027 vss.n5616 vss.n5594 0.0661418
R24028 vss.n5619 vss.n5618 0.0661418
R24029 vss.n5619 vss.n3662 0.0661418
R24030 vss.n5699 vss.n5698 0.0661418
R24031 vss.n5686 vss.n5540 0.0661418
R24032 vss.n5686 vss.n5684 0.0661418
R24033 vss.n5691 vss.n5690 0.0661418
R24034 vss.n5690 vss.n5685 0.0661418
R24035 vss.n5697 vss.n5696 0.0661418
R24036 vss.n5696 vss.n5694 0.0661418
R24037 vss.n5721 vss.n5720 0.0661418
R24038 vss.n5722 vss.n5721 0.0661418
R24039 vss.n5560 vss.n5555 0.0661418
R24040 vss.n5561 vss.n5554 0.0661418
R24041 vss.n5554 vss.n5553 0.0661418
R24042 vss.n5548 vss.n5541 0.0661418
R24043 vss.n5548 vss.n5546 0.0661418
R24044 vss.n5572 vss.n5571 0.0661418
R24045 vss.n5571 vss.n5547 0.0661418
R24046 vss.n5574 vss.n5573 0.0661418
R24047 vss.n5574 vss.n3730 0.0661418
R24048 vss.n5937 vss.n5936 0.0661418
R24049 vss.n5924 vss.n5917 0.0661418
R24050 vss.n5924 vss.n5922 0.0661418
R24051 vss.n5929 vss.n5928 0.0661418
R24052 vss.n5928 vss.n5923 0.0661418
R24053 vss.n5935 vss.n5934 0.0661418
R24054 vss.n5934 vss.n5932 0.0661418
R24055 vss.n5959 vss.n5958 0.0661418
R24056 vss.n5960 vss.n5959 0.0661418
R24057 vss.n5727 vss.n4003 0.0661418
R24058 vss.n5876 vss.n5728 0.0661418
R24059 vss.n5876 vss.n5874 0.0661418
R24060 vss.n5883 vss.n5882 0.0661418
R24061 vss.n5882 vss.n5875 0.0661418
R24062 vss.n5889 vss.n5888 0.0661418
R24063 vss.n5888 vss.n5886 0.0661418
R24064 vss.n5891 vss.n5890 0.0661418
R24065 vss.n5891 vss.n3781 0.0661418
R24066 vss.n5808 vss.n5807 0.0661418
R24067 vss.n5791 vss.n5789 0.0661418
R24068 vss.n5789 vss.n5788 0.0661418
R24069 vss.n5783 vss.n5776 0.0661418
R24070 vss.n5783 vss.n5781 0.0661418
R24071 vss.n5806 vss.n5805 0.0661418
R24072 vss.n5805 vss.n5782 0.0661418
R24073 vss.n5794 vss.n5790 0.0661418
R24074 vss.n5790 vss.n3999 0.0661418
R24075 vss.n5748 vss.n5743 0.0661418
R24076 vss.n5749 vss.n5742 0.0661418
R24077 vss.n5742 vss.n5741 0.0661418
R24078 vss.n5736 vss.n5729 0.0661418
R24079 vss.n5736 vss.n5734 0.0661418
R24080 vss.n5760 vss.n5759 0.0661418
R24081 vss.n5759 vss.n5735 0.0661418
R24082 vss.n5762 vss.n5761 0.0661418
R24083 vss.n5762 vss.n3849 0.0661418
R24084 vss.n6176 vss.n6175 0.0661418
R24085 vss.n6163 vss.n6156 0.0661418
R24086 vss.n6163 vss.n6161 0.0661418
R24087 vss.n6168 vss.n6167 0.0661418
R24088 vss.n6167 vss.n6162 0.0661418
R24089 vss.n6174 vss.n6173 0.0661418
R24090 vss.n6173 vss.n6171 0.0661418
R24091 vss.n6198 vss.n6197 0.0661418
R24092 vss.n6199 vss.n6198 0.0661418
R24093 vss.n5967 vss.n3995 0.0661418
R24094 vss.n6115 vss.n5968 0.0661418
R24095 vss.n6115 vss.n6113 0.0661418
R24096 vss.n6122 vss.n6121 0.0661418
R24097 vss.n6121 vss.n6114 0.0661418
R24098 vss.n6128 vss.n6127 0.0661418
R24099 vss.n6127 vss.n6125 0.0661418
R24100 vss.n6130 vss.n6129 0.0661418
R24101 vss.n6130 vss.n3900 0.0661418
R24102 vss.n6048 vss.n6047 0.0661418
R24103 vss.n6031 vss.n6029 0.0661418
R24104 vss.n6029 vss.n6028 0.0661418
R24105 vss.n6023 vss.n6016 0.0661418
R24106 vss.n6023 vss.n6021 0.0661418
R24107 vss.n6046 vss.n6045 0.0661418
R24108 vss.n6045 vss.n6022 0.0661418
R24109 vss.n6034 vss.n6030 0.0661418
R24110 vss.n6030 vss.n3991 0.0661418
R24111 vss.n5989 vss.n5982 0.0661418
R24112 vss.n5982 vss.n5981 0.0661418
R24113 vss.n5976 vss.n5969 0.0661418
R24114 vss.n5976 vss.n5974 0.0661418
R24115 vss.n6000 vss.n5999 0.0661418
R24116 vss.n5999 vss.n5975 0.0661418
R24117 vss.n6002 vss.n6001 0.0661418
R24118 vss.n6002 vss.n3968 0.0661418
R24119 vss.n5988 vss.n5983 0.0661418
R24120 vss.n4381 vss.n4380 0.0661418
R24121 vss.n4380 vss.n4375 0.0661418
R24122 vss.n4376 vss.n4370 0.0661418
R24123 vss.n4376 vss.n4374 0.0661418
R24124 vss.n4387 vss.n4386 0.0661418
R24125 vss.n4386 vss.n4384 0.0661418
R24126 vss.n4389 vss.n4388 0.0661418
R24127 vss.n4389 vss.n3309 0.0661418
R24128 vss.n4552 vss.n4551 0.0661418
R24129 vss.n4553 vss.n4552 0.0661418
R24130 vss.n6622 vss.n6615 0.0661418
R24131 vss.n6622 vss.n6620 0.0661418
R24132 vss.n6630 vss.n6628 0.0661418
R24133 vss.n6628 vss.n6627 0.0661418
R24134 vss.n6645 vss.n6644 0.0661418
R24135 vss.n6644 vss.n6621 0.0661418
R24136 vss.n6647 vss.n6646 0.0661418
R24137 vss.n6647 vss.n3333 0.0661418
R24138 vss.n6633 vss.n6629 0.0661418
R24139 vss.n6629 vss.n1075 0.0661418
R24140 vss.n6504 vss.n6497 0.0661418
R24141 vss.n6504 vss.n6502 0.0661418
R24142 vss.n6512 vss.n6510 0.0661418
R24143 vss.n6510 vss.n6509 0.0661418
R24144 vss.n6596 vss.n6595 0.0661418
R24145 vss.n6595 vss.n6503 0.0661418
R24146 vss.n6598 vss.n6597 0.0661418
R24147 vss.n6599 vss.n6598 0.0661418
R24148 vss.n6584 vss.n6511 0.0661418
R24149 vss.n6583 vss.n6511 0.0661418
R24150 vss.n5220 vss.n5213 0.0661418
R24151 vss.n5220 vss.n5218 0.0661418
R24152 vss.n5228 vss.n5226 0.0661418
R24153 vss.n5226 vss.n5225 0.0661418
R24154 vss.n5243 vss.n5242 0.0661418
R24155 vss.n5242 vss.n5219 0.0661418
R24156 vss.n5245 vss.n5244 0.0661418
R24157 vss.n5245 vss.n3325 0.0661418
R24158 vss.n5231 vss.n5227 0.0661418
R24159 vss.n5227 vss.n795 0.0661418
R24160 vss.n4071 vss.n4002 0.0661418
R24161 vss.n5432 vss.n5425 0.0661418
R24162 vss.n5432 vss.n5430 0.0661418
R24163 vss.n5440 vss.n5438 0.0661418
R24164 vss.n5438 vss.n5437 0.0661418
R24165 vss.n5455 vss.n5454 0.0661418
R24166 vss.n5454 vss.n5431 0.0661418
R24167 vss.n5457 vss.n5456 0.0661418
R24168 vss.n5457 vss.n3321 0.0661418
R24169 vss.n5443 vss.n5439 0.0661418
R24170 vss.n5439 vss.n742 0.0661418
R24171 vss.n5317 vss.n5310 0.0661418
R24172 vss.n5317 vss.n5315 0.0661418
R24173 vss.n5325 vss.n5323 0.0661418
R24174 vss.n5323 vss.n5322 0.0661418
R24175 vss.n5408 vss.n5407 0.0661418
R24176 vss.n5407 vss.n5316 0.0661418
R24177 vss.n5410 vss.n5409 0.0661418
R24178 vss.n5410 vss.n3324 0.0661418
R24179 vss.n5396 vss.n5324 0.0661418
R24180 vss.n5395 vss.n5324 0.0661418
R24181 vss.n4135 vss.n4128 0.0661418
R24182 vss.n4135 vss.n4133 0.0661418
R24183 vss.n4143 vss.n4141 0.0661418
R24184 vss.n4141 vss.n4140 0.0661418
R24185 vss.n4158 vss.n4157 0.0661418
R24186 vss.n4157 vss.n4134 0.0661418
R24187 vss.n4160 vss.n4159 0.0661418
R24188 vss.n4160 vss.n3317 0.0661418
R24189 vss.n4146 vss.n4142 0.0661418
R24190 vss.n4142 vss.n643 0.0661418
R24191 vss.n4252 vss.n3994 0.0661418
R24192 vss.n4958 vss.n4951 0.0661418
R24193 vss.n4958 vss.n4956 0.0661418
R24194 vss.n4966 vss.n4964 0.0661418
R24195 vss.n4964 vss.n4963 0.0661418
R24196 vss.n4981 vss.n4980 0.0661418
R24197 vss.n4980 vss.n4957 0.0661418
R24198 vss.n4983 vss.n4982 0.0661418
R24199 vss.n4983 vss.n3313 0.0661418
R24200 vss.n4969 vss.n4965 0.0661418
R24201 vss.n4965 vss.n537 0.0661418
R24202 vss.n4089 vss.n4082 0.0661418
R24203 vss.n4089 vss.n4087 0.0661418
R24204 vss.n4097 vss.n4095 0.0661418
R24205 vss.n4095 vss.n4094 0.0661418
R24206 vss.n4112 vss.n4111 0.0661418
R24207 vss.n4111 vss.n4088 0.0661418
R24208 vss.n4114 vss.n4113 0.0661418
R24209 vss.n4114 vss.n3316 0.0661418
R24210 vss.n4100 vss.n4096 0.0661418
R24211 vss.n4096 vss.n628 0.0661418
R24212 vss.n4272 vss.n4265 0.0661418
R24213 vss.n4272 vss.n4270 0.0661418
R24214 vss.n4280 vss.n4278 0.0661418
R24215 vss.n4278 vss.n4277 0.0661418
R24216 vss.n4933 vss.n4932 0.0661418
R24217 vss.n4932 vss.n4271 0.0661418
R24218 vss.n4935 vss.n4934 0.0661418
R24219 vss.n4935 vss.n3312 0.0661418
R24220 vss.n4921 vss.n4279 0.0661418
R24221 vss.n4920 vss.n4279 0.0661418
R24222 vss.n5105 vss.n5098 0.0661418
R24223 vss.n5105 vss.n5103 0.0661418
R24224 vss.n5113 vss.n5111 0.0661418
R24225 vss.n5111 vss.n5110 0.0661418
R24226 vss.n5196 vss.n5195 0.0661418
R24227 vss.n5195 vss.n5104 0.0661418
R24228 vss.n5198 vss.n5197 0.0661418
R24229 vss.n5198 vss.n3320 0.0661418
R24230 vss.n5184 vss.n5112 0.0661418
R24231 vss.n5183 vss.n5112 0.0661418
R24232 vss.n3348 vss.n3341 0.0661418
R24233 vss.n3348 vss.n3346 0.0661418
R24234 vss.n3356 vss.n3354 0.0661418
R24235 vss.n3354 vss.n3353 0.0661418
R24236 vss.n3371 vss.n3370 0.0661418
R24237 vss.n3370 vss.n3347 0.0661418
R24238 vss.n3373 vss.n3372 0.0661418
R24239 vss.n3373 vss.n3328 0.0661418
R24240 vss.n3359 vss.n3355 0.0661418
R24241 vss.n3355 vss.n885 0.0661418
R24242 vss.n3395 vss.n3388 0.0661418
R24243 vss.n3395 vss.n3393 0.0661418
R24244 vss.n3403 vss.n3401 0.0661418
R24245 vss.n3401 vss.n3400 0.0661418
R24246 vss.n3418 vss.n3417 0.0661418
R24247 vss.n3417 vss.n3394 0.0661418
R24248 vss.n3420 vss.n3419 0.0661418
R24249 vss.n3420 vss.n3329 0.0661418
R24250 vss.n3406 vss.n3402 0.0661418
R24251 vss.n3402 vss.n900 0.0661418
R24252 vss.n3533 vss.n3532 0.0661418
R24253 vss.n6389 vss.n6382 0.0661418
R24254 vss.n6389 vss.n6387 0.0661418
R24255 vss.n6397 vss.n6395 0.0661418
R24256 vss.n6395 vss.n6394 0.0661418
R24257 vss.n6480 vss.n6479 0.0661418
R24258 vss.n6479 vss.n6388 0.0661418
R24259 vss.n6482 vss.n6481 0.0661418
R24260 vss.n6482 vss.n3332 0.0661418
R24261 vss.n6468 vss.n6396 0.0661418
R24262 vss.n6467 vss.n6396 0.0661418
R24263 vss.n6688 vss.n6687 0.0661418
R24264 vss.n6689 vss.n6688 0.0661418
R24265 vss.n6673 vss.n6672 0.0661418
R24266 vss.n6672 vss.n6665 0.0661418
R24267 vss.n6666 vss.n3340 0.0661418
R24268 vss.n6666 vss.n3335 0.0661418
R24269 vss.n6683 vss.n6680 0.0661418
R24270 vss.n6683 vss.n378 0.0661418
R24271 vss.n3339 vss.n3337 0.0661418
R24272 vss.n6336 vss.n3437 0.0661418
R24273 vss.n6336 vss.n6335 0.0661418
R24274 vss.n6359 vss.n3434 0.0661418
R24275 vss.n6360 vss.n6359 0.0661418
R24276 vss.n6348 vss.n6341 0.0661418
R24277 vss.n6344 vss.n6341 0.0661418
R24278 vss.n6346 vss.n6342 0.0661418
R24279 vss.n6342 vss.n3334 0.0661418
R24280 vss.n3440 vss.n3438 0.0661418
R24281 vss.n3477 vss.n3445 0.0661418
R24282 vss.n3478 vss.n3477 0.0661418
R24283 vss.n3451 vss.n3450 0.0661418
R24284 vss.n3451 vss.n3449 0.0661418
R24285 vss.n3457 vss.n3456 0.0661418
R24286 vss.n3456 vss.n3454 0.0661418
R24287 vss.n3485 vss.n3484 0.0661418
R24288 vss.n3486 vss.n3485 0.0661418
R24289 vss.n3459 vss.n3458 0.0661418
R24290 vss.n3525 vss.n3492 0.0661418
R24291 vss.n3526 vss.n3525 0.0661418
R24292 vss.n3499 vss.n3498 0.0661418
R24293 vss.n3498 vss.n3496 0.0661418
R24294 vss.n3505 vss.n3504 0.0661418
R24295 vss.n3504 vss.n3502 0.0661418
R24296 vss.n3507 vss.n3506 0.0661418
R24297 vss.n3507 vss.n3330 0.0661418
R24298 vss.n5289 vss.n5288 0.0661418
R24299 vss.n5288 vss.n5264 0.0661418
R24300 vss.n5265 vss.n5258 0.0661418
R24301 vss.n5265 vss.n5263 0.0661418
R24302 vss.n5273 vss.n5271 0.0661418
R24303 vss.n5271 vss.n5270 0.0661418
R24304 vss.n5291 vss.n5290 0.0661418
R24305 vss.n5294 vss.n5291 0.0661418
R24306 vss.n5276 vss.n5272 0.0661418
R24307 vss.n4011 vss.n4010 0.0661418
R24308 vss.n5524 vss.n4011 0.0661418
R24309 vss.n4017 vss.n4016 0.0661418
R24310 vss.n4016 vss.n4014 0.0661418
R24311 vss.n4023 vss.n4022 0.0661418
R24312 vss.n4022 vss.n4020 0.0661418
R24313 vss.n4025 vss.n4024 0.0661418
R24314 vss.n4025 vss.n3326 0.0661418
R24315 vss.n5531 vss.n4007 0.0661418
R24316 vss.n5504 vss.n5503 0.0661418
R24317 vss.n5503 vss.n5479 0.0661418
R24318 vss.n5480 vss.n5473 0.0661418
R24319 vss.n5480 vss.n5478 0.0661418
R24320 vss.n5488 vss.n5486 0.0661418
R24321 vss.n5486 vss.n5485 0.0661418
R24322 vss.n5506 vss.n5505 0.0661418
R24323 vss.n5506 vss.n4004 0.0661418
R24324 vss.n5491 vss.n5487 0.0661418
R24325 vss.n4068 vss.n4067 0.0661418
R24326 vss.n4067 vss.n4044 0.0661418
R24327 vss.n4045 vss.n4038 0.0661418
R24328 vss.n4045 vss.n4043 0.0661418
R24329 vss.n4053 vss.n4051 0.0661418
R24330 vss.n4051 vss.n4050 0.0661418
R24331 vss.n4056 vss.n4052 0.0661418
R24332 vss.n4052 vss.n3322 0.0661418
R24333 vss.n5078 vss.n5077 0.0661418
R24334 vss.n5077 vss.n5053 0.0661418
R24335 vss.n5054 vss.n5047 0.0661418
R24336 vss.n5054 vss.n5052 0.0661418
R24337 vss.n5062 vss.n5060 0.0661418
R24338 vss.n5060 vss.n5059 0.0661418
R24339 vss.n5080 vss.n5079 0.0661418
R24340 vss.n5080 vss.n4001 0.0661418
R24341 vss.n5065 vss.n5061 0.0661418
R24342 vss.n4209 vss.n4176 0.0661418
R24343 vss.n4210 vss.n4209 0.0661418
R24344 vss.n4198 vss.n4173 0.0661418
R24345 vss.n4199 vss.n4198 0.0661418
R24346 vss.n4187 vss.n4185 0.0661418
R24347 vss.n4185 vss.n4184 0.0661418
R24348 vss.n4190 vss.n4186 0.0661418
R24349 vss.n4186 vss.n3318 0.0661418
R24350 vss.n4213 vss.n4177 0.0661418
R24351 vss.n5030 vss.n5029 0.0661418
R24352 vss.n5029 vss.n5005 0.0661418
R24353 vss.n5006 vss.n4999 0.0661418
R24354 vss.n5006 vss.n5004 0.0661418
R24355 vss.n5014 vss.n5012 0.0661418
R24356 vss.n5012 vss.n5011 0.0661418
R24357 vss.n5032 vss.n5031 0.0661418
R24358 vss.n5032 vss.n3996 0.0661418
R24359 vss.n5017 vss.n5013 0.0661418
R24360 vss.n4249 vss.n4248 0.0661418
R24361 vss.n4248 vss.n4225 0.0661418
R24362 vss.n4226 vss.n4219 0.0661418
R24363 vss.n4226 vss.n4224 0.0661418
R24364 vss.n4234 vss.n4232 0.0661418
R24365 vss.n4232 vss.n4231 0.0661418
R24366 vss.n4237 vss.n4233 0.0661418
R24367 vss.n4233 vss.n3314 0.0661418
R24368 vss.n4525 vss.n4524 0.0661418
R24369 vss.n4524 vss.n4500 0.0661418
R24370 vss.n4501 vss.n4494 0.0661418
R24371 vss.n4501 vss.n4499 0.0661418
R24372 vss.n4509 vss.n4507 0.0661418
R24373 vss.n4507 vss.n4506 0.0661418
R24374 vss.n4527 vss.n4526 0.0661418
R24375 vss.n4527 vss.n3993 0.0661418
R24376 vss.n4512 vss.n4508 0.0661418
R24377 vss.n4477 vss.n4476 0.0661418
R24378 vss.n4476 vss.n4453 0.0661418
R24379 vss.n4454 vss.n4447 0.0661418
R24380 vss.n4454 vss.n4452 0.0661418
R24381 vss.n4462 vss.n4460 0.0661418
R24382 vss.n4460 vss.n4459 0.0661418
R24383 vss.n4465 vss.n4461 0.0661418
R24384 vss.n4461 vss.n3310 0.0661418
R24385 vss.n4482 vss.n4478 0.0661418
R24386 vss.n4408 vss.n4401 0.0661418
R24387 vss.n4408 vss.n4406 0.0661418
R24388 vss.n4416 vss.n4414 0.0661418
R24389 vss.n4414 vss.n4413 0.0661418
R24390 vss.n4431 vss.n4430 0.0661418
R24391 vss.n4430 vss.n4407 0.0661418
R24392 vss.n4433 vss.n4432 0.0661418
R24393 vss.n4433 vss.n3988 0.0661418
R24394 vss.n4419 vss.n4415 0.0661418
R24395 vss.n4415 vss.n3307 0.0661418
R24396 vss.n4768 vss.n4767 0.0661418
R24397 vss.n4767 vss.n4762 0.0661418
R24398 vss.n4763 vss.n4757 0.0661418
R24399 vss.n4763 vss.n4761 0.0661418
R24400 vss.n4774 vss.n4773 0.0661418
R24401 vss.n4773 vss.n4771 0.0661418
R24402 vss.n4776 vss.n4775 0.0661418
R24403 vss.n4776 vss.n3308 0.0661418
R24404 vss.n4798 vss.n4797 0.0661418
R24405 vss.n4799 vss.n4798 0.0661418
R24406 vss.n3304 vss.n3303 0.0661418
R24407 vss.n3303 vss.n3280 0.0661418
R24408 vss.n3281 vss.n3274 0.0661418
R24409 vss.n3281 vss.n3279 0.0661418
R24410 vss.n3289 vss.n3287 0.0661418
R24411 vss.n3287 vss.n3286 0.0661418
R24412 vss.n3306 vss.n3305 0.0661418
R24413 vss.n6726 vss.n3306 0.0661418
R24414 vss.n3292 vss.n3288 0.0661418
R24415 vss.n3288 vss.n436 0.0661418
R24416 vss.n15516 vss.n15515 0.0661418
R24417 vss.n15515 vss.n15513 0.0661418
R24418 vss.n15510 vss.n15509 0.0661418
R24419 vss.n15509 vss.n15504 0.0661418
R24420 vss.n15518 vss.n15517 0.0661418
R24421 vss.n15518 vss.n382 0.0661418
R24422 vss.n1048 vss.n1041 0.0661418
R24423 vss.n1048 vss.n1046 0.0661418
R24424 vss.n1071 vss.n1070 0.0661418
R24425 vss.n1070 vss.n1047 0.0661418
R24426 vss.n1056 vss.n1054 0.0661418
R24427 vss.n1054 vss.n1053 0.0661418
R24428 vss.n1059 vss.n1055 0.0661418
R24429 vss.n1055 vss.n407 0.0661418
R24430 vss.n1073 vss.n1072 0.0661418
R24431 vss.n15036 vss.n1073 0.0661418
R24432 vss.n14903 vss.n14901 0.0661418
R24433 vss.n14901 vss.n14900 0.0661418
R24434 vss.n14895 vss.n14888 0.0661418
R24435 vss.n14895 vss.n14893 0.0661418
R24436 vss.n14920 vss.n14919 0.0661418
R24437 vss.n14919 vss.n14894 0.0661418
R24438 vss.n14922 vss.n14921 0.0661418
R24439 vss.n14922 vss.n409 0.0661418
R24440 vss.n14906 vss.n14902 0.0661418
R24441 vss.n510 vss.n503 0.0661418
R24442 vss.n510 vss.n508 0.0661418
R24443 vss.n533 vss.n532 0.0661418
R24444 vss.n532 vss.n509 0.0661418
R24445 vss.n518 vss.n516 0.0661418
R24446 vss.n516 vss.n515 0.0661418
R24447 vss.n521 vss.n517 0.0661418
R24448 vss.n517 vss.n427 0.0661418
R24449 vss.n535 vss.n534 0.0661418
R24450 vss.n15430 vss.n535 0.0661418
R24451 vss.n7308 vss.n7301 0.0661418
R24452 vss.n7308 vss.n7306 0.0661418
R24453 vss.n7331 vss.n7330 0.0661418
R24454 vss.n7330 vss.n7307 0.0661418
R24455 vss.n7316 vss.n7314 0.0661418
R24456 vss.n7314 vss.n7313 0.0661418
R24457 vss.n7319 vss.n7315 0.0661418
R24458 vss.n7315 vss.n423 0.0661418
R24459 vss.n7333 vss.n7332 0.0661418
R24460 vss.n7333 vss.n642 0.0661418
R24461 vss.n715 vss.n708 0.0661418
R24462 vss.n715 vss.n713 0.0661418
R24463 vss.n738 vss.n737 0.0661418
R24464 vss.n737 vss.n714 0.0661418
R24465 vss.n723 vss.n721 0.0661418
R24466 vss.n721 vss.n720 0.0661418
R24467 vss.n726 vss.n722 0.0661418
R24468 vss.n722 vss.n419 0.0661418
R24469 vss.n740 vss.n739 0.0661418
R24470 vss.n15357 vss.n740 0.0661418
R24471 vss.n768 vss.n761 0.0661418
R24472 vss.n768 vss.n766 0.0661418
R24473 vss.n791 vss.n790 0.0661418
R24474 vss.n790 vss.n767 0.0661418
R24475 vss.n776 vss.n774 0.0661418
R24476 vss.n774 vss.n773 0.0661418
R24477 vss.n779 vss.n775 0.0661418
R24478 vss.n775 vss.n415 0.0661418
R24479 vss.n793 vss.n792 0.0661418
R24480 vss.n15280 vss.n793 0.0661418
R24481 vss.n15182 vss.n15175 0.0661418
R24482 vss.n15182 vss.n15180 0.0661418
R24483 vss.n15205 vss.n15204 0.0661418
R24484 vss.n15204 vss.n15181 0.0661418
R24485 vss.n15190 vss.n15188 0.0661418
R24486 vss.n15188 vss.n15187 0.0661418
R24487 vss.n15193 vss.n15189 0.0661418
R24488 vss.n15189 vss.n411 0.0661418
R24489 vss.n15207 vss.n15206 0.0661418
R24490 vss.n15207 vss.n899 0.0661418
R24491 vss.n925 vss.n918 0.0661418
R24492 vss.n925 vss.n923 0.0661418
R24493 vss.n948 vss.n947 0.0661418
R24494 vss.n947 vss.n924 0.0661418
R24495 vss.n933 vss.n931 0.0661418
R24496 vss.n931 vss.n930 0.0661418
R24497 vss.n936 vss.n932 0.0661418
R24498 vss.n932 vss.n410 0.0661418
R24499 vss.n950 vss.n949 0.0661418
R24500 vss.n951 vss.n950 0.0661418
R24501 vss.n819 vss.n818 0.0661418
R24502 vss.n818 vss.n813 0.0661418
R24503 vss.n816 vss.n809 0.0661418
R24504 vss.n816 vss.n814 0.0661418
R24505 vss.n825 vss.n824 0.0661418
R24506 vss.n824 vss.n822 0.0661418
R24507 vss.n827 vss.n826 0.0661418
R24508 vss.n827 vss.n414 0.0661418
R24509 vss.n849 vss.n848 0.0661418
R24510 vss.n850 vss.n849 0.0661418
R24511 vss.n15104 vss.n15099 0.0661418
R24512 vss.n15104 vss.n15102 0.0661418
R24513 vss.n15112 vss.n15111 0.0661418
R24514 vss.n15111 vss.n15103 0.0661418
R24515 vss.n15118 vss.n15117 0.0661418
R24516 vss.n15117 vss.n15115 0.0661418
R24517 vss.n15120 vss.n15119 0.0661418
R24518 vss.n15120 vss.n417 0.0661418
R24519 vss.n7456 vss.n7455 0.0661418
R24520 vss.n7455 vss.n7449 0.0661418
R24521 vss.n7462 vss.n7461 0.0661418
R24522 vss.n7461 vss.n7459 0.0661418
R24523 vss.n7450 vss.n7445 0.0661418
R24524 vss.n7450 vss.n7441 0.0661418
R24525 vss.n7444 vss.n7440 0.0661418
R24526 vss.n7487 vss.n7440 0.0661418
R24527 vss.n7464 vss.n7463 0.0661418
R24528 vss.n15302 vss.n15295 0.0661418
R24529 vss.n15302 vss.n15300 0.0661418
R24530 vss.n15325 vss.n15324 0.0661418
R24531 vss.n15324 vss.n15301 0.0661418
R24532 vss.n15310 vss.n15308 0.0661418
R24533 vss.n15308 vss.n15307 0.0661418
R24534 vss.n15313 vss.n15309 0.0661418
R24535 vss.n15309 vss.n418 0.0661418
R24536 vss.n15327 vss.n15326 0.0661418
R24537 vss.n15328 vss.n15327 0.0661418
R24538 vss.n668 vss.n661 0.0661418
R24539 vss.n668 vss.n666 0.0661418
R24540 vss.n691 vss.n690 0.0661418
R24541 vss.n690 vss.n667 0.0661418
R24542 vss.n676 vss.n674 0.0661418
R24543 vss.n674 vss.n673 0.0661418
R24544 vss.n679 vss.n675 0.0661418
R24545 vss.n675 vss.n422 0.0661418
R24546 vss.n693 vss.n692 0.0661418
R24547 vss.n694 vss.n693 0.0661418
R24548 vss.n7397 vss.n7394 0.0661418
R24549 vss.n7403 vss.n7398 0.0661418
R24550 vss.n7403 vss.n7401 0.0661418
R24551 vss.n7410 vss.n7409 0.0661418
R24552 vss.n7409 vss.n7402 0.0661418
R24553 vss.n7416 vss.n7415 0.0661418
R24554 vss.n7415 vss.n7413 0.0661418
R24555 vss.n7418 vss.n7417 0.0661418
R24556 vss.n7418 vss.n421 0.0661418
R24557 vss.n7374 vss.n7373 0.0661418
R24558 vss.n7356 vss.n3063 0.0661418
R24559 vss.n7356 vss.n7354 0.0661418
R24560 vss.n7361 vss.n7360 0.0661418
R24561 vss.n7360 vss.n7355 0.0661418
R24562 vss.n7367 vss.n7366 0.0661418
R24563 vss.n7366 vss.n7364 0.0661418
R24564 vss.n7391 vss.n7390 0.0661418
R24565 vss.n7392 vss.n7391 0.0661418
R24566 vss.n3083 vss.n3078 0.0661418
R24567 vss.n3084 vss.n3077 0.0661418
R24568 vss.n3077 vss.n3076 0.0661418
R24569 vss.n3071 vss.n3064 0.0661418
R24570 vss.n3071 vss.n3069 0.0661418
R24571 vss.n3095 vss.n3094 0.0661418
R24572 vss.n3094 vss.n3070 0.0661418
R24573 vss.n3097 vss.n3096 0.0661418
R24574 vss.n3097 vss.n425 0.0661418
R24575 vss.n3117 vss.n3110 0.0661418
R24576 vss.n3117 vss.n3115 0.0661418
R24577 vss.n7284 vss.n7283 0.0661418
R24578 vss.n7283 vss.n3116 0.0661418
R24579 vss.n3125 vss.n3123 0.0661418
R24580 vss.n3123 vss.n3122 0.0661418
R24581 vss.n7272 vss.n3124 0.0661418
R24582 vss.n7271 vss.n3124 0.0661418
R24583 vss.n7289 vss.n7285 0.0661418
R24584 vss.n562 vss.n561 0.0661418
R24585 vss.n561 vss.n556 0.0661418
R24586 vss.n559 vss.n551 0.0661418
R24587 vss.n559 vss.n557 0.0661418
R24588 vss.n568 vss.n567 0.0661418
R24589 vss.n567 vss.n565 0.0661418
R24590 vss.n570 vss.n569 0.0661418
R24591 vss.n570 vss.n426 0.0661418
R24592 vss.n592 vss.n591 0.0661418
R24593 vss.n593 vss.n592 0.0661418
R24594 vss.n460 vss.n453 0.0661418
R24595 vss.n460 vss.n458 0.0661418
R24596 vss.n483 vss.n482 0.0661418
R24597 vss.n482 vss.n459 0.0661418
R24598 vss.n468 vss.n466 0.0661418
R24599 vss.n466 vss.n465 0.0661418
R24600 vss.n471 vss.n467 0.0661418
R24601 vss.n467 vss.n434 0.0661418
R24602 vss.n485 vss.n484 0.0661418
R24603 vss.n486 vss.n485 0.0661418
R24604 vss.n4713 vss.n4712 0.0661418
R24605 vss.n4712 vss.n4707 0.0661418
R24606 vss.n4710 vss.n4558 0.0661418
R24607 vss.n4710 vss.n4708 0.0661418
R24608 vss.n4719 vss.n4718 0.0661418
R24609 vss.n4718 vss.n4716 0.0661418
R24610 vss.n4721 vss.n4720 0.0661418
R24611 vss.n4721 vss.n431 0.0661418
R24612 vss.n4743 vss.n4742 0.0661418
R24613 vss.n4744 vss.n4743 0.0661418
R24614 vss.n4328 vss.n4327 0.0661418
R24615 vss.n4327 vss.n4322 0.0661418
R24616 vss.n4325 vss.n4318 0.0661418
R24617 vss.n4325 vss.n4323 0.0661418
R24618 vss.n4334 vss.n4333 0.0661418
R24619 vss.n4333 vss.n4331 0.0661418
R24620 vss.n4336 vss.n4335 0.0661418
R24621 vss.n4336 vss.n430 0.0661418
R24622 vss.n4358 vss.n4357 0.0661418
R24623 vss.n4359 vss.n4358 0.0661418
R24624 vss.n7227 vss.n3128 0.0661418
R24625 vss.n7233 vss.n7228 0.0661418
R24626 vss.n7233 vss.n7231 0.0661418
R24627 vss.n7240 vss.n7239 0.0661418
R24628 vss.n7239 vss.n7232 0.0661418
R24629 vss.n7246 vss.n7245 0.0661418
R24630 vss.n7245 vss.n7243 0.0661418
R24631 vss.n7248 vss.n7247 0.0661418
R24632 vss.n7248 vss.n429 0.0661418
R24633 vss.n4639 vss.n4638 0.0661418
R24634 vss.n4622 vss.n4620 0.0661418
R24635 vss.n4620 vss.n4619 0.0661418
R24636 vss.n4614 vss.n4607 0.0661418
R24637 vss.n4614 vss.n4612 0.0661418
R24638 vss.n4637 vss.n4636 0.0661418
R24639 vss.n4636 vss.n4613 0.0661418
R24640 vss.n4625 vss.n4621 0.0661418
R24641 vss.n4621 vss.n3133 0.0661418
R24642 vss.n4674 vss.n4669 0.0661418
R24643 vss.n4675 vss.n4668 0.0661418
R24644 vss.n4668 vss.n4667 0.0661418
R24645 vss.n4662 vss.n4655 0.0661418
R24646 vss.n4662 vss.n4660 0.0661418
R24647 vss.n4686 vss.n4685 0.0661418
R24648 vss.n4685 vss.n4661 0.0661418
R24649 vss.n4688 vss.n4687 0.0661418
R24650 vss.n4688 vss.n433 0.0661418
R24651 vss.n4592 vss.n4591 0.0661418
R24652 vss.n4574 vss.n4572 0.0661418
R24653 vss.n4572 vss.n4571 0.0661418
R24654 vss.n4566 vss.n4559 0.0661418
R24655 vss.n4566 vss.n4564 0.0661418
R24656 vss.n4590 vss.n4589 0.0661418
R24657 vss.n4589 vss.n4565 0.0661418
R24658 vss.n4578 vss.n4573 0.0661418
R24659 vss.n4577 vss.n4573 0.0661418
R24660 vss.n6838 vss.n6831 0.0661418
R24661 vss.n6838 vss.n6836 0.0661418
R24662 vss.n6846 vss.n6844 0.0661418
R24663 vss.n6844 vss.n6843 0.0661418
R24664 vss.n6861 vss.n6860 0.0661418
R24665 vss.n6860 vss.n6837 0.0661418
R24666 vss.n6863 vss.n6862 0.0661418
R24667 vss.n6863 vss.n6804 0.0661418
R24668 vss.n6849 vss.n6845 0.0661418
R24669 vss.n6845 vss.n2359 0.0661418
R24670 vss.n2609 vss.n2608 0.0661418
R24671 vss.n2609 vss.n2606 0.0661418
R24672 vss.n2615 vss.n2614 0.0661418
R24673 vss.n2614 vss.n2612 0.0661418
R24674 vss.n2630 vss.n2602 0.0661418
R24675 vss.n2630 vss.n2607 0.0661418
R24676 vss.n2641 vss.n2640 0.0661418
R24677 vss.n2642 vss.n2641 0.0661418
R24678 vss.n2617 vss.n2616 0.0661418
R24679 vss.n2617 vss.n1854 0.0661418
R24680 vss.n1912 vss.n1911 0.0661418
R24681 vss.n1911 vss.n1906 0.0661418
R24682 vss.n1907 vss.n1901 0.0661418
R24683 vss.n1907 vss.n1905 0.0661418
R24684 vss.n1918 vss.n1917 0.0661418
R24685 vss.n1917 vss.n1915 0.0661418
R24686 vss.n1920 vss.n1919 0.0661418
R24687 vss.n1921 vss.n1920 0.0661418
R24688 vss.n1943 vss.n1942 0.0661418
R24689 vss.n1944 vss.n1943 0.0661418
R24690 vss.n2845 vss.n2838 0.0661418
R24691 vss.n2845 vss.n2843 0.0661418
R24692 vss.n2853 vss.n2851 0.0661418
R24693 vss.n2851 vss.n2850 0.0661418
R24694 vss.n2868 vss.n2867 0.0661418
R24695 vss.n2867 vss.n2844 0.0661418
R24696 vss.n2870 vss.n2869 0.0661418
R24697 vss.n2870 vss.n2476 0.0661418
R24698 vss.n2856 vss.n2852 0.0661418
R24699 vss.n2852 vss.n1574 0.0661418
R24700 vss.n3057 vss.n3056 0.0661418
R24701 vss.n7629 vss.n7622 0.0661418
R24702 vss.n7629 vss.n7627 0.0661418
R24703 vss.n7637 vss.n7635 0.0661418
R24704 vss.n7635 vss.n7634 0.0661418
R24705 vss.n7652 vss.n7651 0.0661418
R24706 vss.n7651 vss.n7628 0.0661418
R24707 vss.n7654 vss.n7653 0.0661418
R24708 vss.n7654 vss.n2472 0.0661418
R24709 vss.n7640 vss.n7636 0.0661418
R24710 vss.n7636 vss.n1521 0.0661418
R24711 vss.n2731 vss.n2724 0.0661418
R24712 vss.n2731 vss.n2729 0.0661418
R24713 vss.n2739 vss.n2737 0.0661418
R24714 vss.n2737 vss.n2736 0.0661418
R24715 vss.n2822 vss.n2821 0.0661418
R24716 vss.n2821 vss.n2730 0.0661418
R24717 vss.n2824 vss.n2823 0.0661418
R24718 vss.n2824 vss.n2475 0.0661418
R24719 vss.n2810 vss.n2738 0.0661418
R24720 vss.n2809 vss.n2738 0.0661418
R24721 vss.n2937 vss.n2930 0.0661418
R24722 vss.n2937 vss.n2935 0.0661418
R24723 vss.n2945 vss.n2943 0.0661418
R24724 vss.n2943 vss.n2942 0.0661418
R24725 vss.n2960 vss.n2959 0.0661418
R24726 vss.n2959 vss.n2936 0.0661418
R24727 vss.n2962 vss.n2961 0.0661418
R24728 vss.n2963 vss.n2962 0.0661418
R24729 vss.n2948 vss.n2944 0.0661418
R24730 vss.n2944 vss.n1422 0.0661418
R24731 vss.n7056 vss.n3131 0.0661418
R24732 vss.n6998 vss.n6997 0.0661418
R24733 vss.n6998 vss.n6995 0.0661418
R24734 vss.n7004 vss.n7003 0.0661418
R24735 vss.n7003 vss.n7001 0.0661418
R24736 vss.n7019 vss.n6991 0.0661418
R24737 vss.n7019 vss.n6996 0.0661418
R24738 vss.n7030 vss.n7029 0.0661418
R24739 vss.n7031 vss.n7030 0.0661418
R24740 vss.n7006 vss.n7005 0.0661418
R24741 vss.n7006 vss.n1316 0.0661418
R24742 vss.n7138 vss.n7137 0.0661418
R24743 vss.n7137 vss.n7132 0.0661418
R24744 vss.n7144 vss.n7143 0.0661418
R24745 vss.n7143 vss.n7141 0.0661418
R24746 vss.n7135 vss.n7128 0.0661418
R24747 vss.n7135 vss.n7133 0.0661418
R24748 vss.n7168 vss.n7167 0.0661418
R24749 vss.n7169 vss.n7168 0.0661418
R24750 vss.n7146 vss.n7145 0.0661418
R24751 vss.n7146 vss.n1407 0.0661418
R24752 vss.n6934 vss.n6933 0.0661418
R24753 vss.n6933 vss.n6928 0.0661418
R24754 vss.n6940 vss.n6939 0.0661418
R24755 vss.n6939 vss.n6937 0.0661418
R24756 vss.n6931 vss.n6924 0.0661418
R24757 vss.n6931 vss.n6929 0.0661418
R24758 vss.n6985 vss.n6984 0.0661418
R24759 vss.n6986 vss.n6985 0.0661418
R24760 vss.n6942 vss.n6941 0.0661418
R24761 vss.n6962 vss.n6942 0.0661418
R24762 vss.n7513 vss.n7506 0.0661418
R24763 vss.n7513 vss.n7511 0.0661418
R24764 vss.n7521 vss.n7519 0.0661418
R24765 vss.n7519 vss.n7518 0.0661418
R24766 vss.n7604 vss.n7603 0.0661418
R24767 vss.n7603 vss.n7512 0.0661418
R24768 vss.n7606 vss.n7605 0.0661418
R24769 vss.n7606 vss.n2471 0.0661418
R24770 vss.n7592 vss.n7520 0.0661418
R24771 vss.n7591 vss.n7520 0.0661418
R24772 vss.n7776 vss.n7769 0.0661418
R24773 vss.n7776 vss.n7774 0.0661418
R24774 vss.n7784 vss.n7782 0.0661418
R24775 vss.n7782 vss.n7781 0.0661418
R24776 vss.n7799 vss.n7798 0.0661418
R24777 vss.n7798 vss.n7775 0.0661418
R24778 vss.n7801 vss.n7800 0.0661418
R24779 vss.n7801 vss.n2479 0.0661418
R24780 vss.n7787 vss.n7783 0.0661418
R24781 vss.n7783 vss.n1664 0.0661418
R24782 vss.n7824 vss.n7817 0.0661418
R24783 vss.n7824 vss.n7822 0.0661418
R24784 vss.n7832 vss.n7830 0.0661418
R24785 vss.n7830 vss.n7829 0.0661418
R24786 vss.n7847 vss.n7846 0.0661418
R24787 vss.n7846 vss.n7823 0.0661418
R24788 vss.n7849 vss.n7848 0.0661418
R24789 vss.n7849 vss.n2480 0.0661418
R24790 vss.n7835 vss.n7831 0.0661418
R24791 vss.n7831 vss.n1679 0.0661418
R24792 vss.n2712 vss.n987 0.0661418
R24793 vss.n2497 vss.n2496 0.0661418
R24794 vss.n2496 vss.n2491 0.0661418
R24795 vss.n2503 vss.n2502 0.0661418
R24796 vss.n2502 vss.n2500 0.0661418
R24797 vss.n2494 vss.n2487 0.0661418
R24798 vss.n2494 vss.n2492 0.0661418
R24799 vss.n2596 vss.n2595 0.0661418
R24800 vss.n2597 vss.n2596 0.0661418
R24801 vss.n2505 vss.n2504 0.0661418
R24802 vss.n2574 vss.n2505 0.0661418
R24803 vss.n1153 vss.n1152 0.0661418
R24804 vss.n1152 vss.n1147 0.0661418
R24805 vss.n1148 vss.n1141 0.0661418
R24806 vss.n1148 vss.n1146 0.0661418
R24807 vss.n7940 vss.n7939 0.0661418
R24808 vss.n7939 vss.n7926 0.0661418
R24809 vss.n1155 vss.n1154 0.0661418
R24810 vss.n14871 vss.n1155 0.0661418
R24811 vss.n7930 vss.n7928 0.0661418
R24812 vss.n2665 vss.n2660 0.0661418
R24813 vss.n2665 vss.n2664 0.0661418
R24814 vss.n7916 vss.n7915 0.0661418
R24815 vss.n7917 vss.n7916 0.0661418
R24816 vss.n2652 vss.n2647 0.0661418
R24817 vss.n2652 vss.n2651 0.0661418
R24818 vss.n7924 vss.n7923 0.0661418
R24819 vss.n7925 vss.n7924 0.0661418
R24820 vss.n2663 vss.n2661 0.0661418
R24821 vss.n7896 vss.n7895 0.0661418
R24822 vss.n7895 vss.n7871 0.0661418
R24823 vss.n7872 vss.n7865 0.0661418
R24824 vss.n7872 vss.n7870 0.0661418
R24825 vss.n7880 vss.n7878 0.0661418
R24826 vss.n7878 vss.n7877 0.0661418
R24827 vss.n7898 vss.n7897 0.0661418
R24828 vss.n7901 vss.n7898 0.0661418
R24829 vss.n7883 vss.n7879 0.0661418
R24830 vss.n2709 vss.n2708 0.0661418
R24831 vss.n2708 vss.n2685 0.0661418
R24832 vss.n2686 vss.n2679 0.0661418
R24833 vss.n2686 vss.n2684 0.0661418
R24834 vss.n2694 vss.n2692 0.0661418
R24835 vss.n2692 vss.n2691 0.0661418
R24836 vss.n2697 vss.n2693 0.0661418
R24837 vss.n2693 vss.n2481 0.0661418
R24838 vss.n7750 vss.n7749 0.0661418
R24839 vss.n7749 vss.n7725 0.0661418
R24840 vss.n7726 vss.n7719 0.0661418
R24841 vss.n7726 vss.n7724 0.0661418
R24842 vss.n7734 vss.n7732 0.0661418
R24843 vss.n7732 vss.n7731 0.0661418
R24844 vss.n7752 vss.n7751 0.0661418
R24845 vss.n7752 vss.n986 0.0661418
R24846 vss.n7737 vss.n7733 0.0661418
R24847 vss.n2891 vss.n2886 0.0661418
R24848 vss.n2891 vss.n2890 0.0661418
R24849 vss.n2914 vss.n2883 0.0661418
R24850 vss.n2915 vss.n2914 0.0661418
R24851 vss.n2903 vss.n2896 0.0661418
R24852 vss.n2899 vss.n2896 0.0661418
R24853 vss.n2901 vss.n2897 0.0661418
R24854 vss.n2897 vss.n2477 0.0661418
R24855 vss.n2889 vss.n2887 0.0661418
R24856 vss.n7701 vss.n7700 0.0661418
R24857 vss.n7700 vss.n7676 0.0661418
R24858 vss.n7677 vss.n7670 0.0661418
R24859 vss.n7677 vss.n7675 0.0661418
R24860 vss.n7685 vss.n7683 0.0661418
R24861 vss.n7683 vss.n7682 0.0661418
R24862 vss.n7703 vss.n7702 0.0661418
R24863 vss.n7706 vss.n7703 0.0661418
R24864 vss.n7688 vss.n7684 0.0661418
R24865 vss.n3049 vss.n3016 0.0661418
R24866 vss.n3050 vss.n3049 0.0661418
R24867 vss.n3023 vss.n3022 0.0661418
R24868 vss.n3022 vss.n3020 0.0661418
R24869 vss.n3029 vss.n3028 0.0661418
R24870 vss.n3028 vss.n3026 0.0661418
R24871 vss.n3031 vss.n3030 0.0661418
R24872 vss.n3031 vss.n2473 0.0661418
R24873 vss.n3007 vss.n3006 0.0661418
R24874 vss.n3006 vss.n2982 0.0661418
R24875 vss.n2983 vss.n2976 0.0661418
R24876 vss.n2983 vss.n2981 0.0661418
R24877 vss.n2991 vss.n2989 0.0661418
R24878 vss.n2989 vss.n2988 0.0661418
R24879 vss.n3009 vss.n3008 0.0661418
R24880 vss.n7490 vss.n3009 0.0661418
R24881 vss.n2994 vss.n2990 0.0661418
R24882 vss.n2461 vss.n2455 0.0661418
R24883 vss.n2461 vss.n2460 0.0661418
R24884 vss.n7975 vss.n2452 0.0661418
R24885 vss.n7976 vss.n7975 0.0661418
R24886 vss.n7964 vss.n2466 0.0661418
R24887 vss.n7960 vss.n2466 0.0661418
R24888 vss.n7962 vss.n2467 0.0661418
R24889 vss.n7959 vss.n2467 0.0661418
R24890 vss.n2458 vss.n2456 0.0661418
R24891 vss.n7108 vss.n7107 0.0661418
R24892 vss.n7109 vss.n7108 0.0661418
R24893 vss.n7092 vss.n7091 0.0661418
R24894 vss.n7091 vss.n7084 0.0661418
R24895 vss.n7085 vss.n7082 0.0661418
R24896 vss.n7085 vss.n7077 0.0661418
R24897 vss.n7104 vss.n7103 0.0661418
R24898 vss.n7103 vss.n7102 0.0661418
R24899 vss.n7081 vss.n7079 0.0661418
R24900 vss.n7061 vss.n7051 0.0661418
R24901 vss.n7061 vss.n7060 0.0661418
R24902 vss.n7067 vss.n7066 0.0661418
R24903 vss.n7068 vss.n7067 0.0661418
R24904 vss.n7041 vss.n7036 0.0661418
R24905 vss.n7041 vss.n7040 0.0661418
R24906 vss.n7075 vss.n7074 0.0661418
R24907 vss.n7076 vss.n7075 0.0661418
R24908 vss.n6904 vss.n6903 0.0661418
R24909 vss.n6905 vss.n6904 0.0661418
R24910 vss.n6889 vss.n6888 0.0661418
R24911 vss.n6888 vss.n6881 0.0661418
R24912 vss.n6882 vss.n6830 0.0661418
R24913 vss.n6882 vss.n6825 0.0661418
R24914 vss.n6899 vss.n6896 0.0661418
R24915 vss.n6899 vss.n3130 0.0661418
R24916 vss.n6829 vss.n6827 0.0661418
R24917 vss.n3141 vss.n3140 0.0661418
R24918 vss.n7211 vss.n3141 0.0661418
R24919 vss.n3147 vss.n3146 0.0661418
R24920 vss.n3146 vss.n3144 0.0661418
R24921 vss.n6814 vss.n6810 0.0661418
R24922 vss.n6814 vss.n6813 0.0661418
R24923 vss.n6823 vss.n6822 0.0661418
R24924 vss.n6824 vss.n6823 0.0661418
R24925 vss.n7218 vss.n3137 0.0661418
R24926 vss.n3157 vss.n3150 0.0661418
R24927 vss.n3157 vss.n3155 0.0661418
R24928 vss.n3165 vss.n3163 0.0661418
R24929 vss.n3163 vss.n3162 0.0661418
R24930 vss.n7191 vss.n7190 0.0661418
R24931 vss.n7190 vss.n3156 0.0661418
R24932 vss.n7193 vss.n7192 0.0661418
R24933 vss.n7193 vss.n3134 0.0661418
R24934 vss.n7179 vss.n3164 0.0661418
R24935 vss.n7178 vss.n3164 0.0661418
R24936 vss.n3183 vss.n3182 0.0661418
R24937 vss.n3182 vss.n3177 0.0661418
R24938 vss.n3199 vss.n3196 0.0661418
R24939 vss.n3199 vss.n3198 0.0661418
R24940 vss.n3180 vss.n3173 0.0661418
R24941 vss.n3180 vss.n3178 0.0661418
R24942 vss.n6802 vss.n6801 0.0661418
R24943 vss.n6803 vss.n6802 0.0661418
R24944 vss.n3208 vss.n3207 0.0661418
R24945 vss.n3209 vss.n3208 0.0661418
R24946 vss.n6775 vss.n6774 0.0661418
R24947 vss.n6774 vss.n6751 0.0661418
R24948 vss.n6752 vss.n6745 0.0661418
R24949 vss.n6752 vss.n6750 0.0661418
R24950 vss.n6760 vss.n6758 0.0661418
R24951 vss.n6758 vss.n6757 0.0661418
R24952 vss.n6763 vss.n6759 0.0661418
R24953 vss.n6759 vss.n1215 0.0661418
R24954 vss.n6777 vss.n6776 0.0661418
R24955 vss.n6777 vss.n3168 0.0661418
R24956 vss.n14821 vss.n14820 0.0661418
R24957 vss.n14820 vss.n14818 0.0661418
R24958 vss.n14823 vss.n14822 0.0661418
R24959 vss.n14823 vss.n1161 0.0661418
R24960 vss.n1827 vss.n1820 0.0661418
R24961 vss.n1827 vss.n1825 0.0661418
R24962 vss.n1850 vss.n1849 0.0661418
R24963 vss.n1849 vss.n1826 0.0661418
R24964 vss.n1835 vss.n1833 0.0661418
R24965 vss.n1833 vss.n1832 0.0661418
R24966 vss.n1838 vss.n1834 0.0661418
R24967 vss.n1834 vss.n1186 0.0661418
R24968 vss.n1852 vss.n1851 0.0661418
R24969 vss.n14341 vss.n1852 0.0661418
R24970 vss.n14208 vss.n14206 0.0661418
R24971 vss.n14206 vss.n14205 0.0661418
R24972 vss.n14200 vss.n14193 0.0661418
R24973 vss.n14200 vss.n14198 0.0661418
R24974 vss.n14225 vss.n14224 0.0661418
R24975 vss.n14224 vss.n14199 0.0661418
R24976 vss.n14227 vss.n14226 0.0661418
R24977 vss.n14227 vss.n1188 0.0661418
R24978 vss.n14211 vss.n14207 0.0661418
R24979 vss.n1289 vss.n1282 0.0661418
R24980 vss.n1289 vss.n1287 0.0661418
R24981 vss.n1312 vss.n1311 0.0661418
R24982 vss.n1311 vss.n1288 0.0661418
R24983 vss.n1297 vss.n1295 0.0661418
R24984 vss.n1295 vss.n1294 0.0661418
R24985 vss.n1300 vss.n1296 0.0661418
R24986 vss.n1296 vss.n1206 0.0661418
R24987 vss.n1314 vss.n1313 0.0661418
R24988 vss.n14735 vss.n1314 0.0661418
R24989 vss.n13988 vss.n13981 0.0661418
R24990 vss.n13988 vss.n13986 0.0661418
R24991 vss.n14011 vss.n14010 0.0661418
R24992 vss.n14010 vss.n13987 0.0661418
R24993 vss.n13996 vss.n13994 0.0661418
R24994 vss.n13994 vss.n13993 0.0661418
R24995 vss.n13999 vss.n13995 0.0661418
R24996 vss.n13995 vss.n1202 0.0661418
R24997 vss.n14013 vss.n14012 0.0661418
R24998 vss.n14013 vss.n1421 0.0661418
R24999 vss.n1494 vss.n1487 0.0661418
R25000 vss.n1494 vss.n1492 0.0661418
R25001 vss.n1517 vss.n1516 0.0661418
R25002 vss.n1516 vss.n1493 0.0661418
R25003 vss.n1502 vss.n1500 0.0661418
R25004 vss.n1500 vss.n1499 0.0661418
R25005 vss.n1505 vss.n1501 0.0661418
R25006 vss.n1501 vss.n1198 0.0661418
R25007 vss.n1519 vss.n1518 0.0661418
R25008 vss.n14662 vss.n1519 0.0661418
R25009 vss.n1547 vss.n1540 0.0661418
R25010 vss.n1547 vss.n1545 0.0661418
R25011 vss.n1570 vss.n1569 0.0661418
R25012 vss.n1569 vss.n1546 0.0661418
R25013 vss.n1555 vss.n1553 0.0661418
R25014 vss.n1553 vss.n1552 0.0661418
R25015 vss.n1558 vss.n1554 0.0661418
R25016 vss.n1554 vss.n1194 0.0661418
R25017 vss.n1572 vss.n1571 0.0661418
R25018 vss.n14585 vss.n1572 0.0661418
R25019 vss.n14487 vss.n14480 0.0661418
R25020 vss.n14487 vss.n14485 0.0661418
R25021 vss.n14510 vss.n14509 0.0661418
R25022 vss.n14509 vss.n14486 0.0661418
R25023 vss.n14495 vss.n14493 0.0661418
R25024 vss.n14493 vss.n14492 0.0661418
R25025 vss.n14498 vss.n14494 0.0661418
R25026 vss.n14494 vss.n1190 0.0661418
R25027 vss.n14512 vss.n14511 0.0661418
R25028 vss.n14512 vss.n1678 0.0661418
R25029 vss.n1704 vss.n1697 0.0661418
R25030 vss.n1704 vss.n1702 0.0661418
R25031 vss.n1727 vss.n1726 0.0661418
R25032 vss.n1726 vss.n1703 0.0661418
R25033 vss.n1712 vss.n1710 0.0661418
R25034 vss.n1710 vss.n1709 0.0661418
R25035 vss.n1715 vss.n1711 0.0661418
R25036 vss.n1711 vss.n1189 0.0661418
R25037 vss.n1729 vss.n1728 0.0661418
R25038 vss.n1730 vss.n1729 0.0661418
R25039 vss.n1598 vss.n1597 0.0661418
R25040 vss.n1597 vss.n1592 0.0661418
R25041 vss.n1595 vss.n1588 0.0661418
R25042 vss.n1595 vss.n1593 0.0661418
R25043 vss.n1604 vss.n1603 0.0661418
R25044 vss.n1603 vss.n1601 0.0661418
R25045 vss.n1606 vss.n1605 0.0661418
R25046 vss.n1606 vss.n1193 0.0661418
R25047 vss.n1628 vss.n1627 0.0661418
R25048 vss.n1629 vss.n1628 0.0661418
R25049 vss.n14409 vss.n14404 0.0661418
R25050 vss.n14409 vss.n14407 0.0661418
R25051 vss.n14417 vss.n14416 0.0661418
R25052 vss.n14416 vss.n14408 0.0661418
R25053 vss.n14423 vss.n14422 0.0661418
R25054 vss.n14422 vss.n14420 0.0661418
R25055 vss.n14425 vss.n14424 0.0661418
R25056 vss.n14425 vss.n1196 0.0661418
R25057 vss.n13921 vss.n13920 0.0661418
R25058 vss.n13920 vss.n13914 0.0661418
R25059 vss.n13927 vss.n13926 0.0661418
R25060 vss.n13926 vss.n13924 0.0661418
R25061 vss.n13915 vss.n13910 0.0661418
R25062 vss.n13915 vss.n13906 0.0661418
R25063 vss.n13909 vss.n13905 0.0661418
R25064 vss.n13952 vss.n13905 0.0661418
R25065 vss.n13929 vss.n13928 0.0661418
R25066 vss.n14607 vss.n14600 0.0661418
R25067 vss.n14607 vss.n14605 0.0661418
R25068 vss.n14630 vss.n14629 0.0661418
R25069 vss.n14629 vss.n14606 0.0661418
R25070 vss.n14615 vss.n14613 0.0661418
R25071 vss.n14613 vss.n14612 0.0661418
R25072 vss.n14618 vss.n14614 0.0661418
R25073 vss.n14614 vss.n1197 0.0661418
R25074 vss.n14632 vss.n14631 0.0661418
R25075 vss.n14633 vss.n14632 0.0661418
R25076 vss.n1447 vss.n1440 0.0661418
R25077 vss.n1447 vss.n1445 0.0661418
R25078 vss.n1470 vss.n1469 0.0661418
R25079 vss.n1469 vss.n1446 0.0661418
R25080 vss.n1455 vss.n1453 0.0661418
R25081 vss.n1453 vss.n1452 0.0661418
R25082 vss.n1458 vss.n1454 0.0661418
R25083 vss.n1454 vss.n1201 0.0661418
R25084 vss.n1472 vss.n1471 0.0661418
R25085 vss.n1473 vss.n1472 0.0661418
R25086 vss.n13862 vss.n13859 0.0661418
R25087 vss.n13868 vss.n13863 0.0661418
R25088 vss.n13868 vss.n13866 0.0661418
R25089 vss.n13875 vss.n13874 0.0661418
R25090 vss.n13874 vss.n13867 0.0661418
R25091 vss.n13881 vss.n13880 0.0661418
R25092 vss.n13880 vss.n13878 0.0661418
R25093 vss.n13883 vss.n13882 0.0661418
R25094 vss.n13883 vss.n1200 0.0661418
R25095 vss.n8203 vss.n8202 0.0661418
R25096 vss.n8185 vss.n8179 0.0661418
R25097 vss.n8185 vss.n8183 0.0661418
R25098 vss.n8190 vss.n8189 0.0661418
R25099 vss.n8189 vss.n8184 0.0661418
R25100 vss.n8196 vss.n8195 0.0661418
R25101 vss.n8195 vss.n8193 0.0661418
R25102 vss.n8220 vss.n8219 0.0661418
R25103 vss.n8221 vss.n8220 0.0661418
R25104 vss.n8170 vss.n8166 0.0661418
R25105 vss.n8167 vss.n8165 0.0661418
R25106 vss.n8165 vss.n8164 0.0661418
R25107 vss.n8159 vss.n8152 0.0661418
R25108 vss.n8159 vss.n8157 0.0661418
R25109 vss.n13965 vss.n13964 0.0661418
R25110 vss.n13964 vss.n8158 0.0661418
R25111 vss.n13967 vss.n13966 0.0661418
R25112 vss.n13967 vss.n1204 0.0661418
R25113 vss.n14038 vss.n14037 0.0661418
R25114 vss.n14037 vss.n14031 0.0661418
R25115 vss.n14044 vss.n14043 0.0661418
R25116 vss.n14043 vss.n14041 0.0661418
R25117 vss.n14032 vss.n8149 0.0661418
R25118 vss.n14032 vss.n8145 0.0661418
R25119 vss.n8148 vss.n8144 0.0661418
R25120 vss.n14069 vss.n8144 0.0661418
R25121 vss.n14046 vss.n14045 0.0661418
R25122 vss.n1341 vss.n1340 0.0661418
R25123 vss.n1340 vss.n1335 0.0661418
R25124 vss.n1338 vss.n1330 0.0661418
R25125 vss.n1338 vss.n1336 0.0661418
R25126 vss.n1347 vss.n1346 0.0661418
R25127 vss.n1346 vss.n1344 0.0661418
R25128 vss.n1349 vss.n1348 0.0661418
R25129 vss.n1349 vss.n1205 0.0661418
R25130 vss.n1371 vss.n1370 0.0661418
R25131 vss.n1372 vss.n1371 0.0661418
R25132 vss.n1239 vss.n1232 0.0661418
R25133 vss.n1239 vss.n1237 0.0661418
R25134 vss.n1262 vss.n1261 0.0661418
R25135 vss.n1261 vss.n1238 0.0661418
R25136 vss.n1247 vss.n1245 0.0661418
R25137 vss.n1245 vss.n1244 0.0661418
R25138 vss.n1250 vss.n1246 0.0661418
R25139 vss.n1246 vss.n1213 0.0661418
R25140 vss.n1264 vss.n1263 0.0661418
R25141 vss.n1265 vss.n1264 0.0661418
R25142 vss.n2332 vss.n2325 0.0661418
R25143 vss.n2332 vss.n2330 0.0661418
R25144 vss.n2355 vss.n2354 0.0661418
R25145 vss.n2354 vss.n2331 0.0661418
R25146 vss.n2340 vss.n2338 0.0661418
R25147 vss.n2338 vss.n2337 0.0661418
R25148 vss.n2343 vss.n2339 0.0661418
R25149 vss.n2339 vss.n1210 0.0661418
R25150 vss.n2357 vss.n2356 0.0661418
R25151 vss.n8034 vss.n2357 0.0661418
R25152 vss.n2383 vss.n2382 0.0661418
R25153 vss.n2382 vss.n2377 0.0661418
R25154 vss.n2380 vss.n2373 0.0661418
R25155 vss.n2380 vss.n2378 0.0661418
R25156 vss.n2389 vss.n2388 0.0661418
R25157 vss.n2388 vss.n2386 0.0661418
R25158 vss.n2391 vss.n2390 0.0661418
R25159 vss.n2391 vss.n1209 0.0661418
R25160 vss.n2413 vss.n2412 0.0661418
R25161 vss.n2414 vss.n2413 0.0661418
R25162 vss.n8101 vss.n8097 0.0661418
R25163 vss.n8107 vss.n8102 0.0661418
R25164 vss.n8107 vss.n8105 0.0661418
R25165 vss.n8114 vss.n8113 0.0661418
R25166 vss.n8113 vss.n8106 0.0661418
R25167 vss.n8120 vss.n8119 0.0661418
R25168 vss.n8119 vss.n8117 0.0661418
R25169 vss.n8122 vss.n8121 0.0661418
R25170 vss.n8122 vss.n1208 0.0661418
R25171 vss.n8075 vss.n8074 0.0661418
R25172 vss.n8057 vss.n2230 0.0661418
R25173 vss.n8057 vss.n8055 0.0661418
R25174 vss.n8062 vss.n8061 0.0661418
R25175 vss.n8061 vss.n8056 0.0661418
R25176 vss.n8068 vss.n8067 0.0661418
R25177 vss.n8067 vss.n8065 0.0661418
R25178 vss.n8092 vss.n8091 0.0661418
R25179 vss.n8093 vss.n8092 0.0661418
R25180 vss.n2250 vss.n2245 0.0661418
R25181 vss.n2251 vss.n2244 0.0661418
R25182 vss.n2244 vss.n2243 0.0661418
R25183 vss.n2238 vss.n2231 0.0661418
R25184 vss.n2238 vss.n2236 0.0661418
R25185 vss.n2262 vss.n2261 0.0661418
R25186 vss.n2261 vss.n2237 0.0661418
R25187 vss.n2264 vss.n2263 0.0661418
R25188 vss.n2264 vss.n1212 0.0661418
R25189 vss.n2310 vss.n2309 0.0661418
R25190 vss.n2292 vss.n2290 0.0661418
R25191 vss.n2290 vss.n2289 0.0661418
R25192 vss.n2284 vss.n2277 0.0661418
R25193 vss.n2284 vss.n2282 0.0661418
R25194 vss.n2308 vss.n2307 0.0661418
R25195 vss.n2307 vss.n2283 0.0661418
R25196 vss.n2296 vss.n2291 0.0661418
R25197 vss.n2295 vss.n2291 0.0661418
R25198 vss.n2094 vss.n2087 0.0661418
R25199 vss.n2094 vss.n2092 0.0661418
R25200 vss.n11952 vss.n11949 0.0661418
R25201 vss.n11952 vss.n11951 0.0661418
R25202 vss.n2099 vss.n2098 0.0661418
R25203 vss.n2098 vss.n2093 0.0661418
R25204 vss.n2101 vss.n2100 0.0661418
R25205 vss.n14125 vss.n2101 0.0661418
R25206 vss.n11961 vss.n11960 0.0661418
R25207 vss.n11962 vss.n11961 0.0661418
R25208 vss.n13474 vss.n13467 0.0661418
R25209 vss.n13474 vss.n13472 0.0661418
R25210 vss.n13482 vss.n13480 0.0661418
R25211 vss.n13480 vss.n13479 0.0661418
R25212 vss.n13497 vss.n13496 0.0661418
R25213 vss.n13496 vss.n13473 0.0661418
R25214 vss.n13499 vss.n13498 0.0661418
R25215 vss.n13499 vss.n2105 0.0661418
R25216 vss.n13485 vss.n13481 0.0661418
R25217 vss.n13481 vss.n8356 0.0661418
R25218 vss.n12030 vss.n12029 0.0661418
R25219 vss.n12029 vss.n12024 0.0661418
R25220 vss.n12025 vss.n12019 0.0661418
R25221 vss.n12025 vss.n12023 0.0661418
R25222 vss.n12036 vss.n12035 0.0661418
R25223 vss.n12035 vss.n12033 0.0661418
R25224 vss.n12038 vss.n12037 0.0661418
R25225 vss.n12038 vss.n2102 0.0661418
R25226 vss.n12059 vss.n12058 0.0661418
R25227 vss.n12060 vss.n12059 0.0661418
R25228 vss.n8309 vss.n8302 0.0661418
R25229 vss.n8309 vss.n8307 0.0661418
R25230 vss.n8317 vss.n8315 0.0661418
R25231 vss.n8315 vss.n8314 0.0661418
R25232 vss.n13729 vss.n13728 0.0661418
R25233 vss.n13728 vss.n8308 0.0661418
R25234 vss.n13731 vss.n13730 0.0661418
R25235 vss.n13731 vss.n2109 0.0661418
R25236 vss.n13717 vss.n8316 0.0661418
R25237 vss.n13716 vss.n8316 0.0661418
R25238 vss.n8456 vss.n8455 0.0661418
R25239 vss.n8455 vss.n8450 0.0661418
R25240 vss.n8451 vss.n8445 0.0661418
R25241 vss.n8451 vss.n8449 0.0661418
R25242 vss.n8462 vss.n8461 0.0661418
R25243 vss.n8461 vss.n8459 0.0661418
R25244 vss.n8464 vss.n8463 0.0661418
R25245 vss.n8464 vss.n2113 0.0661418
R25246 vss.n8485 vss.n8484 0.0661418
R25247 vss.n8486 vss.n8485 0.0661418
R25248 vss.n8533 vss.n8532 0.0661418
R25249 vss.n8532 vss.n8527 0.0661418
R25250 vss.n8528 vss.n8522 0.0661418
R25251 vss.n8528 vss.n8526 0.0661418
R25252 vss.n8539 vss.n8538 0.0661418
R25253 vss.n8538 vss.n8536 0.0661418
R25254 vss.n8541 vss.n8540 0.0661418
R25255 vss.n8541 vss.n2110 0.0661418
R25256 vss.n8562 vss.n8561 0.0661418
R25257 vss.n8563 vss.n8562 0.0661418
R25258 vss.n9095 vss.n9088 0.0661418
R25259 vss.n9095 vss.n9093 0.0661418
R25260 vss.n9103 vss.n9101 0.0661418
R25261 vss.n9101 vss.n9100 0.0661418
R25262 vss.n13017 vss.n13016 0.0661418
R25263 vss.n13016 vss.n9094 0.0661418
R25264 vss.n13019 vss.n13018 0.0661418
R25265 vss.n13019 vss.n2117 0.0661418
R25266 vss.n13005 vss.n9102 0.0661418
R25267 vss.n13004 vss.n9102 0.0661418
R25268 vss.n8959 vss.n8952 0.0661418
R25269 vss.n8959 vss.n8957 0.0661418
R25270 vss.n8967 vss.n8965 0.0661418
R25271 vss.n8965 vss.n8964 0.0661418
R25272 vss.n8982 vss.n8981 0.0661418
R25273 vss.n8981 vss.n8958 0.0661418
R25274 vss.n8984 vss.n8983 0.0661418
R25275 vss.n8984 vss.n2121 0.0661418
R25276 vss.n8970 vss.n8966 0.0661418
R25277 vss.n8966 vss.n8900 0.0661418
R25278 vss.n9128 vss.n9127 0.0661418
R25279 vss.n9127 vss.n9122 0.0661418
R25280 vss.n9123 vss.n9117 0.0661418
R25281 vss.n9123 vss.n9121 0.0661418
R25282 vss.n9134 vss.n9133 0.0661418
R25283 vss.n9133 vss.n9131 0.0661418
R25284 vss.n9136 vss.n9135 0.0661418
R25285 vss.n9136 vss.n2118 0.0661418
R25286 vss.n9157 vss.n9156 0.0661418
R25287 vss.n9158 vss.n9157 0.0661418
R25288 vss.n12559 vss.n12558 0.0661418
R25289 vss.n12558 vss.n12553 0.0661418
R25290 vss.n12554 vss.n12548 0.0661418
R25291 vss.n12554 vss.n12552 0.0661418
R25292 vss.n12565 vss.n12564 0.0661418
R25293 vss.n12564 vss.n12562 0.0661418
R25294 vss.n12567 vss.n12566 0.0661418
R25295 vss.n12567 vss.n2125 0.0661418
R25296 vss.n12637 vss.n12636 0.0661418
R25297 vss.n12638 vss.n12637 0.0661418
R25298 vss.n9030 vss.n8096 0.0661418
R25299 vss.n13858 vss.n13857 0.0661418
R25300 vss.n13545 vss.n1766 0.0661418
R25301 vss.n14146 vss.n2058 0.0661418
R25302 vss.n14147 vss.n14146 0.0661418
R25303 vss.n2065 vss.n2064 0.0661418
R25304 vss.n2064 vss.n2062 0.0661418
R25305 vss.n2071 vss.n2070 0.0661418
R25306 vss.n2070 vss.n2068 0.0661418
R25307 vss.n14154 vss.n14153 0.0661418
R25308 vss.n14155 vss.n14154 0.0661418
R25309 vss.n2073 vss.n2072 0.0661418
R25310 vss.n13587 vss.n13586 0.0661418
R25311 vss.n13586 vss.n13562 0.0661418
R25312 vss.n13563 vss.n13556 0.0661418
R25313 vss.n13563 vss.n13561 0.0661418
R25314 vss.n13571 vss.n13569 0.0661418
R25315 vss.n13569 vss.n13568 0.0661418
R25316 vss.n13575 vss.n13570 0.0661418
R25317 vss.n13574 vss.n13570 0.0661418
R25318 vss.n13593 vss.n13588 0.0661418
R25319 vss.n13636 vss.n13635 0.0661418
R25320 vss.n13635 vss.n13611 0.0661418
R25321 vss.n13612 vss.n13605 0.0661418
R25322 vss.n13612 vss.n13610 0.0661418
R25323 vss.n13620 vss.n13618 0.0661418
R25324 vss.n13618 vss.n13617 0.0661418
R25325 vss.n13638 vss.n13637 0.0661418
R25326 vss.n13641 vss.n13638 0.0661418
R25327 vss.n13623 vss.n13619 0.0661418
R25328 vss.n13542 vss.n13541 0.0661418
R25329 vss.n13541 vss.n13518 0.0661418
R25330 vss.n13519 vss.n13512 0.0661418
R25331 vss.n13519 vss.n13517 0.0661418
R25332 vss.n13527 vss.n13525 0.0661418
R25333 vss.n13525 vss.n13524 0.0661418
R25334 vss.n13530 vss.n13526 0.0661418
R25335 vss.n13526 vss.n2103 0.0661418
R25336 vss.n8286 vss.n8285 0.0661418
R25337 vss.n8285 vss.n8261 0.0661418
R25338 vss.n8262 vss.n8255 0.0661418
R25339 vss.n8262 vss.n8260 0.0661418
R25340 vss.n8270 vss.n8268 0.0661418
R25341 vss.n8268 vss.n8267 0.0661418
R25342 vss.n8288 vss.n8287 0.0661418
R25343 vss.n8288 vss.n1765 0.0661418
R25344 vss.n8273 vss.n8269 0.0661418
R25345 vss.n13776 vss.n13775 0.0661418
R25346 vss.n13775 vss.n13752 0.0661418
R25347 vss.n13753 vss.n13746 0.0661418
R25348 vss.n13753 vss.n13751 0.0661418
R25349 vss.n13761 vss.n13759 0.0661418
R25350 vss.n13759 vss.n13758 0.0661418
R25351 vss.n13764 vss.n13760 0.0661418
R25352 vss.n13760 vss.n2107 0.0661418
R25353 vss.n13782 vss.n13777 0.0661418
R25354 vss.n13825 vss.n13824 0.0661418
R25355 vss.n13824 vss.n13800 0.0661418
R25356 vss.n13801 vss.n13794 0.0661418
R25357 vss.n13801 vss.n13799 0.0661418
R25358 vss.n13809 vss.n13807 0.0661418
R25359 vss.n13807 vss.n13806 0.0661418
R25360 vss.n13827 vss.n13826 0.0661418
R25361 vss.n13830 vss.n13827 0.0661418
R25362 vss.n13812 vss.n13808 0.0661418
R25363 vss.n13850 vss.n8227 0.0661418
R25364 vss.n13851 vss.n13850 0.0661418
R25365 vss.n8234 vss.n8233 0.0661418
R25366 vss.n8233 vss.n8231 0.0661418
R25367 vss.n8240 vss.n8239 0.0661418
R25368 vss.n8239 vss.n8237 0.0661418
R25369 vss.n8242 vss.n8241 0.0661418
R25370 vss.n8242 vss.n2111 0.0661418
R25371 vss.n9072 vss.n9071 0.0661418
R25372 vss.n9071 vss.n9047 0.0661418
R25373 vss.n9048 vss.n9041 0.0661418
R25374 vss.n9048 vss.n9046 0.0661418
R25375 vss.n9056 vss.n9054 0.0661418
R25376 vss.n9054 vss.n9053 0.0661418
R25377 vss.n9074 vss.n9073 0.0661418
R25378 vss.n9074 vss.n8223 0.0661418
R25379 vss.n9059 vss.n9055 0.0661418
R25380 vss.n13064 vss.n13063 0.0661418
R25381 vss.n13063 vss.n13040 0.0661418
R25382 vss.n13041 vss.n13034 0.0661418
R25383 vss.n13041 vss.n13039 0.0661418
R25384 vss.n13049 vss.n13047 0.0661418
R25385 vss.n13047 vss.n13046 0.0661418
R25386 vss.n13052 vss.n13048 0.0661418
R25387 vss.n13048 vss.n2115 0.0661418
R25388 vss.n13070 vss.n13065 0.0661418
R25389 vss.n13113 vss.n13112 0.0661418
R25390 vss.n13112 vss.n13088 0.0661418
R25391 vss.n13089 vss.n13082 0.0661418
R25392 vss.n13089 vss.n13087 0.0661418
R25393 vss.n13097 vss.n13095 0.0661418
R25394 vss.n13095 vss.n13094 0.0661418
R25395 vss.n13115 vss.n13114 0.0661418
R25396 vss.n13118 vss.n13115 0.0661418
R25397 vss.n13100 vss.n13096 0.0661418
R25398 vss.n9027 vss.n9026 0.0661418
R25399 vss.n9026 vss.n9003 0.0661418
R25400 vss.n9004 vss.n8997 0.0661418
R25401 vss.n9004 vss.n9002 0.0661418
R25402 vss.n9012 vss.n9010 0.0661418
R25403 vss.n9010 vss.n9009 0.0661418
R25404 vss.n9015 vss.n9011 0.0661418
R25405 vss.n9011 vss.n2119 0.0661418
R25406 vss.n12610 vss.n12609 0.0661418
R25407 vss.n12609 vss.n12585 0.0661418
R25408 vss.n12586 vss.n12579 0.0661418
R25409 vss.n12586 vss.n12584 0.0661418
R25410 vss.n12594 vss.n12592 0.0661418
R25411 vss.n12592 vss.n12591 0.0661418
R25412 vss.n12612 vss.n12611 0.0661418
R25413 vss.n12612 vss.n8095 0.0661418
R25414 vss.n12597 vss.n12593 0.0661418
R25415 vss.n2176 vss.n2175 0.0661418
R25416 vss.n2175 vss.n2152 0.0661418
R25417 vss.n2153 vss.n2146 0.0661418
R25418 vss.n2153 vss.n2151 0.0661418
R25419 vss.n2161 vss.n2159 0.0661418
R25420 vss.n2159 vss.n2158 0.0661418
R25421 vss.n2164 vss.n2160 0.0661418
R25422 vss.n2160 vss.n2123 0.0661418
R25423 vss.n14076 vss.n2177 0.0661418
R25424 vss.n2191 vss.n2190 0.0661418
R25425 vss.n2191 vss.n2188 0.0661418
R25426 vss.n2197 vss.n2196 0.0661418
R25427 vss.n2196 vss.n2194 0.0661418
R25428 vss.n2212 vss.n2184 0.0661418
R25429 vss.n2212 vss.n2189 0.0661418
R25430 vss.n2223 vss.n2222 0.0661418
R25431 vss.n2224 vss.n2223 0.0661418
R25432 vss.n2199 vss.n2198 0.0661418
R25433 vss.n2199 vss.n2127 0.0661418
R25434 vss.n2142 vss.n2141 0.0661418
R25435 vss.n2141 vss.n2136 0.0661418
R25436 vss.n9291 vss.n9288 0.0661418
R25437 vss.n9291 vss.n9290 0.0661418
R25438 vss.n2139 vss.n2132 0.0661418
R25439 vss.n2139 vss.n2137 0.0661418
R25440 vss.n14102 vss.n14101 0.0661418
R25441 vss.n14103 vss.n14102 0.0661418
R25442 vss.n9300 vss.n9299 0.0661418
R25443 vss.n9301 vss.n9300 0.0661418
R25444 vss.n9399 vss.n9392 0.0661418
R25445 vss.n9399 vss.n9397 0.0661418
R25446 vss.n9407 vss.n9405 0.0661418
R25447 vss.n9405 vss.n9404 0.0661418
R25448 vss.n12854 vss.n12853 0.0661418
R25449 vss.n12853 vss.n9398 0.0661418
R25450 vss.n12856 vss.n12855 0.0661418
R25451 vss.n12856 vss.n2126 0.0661418
R25452 vss.n12842 vss.n9406 0.0661418
R25453 vss.n12841 vss.n9406 0.0661418
R25454 vss.n12743 vss.n12742 0.0661418
R25455 vss.n12742 vss.n12737 0.0661418
R25456 vss.n12738 vss.n12732 0.0661418
R25457 vss.n12738 vss.n12736 0.0661418
R25458 vss.n12749 vss.n12748 0.0661418
R25459 vss.n12748 vss.n12746 0.0661418
R25460 vss.n12751 vss.n12750 0.0661418
R25461 vss.n12751 vss.n2122 0.0661418
R25462 vss.n12773 vss.n12772 0.0661418
R25463 vss.n12774 vss.n12773 0.0661418
R25464 vss.n8417 vss.n8410 0.0661418
R25465 vss.n8417 vss.n8415 0.0661418
R25466 vss.n8425 vss.n8423 0.0661418
R25467 vss.n8423 vss.n8422 0.0661418
R25468 vss.n13331 vss.n13330 0.0661418
R25469 vss.n13330 vss.n8416 0.0661418
R25470 vss.n13333 vss.n13332 0.0661418
R25471 vss.n13333 vss.n2114 0.0661418
R25472 vss.n13319 vss.n8424 0.0661418
R25473 vss.n13318 vss.n8424 0.0661418
R25474 vss.n13359 vss.n13352 0.0661418
R25475 vss.n13359 vss.n13357 0.0661418
R25476 vss.n13367 vss.n13365 0.0661418
R25477 vss.n13365 vss.n13364 0.0661418
R25478 vss.n13450 vss.n13449 0.0661418
R25479 vss.n13449 vss.n13358 0.0661418
R25480 vss.n13452 vss.n13451 0.0661418
R25481 vss.n13452 vss.n2106 0.0661418
R25482 vss.n13438 vss.n13366 0.0661418
R25483 vss.n13437 vss.n13366 0.0661418
R25484 vss.n2047 vss.n2046 0.0661418
R25485 vss.n2046 vss.n2041 0.0661418
R25486 vss.n2042 vss.n2035 0.0661418
R25487 vss.n2042 vss.n2040 0.0661418
R25488 vss.n11855 vss.n11852 0.0661418
R25489 vss.n11855 vss.n11854 0.0661418
R25490 vss.n11864 vss.n11863 0.0661418
R25491 vss.n11865 vss.n11864 0.0661418
R25492 vss.n2049 vss.n2048 0.0661418
R25493 vss.n14179 vss.n2049 0.0661418
R25494 vss.n14403 vss.n14401 0.0661418
R25495 vss.n1760 vss.n1758 0.0661418
R25496 vss.n1758 vss.n1757 0.0661418
R25497 vss.n1752 vss.n1745 0.0661418
R25498 vss.n1752 vss.n1750 0.0661418
R25499 vss.n14461 vss.n14460 0.0661418
R25500 vss.n14460 vss.n1751 0.0661418
R25501 vss.n14449 vss.n1759 0.0661418
R25502 vss.n14448 vss.n1759 0.0661418
R25503 vss.n14463 vss.n14462 0.0661418
R25504 vss.n1790 vss.n1789 0.0661418
R25505 vss.n1789 vss.n1787 0.0661418
R25506 vss.n1784 vss.n1783 0.0661418
R25507 vss.n1783 vss.n1776 0.0661418
R25508 vss.n1777 vss.n1772 0.0661418
R25509 vss.n1777 vss.n1775 0.0661418
R25510 vss.n1792 vss.n1791 0.0661418
R25511 vss.n1792 vss.n1192 0.0661418
R25512 vss.n1771 vss.n1768 0.0661418
R25513 vss.n14366 vss.n14365 0.0661418
R25514 vss.n14365 vss.n14359 0.0661418
R25515 vss.n14372 vss.n14371 0.0661418
R25516 vss.n14371 vss.n14369 0.0661418
R25517 vss.n14360 vss.n1819 0.0661418
R25518 vss.n14360 vss.n1815 0.0661418
R25519 vss.n1818 vss.n1814 0.0661418
R25520 vss.n14397 vss.n1814 0.0661418
R25521 vss.n14374 vss.n14373 0.0661418
R25522 vss.n1994 vss.n1987 0.0661418
R25523 vss.n1994 vss.n1992 0.0661418
R25524 vss.n2017 vss.n2016 0.0661418
R25525 vss.n2016 vss.n1993 0.0661418
R25526 vss.n2002 vss.n2000 0.0661418
R25527 vss.n2000 vss.n1999 0.0661418
R25528 vss.n2005 vss.n2001 0.0661418
R25529 vss.n2001 vss.n1185 0.0661418
R25530 vss.n2019 vss.n2018 0.0661418
R25531 vss.n2020 vss.n2019 0.0661418
R25532 vss.n14259 vss.n14255 0.0661418
R25533 vss.n14259 vss.n14250 0.0661418
R25534 vss.n14253 vss.n14241 0.0661418
R25535 vss.n14253 vss.n14250 0.0661418
R25536 vss.n14247 vss.n14245 0.0661418
R25537 vss.n14250 vss.n14245 0.0661418
R25538 vss.n14274 vss.n14246 0.0661418
R25539 vss.n14250 vss.n14246 0.0661418
R25540 vss.n14264 vss.n14263 0.0661418
R25541 vss.n14263 vss.n14250 0.0661418
R25542 vss.n14169 vss.n14168 0.0661418
R25543 vss.n14168 vss.n14167 0.0661418
R25544 vss.n1175 vss.n1168 0.0661418
R25545 vss.n1175 vss.n1173 0.0661418
R25546 vss.n1180 vss.n1179 0.0661418
R25547 vss.n1179 vss.n1174 0.0661418
R25548 vss.n1182 vss.n1181 0.0661418
R25549 vss.n14791 vss.n1182 0.0661418
R25550 vss.n14173 vss.n14172 0.0661418
R25551 vss.n14174 vss.n14173 0.0661418
R25552 vss.n14316 vss.n14315 0.0661418
R25553 vss.n14315 vss.n14288 0.0661418
R25554 vss.n14297 vss.n14283 0.0661418
R25555 vss.n14297 vss.n14288 0.0661418
R25556 vss.n14304 vss.n14303 0.0661418
R25557 vss.n14303 vss.n14288 0.0661418
R25558 vss.n14309 vss.n14302 0.0661418
R25559 vss.n14302 vss.n14288 0.0661418
R25560 vss.n14293 vss.n14291 0.0661418
R25561 vss.n14291 vss.n14288 0.0661418
R25562 vss.n14815 vss.n14814 0.0661418
R25563 vss.n14814 vss.n14809 0.0661418
R25564 vss.n14812 vss.n1166 0.0661418
R25565 vss.n14812 vss.n14810 0.0661418
R25566 vss.n14845 vss.n14844 0.0661418
R25567 vss.n14846 vss.n14845 0.0661418
R25568 vss.n15098 vss.n15096 0.0661418
R25569 vss.n981 vss.n979 0.0661418
R25570 vss.n979 vss.n978 0.0661418
R25571 vss.n973 vss.n966 0.0661418
R25572 vss.n973 vss.n971 0.0661418
R25573 vss.n15156 vss.n15155 0.0661418
R25574 vss.n15155 vss.n972 0.0661418
R25575 vss.n15144 vss.n980 0.0661418
R25576 vss.n15143 vss.n980 0.0661418
R25577 vss.n15158 vss.n15157 0.0661418
R25578 vss.n1011 vss.n1010 0.0661418
R25579 vss.n1010 vss.n1008 0.0661418
R25580 vss.n1005 vss.n1004 0.0661418
R25581 vss.n1004 vss.n997 0.0661418
R25582 vss.n998 vss.n993 0.0661418
R25583 vss.n998 vss.n996 0.0661418
R25584 vss.n1013 vss.n1012 0.0661418
R25585 vss.n1013 vss.n413 0.0661418
R25586 vss.n992 vss.n989 0.0661418
R25587 vss.n15061 vss.n15060 0.0661418
R25588 vss.n15060 vss.n15054 0.0661418
R25589 vss.n15067 vss.n15066 0.0661418
R25590 vss.n15066 vss.n15064 0.0661418
R25591 vss.n15055 vss.n1040 0.0661418
R25592 vss.n15055 vss.n1036 0.0661418
R25593 vss.n1039 vss.n1035 0.0661418
R25594 vss.n15092 vss.n1035 0.0661418
R25595 vss.n15069 vss.n15068 0.0661418
R25596 vss.n1099 vss.n1092 0.0661418
R25597 vss.n1099 vss.n1097 0.0661418
R25598 vss.n1122 vss.n1121 0.0661418
R25599 vss.n1121 vss.n1098 0.0661418
R25600 vss.n1107 vss.n1105 0.0661418
R25601 vss.n1105 vss.n1104 0.0661418
R25602 vss.n1110 vss.n1106 0.0661418
R25603 vss.n1106 vss.n406 0.0661418
R25604 vss.n1124 vss.n1123 0.0661418
R25605 vss.n1125 vss.n1124 0.0661418
R25606 vss.n14954 vss.n14950 0.0661418
R25607 vss.n14954 vss.n14945 0.0661418
R25608 vss.n14948 vss.n14936 0.0661418
R25609 vss.n14948 vss.n14945 0.0661418
R25610 vss.n14942 vss.n14940 0.0661418
R25611 vss.n14945 vss.n14940 0.0661418
R25612 vss.n14969 vss.n14941 0.0661418
R25613 vss.n14945 vss.n14941 0.0661418
R25614 vss.n14959 vss.n14958 0.0661418
R25615 vss.n14958 vss.n14945 0.0661418
R25616 vss.n14863 vss.n14862 0.0661418
R25617 vss.n14862 vss.n14861 0.0661418
R25618 vss.n396 vss.n389 0.0661418
R25619 vss.n396 vss.n394 0.0661418
R25620 vss.n401 vss.n400 0.0661418
R25621 vss.n400 vss.n395 0.0661418
R25622 vss.n403 vss.n402 0.0661418
R25623 vss.n15486 vss.n403 0.0661418
R25624 vss.n14867 vss.n14866 0.0661418
R25625 vss.n14868 vss.n14867 0.0661418
R25626 vss.n15011 vss.n15010 0.0661418
R25627 vss.n15010 vss.n14983 0.0661418
R25628 vss.n14992 vss.n14978 0.0661418
R25629 vss.n14992 vss.n14983 0.0661418
R25630 vss.n14999 vss.n14998 0.0661418
R25631 vss.n14998 vss.n14983 0.0661418
R25632 vss.n15004 vss.n14997 0.0661418
R25633 vss.n14997 vss.n14983 0.0661418
R25634 vss.n14988 vss.n14986 0.0661418
R25635 vss.n14986 vss.n14983 0.0661418
R25636 vss.n15507 vss.n387 0.0661418
R25637 vss.n15507 vss.n15505 0.0661418
R25638 vss.n15540 vss.n15539 0.0661418
R25639 vss.n15541 vss.n15540 0.0661418
R25640 vss.n6220 vss.n6219 0.0661418
R25641 vss.n6219 vss.n6213 0.0661418
R25642 vss.n6226 vss.n6225 0.0661418
R25643 vss.n6225 vss.n6223 0.0661418
R25644 vss.n6214 vss.n6209 0.0661418
R25645 vss.n6214 vss.n6205 0.0661418
R25646 vss.n6208 vss.n6204 0.0661418
R25647 vss.n6251 vss.n6204 0.0661418
R25648 vss.n6228 vss.n6227 0.0661418
R25649 vss.n36 vss.n29 0.0661418
R25650 vss.n36 vss.n34 0.0661418
R25651 vss.n41 vss.n40 0.0661418
R25652 vss.n40 vss.n35 0.0661418
R25653 vss.n3961 vss.n3960 0.0661418
R25654 vss.n3960 vss.n3949 0.0661418
R25655 vss.n3952 vss.n3948 0.0661418
R25656 vss.n3966 vss.n3948 0.0661418
R25657 vss.n43 vss.n42 0.0661418
R25658 vss.n15856 vss.n43 0.0661418
R25659 vss.n3866 vss.n3865 0.0661418
R25660 vss.n3865 vss.n3859 0.0661418
R25661 vss.n3872 vss.n3871 0.0661418
R25662 vss.n3871 vss.n3869 0.0661418
R25663 vss.n3860 vss.n3855 0.0661418
R25664 vss.n3860 vss.n3851 0.0661418
R25665 vss.n3854 vss.n3850 0.0661418
R25666 vss.n3897 vss.n3850 0.0661418
R25667 vss.n3874 vss.n3873 0.0661418
R25668 vss.n3875 vss.n3874 0.0661418
R25669 vss.n3747 vss.n3746 0.0661418
R25670 vss.n3746 vss.n3740 0.0661418
R25671 vss.n3753 vss.n3752 0.0661418
R25672 vss.n3752 vss.n3750 0.0661418
R25673 vss.n3741 vss.n3736 0.0661418
R25674 vss.n3741 vss.n3732 0.0661418
R25675 vss.n3735 vss.n3731 0.0661418
R25676 vss.n3778 vss.n3731 0.0661418
R25677 vss.n3755 vss.n3754 0.0661418
R25678 vss.n3756 vss.n3755 0.0661418
R25679 vss.n3628 vss.n3627 0.0661418
R25680 vss.n3627 vss.n3621 0.0661418
R25681 vss.n3634 vss.n3633 0.0661418
R25682 vss.n3633 vss.n3631 0.0661418
R25683 vss.n3622 vss.n3617 0.0661418
R25684 vss.n3622 vss.n3613 0.0661418
R25685 vss.n3616 vss.n3612 0.0661418
R25686 vss.n3659 vss.n3612 0.0661418
R25687 vss.n3636 vss.n3635 0.0661418
R25688 vss.n3637 vss.n3636 0.0661418
R25689 vss.n6304 vss.n6303 0.0661418
R25690 vss.n6303 vss.n6302 0.0661418
R25691 vss.n251 vss.n244 0.0661418
R25692 vss.n251 vss.n249 0.0661418
R25693 vss.n256 vss.n255 0.0661418
R25694 vss.n255 vss.n250 0.0661418
R25695 vss.n258 vss.n257 0.0661418
R25696 vss.n15688 vss.n258 0.0661418
R25697 vss.n6308 vss.n6307 0.0661418
R25698 vss.n6309 vss.n6308 0.0661418
R25699 vss.n15597 vss.n15593 0.0661418
R25700 vss.n15597 vss.n15588 0.0661418
R25701 vss.n15591 vss.n15579 0.0661418
R25702 vss.n15591 vss.n15588 0.0661418
R25703 vss.n15585 vss.n15583 0.0661418
R25704 vss.n15588 vss.n15583 0.0661418
R25705 vss.n15612 vss.n15584 0.0661418
R25706 vss.n15588 vss.n15584 0.0661418
R25707 vss.n15602 vss.n15601 0.0661418
R25708 vss.n15601 vss.n15588 0.0661418
R25709 vss.n319 vss.n318 0.0661418
R25710 vss.n318 vss.n312 0.0661418
R25711 vss.n325 vss.n324 0.0661418
R25712 vss.n324 vss.n322 0.0661418
R25713 vss.n313 vss.n309 0.0661418
R25714 vss.n313 vss.n305 0.0661418
R25715 vss.n308 vss.n304 0.0661418
R25716 vss.n350 vss.n304 0.0661418
R25717 vss.n327 vss.n326 0.0661418
R25718 vss.n328 vss.n327 0.0661418
R25719 vss.n3584 vss.n3583 0.0661418
R25720 vss.n3583 vss.n3581 0.0661418
R25721 vss.n3578 vss.n3577 0.0661418
R25722 vss.n3577 vss.n3572 0.0661418
R25723 vss.n3575 vss.n3568 0.0661418
R25724 vss.n3575 vss.n3573 0.0661418
R25725 vss.n3610 vss.n3609 0.0661418
R25726 vss.n3611 vss.n3610 0.0661418
R25727 vss.n3560 vss.n3559 0.0661418
R25728 vss.n3586 vss.n3585 0.0661418
R25729 vss.n15635 vss.n15634 0.0661418
R25730 vss.n15634 vss.n353 0.0661418
R25731 vss.n15631 vss.n15630 0.0661418
R25732 vss.n15630 vss.n353 0.0661418
R25733 vss.n15625 vss.n15623 0.0661418
R25734 vss.n15625 vss.n353 0.0661418
R25735 vss.n15651 vss.n15650 0.0661418
R25736 vss.n15650 vss.n353 0.0661418
R25737 vss.n15640 vss.n15639 0.0661418
R25738 vss.n15639 vss.n353 0.0661418
R25739 vss.n367 vss.n360 0.0661418
R25740 vss.n367 vss.n365 0.0661418
R25741 vss.n15560 vss.n15559 0.0661418
R25742 vss.n15559 vss.n366 0.0661418
R25743 vss.n375 vss.n373 0.0661418
R25744 vss.n373 vss.n372 0.0661418
R25745 vss.n15548 vss.n374 0.0661418
R25746 vss.n15547 vss.n374 0.0661418
R25747 vss.n15562 vss.n15561 0.0661418
R25748 vss.n15562 vss.n303 0.0661418
R25749 vss.n12145 vss.n12137 0.0661418
R25750 vss.n12145 vss.n12143 0.0661418
R25751 vss.n12150 vss.n12149 0.0661418
R25752 vss.n12149 vss.n12144 0.0661418
R25753 vss.n12156 vss.n12155 0.0661418
R25754 vss.n12155 vss.n12153 0.0661418
R25755 vss.n12158 vss.n12157 0.0661418
R25756 vss.n12158 vss.n12132 0.0661418
R25757 vss.n12179 vss.n12178 0.0661418
R25758 vss.n12180 vss.n12179 0.0661418
R25759 vss.n11769 vss.n11766 0.0661418
R25760 vss.n11771 vss.n11765 0.0661418
R25761 vss.n11765 vss.n11763 0.0661418
R25762 vss.n11773 vss.n11758 0.0661418
R25763 vss.n11773 vss.n11763 0.0661418
R25764 vss.n11779 vss.n11778 0.0661418
R25765 vss.n11778 vss.n11763 0.0661418
R25766 vss.n11783 vss.n11777 0.0661418
R25767 vss.n11777 vss.n11763 0.0661418
R25768 vss.n8831 vss.n8830 0.0661418
R25769 vss.n8830 vss.n8828 0.0661418
R25770 vss.n8825 vss.n8824 0.0661418
R25771 vss.n8824 vss.n8819 0.0661418
R25772 vss.n8822 vss.n8815 0.0661418
R25773 vss.n8822 vss.n8820 0.0661418
R25774 vss.n13247 vss.n13246 0.0661418
R25775 vss.n13248 vss.n13247 0.0661418
R25776 vss.n8833 vss.n8832 0.0661418
R25777 vss.n13225 vss.n8833 0.0661418
R25778 vss.n11716 vss.n9883 0.0661418
R25779 vss.n11717 vss.n11716 0.0661418
R25780 vss.n9890 vss.n9889 0.0661418
R25781 vss.n9889 vss.n9887 0.0661418
R25782 vss.n9896 vss.n9895 0.0661418
R25783 vss.n9895 vss.n9893 0.0661418
R25784 vss.n11724 vss.n11723 0.0661418
R25785 vss.n11725 vss.n11724 0.0661418
R25786 vss.n9898 vss.n9897 0.0661418
R25787 vss.n11545 vss.n11544 0.0661418
R25788 vss.n11544 vss.n11521 0.0661418
R25789 vss.n11522 vss.n11515 0.0661418
R25790 vss.n11522 vss.n11520 0.0661418
R25791 vss.n11530 vss.n11528 0.0661418
R25792 vss.n11528 vss.n11527 0.0661418
R25793 vss.n11533 vss.n11529 0.0661418
R25794 vss.n11529 vss.n8837 0.0661418
R25795 vss.n11551 vss.n11546 0.0661418
R25796 vss.n11594 vss.n11593 0.0661418
R25797 vss.n11593 vss.n11569 0.0661418
R25798 vss.n11570 vss.n11563 0.0661418
R25799 vss.n11570 vss.n11568 0.0661418
R25800 vss.n11578 vss.n11576 0.0661418
R25801 vss.n11576 vss.n11575 0.0661418
R25802 vss.n11596 vss.n11595 0.0661418
R25803 vss.n11599 vss.n11596 0.0661418
R25804 vss.n11581 vss.n11577 0.0661418
R25805 vss.n11501 vss.n11500 0.0661418
R25806 vss.n11500 vss.n11477 0.0661418
R25807 vss.n11478 vss.n11471 0.0661418
R25808 vss.n11478 vss.n11476 0.0661418
R25809 vss.n11486 vss.n11484 0.0661418
R25810 vss.n11484 vss.n11483 0.0661418
R25811 vss.n11489 vss.n11485 0.0661418
R25812 vss.n11485 vss.n8841 0.0661418
R25813 vss.n11141 vss.n11140 0.0661418
R25814 vss.n11140 vss.n11116 0.0661418
R25815 vss.n11117 vss.n11110 0.0661418
R25816 vss.n11117 vss.n11115 0.0661418
R25817 vss.n11125 vss.n11123 0.0661418
R25818 vss.n11123 vss.n11122 0.0661418
R25819 vss.n11143 vss.n11142 0.0661418
R25820 vss.n11143 vss.n9803 0.0661418
R25821 vss.n11128 vss.n11124 0.0661418
R25822 vss.n11234 vss.n11233 0.0661418
R25823 vss.n11233 vss.n11210 0.0661418
R25824 vss.n11211 vss.n11204 0.0661418
R25825 vss.n11211 vss.n11209 0.0661418
R25826 vss.n11219 vss.n11217 0.0661418
R25827 vss.n11217 vss.n11216 0.0661418
R25828 vss.n11222 vss.n11218 0.0661418
R25829 vss.n11218 vss.n8845 0.0661418
R25830 vss.n11240 vss.n11235 0.0661418
R25831 vss.n11283 vss.n11282 0.0661418
R25832 vss.n11282 vss.n11258 0.0661418
R25833 vss.n11259 vss.n11252 0.0661418
R25834 vss.n11259 vss.n11257 0.0661418
R25835 vss.n11267 vss.n11265 0.0661418
R25836 vss.n11265 vss.n11264 0.0661418
R25837 vss.n11285 vss.n11284 0.0661418
R25838 vss.n11288 vss.n11285 0.0661418
R25839 vss.n11270 vss.n11266 0.0661418
R25840 vss.n11096 vss.n11095 0.0661418
R25841 vss.n11095 vss.n11072 0.0661418
R25842 vss.n11073 vss.n11066 0.0661418
R25843 vss.n11073 vss.n11071 0.0661418
R25844 vss.n11081 vss.n11079 0.0661418
R25845 vss.n11079 vss.n11078 0.0661418
R25846 vss.n11084 vss.n11080 0.0661418
R25847 vss.n11080 vss.n8849 0.0661418
R25848 vss.n10944 vss.n10943 0.0661418
R25849 vss.n10943 vss.n10919 0.0661418
R25850 vss.n10920 vss.n10913 0.0661418
R25851 vss.n10920 vss.n10918 0.0661418
R25852 vss.n10928 vss.n10926 0.0661418
R25853 vss.n10926 vss.n10925 0.0661418
R25854 vss.n10946 vss.n10945 0.0661418
R25855 vss.n10946 vss.n9674 0.0661418
R25856 vss.n10931 vss.n10927 0.0661418
R25857 vss.n10895 vss.n10894 0.0661418
R25858 vss.n10894 vss.n10871 0.0661418
R25859 vss.n10872 vss.n10865 0.0661418
R25860 vss.n10872 vss.n10870 0.0661418
R25861 vss.n10880 vss.n10878 0.0661418
R25862 vss.n10878 vss.n10877 0.0661418
R25863 vss.n10883 vss.n10879 0.0661418
R25864 vss.n10879 vss.n8853 0.0661418
R25865 vss.n10901 vss.n10896 0.0661418
R25866 vss.n10848 vss.n10847 0.0661418
R25867 vss.n10847 vss.n10823 0.0661418
R25868 vss.n10824 vss.n10817 0.0661418
R25869 vss.n10824 vss.n10822 0.0661418
R25870 vss.n10832 vss.n10830 0.0661418
R25871 vss.n10830 vss.n10829 0.0661418
R25872 vss.n10850 vss.n10849 0.0661418
R25873 vss.n10853 vss.n10850 0.0661418
R25874 vss.n10835 vss.n10831 0.0661418
R25875 vss.n10199 vss.n10198 0.0661418
R25876 vss.n10198 vss.n10175 0.0661418
R25877 vss.n10176 vss.n10169 0.0661418
R25878 vss.n10176 vss.n10174 0.0661418
R25879 vss.n10184 vss.n10182 0.0661418
R25880 vss.n10182 vss.n10181 0.0661418
R25881 vss.n10187 vss.n10183 0.0661418
R25882 vss.n10183 vss.n8857 0.0661418
R25883 vss.n10550 vss.n10549 0.0661418
R25884 vss.n10549 vss.n10525 0.0661418
R25885 vss.n10526 vss.n10519 0.0661418
R25886 vss.n10526 vss.n10524 0.0661418
R25887 vss.n10534 vss.n10532 0.0661418
R25888 vss.n10532 vss.n10531 0.0661418
R25889 vss.n10552 vss.n10551 0.0661418
R25890 vss.n10552 vss.n9545 0.0661418
R25891 vss.n10537 vss.n10533 0.0661418
R25892 vss.n10501 vss.n10500 0.0661418
R25893 vss.n10500 vss.n10477 0.0661418
R25894 vss.n10478 vss.n10471 0.0661418
R25895 vss.n10478 vss.n10476 0.0661418
R25896 vss.n10486 vss.n10484 0.0661418
R25897 vss.n10484 vss.n10483 0.0661418
R25898 vss.n10489 vss.n10485 0.0661418
R25899 vss.n10485 vss.n8861 0.0661418
R25900 vss.n10507 vss.n10502 0.0661418
R25901 vss.n10431 vss.n10424 0.0661418
R25902 vss.n10431 vss.n10429 0.0661418
R25903 vss.n10439 vss.n10437 0.0661418
R25904 vss.n10437 vss.n10436 0.0661418
R25905 vss.n10454 vss.n10453 0.0661418
R25906 vss.n10453 vss.n10430 0.0661418
R25907 vss.n10456 vss.n10455 0.0661418
R25908 vss.n10457 vss.n10456 0.0661418
R25909 vss.n10442 vss.n10438 0.0661418
R25910 vss.n10438 vss.n8865 0.0661418
R25911 vss.n10576 vss.n10569 0.0661418
R25912 vss.n10576 vss.n10574 0.0661418
R25913 vss.n10584 vss.n10582 0.0661418
R25914 vss.n10582 vss.n10581 0.0661418
R25915 vss.n10600 vss.n10599 0.0661418
R25916 vss.n10599 vss.n10575 0.0661418
R25917 vss.n10602 vss.n10601 0.0661418
R25918 vss.n10602 vss.n8860 0.0661418
R25919 vss.n10588 vss.n10583 0.0661418
R25920 vss.n10587 vss.n10583 0.0661418
R25921 vss.n10970 vss.n10963 0.0661418
R25922 vss.n10970 vss.n10968 0.0661418
R25923 vss.n10978 vss.n10976 0.0661418
R25924 vss.n10976 vss.n10975 0.0661418
R25925 vss.n10994 vss.n10993 0.0661418
R25926 vss.n10993 vss.n10969 0.0661418
R25927 vss.n10996 vss.n10995 0.0661418
R25928 vss.n10996 vss.n8852 0.0661418
R25929 vss.n10982 vss.n10977 0.0661418
R25930 vss.n10981 vss.n10977 0.0661418
R25931 vss.n10007 vss.n10006 0.0661418
R25932 vss.n10006 vss.n10001 0.0661418
R25933 vss.n10002 vss.n9996 0.0661418
R25934 vss.n10002 vss.n10000 0.0661418
R25935 vss.n10013 vss.n10012 0.0661418
R25936 vss.n10012 vss.n10010 0.0661418
R25937 vss.n10015 vss.n10014 0.0661418
R25938 vss.n10015 vss.n8844 0.0661418
R25939 vss.n10037 vss.n10036 0.0661418
R25940 vss.n10038 vss.n10037 0.0661418
R25941 vss.n11625 vss.n11620 0.0661418
R25942 vss.n11623 vss.n11620 0.0661418
R25943 vss.n11639 vss.n11638 0.0661418
R25944 vss.n11640 vss.n11639 0.0661418
R25945 vss.n9957 vss.n9952 0.0661418
R25946 vss.n9957 vss.n9956 0.0661418
R25947 vss.n11647 vss.n11646 0.0661418
R25948 vss.n11648 vss.n11647 0.0661418
R25949 vss.n11629 vss.n11621 0.0661418
R25950 vss.n11621 vss.n8836 0.0661418
R25951 vss.n9600 vss 0.0465526
R25952 vss.n9730 vss 0.0465526
R25953 vss.n12194 vss 0.0465526
R25954 vss.n12312 vss 0.0465526
R25955 vss.n12431 vss 0.0465526
R25956 vss.n9471 vss 0.0465526
R25957 vss.n9470 vss 0.0465526
R25958 vss.n6157 vss 0.0465526
R25959 vss.n5918 vss 0.0465526
R25960 vss.n3541 vss 0.0465526
R25961 vss.n7349 vss 0.0465526
R25962 vss.n15173 vss 0.0465526
R25963 vss.n7446 vss 0.0465526
R25964 vss.n7300 vss 0.0465526
R25965 vss.n4653 vss 0.0465526
R25966 vss.n4606 vss 0.0465526
R25967 vss.n8150 vss 0.0465526
R25968 vss.n14478 vss 0.0465526
R25969 vss.n13911 vss 0.0465526
R25970 vss.n14028 vss 0.0465526
R25971 vss.n8050 vss 0.0465526
R25972 vss.n2324 vss 0.0465526
R25973 vss.n14356 vss 0.0465526
R25974 vss.n14282 vss 0.0465526
R25975 vss.n15051 vss 0.0465526
R25976 vss.n14977 vss 0.0465526
R25977 vss.n6210 vss 0.0465526
R25978 vss.n6063 vss 0.0465526
R25979 vss.n5823 vss 0.0465526
R25980 vss.n5679 vss 0.0465526
R25981 vss.n15620 vss 0.0465526
R25982 vss.n11802 vss 0.0465526
R25983 vss.n11792 vss.n11766 0.033698
R25984 vss.n10508 vss.n10507 0.0290121
R25985 vss.n10902 vss.n10901 0.0290121
R25986 vss.n11241 vss.n11240 0.0290121
R25987 vss.n11552 vss.n11551 0.0290121
R25988 vss.n9782 vss.n9781 0.0290121
R25989 vss.n9753 vss.n9746 0.0290121
R25990 vss.n12333 vss.n12330 0.0290121
R25991 vss.n9653 vss.n9652 0.0290121
R25992 vss.n9623 vss.n9616 0.0290121
R25993 vss.n12452 vss.n12449 0.0290121
R25994 vss.n9523 vss.n9522 0.0290121
R25995 vss.n9494 vss.n9487 0.0290121
R25996 vss.n9460 vss.n9456 0.0290121
R25997 vss.n12215 vss.n12212 0.0290121
R25998 vss.n5702 vss.n5699 0.0290121
R25999 vss.n5557 vss.n5555 0.0290121
R26000 vss.n5940 vss.n5937 0.0290121
R26001 vss.n5812 vss.n5808 0.0290121
R26002 vss.n5745 vss.n5743 0.0290121
R26003 vss.n6179 vss.n6176 0.0290121
R26004 vss.n6052 vss.n6048 0.0290121
R26005 vss.n5985 vss.n5983 0.0290121
R26006 vss.n4483 vss.n4482 0.0290121
R26007 vss.n4213 vss.n4212 0.0290121
R26008 vss.n5528 vss.n4007 0.0290121
R26009 vss.n6367 vss.n3440 0.0290121
R26010 vss.n3337 vss.n3336 0.0290121
R26011 vss.n3464 vss.n3459 0.0290121
R26012 vss.n5279 vss.n5272 0.0290121
R26013 vss.n5494 vss.n5487 0.0290121
R26014 vss.n5068 vss.n5061 0.0290121
R26015 vss.n5020 vss.n5013 0.0290121
R26016 vss.n4515 vss.n4508 0.0290121
R26017 vss.n14909 vss.n14902 0.0290121
R26018 vss.n7467 vss.n7464 0.0290121
R26019 vss.n7373 vss.n7372 0.0290121
R26020 vss.n3080 vss.n3078 0.0290121
R26021 vss.n7290 vss.n7289 0.0290121
R26022 vss.n4643 vss.n4639 0.0290121
R26023 vss.n4671 vss.n4669 0.0290121
R26024 vss.n4596 vss.n4592 0.0290121
R26025 vss.n7215 vss.n3137 0.0290121
R26026 vss.n7983 vss.n2458 0.0290121
R26027 vss.n2922 vss.n2889 0.0290121
R26028 vss.n2672 vss.n2663 0.0290121
R26029 vss.n7928 vss.n7927 0.0290121
R26030 vss.n7886 vss.n7879 0.0290121
R26031 vss.n7740 vss.n7733 0.0290121
R26032 vss.n7691 vss.n7684 0.0290121
R26033 vss.n2997 vss.n2990 0.0290121
R26034 vss.n7079 vss.n7078 0.0290121
R26035 vss.n6827 vss.n6826 0.0290121
R26036 vss.n14214 vss.n14207 0.0290121
R26037 vss.n13932 vss.n13929 0.0290121
R26038 vss.n8202 vss.n8201 0.0290121
R26039 vss.n8173 vss.n8166 0.0290121
R26040 vss.n14049 vss.n14046 0.0290121
R26041 vss.n8074 vss.n8073 0.0290121
R26042 vss.n2247 vss.n2245 0.0290121
R26043 vss.n2314 vss.n2310 0.0290121
R26044 vss.n14077 vss.n14076 0.0290121
R26045 vss.n13071 vss.n13070 0.0290121
R26046 vss.n13783 vss.n13782 0.0290121
R26047 vss.n13594 vss.n13593 0.0290121
R26048 vss.n2078 vss.n2073 0.0290121
R26049 vss.n13626 vss.n13619 0.0290121
R26050 vss.n8276 vss.n8269 0.0290121
R26051 vss.n13815 vss.n13808 0.0290121
R26052 vss.n9062 vss.n9055 0.0290121
R26053 vss.n13103 vss.n13096 0.0290121
R26054 vss.n12600 vss.n12593 0.0290121
R26055 vss.n14412 vss.n14401 0.0290121
R26056 vss.n14467 vss.n14463 0.0290121
R26057 vss.n14377 vss.n14374 0.0290121
R26058 vss.n15107 vss.n15096 0.0290121
R26059 vss.n15162 vss.n15158 0.0290121
R26060 vss.n15072 vss.n15069 0.0290121
R26061 vss.n6231 vss.n6228 0.0290121
R26062 vss.n3563 vss.n3560 0.0290121
R26063 vss.n3589 vss.n3586 0.0290121
R26064 vss.n9902 vss.n9898 0.0290121
R26065 vss.n11584 vss.n11577 0.0290121
R26066 vss.n11131 vss.n11124 0.0290121
R26067 vss.n11273 vss.n11266 0.0290121
R26068 vss.n10934 vss.n10927 0.0290121
R26069 vss.n10838 vss.n10831 0.0290121
R26070 vss.n10540 vss.n10533 0.0290121
R26071 vss.n11615 vss.n9964 0.021882
R26072 vss.n11305 vss.n11304 0.021882
R26073 vss.n10641 vss.n10167 0.021882
R26074 vss.n13673 vss.n8338 0.021882
R26075 vss.n13703 vss.n13702 0.021882
R26076 vss.n13292 vss.n13291 0.021882
R26077 vss.n12991 vss.n8617 0.021882
R26078 vss.n13150 vss.n8882 0.021882
R26079 vss.n13181 vss.n8880 0.021882
R26080 vss.n13179 vss.n8881 0.021882
R26081 vss.n15731 vss.n163 0.021882
R26082 vss.n15787 vss.n85 0.021882
R26083 vss.n15843 vss.n27 0.021882
R26084 vss.n15223 vss.n15222 0.021882
R26085 vss.n15266 vss.n759 0.021882
R26086 vss.n15343 vss.n15342 0.021882
R26087 vss.n15373 vss.n15372 0.021882
R26088 vss.n15416 vss.n501 0.021882
R26089 vss.n15448 vss.n15447 0.021882
R26090 vss.n15445 vss.n500 0.021882
R26091 vss.n14528 vss.n14527 0.021882
R26092 vss.n14571 vss.n1538 0.021882
R26093 vss.n14648 vss.n14647 0.021882
R26094 vss.n14678 vss.n14677 0.021882
R26095 vss.n14721 vss.n1280 0.021882
R26096 vss.n14753 vss.n14752 0.021882
R26097 vss.n14750 vss.n1279 0.021882
R26098 vss.n14327 vss.n14326 0.021882
R26099 vss.n15022 vss.n15021 0.021882
R26100 vss.n15816 vss.n15815 0.021882
R26101 vss.n15760 vss.n15759 0.021882
R26102 vss.n15704 vss.n15703 0.021882
R26103 vss.n15674 vss.n242 0.021882
R26104 vss.n12190 vss.n9859 0.021882
R26105 vss.n10618 vss.n10617 0.021882
R26106 vss.n11011 vss.n11010 0.021882
R26107 vss.n11331 vss.n9965 0.021882
R26108 vss.n11617 vss.n9935 0.021882
R26109 vss.n10369 vss.n10254 0.021882
R26110 vss.n15872 vss.n15871 0.021882
R26111 vss vss 0.0202368
R26112 vss vss 0.0202368
R26113 vss vss 0.0202368
R26114 vss vss 0.0202368
R26115 vss vss 0.0185921
R26116 vss vss 0.0185921
R26117 vss vss 0.0169474
R26118 vss vss 0.0169474
R26119 vss.n10565 vss 0.0136579
R26120 vss.n10959 vss 0.0136579
R26121 vss.n11156 vss 0.0136579
R26122 vss.n11710 vss 0.0136579
R26123 vss.n4540 vss 0.0136579
R26124 vss vss 0.0136579
R26125 vss.n5305 vss 0.0136579
R26126 vss.n5093 vss 0.0136579
R26127 vss.n4998 vss 0.0136579
R26128 vss.n5472 vss 0.0136579
R26129 vss.n6377 vss 0.0136579
R26130 vss.n6662 vss 0.0136579
R26131 vss.n3273 vss 0.0136579
R26132 vss.n6878 vss 0.0136579
R26133 vss vss 0.0136579
R26134 vss.n7765 vss 0.0136579
R26135 vss.n7501 vss 0.0136579
R26136 vss.n7993 vss 0.0136579
R26137 vss.n7669 vss 0.0136579
R26138 vss.n7864 vss 0.0136579
R26139 vss.n14882 vss 0.0136579
R26140 vss.n3149 vss 0.0136579
R26141 vss.n12625 vss 0.0136579
R26142 vss.n9087 vss 0.0136579
R26143 vss.n8301 vss 0.0136579
R26144 vss.n14140 vss 0.0136579
R26145 vss.n14089 vss 0.0136579
R26146 vss.n13130 vss 0.0136579
R26147 vss.n13842 vss 0.0136579
R26148 vss.n13653 vss 0.0136579
R26149 vss vss 0.0136579
R26150 vss.n8879 vss 0.0136579
R26151 vss.n10816 vss 0.0136579
R26152 vss.n11300 vss 0.0136579
R26153 vss.n11611 vss 0.0136579
R26154 vss vss 0.0136579
R26155 vss.n3242 vss.n3241 0.0126193
R26156 vss.n3244 vss.n3241 0.0126193
R26157 vss.n3255 vss.n3254 0.0126193
R26158 vss.n3254 vss.n3236 0.0126193
R26159 vss.n3270 vss.n3269 0.0126193
R26160 vss.n3269 vss.n3268 0.0126193
R26161 vss.n3223 vss.n3222 0.0126193
R26162 vss.n3222 vss.n3210 0.0126193
R26163 vss.n3216 vss.n3215 0.0126193
R26164 vss.n3215 vss.n2358 0.0126193
R26165 vss.n2425 vss.n2423 0.0126193
R26166 vss.n2423 vss.n2420 0.0126193
R26167 vss.n8013 vss.n8012 0.0126193
R26168 vss.n8012 vss.n8011 0.0126193
R26169 vss.n8000 vss.n7999 0.0126193
R26170 vss.n8001 vss.n8000 0.0126193
R26171 vss.n6956 vss.n6955 0.0126193
R26172 vss.n6955 vss.n6943 0.0126193
R26173 vss.n6949 vss.n6948 0.0126193
R26174 vss.n6948 vss.n1315 0.0126193
R26175 vss.n1398 vss.n1394 0.0126193
R26176 vss.n1398 vss.n1397 0.0126193
R26177 vss.n1402 vss.n1401 0.0126193
R26178 vss.n1401 vss.n1382 0.0126193
R26179 vss.n14707 vss.n14706 0.0126193
R26180 vss.n14706 vss.n14705 0.0126193
R26181 vss.n1415 vss.n1410 0.0126193
R26182 vss.n1410 vss.n1408 0.0126193
R26183 vss.n1418 vss.n1411 0.0126193
R26184 vss.n14692 vss.n1411 0.0126193
R26185 vss.n7546 vss.n7545 0.0126193
R26186 vss.n7547 vss.n7546 0.0126193
R26187 vss.n7559 vss.n7558 0.0126193
R26188 vss.n7560 vss.n7559 0.0126193
R26189 vss.n7572 vss.n7571 0.0126193
R26190 vss.n7571 vss.n7570 0.0126193
R26191 vss.n7585 vss.n7584 0.0126193
R26192 vss.n7584 vss.n7525 0.0126193
R26193 vss.n7578 vss.n7577 0.0126193
R26194 vss.n7577 vss.n1520 0.0126193
R26195 vss.n2764 vss.n2763 0.0126193
R26196 vss.n2765 vss.n2764 0.0126193
R26197 vss.n2777 vss.n2776 0.0126193
R26198 vss.n2778 vss.n2777 0.0126193
R26199 vss.n2790 vss.n2789 0.0126193
R26200 vss.n2789 vss.n2788 0.0126193
R26201 vss.n2803 vss.n2802 0.0126193
R26202 vss.n2802 vss.n2743 0.0126193
R26203 vss.n2796 vss.n2795 0.0126193
R26204 vss.n2795 vss.n1573 0.0126193
R26205 vss.n1655 vss.n1651 0.0126193
R26206 vss.n1655 vss.n1654 0.0126193
R26207 vss.n1659 vss.n1658 0.0126193
R26208 vss.n1658 vss.n1639 0.0126193
R26209 vss.n14557 vss.n14556 0.0126193
R26210 vss.n14556 vss.n14555 0.0126193
R26211 vss.n1672 vss.n1667 0.0126193
R26212 vss.n1667 vss.n1665 0.0126193
R26213 vss.n1675 vss.n1668 0.0126193
R26214 vss.n14542 vss.n1668 0.0126193
R26215 vss.n2532 vss.n2531 0.0126193
R26216 vss.n2533 vss.n2532 0.0126193
R26217 vss.n2543 vss.n2542 0.0126193
R26218 vss.n2544 vss.n2543 0.0126193
R26219 vss.n2556 vss.n2555 0.0126193
R26220 vss.n2555 vss.n2554 0.0126193
R26221 vss.n2568 vss.n2567 0.0126193
R26222 vss.n2567 vss.n2507 0.0126193
R26223 vss.n2561 vss.n2560 0.0126193
R26224 vss.n2560 vss.n1853 0.0126193
R26225 vss.n1888 vss.n1887 0.0126193
R26226 vss.n1887 vss.n1886 0.0126193
R26227 vss.n1893 vss.n1892 0.0126193
R26228 vss.n1892 vss.n1873 0.0126193
R26229 vss.n1973 vss.n1972 0.0126193
R26230 vss.n1972 vss.n1971 0.0126193
R26231 vss.n1952 vss.n1947 0.0126193
R26232 vss.n1947 vss.n1945 0.0126193
R26233 vss.n1955 vss.n1948 0.0126193
R26234 vss.n1958 vss.n1948 0.0126193
R26235 vss.n1865 vss.n1859 0.0126193
R26236 vss.n1865 vss.n1863 0.0126193
R26237 vss.n1884 vss.n1869 0.0126193
R26238 vss.n1885 vss.n1884 0.0126193
R26239 vss.n1980 vss.n1979 0.0126193
R26240 vss.n1979 vss.n1978 0.0126193
R26241 vss.n1969 vss.n1968 0.0126193
R26242 vss.n1970 vss.n1969 0.0126193
R26243 vss.n14337 vss.n14336 0.0126193
R26244 vss.n14338 vss.n14337 0.0126193
R26245 vss.n1690 vss.n1684 0.0126193
R26246 vss.n1690 vss.n1688 0.0126193
R26247 vss.n2534 vss.n1694 0.0126193
R26248 vss.n2535 vss.n2534 0.0126193
R26249 vss.n2547 vss.n2546 0.0126193
R26250 vss.n2546 vss.n2545 0.0126193
R26251 vss.n2550 vss.n2518 0.0126193
R26252 vss.n2518 vss.n2506 0.0126193
R26253 vss.n14538 vss.n14537 0.0126193
R26254 vss.n14539 vss.n14538 0.0126193
R26255 vss.n1631 vss.n1579 0.0126193
R26256 vss.n1631 vss.n1583 0.0126193
R26257 vss.n1652 vss.n1635 0.0126193
R26258 vss.n1653 vss.n1652 0.0126193
R26259 vss.n14564 vss.n14563 0.0126193
R26260 vss.n14563 vss.n14562 0.0126193
R26261 vss.n14553 vss.n14552 0.0126193
R26262 vss.n14554 vss.n14553 0.0126193
R26263 vss.n14581 vss.n14580 0.0126193
R26264 vss.n14582 vss.n14581 0.0126193
R26265 vss.n1532 vss.n1526 0.0126193
R26266 vss.n1532 vss.n1530 0.0126193
R26267 vss.n2766 vss.n1536 0.0126193
R26268 vss.n2767 vss.n2766 0.0126193
R26269 vss.n2781 vss.n2780 0.0126193
R26270 vss.n2780 vss.n2779 0.0126193
R26271 vss.n2784 vss.n2752 0.0126193
R26272 vss.n2752 vss.n2742 0.0126193
R26273 vss.n14658 vss.n14657 0.0126193
R26274 vss.n14659 vss.n14658 0.0126193
R26275 vss.n1433 vss.n1427 0.0126193
R26276 vss.n1433 vss.n1431 0.0126193
R26277 vss.n7548 vss.n1437 0.0126193
R26278 vss.n7549 vss.n7548 0.0126193
R26279 vss.n7563 vss.n7562 0.0126193
R26280 vss.n7562 vss.n7561 0.0126193
R26281 vss.n7566 vss.n7534 0.0126193
R26282 vss.n7534 vss.n7524 0.0126193
R26283 vss.n14688 vss.n14687 0.0126193
R26284 vss.n14689 vss.n14688 0.0126193
R26285 vss.n1374 vss.n1321 0.0126193
R26286 vss.n1374 vss.n1325 0.0126193
R26287 vss.n1395 vss.n1378 0.0126193
R26288 vss.n1396 vss.n1395 0.0126193
R26289 vss.n14714 vss.n14713 0.0126193
R26290 vss.n14713 vss.n14712 0.0126193
R26291 vss.n14703 vss.n14702 0.0126193
R26292 vss.n14704 vss.n14703 0.0126193
R26293 vss.n14731 vss.n14730 0.0126193
R26294 vss.n14732 vss.n14731 0.0126193
R26295 vss.n2416 vss.n2364 0.0126193
R26296 vss.n2416 vss.n2368 0.0126193
R26297 vss.n8020 vss.n8019 0.0126193
R26298 vss.n8019 vss.n8018 0.0126193
R26299 vss.n8009 vss.n8008 0.0126193
R26300 vss.n8010 vss.n8009 0.0126193
R26301 vss.n2439 vss.n2438 0.0126193
R26302 vss.n2440 vss.n2439 0.0126193
R26303 vss.n8030 vss.n8029 0.0126193
R26304 vss.n8031 vss.n8030 0.0126193
R26305 vss.n1226 vss.n1220 0.0126193
R26306 vss.n1226 vss.n1224 0.0126193
R26307 vss.n3245 vss.n1230 0.0126193
R26308 vss.n3246 vss.n3245 0.0126193
R26309 vss.n3262 vss.n3261 0.0126193
R26310 vss.n3261 vss.n3260 0.0126193
R26311 vss.n3266 vss.n3265 0.0126193
R26312 vss.n3267 vss.n3266 0.0126193
R26313 vss.n14763 vss.n14762 0.0126193
R26314 vss.n14764 vss.n14763 0.0126193
R26315 vss.n4821 vss.n4820 0.0126193
R26316 vss.n4822 vss.n4821 0.0126193
R26317 vss.n4834 vss.n4833 0.0126193
R26318 vss.n4834 vss.n4814 0.0126193
R26319 vss.n4848 vss.n4847 0.0126193
R26320 vss.n4847 vss.n4846 0.0126193
R26321 vss.n4803 vss.n4749 0.0126193
R26322 vss.n4803 vss.n4801 0.0126193
R26323 vss.n4859 vss.n4858 0.0126193
R26324 vss.n4860 vss.n4859 0.0126193
R26325 vss.n4303 vss.n4302 0.0126193
R26326 vss.n4304 vss.n4303 0.0126193
R26327 vss.n4888 vss.n4887 0.0126193
R26328 vss.n4889 vss.n4888 0.0126193
R26329 vss.n4901 vss.n4900 0.0126193
R26330 vss.n4900 vss.n4899 0.0126193
R26331 vss.n4914 vss.n4913 0.0126193
R26332 vss.n4913 vss.n4284 0.0126193
R26333 vss.n4907 vss.n4906 0.0126193
R26334 vss.n4906 vss.n536 0.0126193
R26335 vss.n619 vss.n615 0.0126193
R26336 vss.n619 vss.n618 0.0126193
R26337 vss.n623 vss.n622 0.0126193
R26338 vss.n622 vss.n603 0.0126193
R26339 vss.n15402 vss.n15401 0.0126193
R26340 vss.n15401 vss.n15400 0.0126193
R26341 vss.n636 vss.n631 0.0126193
R26342 vss.n631 vss.n629 0.0126193
R26343 vss.n639 vss.n632 0.0126193
R26344 vss.n15387 vss.n632 0.0126193
R26345 vss.n5138 vss.n5137 0.0126193
R26346 vss.n5139 vss.n5138 0.0126193
R26347 vss.n5151 vss.n5150 0.0126193
R26348 vss.n5152 vss.n5151 0.0126193
R26349 vss.n5164 vss.n5163 0.0126193
R26350 vss.n5163 vss.n5162 0.0126193
R26351 vss.n5177 vss.n5176 0.0126193
R26352 vss.n5176 vss.n5117 0.0126193
R26353 vss.n5170 vss.n5169 0.0126193
R26354 vss.n5169 vss.n741 0.0126193
R26355 vss.n5350 vss.n5349 0.0126193
R26356 vss.n5351 vss.n5350 0.0126193
R26357 vss.n5363 vss.n5362 0.0126193
R26358 vss.n5364 vss.n5363 0.0126193
R26359 vss.n5376 vss.n5375 0.0126193
R26360 vss.n5375 vss.n5374 0.0126193
R26361 vss.n5389 vss.n5388 0.0126193
R26362 vss.n5388 vss.n5329 0.0126193
R26363 vss.n5382 vss.n5381 0.0126193
R26364 vss.n5381 vss.n794 0.0126193
R26365 vss.n876 vss.n872 0.0126193
R26366 vss.n876 vss.n875 0.0126193
R26367 vss.n880 vss.n879 0.0126193
R26368 vss.n879 vss.n860 0.0126193
R26369 vss.n15252 vss.n15251 0.0126193
R26370 vss.n15251 vss.n15250 0.0126193
R26371 vss.n893 vss.n888 0.0126193
R26372 vss.n888 vss.n886 0.0126193
R26373 vss.n896 vss.n889 0.0126193
R26374 vss.n15237 vss.n889 0.0126193
R26375 vss.n6422 vss.n6421 0.0126193
R26376 vss.n6423 vss.n6422 0.0126193
R26377 vss.n6435 vss.n6434 0.0126193
R26378 vss.n6436 vss.n6435 0.0126193
R26379 vss.n6448 vss.n6447 0.0126193
R26380 vss.n6447 vss.n6446 0.0126193
R26381 vss.n6461 vss.n6460 0.0126193
R26382 vss.n6460 vss.n6401 0.0126193
R26383 vss.n6454 vss.n6453 0.0126193
R26384 vss.n6453 vss.n1074 0.0126193
R26385 vss.n6537 vss.n6536 0.0126193
R26386 vss.n6538 vss.n6537 0.0126193
R26387 vss.n6550 vss.n6549 0.0126193
R26388 vss.n6551 vss.n6550 0.0126193
R26389 vss.n6563 vss.n6562 0.0126193
R26390 vss.n6562 vss.n6561 0.0126193
R26391 vss.n6577 vss.n6576 0.0126193
R26392 vss.n6576 vss.n6516 0.0126193
R26393 vss.n6569 vss.n6568 0.0126193
R26394 vss.n6571 vss.n6568 0.0126193
R26395 vss.n1086 vss.n1080 0.0126193
R26396 vss.n1086 vss.n1084 0.0126193
R26397 vss.n6539 vss.n1090 0.0126193
R26398 vss.n6540 vss.n6539 0.0126193
R26399 vss.n6554 vss.n6553 0.0126193
R26400 vss.n6553 vss.n6552 0.0126193
R26401 vss.n6557 vss.n6525 0.0126193
R26402 vss.n6525 vss.n6515 0.0126193
R26403 vss.n15032 vss.n15031 0.0126193
R26404 vss.n15033 vss.n15032 0.0126193
R26405 vss.n911 vss.n905 0.0126193
R26406 vss.n911 vss.n909 0.0126193
R26407 vss.n6424 vss.n915 0.0126193
R26408 vss.n6425 vss.n6424 0.0126193
R26409 vss.n6439 vss.n6438 0.0126193
R26410 vss.n6438 vss.n6437 0.0126193
R26411 vss.n6442 vss.n6410 0.0126193
R26412 vss.n6410 vss.n6400 0.0126193
R26413 vss.n15233 vss.n15232 0.0126193
R26414 vss.n15234 vss.n15233 0.0126193
R26415 vss.n852 vss.n800 0.0126193
R26416 vss.n852 vss.n804 0.0126193
R26417 vss.n873 vss.n856 0.0126193
R26418 vss.n874 vss.n873 0.0126193
R26419 vss.n15259 vss.n15258 0.0126193
R26420 vss.n15258 vss.n15257 0.0126193
R26421 vss.n15248 vss.n15247 0.0126193
R26422 vss.n15249 vss.n15248 0.0126193
R26423 vss.n15276 vss.n15275 0.0126193
R26424 vss.n15277 vss.n15276 0.0126193
R26425 vss.n753 vss.n747 0.0126193
R26426 vss.n753 vss.n751 0.0126193
R26427 vss.n5352 vss.n757 0.0126193
R26428 vss.n5353 vss.n5352 0.0126193
R26429 vss.n5367 vss.n5366 0.0126193
R26430 vss.n5366 vss.n5365 0.0126193
R26431 vss.n5370 vss.n5338 0.0126193
R26432 vss.n5338 vss.n5328 0.0126193
R26433 vss.n15353 vss.n15352 0.0126193
R26434 vss.n15354 vss.n15353 0.0126193
R26435 vss.n654 vss.n648 0.0126193
R26436 vss.n654 vss.n652 0.0126193
R26437 vss.n5140 vss.n658 0.0126193
R26438 vss.n5141 vss.n5140 0.0126193
R26439 vss.n5155 vss.n5154 0.0126193
R26440 vss.n5154 vss.n5153 0.0126193
R26441 vss.n5158 vss.n5126 0.0126193
R26442 vss.n5126 vss.n5116 0.0126193
R26443 vss.n15383 vss.n15382 0.0126193
R26444 vss.n15384 vss.n15383 0.0126193
R26445 vss.n595 vss.n542 0.0126193
R26446 vss.n595 vss.n546 0.0126193
R26447 vss.n616 vss.n599 0.0126193
R26448 vss.n617 vss.n616 0.0126193
R26449 vss.n15409 vss.n15408 0.0126193
R26450 vss.n15408 vss.n15407 0.0126193
R26451 vss.n15398 vss.n15397 0.0126193
R26452 vss.n15399 vss.n15398 0.0126193
R26453 vss.n15426 vss.n15425 0.0126193
R26454 vss.n15427 vss.n15426 0.0126193
R26455 vss.n4363 vss.n4362 0.0126193
R26456 vss.n4362 vss.n4313 0.0126193
R26457 vss.n4877 vss.n4876 0.0126193
R26458 vss.n4878 vss.n4877 0.0126193
R26459 vss.n4892 vss.n4891 0.0126193
R26460 vss.n4891 vss.n4890 0.0126193
R26461 vss.n4895 vss.n4293 0.0126193
R26462 vss.n4293 vss.n4283 0.0126193
R26463 vss.n4365 vss.n4364 0.0126193
R26464 vss.n4863 vss.n4365 0.0126193
R26465 vss.n447 vss.n441 0.0126193
R26466 vss.n447 vss.n445 0.0126193
R26467 vss.n4823 vss.n451 0.0126193
R26468 vss.n4824 vss.n4823 0.0126193
R26469 vss.n4840 vss.n4839 0.0126193
R26470 vss.n4839 vss.n4838 0.0126193
R26471 vss.n4844 vss.n4843 0.0126193
R26472 vss.n4845 vss.n4844 0.0126193
R26473 vss.n15458 vss.n15457 0.0126193
R26474 vss.n15459 vss.n15458 0.0126193
R26475 vss.n6265 vss.n6264 0.0126193
R26476 vss.n6264 vss.n6263 0.0126193
R26477 vss.n15888 vss.n15887 0.0126193
R26478 vss.n15889 vss.n15888 0.0126193
R26479 vss.n15882 vss.n24 0.0126193
R26480 vss.n15882 vss.n15881 0.0126193
R26481 vss.n15877 vss.n26 0.0126193
R26482 vss.n26 vss.n25 0.0126193
R26483 vss.n6269 vss.n6268 0.0126193
R26484 vss.n6270 vss.n6269 0.0126193
R26485 vss.n54 vss.n48 0.0126193
R26486 vss.n54 vss.n52 0.0126193
R26487 vss.n61 vss.n58 0.0126193
R26488 vss.n62 vss.n61 0.0126193
R26489 vss.n15836 vss.n15835 0.0126193
R26490 vss.n15835 vss.n63 0.0126193
R26491 vss.n66 vss.n65 0.0126193
R26492 vss.n15829 vss.n66 0.0126193
R26493 vss.n15853 vss.n15852 0.0126193
R26494 vss.n15854 vss.n15853 0.0126193
R26495 vss.n78 vss.n72 0.0126193
R26496 vss.n78 vss.n76 0.0126193
R26497 vss.n110 vss.n82 0.0126193
R26498 vss.n111 vss.n110 0.0126193
R26499 vss.n117 vss.n116 0.0126193
R26500 vss.n116 vss.n115 0.0126193
R26501 vss.n121 vss.n120 0.0126193
R26502 vss.n122 vss.n121 0.0126193
R26503 vss.n15826 vss.n15825 0.0126193
R26504 vss.n15827 vss.n15826 0.0126193
R26505 vss.n133 vss.n127 0.0126193
R26506 vss.n133 vss.n131 0.0126193
R26507 vss.n140 vss.n137 0.0126193
R26508 vss.n141 vss.n140 0.0126193
R26509 vss.n15780 vss.n15779 0.0126193
R26510 vss.n15779 vss.n142 0.0126193
R26511 vss.n145 vss.n144 0.0126193
R26512 vss.n15773 vss.n145 0.0126193
R26513 vss.n15797 vss.n15796 0.0126193
R26514 vss.n15798 vss.n15797 0.0126193
R26515 vss.n157 vss.n151 0.0126193
R26516 vss.n157 vss.n155 0.0126193
R26517 vss.n188 vss.n161 0.0126193
R26518 vss.n189 vss.n188 0.0126193
R26519 vss.n195 vss.n194 0.0126193
R26520 vss.n194 vss.n193 0.0126193
R26521 vss.n199 vss.n198 0.0126193
R26522 vss.n200 vss.n199 0.0126193
R26523 vss.n15770 vss.n15769 0.0126193
R26524 vss.n15771 vss.n15770 0.0126193
R26525 vss.n211 vss.n205 0.0126193
R26526 vss.n211 vss.n209 0.0126193
R26527 vss.n218 vss.n215 0.0126193
R26528 vss.n219 vss.n218 0.0126193
R26529 vss.n15724 vss.n15723 0.0126193
R26530 vss.n15723 vss.n220 0.0126193
R26531 vss.n223 vss.n222 0.0126193
R26532 vss.n15717 vss.n223 0.0126193
R26533 vss.n15741 vss.n15740 0.0126193
R26534 vss.n15742 vss.n15741 0.0126193
R26535 vss.n235 vss.n229 0.0126193
R26536 vss.n235 vss.n233 0.0126193
R26537 vss.n267 vss.n239 0.0126193
R26538 vss.n268 vss.n267 0.0126193
R26539 vss.n274 vss.n273 0.0126193
R26540 vss.n273 vss.n272 0.0126193
R26541 vss.n278 vss.n277 0.0126193
R26542 vss.n279 vss.n278 0.0126193
R26543 vss.n15714 vss.n15713 0.0126193
R26544 vss.n15715 vss.n15714 0.0126193
R26545 vss.n15681 vss.n15680 0.0126193
R26546 vss.n15680 vss.n15679 0.0126193
R26547 vss.n296 vss.n291 0.0126193
R26548 vss.n296 vss.n294 0.0126193
R26549 vss.n15667 vss.n15666 0.0126193
R26550 vss.n15666 vss.n295 0.0126193
R26551 vss.n301 vss.n300 0.0126193
R26552 vss.n15660 vss.n301 0.0126193
R26553 vss.n15685 vss.n15684 0.0126193
R26554 vss.n15686 vss.n15685 0.0126193
R26555 vss.n8367 vss.n8361 0.0126193
R26556 vss.n8367 vss.n8365 0.0126193
R26557 vss.n8392 vss.n8371 0.0126193
R26558 vss.n8393 vss.n8392 0.0126193
R26559 vss.n8380 vss.n8377 0.0126193
R26560 vss.n8381 vss.n8380 0.0126193
R26561 vss.n8379 vss.n8378 0.0126193
R26562 vss.n8383 vss.n8379 0.0126193
R26563 vss.n13683 vss.n13682 0.0126193
R26564 vss.n13684 vss.n13683 0.0126193
R26565 vss.n8331 vss.n8325 0.0126193
R26566 vss.n8331 vss.n8329 0.0126193
R26567 vss.n13394 vss.n8335 0.0126193
R26568 vss.n13395 vss.n13394 0.0126193
R26569 vss.n13385 vss.n13382 0.0126193
R26570 vss.n13386 vss.n13385 0.0126193
R26571 vss.n13412 vss.n13380 0.0126193
R26572 vss.n13380 vss.n13370 0.0126193
R26573 vss.n13713 vss.n13712 0.0126193
R26574 vss.n13714 vss.n13713 0.0126193
R26575 vss.n8497 vss.n8491 0.0126193
R26576 vss.n8497 vss.n8495 0.0126193
R26577 vss.n8588 vss.n8501 0.0126193
R26578 vss.n8589 vss.n8588 0.0126193
R26579 vss.n8510 vss.n8507 0.0126193
R26580 vss.n8511 vss.n8510 0.0126193
R26581 vss.n8509 vss.n8508 0.0126193
R26582 vss.n8513 vss.n8509 0.0126193
R26583 vss.n13302 vss.n13301 0.0126193
R26584 vss.n13303 vss.n13302 0.0126193
R26585 vss.n12941 vss.n9177 0.0126193
R26586 vss.n12941 vss.n9181 0.0126193
R26587 vss.n12961 vss.n12945 0.0126193
R26588 vss.n12962 vss.n12961 0.0126193
R26589 vss.n12954 vss.n12951 0.0126193
R26590 vss.n12955 vss.n12954 0.0126193
R26591 vss.n12953 vss.n12952 0.0126193
R26592 vss.n12953 vss.n8428 0.0126193
R26593 vss.n13001 vss.n13000 0.0126193
R26594 vss.n13002 vss.n13001 0.0126193
R26595 vss.n8911 vss.n8905 0.0126193
R26596 vss.n8911 vss.n8909 0.0126193
R26597 vss.n8936 vss.n8915 0.0126193
R26598 vss.n8937 vss.n8936 0.0126193
R26599 vss.n8924 vss.n8921 0.0126193
R26600 vss.n8925 vss.n8924 0.0126193
R26601 vss.n8923 vss.n8922 0.0126193
R26602 vss.n8927 vss.n8923 0.0126193
R26603 vss.n13160 vss.n13159 0.0126193
R26604 vss.n13161 vss.n13160 0.0126193
R26605 vss.n12695 vss.n12643 0.0126193
R26606 vss.n12695 vss.n12647 0.0126193
R26607 vss.n12815 vss.n12814 0.0126193
R26608 vss.n12814 vss.n12813 0.0126193
R26609 vss.n12804 vss.n12803 0.0126193
R26610 vss.n12805 vss.n12804 0.0126193
R26611 vss.n12718 vss.n12717 0.0126193
R26612 vss.n12719 vss.n12718 0.0126193
R26613 vss.n12825 vss.n12824 0.0126193
R26614 vss.n12826 vss.n12825 0.0126193
R26615 vss.n9359 vss.n9306 0.0126193
R26616 vss.n9359 vss.n9310 0.0126193
R26617 vss.n12892 vss.n12891 0.0126193
R26618 vss.n12891 vss.n12890 0.0126193
R26619 vss.n12881 vss.n12880 0.0126193
R26620 vss.n12882 vss.n12881 0.0126193
R26621 vss.n9382 vss.n9381 0.0126193
R26622 vss.n9383 vss.n9382 0.0126193
R26623 vss.n12902 vss.n12901 0.0126193
R26624 vss.n12903 vss.n12902 0.0126193
R26625 vss.n9368 vss.n9366 0.0126193
R26626 vss.n9366 vss.n9363 0.0126193
R26627 vss.n12885 vss.n12884 0.0126193
R26628 vss.n12884 vss.n12883 0.0126193
R26629 vss.n12872 vss.n12871 0.0126193
R26630 vss.n12873 vss.n12872 0.0126193
R26631 vss.n12835 vss.n12834 0.0126193
R26632 vss.n12834 vss.n9410 0.0126193
R26633 vss.n9416 vss.n9415 0.0126193
R26634 vss.n12829 vss.n9415 0.0126193
R26635 vss.n12704 vss.n12702 0.0126193
R26636 vss.n12702 vss.n12699 0.0126193
R26637 vss.n12808 vss.n12807 0.0126193
R26638 vss.n12807 vss.n12806 0.0126193
R26639 vss.n12795 vss.n12794 0.0126193
R26640 vss.n12796 vss.n12795 0.0126193
R26641 vss.n12786 vss.n12785 0.0126193
R26642 vss.n12785 vss.n12776 0.0126193
R26643 vss.n12779 vss.n12778 0.0126193
R26644 vss.n12779 vss.n8899 0.0126193
R26645 vss.n8939 vss.n8935 0.0126193
R26646 vss.n8939 vss.n8938 0.0126193
R26647 vss.n8946 vss.n8945 0.0126193
R26648 vss.n8946 vss.n8919 0.0126193
R26649 vss.n13137 vss.n13136 0.0126193
R26650 vss.n13138 vss.n13137 0.0126193
R26651 vss.n9166 vss.n9165 0.0126193
R26652 vss.n9165 vss.n9164 0.0126193
R26653 vss.n9170 vss.n9169 0.0126193
R26654 vss.n9171 vss.n9170 0.0126193
R26655 vss.n12965 vss.n12964 0.0126193
R26656 vss.n12964 vss.n12963 0.0126193
R26657 vss.n12972 vss.n12971 0.0126193
R26658 vss.n12971 vss.n12949 0.0126193
R26659 vss.n12978 vss.n12977 0.0126193
R26660 vss.n12979 vss.n12978 0.0126193
R26661 vss.n13312 vss.n13311 0.0126193
R26662 vss.n13311 vss.n8429 0.0126193
R26663 vss.n8438 vss.n8437 0.0126193
R26664 vss.n13306 vss.n8437 0.0126193
R26665 vss.n8591 vss.n8587 0.0126193
R26666 vss.n8591 vss.n8590 0.0126193
R26667 vss.n8598 vss.n8597 0.0126193
R26668 vss.n8598 vss.n8505 0.0126193
R26669 vss.n8604 vss.n8603 0.0126193
R26670 vss.n8605 vss.n8604 0.0126193
R26671 vss.n8576 vss.n8575 0.0126193
R26672 vss.n8575 vss.n8565 0.0126193
R26673 vss.n8573 vss.n8572 0.0126193
R26674 vss.n8572 vss.n8571 0.0126193
R26675 vss.n13397 vss.n13391 0.0126193
R26676 vss.n13397 vss.n13396 0.0126193
R26677 vss.n13404 vss.n13403 0.0126193
R26678 vss.n13405 vss.n13404 0.0126193
R26679 vss.n13418 vss.n13417 0.0126193
R26680 vss.n13417 vss.n13416 0.0126193
R26681 vss.n13431 vss.n13430 0.0126193
R26682 vss.n13430 vss.n13371 0.0126193
R26683 vss.n13424 vss.n13423 0.0126193
R26684 vss.n13423 vss.n8355 0.0126193
R26685 vss.n8395 vss.n8391 0.0126193
R26686 vss.n8395 vss.n8394 0.0126193
R26687 vss.n8402 vss.n8401 0.0126193
R26688 vss.n8402 vss.n8375 0.0126193
R26689 vss.n13660 vss.n13659 0.0126193
R26690 vss.n13661 vss.n13660 0.0126193
R26691 vss.n12068 vss.n12067 0.0126193
R26692 vss.n12067 vss.n12066 0.0126193
R26693 vss.n12072 vss.n12071 0.0126193
R26694 vss.n12073 vss.n12072 0.0126193
R26695 vss.n12093 vss.n11888 0.0126193
R26696 vss.n12093 vss.n12092 0.0126193
R26697 vss.n12099 vss.n12098 0.0126193
R26698 vss.n12099 vss.n11881 0.0126193
R26699 vss.n12119 vss.n12118 0.0126193
R26700 vss.n12118 vss.n12117 0.0126193
R26701 vss.n11869 vss.n11844 0.0126193
R26702 vss.n11869 vss.n11867 0.0126193
R26703 vss.n12130 vss.n12129 0.0126193
R26704 vss.n12131 vss.n12130 0.0126193
R26705 vss.n12104 vss.n11876 0.0126193
R26706 vss.n12104 vss.n12103 0.0126193
R26707 vss.n12090 vss.n12089 0.0126193
R26708 vss.n12091 vss.n12090 0.0126193
R26709 vss.n11941 vss.n11940 0.0126193
R26710 vss.n11940 vss.n11938 0.0126193
R26711 vss.n11943 vss.n11942 0.0126193
R26712 vss.n12076 vss.n11943 0.0126193
R26713 vss.n12115 vss.n12114 0.0126193
R26714 vss.n12116 vss.n12115 0.0126193
R26715 vss.n10393 vss.n10392 0.0126193
R26716 vss.n10394 vss.n10393 0.0126193
R26717 vss.n10252 vss.n10251 0.0126193
R26718 vss.n10251 vss.n10247 0.0126193
R26719 vss.n10248 vss.n10244 0.0126193
R26720 vss.n10249 vss.n10248 0.0126193
R26721 vss.n10242 vss.n10235 0.0126193
R26722 vss.n10242 vss.n10240 0.0126193
R26723 vss.n10634 vss.n10633 0.0126193
R26724 vss.n10635 vss.n10634 0.0126193
R26725 vss.n10783 vss.n10782 0.0126193
R26726 vss.n10784 vss.n10783 0.0126193
R26727 vss.n10646 vss.n10640 0.0126193
R26728 vss.n10646 vss.n10644 0.0126193
R26729 vss.n10651 vss.n10650 0.0126193
R26730 vss.n10650 vss.n10645 0.0126193
R26731 vss.n10705 vss.n10704 0.0126193
R26732 vss.n10704 vss.n10701 0.0126193
R26733 vss.n10766 vss.n10765 0.0126193
R26734 vss.n10765 vss.n10764 0.0126193
R26735 vss.n10761 vss.n10760 0.0126193
R26736 vss.n10762 vss.n10761 0.0126193
R26737 vss.n10165 vss.n10164 0.0126193
R26738 vss.n10164 vss.n10160 0.0126193
R26739 vss.n10161 vss.n10157 0.0126193
R26740 vss.n10162 vss.n10161 0.0126193
R26741 vss.n10155 vss.n10148 0.0126193
R26742 vss.n10155 vss.n10153 0.0126193
R26743 vss.n11027 vss.n11026 0.0126193
R26744 vss.n11028 vss.n11027 0.0126193
R26745 vss.n11035 vss.n11034 0.0126193
R26746 vss.n11036 vss.n11035 0.0126193
R26747 vss.n10077 vss.n10076 0.0126193
R26748 vss.n10076 vss.n10072 0.0126193
R26749 vss.n10073 vss.n10069 0.0126193
R26750 vss.n10074 vss.n10073 0.0126193
R26751 vss.n10067 vss.n10060 0.0126193
R26752 vss.n10067 vss.n10065 0.0126193
R26753 vss.n11321 vss.n11320 0.0126193
R26754 vss.n11322 vss.n11321 0.0126193
R26755 vss.n10054 vss.n10053 0.0126193
R26756 vss.n11324 vss.n10054 0.0126193
R26757 vss.n10052 vss.n10051 0.0126193
R26758 vss.n10051 vss.n10047 0.0126193
R26759 vss.n10048 vss.n10044 0.0126193
R26760 vss.n10049 vss.n10048 0.0126193
R26761 vss.n10042 vss.n9988 0.0126193
R26762 vss.n10042 vss.n10040 0.0126193
R26763 vss.n11347 vss.n11346 0.0126193
R26764 vss.n11348 vss.n11347 0.0126193
R26765 vss.n11440 vss.n11439 0.0126193
R26766 vss.n11441 vss.n11440 0.0126193
R26767 vss.n11358 vss.n11353 0.0126193
R26768 vss.n11358 vss.n11356 0.0126193
R26769 vss.n11363 vss.n11362 0.0126193
R26770 vss.n11362 vss.n11357 0.0126193
R26771 vss.n11417 vss.n11416 0.0126193
R26772 vss.n11416 vss.n11413 0.0126193
R26773 vss.n11423 vss.n11422 0.0126193
R26774 vss.n11422 vss.n9929 0.0126193
R26775 vss.n11677 vss.n11676 0.0126193
R26776 vss.n11678 vss.n11677 0.0126193
R26777 vss.n9940 vss.n9934 0.0126193
R26778 vss.n9940 vss.n9938 0.0126193
R26779 vss.n9945 vss.n9944 0.0126193
R26780 vss.n9944 vss.n9939 0.0126193
R26781 vss.n11654 vss.n11653 0.0126193
R26782 vss.n11653 vss.n11650 0.0126193
R26783 vss.n11660 vss.n11659 0.0126193
R26784 vss.n11659 vss.n8834 0.0126193
R26785 vss.n10330 vss.n10277 0.0126193
R26786 vss.n10330 vss.n10328 0.0126193
R26787 vss.n10336 vss.n10332 0.0126193
R26788 vss.n10337 vss.n10336 0.0126193
R26789 vss.n10340 vss.n10339 0.0126193
R26790 vss.n10339 vss.n10335 0.0126193
R26791 vss.n10342 vss.n10341 0.0126193
R26792 vss.n10362 vss.n10342 0.0126193
R26793 vss.n10385 vss.n10384 0.0126193
R26794 vss.n10386 vss.n10385 0.0126193
R26795 vss vss 0.00214474
R26796 vss vss 0.00214474
R26797 vss.n12381 vss.n12380 0.000501408
R26798 vss.n9630 vss.n9601 0.000501408
R26799 vss.n12263 vss.n12262 0.000501408
R26800 vss.n9760 vss.n9731 0.000501408
R26801 vss.n11757 vss.n11756 0.000501408
R26802 vss.n12192 vss.n9858 0.000501408
R26803 vss.n8764 vss.n8763 0.000501408
R26804 vss.n13700 vss.n13699 0.000501408
R26805 vss.n12310 vss.n12309 0.000501408
R26806 vss.n8645 vss.n8644 0.000501408
R26807 vss.n13289 vss.n13288 0.000501408
R26808 vss.n12429 vss.n12427 0.000501408
R26809 vss.n9215 vss.n9214 0.000501408
R26810 vss.n9317 vss.n9316 0.000501408
R26811 vss.n9501 vss.n9472 0.000501408
R26812 vss.n12500 vss.n12499 0.000501408
R26813 vss.n12503 vss.n12502 0.000501408
R26814 vss.n13177 vss.n13176 0.000501408
R26815 vss.n6612 vss.n6611 0.000501408
R26816 vss.n4948 vss.n4947 0.000501408
R26817 vss.n4996 vss.n4995 0.000501408
R26818 vss.n5045 vss.n5044 0.000501408
R26819 vss.n5046 vss.n4218 0.000501408
R26820 vss.n5095 vss.n4172 0.000501408
R26821 vss.n5211 vss.n5210 0.000501408
R26822 vss.n5470 vss.n5469 0.000501408
R26823 vss.n5519 vss.n5518 0.000501408
R26824 vss.n5521 vss.n5520 0.000501408
R26825 vss.n5307 vss.n5257 0.000501408
R26826 vss.n3386 vss.n3385 0.000501408
R26827 vss.n6375 vss.n6374 0.000501408
R26828 vss.n6376 vss.n3433 0.000501408
R26829 vss.n6379 vss.n3432 0.000501408
R26830 vss.n6660 vss.n6659 0.000501408
R26831 vss.n4446 vss.n4445 0.000501408
R26832 vss.n4493 vss.n4492 0.000501408
R26833 vss.n4543 vss.n4542 0.000501408
R26834 vss.n6739 vss.n6738 0.000501408
R26835 vss.n14935 vss.n14934 0.000501408
R26836 vss.n7348 vss.n3109 0.000501408
R26837 vss.n7351 vss.n7350 0.000501408
R26838 vss.n964 vss.n963 0.000501408
R26839 vss.n15220 vss.n15219 0.000501408
R26840 vss.n15172 vss.n15171 0.000501408
R26841 vss.n15100 vss.n965 0.000501408
R26842 vss.n15293 vss.n15292 0.000501408
R26843 vss.n15341 vss.n15340 0.000501408
R26844 vss.n15370 vss.n15369 0.000501408
R26845 vss.n7346 vss.n7345 0.000501408
R26846 vss.n553 vss.n552 0.000501408
R26847 vss.n499 vss.n498 0.000501408
R26848 vss.n4654 vss.n4652 0.000501408
R26849 vss.n4701 vss.n4700 0.000501408
R26850 vss.n4704 vss.n4703 0.000501408
R26851 vss.n15443 vss.n15442 0.000501408
R26852 vss.n1934 vss.n1933 0.000501408
R26853 vss.n6975 vss.n6974 0.000501408
R26854 vss.n7995 vss.n2450 0.000501408
R26855 vss.n7992 vss.n2451 0.000501408
R26856 vss.n7991 vss.n7990 0.000501408
R26857 vss.n7503 vss.n2975 0.000501408
R26858 vss.n7619 vss.n7618 0.000501408
R26859 vss.n7667 vss.n7666 0.000501408
R26860 vss.n7717 vss.n7716 0.000501408
R26861 vss.n7718 vss.n2929 0.000501408
R26862 vss.n7767 vss.n2882 0.000501408
R26863 vss.n7814 vss.n7813 0.000501408
R26864 vss.n7914 vss.n7913 0.000501408
R26865 vss.n7912 vss.n7911 0.000501408
R26866 vss.n7862 vss.n7861 0.000501408
R26867 vss.n14884 vss.n1140 0.000501408
R26868 vss.n7206 vss.n7205 0.000501408
R26869 vss.n7208 vss.n7207 0.000501408
R26870 vss.n6876 vss.n6875 0.000501408
R26871 vss.n6790 vss.n6789 0.000501408
R26872 vss.n14240 vss.n14239 0.000501408
R26873 vss.n13980 vss.n13979 0.000501408
R26874 vss.n8180 vss.n8151 0.000501408
R26875 vss.n1743 vss.n1742 0.000501408
R26876 vss.n14525 vss.n14524 0.000501408
R26877 vss.n14477 vss.n14476 0.000501408
R26878 vss.n14405 vss.n1744 0.000501408
R26879 vss.n14598 vss.n14597 0.000501408
R26880 vss.n14646 vss.n14645 0.000501408
R26881 vss.n14675 vss.n14674 0.000501408
R26882 vss.n14026 vss.n14025 0.000501408
R26883 vss.n1332 vss.n1331 0.000501408
R26884 vss.n1278 vss.n1277 0.000501408
R26885 vss.n8052 vss.n8051 0.000501408
R26886 vss.n8049 vss.n2276 0.000501408
R26887 vss.n8047 vss.n8046 0.000501408
R26888 vss.n14748 vss.n14747 0.000501408
R26889 vss.n14092 vss.n14091 0.000501408
R26890 vss.n14088 vss.n2145 0.000501408
R26891 vss.n14087 vss.n14086 0.000501408
R26892 vss.n12628 vss.n12627 0.000501408
R26893 vss.n12764 vss.n12763 0.000501408
R26894 vss.n13132 vss.n8996 0.000501408
R26895 vss.n13129 vss.n13128 0.000501408
R26896 vss.n13081 vss.n13080 0.000501408
R26897 vss.n13032 vss.n13031 0.000501408
R26898 vss.n13346 vss.n13345 0.000501408
R26899 vss.n8476 vss.n8254 0.000501408
R26900 vss.n13841 vss.n13840 0.000501408
R26901 vss.n13793 vss.n13792 0.000501408
R26902 vss.n13744 vss.n13743 0.000501408
R26903 vss.n13465 vss.n13464 0.000501408
R26904 vss.n13655 vss.n13511 0.000501408
R26905 vss.n13652 vss.n13651 0.000501408
R26906 vss.n13604 vss.n13603 0.000501408
R26907 vss.n14138 vss.n14137 0.000501408
R26908 vss.n14190 vss.n14189 0.000501408
R26909 vss.n14354 vss.n14353 0.000501408
R26910 vss.n14324 vss.n14323 0.000501408
R26911 vss.n14281 vss.n14280 0.000501408
R26912 vss.n15049 vss.n15048 0.000501408
R26913 vss.n15019 vss.n15018 0.000501408
R26914 vss.n14976 vss.n14975 0.000501408
R26915 vss.n15869 vss.n15868 0.000501408
R26916 vss.n6015 vss.n6014 0.000501408
R26917 vss.n6062 vss.n6061 0.000501408
R26918 vss.n6109 vss.n6108 0.000501408
R26919 vss.n3857 vss.n3856 0.000501408
R26920 vss.n15813 vss.n15812 0.000501408
R26921 vss.n5775 vss.n5774 0.000501408
R26922 vss.n5822 vss.n5821 0.000501408
R26923 vss.n5870 vss.n5868 0.000501408
R26924 vss.n3738 vss.n3737 0.000501408
R26925 vss.n15757 vss.n15756 0.000501408
R26926 vss.n5587 vss.n5586 0.000501408
R26927 vss.n5681 vss.n5680 0.000501408
R26928 vss.n5677 vss.n5676 0.000501408
R26929 vss.n3619 vss.n3618 0.000501408
R26930 vss.n15701 vss.n15700 0.000501408
R26931 vss.n15619 vss.n15618 0.000501408
R26932 vss.n15622 vss.n15621 0.000501408
R26933 vss.n3569 vss.n359 0.000501408
R26934 vss.n15575 vss.n15574 0.000501408
R26935 vss.n12138 vss.n8816 0.000501408
R26936 vss.n14804 vss.n14803 0.000501408
R26937 vss.n14806 vss.n14805 0.000501408
R26938 vss.n15499 vss.n15498 0.000501408
R26939 vss.n15501 vss.n15500 0.000501408
R26940 vss.n12140 vss.n12139 0.000501408
R26941 vss.n12188 vss.n12187 0.000501408
R26942 vss.n11801 vss.n11800 0.000501408
R26943 vss.n10470 vss.n10469 0.000501408
R26944 vss.n10518 vss.n10517 0.000501408
R26945 vss.n10567 vss.n10423 0.000501408
R26946 vss.n10615 vss.n10614 0.000501408
R26947 vss.n10814 vss.n10813 0.000501408
R26948 vss.n10864 vss.n10863 0.000501408
R26949 vss.n10912 vss.n10911 0.000501408
R26950 vss.n10961 vss.n10168 0.000501408
R26951 vss.n11009 vss.n11008 0.000501408
R26952 vss.n11302 vss.n11065 0.000501408
R26953 vss.n11299 vss.n11298 0.000501408
R26954 vss.n11251 vss.n11250 0.000501408
R26955 vss.n11202 vss.n11201 0.000501408
R26956 vss.n10028 vss.n10027 0.000501408
R26957 vss.n11613 vss.n11470 0.000501408
R26958 vss.n11610 vss.n11609 0.000501408
R26959 vss.n11562 vss.n11561 0.000501408
R26960 vss.n11708 vss.n11707 0.000501408
R26961 vss.n11637 vss.n11618 0.000501408
R26962 vss.n13185 vss.n13184 0.000501408
R26963 vss.n15904 vss.n15903 0.000501408
R26964 d0.n0 d0.t0 40.0866
R26965 d0.n314 d0.t2 40.0866
R26966 d0.n1 d0.t4 40.0866
R26967 d0.n310 d0.t6 40.0866
R26968 d0.n3 d0.t8 40.0866
R26969 d0.n306 d0.t10 40.0866
R26970 d0.n5 d0.t12 40.0866
R26971 d0.n302 d0.t14 40.0866
R26972 d0.n7 d0.t16 40.0866
R26973 d0.n298 d0.t18 40.0866
R26974 d0.n9 d0.t20 40.0866
R26975 d0.n294 d0.t22 40.0866
R26976 d0.n11 d0.t24 40.0866
R26977 d0.n290 d0.t26 40.0866
R26978 d0.n13 d0.t28 40.0866
R26979 d0.n286 d0.t30 40.0866
R26980 d0.n283 d0.t32 40.0866
R26981 d0.n281 d0.t34 40.0866
R26982 d0.n279 d0.t36 40.0866
R26983 d0.n277 d0.t38 40.0866
R26984 d0.n275 d0.t40 40.0866
R26985 d0.n273 d0.t42 40.0866
R26986 d0.n271 d0.t44 40.0866
R26987 d0.n269 d0.t46 40.0866
R26988 d0.n267 d0.t48 40.0866
R26989 d0.n265 d0.t50 40.0866
R26990 d0.n263 d0.t52 40.0866
R26991 d0.n261 d0.t54 40.0866
R26992 d0.n259 d0.t56 40.0866
R26993 d0.n257 d0.t58 40.0866
R26994 d0.n254 d0.t62 40.0866
R26995 d0.n255 d0.t60 40.0866
R26996 d0.n247 d0.t92 40.0866
R26997 d0.n241 d0.t88 40.0866
R26998 d0.n235 d0.t84 40.0866
R26999 d0.n229 d0.t80 40.0866
R27000 d0.n223 d0.t76 40.0866
R27001 d0.n217 d0.t72 40.0866
R27002 d0.n211 d0.t68 40.0866
R27003 d0.n206 d0.t64 40.0866
R27004 d0.n208 d0.t66 40.0866
R27005 d0.n214 d0.t70 40.0866
R27006 d0.n220 d0.t74 40.0866
R27007 d0.n226 d0.t78 40.0866
R27008 d0.n232 d0.t82 40.0866
R27009 d0.n238 d0.t86 40.0866
R27010 d0.n244 d0.t90 40.0866
R27011 d0.n250 d0.t94 40.0866
R27012 d0.n203 d0.t96 40.0866
R27013 d0.n201 d0.t98 40.0866
R27014 d0.n199 d0.t100 40.0866
R27015 d0.n197 d0.t102 40.0866
R27016 d0.n195 d0.t104 40.0866
R27017 d0.n193 d0.t106 40.0866
R27018 d0.n191 d0.t108 40.0866
R27019 d0.n189 d0.t110 40.0866
R27020 d0.n187 d0.t112 40.0866
R27021 d0.n185 d0.t114 40.0866
R27022 d0.n183 d0.t116 40.0866
R27023 d0.n181 d0.t118 40.0866
R27024 d0.n179 d0.t120 40.0866
R27025 d0.n177 d0.t122 40.0866
R27026 d0.n174 d0.t126 40.0866
R27027 d0.n175 d0.t124 40.0866
R27028 d0.n167 d0.t156 40.0866
R27029 d0.n161 d0.t152 40.0866
R27030 d0.n155 d0.t148 40.0866
R27031 d0.n149 d0.t144 40.0866
R27032 d0.n143 d0.t140 40.0866
R27033 d0.n137 d0.t136 40.0866
R27034 d0.n131 d0.t132 40.0866
R27035 d0.n126 d0.t128 40.0866
R27036 d0.n128 d0.t130 40.0866
R27037 d0.n134 d0.t134 40.0866
R27038 d0.n140 d0.t138 40.0866
R27039 d0.n146 d0.t142 40.0866
R27040 d0.n152 d0.t146 40.0866
R27041 d0.n158 d0.t150 40.0866
R27042 d0.n164 d0.t154 40.0866
R27043 d0.n170 d0.t158 40.0866
R27044 d0.n123 d0.t160 40.0866
R27045 d0.n121 d0.t162 40.0866
R27046 d0.n119 d0.t164 40.0866
R27047 d0.n117 d0.t166 40.0866
R27048 d0.n115 d0.t168 40.0866
R27049 d0.n113 d0.t170 40.0866
R27050 d0.n111 d0.t172 40.0866
R27051 d0.n109 d0.t174 40.0866
R27052 d0.n107 d0.t176 40.0866
R27053 d0.n105 d0.t178 40.0866
R27054 d0.n103 d0.t180 40.0866
R27055 d0.n101 d0.t182 40.0866
R27056 d0.n99 d0.t184 40.0866
R27057 d0.n97 d0.t186 40.0866
R27058 d0.n94 d0.t190 40.0866
R27059 d0.n95 d0.t188 40.0866
R27060 d0.n87 d0.t220 40.0866
R27061 d0.n81 d0.t216 40.0866
R27062 d0.n75 d0.t212 40.0866
R27063 d0.n69 d0.t208 40.0866
R27064 d0.n63 d0.t204 40.0866
R27065 d0.n57 d0.t200 40.0866
R27066 d0.n51 d0.t196 40.0866
R27067 d0.n46 d0.t192 40.0866
R27068 d0.n48 d0.t194 40.0866
R27069 d0.n54 d0.t198 40.0866
R27070 d0.n60 d0.t202 40.0866
R27071 d0.n66 d0.t206 40.0866
R27072 d0.n72 d0.t210 40.0866
R27073 d0.n78 d0.t214 40.0866
R27074 d0.n84 d0.t218 40.0866
R27075 d0.n90 d0.t222 40.0866
R27076 d0.n44 d0.t224 40.0866
R27077 d0.n42 d0.t226 40.0866
R27078 d0.n40 d0.t228 40.0866
R27079 d0.n38 d0.t230 40.0866
R27080 d0.n36 d0.t232 40.0866
R27081 d0.n34 d0.t234 40.0866
R27082 d0.n32 d0.t236 40.0866
R27083 d0.n30 d0.t238 40.0866
R27084 d0.n28 d0.t240 40.0866
R27085 d0.n26 d0.t242 40.0866
R27086 d0.n24 d0.t244 40.0866
R27087 d0.n22 d0.t246 40.0866
R27088 d0.n20 d0.t248 40.0866
R27089 d0.n18 d0.t250 40.0866
R27090 d0.n15 d0.t254 40.0866
R27091 d0.n16 d0.t252 40.0866
R27092 d0.n93 d0.n45 26.0319
R27093 d0.n288 d0.n285 25.885
R27094 d0.n314 d0.t3 23.8528
R27095 d0.n1 d0.t5 23.8528
R27096 d0.n310 d0.t7 23.8528
R27097 d0.n3 d0.t9 23.8528
R27098 d0.n306 d0.t11 23.8528
R27099 d0.n5 d0.t13 23.8528
R27100 d0.n302 d0.t15 23.8528
R27101 d0.n7 d0.t17 23.8528
R27102 d0.n298 d0.t19 23.8528
R27103 d0.n9 d0.t21 23.8528
R27104 d0.n294 d0.t23 23.8528
R27105 d0.n11 d0.t25 23.8528
R27106 d0.n290 d0.t27 23.8528
R27107 d0.n13 d0.t29 23.8528
R27108 d0.n286 d0.t31 23.8528
R27109 d0.n283 d0.t33 23.8528
R27110 d0.n281 d0.t35 23.8528
R27111 d0.n279 d0.t37 23.8528
R27112 d0.n277 d0.t39 23.8528
R27113 d0.n275 d0.t41 23.8528
R27114 d0.n273 d0.t43 23.8528
R27115 d0.n271 d0.t45 23.8528
R27116 d0.n269 d0.t47 23.8528
R27117 d0.n267 d0.t49 23.8528
R27118 d0.n265 d0.t51 23.8528
R27119 d0.n263 d0.t53 23.8528
R27120 d0.n261 d0.t55 23.8528
R27121 d0.n259 d0.t57 23.8528
R27122 d0.n257 d0.t59 23.8528
R27123 d0.n254 d0.t63 23.8528
R27124 d0.n255 d0.t61 23.8528
R27125 d0.n247 d0.t93 23.8528
R27126 d0.n241 d0.t89 23.8528
R27127 d0.n235 d0.t85 23.8528
R27128 d0.n229 d0.t81 23.8528
R27129 d0.n223 d0.t77 23.8528
R27130 d0.n217 d0.t73 23.8528
R27131 d0.n211 d0.t69 23.8528
R27132 d0.n206 d0.t65 23.8528
R27133 d0.n208 d0.t67 23.8528
R27134 d0.n214 d0.t71 23.8528
R27135 d0.n220 d0.t75 23.8528
R27136 d0.n226 d0.t79 23.8528
R27137 d0.n232 d0.t83 23.8528
R27138 d0.n238 d0.t87 23.8528
R27139 d0.n244 d0.t91 23.8528
R27140 d0.n250 d0.t95 23.8528
R27141 d0.n203 d0.t97 23.8528
R27142 d0.n201 d0.t99 23.8528
R27143 d0.n199 d0.t101 23.8528
R27144 d0.n197 d0.t103 23.8528
R27145 d0.n195 d0.t105 23.8528
R27146 d0.n193 d0.t107 23.8528
R27147 d0.n191 d0.t109 23.8528
R27148 d0.n189 d0.t111 23.8528
R27149 d0.n187 d0.t113 23.8528
R27150 d0.n185 d0.t115 23.8528
R27151 d0.n183 d0.t117 23.8528
R27152 d0.n181 d0.t119 23.8528
R27153 d0.n179 d0.t121 23.8528
R27154 d0.n177 d0.t123 23.8528
R27155 d0.n174 d0.t127 23.8528
R27156 d0.n175 d0.t125 23.8528
R27157 d0.n167 d0.t157 23.8528
R27158 d0.n161 d0.t153 23.8528
R27159 d0.n155 d0.t149 23.8528
R27160 d0.n149 d0.t145 23.8528
R27161 d0.n143 d0.t141 23.8528
R27162 d0.n137 d0.t137 23.8528
R27163 d0.n131 d0.t133 23.8528
R27164 d0.n126 d0.t129 23.8528
R27165 d0.n128 d0.t131 23.8528
R27166 d0.n134 d0.t135 23.8528
R27167 d0.n140 d0.t139 23.8528
R27168 d0.n146 d0.t143 23.8528
R27169 d0.n152 d0.t147 23.8528
R27170 d0.n158 d0.t151 23.8528
R27171 d0.n164 d0.t155 23.8528
R27172 d0.n170 d0.t159 23.8528
R27173 d0.n123 d0.t161 23.8528
R27174 d0.n121 d0.t163 23.8528
R27175 d0.n119 d0.t165 23.8528
R27176 d0.n117 d0.t167 23.8528
R27177 d0.n115 d0.t169 23.8528
R27178 d0.n113 d0.t171 23.8528
R27179 d0.n111 d0.t173 23.8528
R27180 d0.n109 d0.t175 23.8528
R27181 d0.n107 d0.t177 23.8528
R27182 d0.n105 d0.t179 23.8528
R27183 d0.n103 d0.t181 23.8528
R27184 d0.n101 d0.t183 23.8528
R27185 d0.n99 d0.t185 23.8528
R27186 d0.n97 d0.t187 23.8528
R27187 d0.n94 d0.t191 23.8528
R27188 d0.n95 d0.t189 23.8528
R27189 d0.n87 d0.t221 23.8528
R27190 d0.n81 d0.t217 23.8528
R27191 d0.n75 d0.t213 23.8528
R27192 d0.n69 d0.t209 23.8528
R27193 d0.n63 d0.t205 23.8528
R27194 d0.n57 d0.t201 23.8528
R27195 d0.n51 d0.t197 23.8528
R27196 d0.n46 d0.t193 23.8528
R27197 d0.n48 d0.t195 23.8528
R27198 d0.n54 d0.t199 23.8528
R27199 d0.n60 d0.t203 23.8528
R27200 d0.n66 d0.t207 23.8528
R27201 d0.n72 d0.t211 23.8528
R27202 d0.n78 d0.t215 23.8528
R27203 d0.n84 d0.t219 23.8528
R27204 d0.n90 d0.t223 23.8528
R27205 d0.n44 d0.t225 23.8528
R27206 d0.n42 d0.t227 23.8528
R27207 d0.n40 d0.t229 23.8528
R27208 d0.n38 d0.t231 23.8528
R27209 d0.n36 d0.t233 23.8528
R27210 d0.n34 d0.t235 23.8528
R27211 d0.n32 d0.t237 23.8528
R27212 d0.n30 d0.t239 23.8528
R27213 d0.n28 d0.t241 23.8528
R27214 d0.n26 d0.t243 23.8528
R27215 d0.n24 d0.t245 23.8528
R27216 d0.n22 d0.t247 23.8528
R27217 d0.n20 d0.t249 23.8528
R27218 d0.n18 d0.t251 23.8528
R27219 d0.n15 d0.t255 23.8528
R27220 d0.n16 d0.t253 23.8528
R27221 d0.n0 d0.t1 23.8528
R27222 d0.n173 d0.n125 20.6255
R27223 d0.n253 d0.n205 20.6255
R27224 d0.n258 d0.n256 7.54113
R27225 d0.n262 d0.n260 7.54113
R27226 d0.n266 d0.n264 7.54113
R27227 d0.n270 d0.n268 7.54113
R27228 d0.n274 d0.n272 7.54113
R27229 d0.n278 d0.n276 7.54113
R27230 d0.n282 d0.n280 7.54113
R27231 d0.n213 d0.n210 7.54113
R27232 d0.n219 d0.n216 7.54113
R27233 d0.n225 d0.n222 7.54113
R27234 d0.n231 d0.n228 7.54113
R27235 d0.n237 d0.n234 7.54113
R27236 d0.n243 d0.n240 7.54113
R27237 d0.n249 d0.n246 7.54113
R27238 d0.n178 d0.n176 7.54113
R27239 d0.n182 d0.n180 7.54113
R27240 d0.n186 d0.n184 7.54113
R27241 d0.n190 d0.n188 7.54113
R27242 d0.n194 d0.n192 7.54113
R27243 d0.n198 d0.n196 7.54113
R27244 d0.n202 d0.n200 7.54113
R27245 d0.n133 d0.n130 7.54113
R27246 d0.n139 d0.n136 7.54113
R27247 d0.n145 d0.n142 7.54113
R27248 d0.n151 d0.n148 7.54113
R27249 d0.n157 d0.n154 7.54113
R27250 d0.n163 d0.n160 7.54113
R27251 d0.n169 d0.n166 7.54113
R27252 d0.n98 d0.n96 7.54113
R27253 d0.n102 d0.n100 7.54113
R27254 d0.n106 d0.n104 7.54113
R27255 d0.n110 d0.n108 7.54113
R27256 d0.n114 d0.n112 7.54113
R27257 d0.n118 d0.n116 7.54113
R27258 d0.n122 d0.n120 7.54113
R27259 d0.n53 d0.n50 7.54113
R27260 d0.n59 d0.n56 7.54113
R27261 d0.n65 d0.n62 7.54113
R27262 d0.n71 d0.n68 7.54113
R27263 d0.n77 d0.n74 7.54113
R27264 d0.n83 d0.n80 7.54113
R27265 d0.n89 d0.n86 7.54113
R27266 d0.n19 d0.n17 7.54113
R27267 d0.n23 d0.n21 7.54113
R27268 d0.n27 d0.n25 7.54113
R27269 d0.n31 d0.n29 7.54113
R27270 d0.n35 d0.n33 7.54113
R27271 d0.n39 d0.n37 7.54113
R27272 d0.n43 d0.n41 7.54113
R27273 d0.n292 d0.n289 7.54113
R27274 d0.n296 d0.n293 7.54113
R27275 d0.n300 d0.n297 7.54113
R27276 d0.n304 d0.n301 7.54113
R27277 d0.n308 d0.n305 7.54113
R27278 d0.n312 d0.n309 7.54113
R27279 d0.n316 d0.n313 7.54113
R27280 d0.n285 d0.n284 5.40687
R27281 d0.n205 d0.n204 5.40687
R27282 d0.n125 d0.n124 5.40687
R27283 d0.n253 d0.n252 5.25999
R27284 d0.n173 d0.n172 5.25999
R27285 d0.n93 d0.n92 5.25999
R27286 d0.n256 d0 2.97874
R27287 d0.n176 d0 2.97874
R27288 d0.n96 d0 2.97874
R27289 d0.n17 d0 2.97874
R27290 d0.n210 d0.n207 2.91624
R27291 d0.n130 d0.n127 2.91624
R27292 d0.n50 d0.n47 2.91624
R27293 d0.n317 d0.n316 2.91624
R27294 d0.n260 d0.n258 2.91613
R27295 d0.n264 d0.n262 2.91613
R27296 d0.n268 d0.n266 2.91613
R27297 d0.n272 d0.n270 2.91613
R27298 d0.n276 d0.n274 2.91613
R27299 d0.n280 d0.n278 2.91613
R27300 d0.n284 d0.n282 2.91613
R27301 d0.n216 d0.n213 2.91613
R27302 d0.n222 d0.n219 2.91613
R27303 d0.n228 d0.n225 2.91613
R27304 d0.n234 d0.n231 2.91613
R27305 d0.n240 d0.n237 2.91613
R27306 d0.n246 d0.n243 2.91613
R27307 d0.n252 d0.n249 2.91613
R27308 d0.n180 d0.n178 2.91613
R27309 d0.n184 d0.n182 2.91613
R27310 d0.n188 d0.n186 2.91613
R27311 d0.n192 d0.n190 2.91613
R27312 d0.n196 d0.n194 2.91613
R27313 d0.n200 d0.n198 2.91613
R27314 d0.n204 d0.n202 2.91613
R27315 d0.n136 d0.n133 2.91613
R27316 d0.n142 d0.n139 2.91613
R27317 d0.n148 d0.n145 2.91613
R27318 d0.n154 d0.n151 2.91613
R27319 d0.n160 d0.n157 2.91613
R27320 d0.n166 d0.n163 2.91613
R27321 d0.n172 d0.n169 2.91613
R27322 d0.n100 d0.n98 2.91613
R27323 d0.n104 d0.n102 2.91613
R27324 d0.n108 d0.n106 2.91613
R27325 d0.n112 d0.n110 2.91613
R27326 d0.n116 d0.n114 2.91613
R27327 d0.n120 d0.n118 2.91613
R27328 d0.n124 d0.n122 2.91613
R27329 d0.n56 d0.n53 2.91613
R27330 d0.n62 d0.n59 2.91613
R27331 d0.n68 d0.n65 2.91613
R27332 d0.n74 d0.n71 2.91613
R27333 d0.n80 d0.n77 2.91613
R27334 d0.n86 d0.n83 2.91613
R27335 d0.n92 d0.n89 2.91613
R27336 d0.n21 d0.n19 2.91613
R27337 d0.n25 d0.n23 2.91613
R27338 d0.n29 d0.n27 2.91613
R27339 d0.n33 d0.n31 2.91613
R27340 d0.n37 d0.n35 2.91613
R27341 d0.n41 d0.n39 2.91613
R27342 d0.n45 d0.n43 2.91613
R27343 d0.n289 d0.n288 2.91613
R27344 d0.n293 d0.n292 2.91613
R27345 d0.n297 d0.n296 2.91613
R27346 d0.n301 d0.n300 2.91613
R27347 d0.n305 d0.n304 2.91613
R27348 d0.n309 d0.n308 2.91613
R27349 d0.n313 d0.n312 2.91613
R27350 d0.n125 d0.n93 2.2505
R27351 d0.n205 d0.n173 2.2505
R27352 d0.n285 d0.n253 2.2505
R27353 d0.n315 d0.n314 0.2505
R27354 d0.n2 d0.n1 0.2505
R27355 d0.n311 d0.n310 0.2505
R27356 d0.n4 d0.n3 0.2505
R27357 d0.n307 d0.n306 0.2505
R27358 d0.n6 d0.n5 0.2505
R27359 d0.n303 d0.n302 0.2505
R27360 d0.n8 d0.n7 0.2505
R27361 d0.n299 d0.n298 0.2505
R27362 d0.n10 d0.n9 0.2505
R27363 d0.n295 d0.n294 0.2505
R27364 d0.n12 d0.n11 0.2505
R27365 d0.n291 d0.n290 0.2505
R27366 d0.n14 d0.n13 0.2505
R27367 d0.n287 d0.n286 0.2505
R27368 d0 d0.n279 0.2505
R27369 d0 d0.n277 0.2505
R27370 d0 d0.n275 0.2505
R27371 d0 d0.n271 0.2505
R27372 d0 d0.n269 0.2505
R27373 d0 d0.n267 0.2505
R27374 d0 d0.n263 0.2505
R27375 d0 d0.n261 0.2505
R27376 d0 d0.n259 0.2505
R27377 d0 d0.n254 0.2505
R27378 d0 d0.n255 0.2505
R27379 d0.n248 d0.n247 0.2505
R27380 d0.n242 d0.n241 0.2505
R27381 d0.n236 d0.n235 0.2505
R27382 d0.n230 d0.n229 0.2505
R27383 d0.n224 d0.n223 0.2505
R27384 d0.n218 d0.n217 0.2505
R27385 d0.n212 d0.n211 0.2505
R27386 d0.n207 d0.n206 0.2505
R27387 d0.n209 d0.n208 0.2505
R27388 d0.n215 d0.n214 0.2505
R27389 d0.n221 d0.n220 0.2505
R27390 d0.n227 d0.n226 0.2505
R27391 d0.n233 d0.n232 0.2505
R27392 d0.n239 d0.n238 0.2505
R27393 d0.n245 d0.n244 0.2505
R27394 d0.n251 d0.n250 0.2505
R27395 d0 d0.n199 0.2505
R27396 d0 d0.n197 0.2505
R27397 d0 d0.n195 0.2505
R27398 d0 d0.n191 0.2505
R27399 d0 d0.n189 0.2505
R27400 d0 d0.n187 0.2505
R27401 d0 d0.n183 0.2505
R27402 d0 d0.n181 0.2505
R27403 d0 d0.n179 0.2505
R27404 d0 d0.n174 0.2505
R27405 d0 d0.n175 0.2505
R27406 d0.n168 d0.n167 0.2505
R27407 d0.n162 d0.n161 0.2505
R27408 d0.n156 d0.n155 0.2505
R27409 d0.n150 d0.n149 0.2505
R27410 d0.n144 d0.n143 0.2505
R27411 d0.n138 d0.n137 0.2505
R27412 d0.n132 d0.n131 0.2505
R27413 d0.n127 d0.n126 0.2505
R27414 d0.n129 d0.n128 0.2505
R27415 d0.n135 d0.n134 0.2505
R27416 d0.n141 d0.n140 0.2505
R27417 d0.n147 d0.n146 0.2505
R27418 d0.n153 d0.n152 0.2505
R27419 d0.n159 d0.n158 0.2505
R27420 d0.n165 d0.n164 0.2505
R27421 d0.n171 d0.n170 0.2505
R27422 d0 d0.n119 0.2505
R27423 d0 d0.n117 0.2505
R27424 d0 d0.n115 0.2505
R27425 d0 d0.n111 0.2505
R27426 d0 d0.n109 0.2505
R27427 d0 d0.n107 0.2505
R27428 d0 d0.n103 0.2505
R27429 d0 d0.n101 0.2505
R27430 d0 d0.n99 0.2505
R27431 d0 d0.n94 0.2505
R27432 d0 d0.n95 0.2505
R27433 d0.n88 d0.n87 0.2505
R27434 d0.n82 d0.n81 0.2505
R27435 d0.n76 d0.n75 0.2505
R27436 d0.n70 d0.n69 0.2505
R27437 d0.n64 d0.n63 0.2505
R27438 d0.n58 d0.n57 0.2505
R27439 d0.n52 d0.n51 0.2505
R27440 d0.n47 d0.n46 0.2505
R27441 d0.n49 d0.n48 0.2505
R27442 d0.n55 d0.n54 0.2505
R27443 d0.n61 d0.n60 0.2505
R27444 d0.n67 d0.n66 0.2505
R27445 d0.n73 d0.n72 0.2505
R27446 d0.n79 d0.n78 0.2505
R27447 d0.n85 d0.n84 0.2505
R27448 d0.n91 d0.n90 0.2505
R27449 d0 d0.n40 0.2505
R27450 d0 d0.n38 0.2505
R27451 d0 d0.n36 0.2505
R27452 d0 d0.n32 0.2505
R27453 d0 d0.n30 0.2505
R27454 d0 d0.n28 0.2505
R27455 d0 d0.n24 0.2505
R27456 d0 d0.n22 0.2505
R27457 d0 d0.n20 0.2505
R27458 d0 d0.n15 0.2505
R27459 d0 d0.n16 0.2505
R27460 d0.n317 d0.n0 0.2505
R27461 d0 d0.n283 0.188
R27462 d0 d0.n281 0.188
R27463 d0 d0.n273 0.188
R27464 d0 d0.n265 0.188
R27465 d0 d0.n257 0.188
R27466 d0 d0.n203 0.188
R27467 d0 d0.n201 0.188
R27468 d0 d0.n193 0.188
R27469 d0 d0.n185 0.188
R27470 d0 d0.n177 0.188
R27471 d0 d0.n123 0.188
R27472 d0 d0.n121 0.188
R27473 d0 d0.n113 0.188
R27474 d0 d0.n105 0.188
R27475 d0 d0.n97 0.188
R27476 d0 d0.n44 0.188
R27477 d0 d0.n42 0.188
R27478 d0 d0.n34 0.188
R27479 d0 d0.n26 0.188
R27480 d0 d0.n18 0.188
R27481 d0.n315 d0 0.063
R27482 d0.n2 d0 0.063
R27483 d0.n311 d0 0.063
R27484 d0.n4 d0 0.063
R27485 d0.n307 d0 0.063
R27486 d0.n6 d0 0.063
R27487 d0.n303 d0 0.063
R27488 d0.n8 d0 0.063
R27489 d0.n299 d0 0.063
R27490 d0.n10 d0 0.063
R27491 d0.n295 d0 0.063
R27492 d0.n12 d0 0.063
R27493 d0.n291 d0 0.063
R27494 d0.n14 d0 0.063
R27495 d0.n287 d0 0.063
R27496 d0 d0 0.063
R27497 d0 d0 0.063
R27498 d0 d0 0.063
R27499 d0 d0 0.063
R27500 d0 d0 0.063
R27501 d0.n248 d0 0.063
R27502 d0.n242 d0 0.063
R27503 d0.n236 d0 0.063
R27504 d0.n230 d0 0.063
R27505 d0.n224 d0 0.063
R27506 d0.n218 d0 0.063
R27507 d0.n212 d0 0.063
R27508 d0.n207 d0 0.063
R27509 d0.n209 d0 0.063
R27510 d0.n215 d0 0.063
R27511 d0.n221 d0 0.063
R27512 d0.n227 d0 0.063
R27513 d0.n233 d0 0.063
R27514 d0.n239 d0 0.063
R27515 d0.n245 d0 0.063
R27516 d0.n251 d0 0.063
R27517 d0 d0 0.063
R27518 d0 d0 0.063
R27519 d0 d0 0.063
R27520 d0 d0 0.063
R27521 d0 d0 0.063
R27522 d0.n168 d0 0.063
R27523 d0.n162 d0 0.063
R27524 d0.n156 d0 0.063
R27525 d0.n150 d0 0.063
R27526 d0.n144 d0 0.063
R27527 d0.n138 d0 0.063
R27528 d0.n132 d0 0.063
R27529 d0.n129 d0 0.063
R27530 d0.n135 d0 0.063
R27531 d0.n141 d0 0.063
R27532 d0.n147 d0 0.063
R27533 d0.n153 d0 0.063
R27534 d0.n159 d0 0.063
R27535 d0.n165 d0 0.063
R27536 d0.n171 d0 0.063
R27537 d0 d0 0.063
R27538 d0 d0 0.063
R27539 d0 d0 0.063
R27540 d0 d0 0.063
R27541 d0 d0 0.063
R27542 d0.n88 d0 0.063
R27543 d0.n82 d0 0.063
R27544 d0.n76 d0 0.063
R27545 d0.n70 d0 0.063
R27546 d0.n64 d0 0.063
R27547 d0.n58 d0 0.063
R27548 d0.n52 d0 0.063
R27549 d0.n47 d0 0.063
R27550 d0.n49 d0 0.063
R27551 d0.n55 d0 0.063
R27552 d0.n61 d0 0.063
R27553 d0.n67 d0 0.063
R27554 d0.n73 d0 0.063
R27555 d0.n79 d0 0.063
R27556 d0.n85 d0 0.063
R27557 d0.n91 d0 0.063
R27558 d0 d0 0.063
R27559 d0 d0 0.063
R27560 d0 d0 0.063
R27561 d0 d0 0.063
R27562 d0 d0 0.063
R27563 d0.n127 d0 0.03175
R27564 d0 d0 0.03175
R27565 d0 d0.n317 0.03175
R27566 d0 d0 0.03175
R27567 d0.n256 d0 0.000617139
R27568 d0.n258 d0 0.000617139
R27569 d0.n260 d0 0.000617139
R27570 d0.n262 d0 0.000617139
R27571 d0.n264 d0 0.000617139
R27572 d0.n266 d0 0.000617139
R27573 d0.n268 d0 0.000617139
R27574 d0.n270 d0 0.000617139
R27575 d0.n272 d0 0.000617139
R27576 d0.n274 d0 0.000617139
R27577 d0.n276 d0 0.000617139
R27578 d0.n278 d0 0.000617139
R27579 d0.n280 d0 0.000617139
R27580 d0.n282 d0 0.000617139
R27581 d0.n284 d0 0.000617139
R27582 d0.n210 d0.n209 0.000617139
R27583 d0.n213 d0.n212 0.000617139
R27584 d0.n216 d0.n215 0.000617139
R27585 d0.n219 d0.n218 0.000617139
R27586 d0.n222 d0.n221 0.000617139
R27587 d0.n225 d0.n224 0.000617139
R27588 d0.n228 d0.n227 0.000617139
R27589 d0.n231 d0.n230 0.000617139
R27590 d0.n234 d0.n233 0.000617139
R27591 d0.n237 d0.n236 0.000617139
R27592 d0.n240 d0.n239 0.000617139
R27593 d0.n243 d0.n242 0.000617139
R27594 d0.n246 d0.n245 0.000617139
R27595 d0.n249 d0.n248 0.000617139
R27596 d0.n252 d0.n251 0.000617139
R27597 d0.n176 d0 0.000617139
R27598 d0.n178 d0 0.000617139
R27599 d0.n180 d0 0.000617139
R27600 d0.n182 d0 0.000617139
R27601 d0.n184 d0 0.000617139
R27602 d0.n186 d0 0.000617139
R27603 d0.n188 d0 0.000617139
R27604 d0.n190 d0 0.000617139
R27605 d0.n192 d0 0.000617139
R27606 d0.n194 d0 0.000617139
R27607 d0.n196 d0 0.000617139
R27608 d0.n198 d0 0.000617139
R27609 d0.n200 d0 0.000617139
R27610 d0.n202 d0 0.000617139
R27611 d0.n204 d0 0.000617139
R27612 d0.n130 d0.n129 0.000617139
R27613 d0.n133 d0.n132 0.000617139
R27614 d0.n136 d0.n135 0.000617139
R27615 d0.n139 d0.n138 0.000617139
R27616 d0.n142 d0.n141 0.000617139
R27617 d0.n145 d0.n144 0.000617139
R27618 d0.n148 d0.n147 0.000617139
R27619 d0.n151 d0.n150 0.000617139
R27620 d0.n154 d0.n153 0.000617139
R27621 d0.n157 d0.n156 0.000617139
R27622 d0.n160 d0.n159 0.000617139
R27623 d0.n163 d0.n162 0.000617139
R27624 d0.n166 d0.n165 0.000617139
R27625 d0.n169 d0.n168 0.000617139
R27626 d0.n172 d0.n171 0.000617139
R27627 d0.n96 d0 0.000617139
R27628 d0.n98 d0 0.000617139
R27629 d0.n100 d0 0.000617139
R27630 d0.n102 d0 0.000617139
R27631 d0.n104 d0 0.000617139
R27632 d0.n106 d0 0.000617139
R27633 d0.n108 d0 0.000617139
R27634 d0.n110 d0 0.000617139
R27635 d0.n112 d0 0.000617139
R27636 d0.n114 d0 0.000617139
R27637 d0.n116 d0 0.000617139
R27638 d0.n118 d0 0.000617139
R27639 d0.n120 d0 0.000617139
R27640 d0.n122 d0 0.000617139
R27641 d0.n124 d0 0.000617139
R27642 d0.n50 d0.n49 0.000617139
R27643 d0.n53 d0.n52 0.000617139
R27644 d0.n56 d0.n55 0.000617139
R27645 d0.n59 d0.n58 0.000617139
R27646 d0.n62 d0.n61 0.000617139
R27647 d0.n65 d0.n64 0.000617139
R27648 d0.n68 d0.n67 0.000617139
R27649 d0.n71 d0.n70 0.000617139
R27650 d0.n74 d0.n73 0.000617139
R27651 d0.n77 d0.n76 0.000617139
R27652 d0.n80 d0.n79 0.000617139
R27653 d0.n83 d0.n82 0.000617139
R27654 d0.n86 d0.n85 0.000617139
R27655 d0.n89 d0.n88 0.000617139
R27656 d0.n92 d0.n91 0.000617139
R27657 d0.n17 d0 0.000617139
R27658 d0.n19 d0 0.000617139
R27659 d0.n21 d0 0.000617139
R27660 d0.n23 d0 0.000617139
R27661 d0.n25 d0 0.000617139
R27662 d0.n27 d0 0.000617139
R27663 d0.n29 d0 0.000617139
R27664 d0.n31 d0 0.000617139
R27665 d0.n33 d0 0.000617139
R27666 d0.n35 d0 0.000617139
R27667 d0.n37 d0 0.000617139
R27668 d0.n39 d0 0.000617139
R27669 d0.n41 d0 0.000617139
R27670 d0.n43 d0 0.000617139
R27671 d0.n45 d0 0.000617139
R27672 d0.n288 d0.n287 0.000617139
R27673 d0.n289 d0.n14 0.000617139
R27674 d0.n292 d0.n291 0.000617139
R27675 d0.n293 d0.n12 0.000617139
R27676 d0.n296 d0.n295 0.000617139
R27677 d0.n297 d0.n10 0.000617139
R27678 d0.n300 d0.n299 0.000617139
R27679 d0.n301 d0.n8 0.000617139
R27680 d0.n304 d0.n303 0.000617139
R27681 d0.n305 d0.n6 0.000617139
R27682 d0.n308 d0.n307 0.000617139
R27683 d0.n309 d0.n4 0.000617139
R27684 d0.n312 d0.n311 0.000617139
R27685 d0.n313 d0.n2 0.000617139
R27686 d0.n316 d0.n315 0.000617139
R27687 vdd.n135 vdd.n130 1560
R27688 vdd.n120 vdd.n111 1560
R27689 vdd.n183 vdd.n178 1560
R27690 vdd.n168 vdd.n159 1560
R27691 vdd.n284 vdd.n279 1560
R27692 vdd.n269 vdd.n260 1560
R27693 vdd.n332 vdd.n327 1560
R27694 vdd.n317 vdd.n308 1560
R27695 vdd.n380 vdd.n375 1560
R27696 vdd.n365 vdd.n356 1560
R27697 vdd.n428 vdd.n423 1560
R27698 vdd.n413 vdd.n404 1560
R27699 vdd.n529 vdd.n524 1560
R27700 vdd.n514 vdd.n505 1560
R27701 vdd.n577 vdd.n572 1560
R27702 vdd.n562 vdd.n553 1560
R27703 vdd.n6985 vdd.n6984 1560
R27704 vdd.n7002 vdd.n7000 1560
R27705 vdd.n7033 vdd.n7032 1560
R27706 vdd.n7050 vdd.n7048 1560
R27707 vdd.n7135 vdd.n7134 1560
R27708 vdd.n7152 vdd.n7150 1560
R27709 vdd.n7183 vdd.n7182 1560
R27710 vdd.n7200 vdd.n7198 1560
R27711 vdd.n7231 vdd.n7230 1560
R27712 vdd.n7248 vdd.n7246 1560
R27713 vdd.n7279 vdd.n7278 1560
R27714 vdd.n7296 vdd.n7294 1560
R27715 vdd.n7381 vdd.n7380 1560
R27716 vdd.n7398 vdd.n7396 1560
R27717 vdd.n8901 vdd.n8900 1560
R27718 vdd.n8918 vdd.n8916 1560
R27719 vdd.n7449 vdd.n7444 1560
R27720 vdd.n7434 vdd.n7425 1560
R27721 vdd.n7497 vdd.n7492 1560
R27722 vdd.n7482 vdd.n7473 1560
R27723 vdd.n7598 vdd.n7593 1560
R27724 vdd.n7583 vdd.n7574 1560
R27725 vdd.n7646 vdd.n7641 1560
R27726 vdd.n7631 vdd.n7622 1560
R27727 vdd.n7694 vdd.n7689 1560
R27728 vdd.n7679 vdd.n7670 1560
R27729 vdd.n7742 vdd.n7737 1560
R27730 vdd.n7727 vdd.n7718 1560
R27731 vdd.n7843 vdd.n7838 1560
R27732 vdd.n7828 vdd.n7819 1560
R27733 vdd.n6956 vdd.n6951 1560
R27734 vdd.n6941 vdd.n6932 1560
R27735 vdd.n7891 vdd.n7886 1560
R27736 vdd.n7876 vdd.n7867 1560
R27737 vdd.n7938 vdd.n7933 1560
R27738 vdd.n7923 vdd.n7914 1560
R27739 vdd.n7988 vdd.n7983 1560
R27740 vdd.n7973 vdd.n7964 1560
R27741 vdd.n8038 vdd.n8033 1560
R27742 vdd.n8023 vdd.n8014 1560
R27743 vdd.n8086 vdd.n8081 1560
R27744 vdd.n8071 vdd.n8062 1560
R27745 vdd.n7778 vdd.n7772 1560
R27746 vdd.n7799 vdd.n7756 1560
R27747 vdd.n8137 vdd.n8132 1560
R27748 vdd.n8122 vdd.n8113 1560
R27749 vdd.n8184 vdd.n8179 1560
R27750 vdd.n8169 vdd.n8160 1560
R27751 vdd.n8232 vdd.n8227 1560
R27752 vdd.n8217 vdd.n8208 1560
R27753 vdd.n8283 vdd.n8278 1560
R27754 vdd.n8268 vdd.n8259 1560
R27755 vdd.n8333 vdd.n8328 1560
R27756 vdd.n8318 vdd.n8309 1560
R27757 vdd.n8381 vdd.n8376 1560
R27758 vdd.n8366 vdd.n8357 1560
R27759 vdd.n8431 vdd.n8426 1560
R27760 vdd.n8416 vdd.n8407 1560
R27761 vdd.n8478 vdd.n8473 1560
R27762 vdd.n8463 vdd.n8454 1560
R27763 vdd.n8528 vdd.n8523 1560
R27764 vdd.n8513 vdd.n8504 1560
R27765 vdd.n8578 vdd.n8573 1560
R27766 vdd.n8563 vdd.n8554 1560
R27767 vdd.n8626 vdd.n8621 1560
R27768 vdd.n8611 vdd.n8602 1560
R27769 vdd.n7533 vdd.n7527 1560
R27770 vdd.n7554 vdd.n7511 1560
R27771 vdd.n8677 vdd.n8672 1560
R27772 vdd.n8662 vdd.n8653 1560
R27773 vdd.n8724 vdd.n8719 1560
R27774 vdd.n8709 vdd.n8700 1560
R27775 vdd.n8774 vdd.n8769 1560
R27776 vdd.n8759 vdd.n8750 1560
R27777 vdd.n8824 vdd.n8819 1560
R27778 vdd.n8809 vdd.n8800 1560
R27779 vdd.n8872 vdd.n8867 1560
R27780 vdd.n8857 vdd.n8848 1560
R27781 vdd.n8998 vdd.n8997 1560
R27782 vdd.n9015 vdd.n9013 1560
R27783 vdd.n8950 vdd.n8949 1560
R27784 vdd.n8967 vdd.n8965 1560
R27785 vdd.n9047 vdd.n9046 1560
R27786 vdd.n9064 vdd.n9062 1560
R27787 vdd.n9097 vdd.n9096 1560
R27788 vdd.n9114 vdd.n9112 1560
R27789 vdd.n9145 vdd.n9144 1560
R27790 vdd.n9162 vdd.n9160 1560
R27791 vdd.n7331 vdd.n7325 1560
R27792 vdd.n7352 vdd.n7312 1560
R27793 vdd.n9293 vdd.n9292 1560
R27794 vdd.n9310 vdd.n9308 1560
R27795 vdd.n9244 vdd.n9243 1560
R27796 vdd.n9261 vdd.n9259 1560
R27797 vdd.n9196 vdd.n9195 1560
R27798 vdd.n9213 vdd.n9211 1560
R27799 vdd.n9342 vdd.n9341 1560
R27800 vdd.n9359 vdd.n9357 1560
R27801 vdd.n9392 vdd.n9391 1560
R27802 vdd.n9409 vdd.n9407 1560
R27803 vdd.n9440 vdd.n9439 1560
R27804 vdd.n9457 vdd.n9455 1560
R27805 vdd.n9538 vdd.n9537 1560
R27806 vdd.n9555 vdd.n9553 1560
R27807 vdd.n9490 vdd.n9489 1560
R27808 vdd.n9507 vdd.n9505 1560
R27809 vdd.n9587 vdd.n9586 1560
R27810 vdd.n9604 vdd.n9602 1560
R27811 vdd.n9637 vdd.n9636 1560
R27812 vdd.n9654 vdd.n9652 1560
R27813 vdd.n9685 vdd.n9684 1560
R27814 vdd.n9702 vdd.n9700 1560
R27815 vdd.n7085 vdd.n7079 1560
R27816 vdd.n7106 vdd.n7066 1560
R27817 vdd.n9784 vdd.n9783 1560
R27818 vdd.n9801 vdd.n9799 1560
R27819 vdd.n9736 vdd.n9735 1560
R27820 vdd.n9753 vdd.n9751 1560
R27821 vdd.n9833 vdd.n9832 1560
R27822 vdd.n9850 vdd.n9848 1560
R27823 vdd.n9883 vdd.n9882 1560
R27824 vdd.n9900 vdd.n9898 1560
R27825 vdd.n9931 vdd.n9930 1560
R27826 vdd.n9948 vdd.n9946 1560
R27827 vdd.n3843 vdd.n3842 1560
R27828 vdd.n3860 vdd.n3858 1560
R27829 vdd.n3891 vdd.n3890 1560
R27830 vdd.n3908 vdd.n3906 1560
R27831 vdd.n3993 vdd.n3992 1560
R27832 vdd.n4010 vdd.n4008 1560
R27833 vdd.n4041 vdd.n4040 1560
R27834 vdd.n4058 vdd.n4056 1560
R27835 vdd.n4089 vdd.n4088 1560
R27836 vdd.n4106 vdd.n4104 1560
R27837 vdd.n4137 vdd.n4136 1560
R27838 vdd.n4154 vdd.n4152 1560
R27839 vdd.n4239 vdd.n4238 1560
R27840 vdd.n4256 vdd.n4254 1560
R27841 vdd.n5759 vdd.n5758 1560
R27842 vdd.n5776 vdd.n5774 1560
R27843 vdd.n4307 vdd.n4302 1560
R27844 vdd.n4292 vdd.n4283 1560
R27845 vdd.n4355 vdd.n4350 1560
R27846 vdd.n4340 vdd.n4331 1560
R27847 vdd.n4456 vdd.n4451 1560
R27848 vdd.n4441 vdd.n4432 1560
R27849 vdd.n4504 vdd.n4499 1560
R27850 vdd.n4489 vdd.n4480 1560
R27851 vdd.n4552 vdd.n4547 1560
R27852 vdd.n4537 vdd.n4528 1560
R27853 vdd.n4600 vdd.n4595 1560
R27854 vdd.n4585 vdd.n4576 1560
R27855 vdd.n4701 vdd.n4696 1560
R27856 vdd.n4686 vdd.n4677 1560
R27857 vdd.n3814 vdd.n3809 1560
R27858 vdd.n3799 vdd.n3790 1560
R27859 vdd.n4749 vdd.n4744 1560
R27860 vdd.n4734 vdd.n4725 1560
R27861 vdd.n4796 vdd.n4791 1560
R27862 vdd.n4781 vdd.n4772 1560
R27863 vdd.n4846 vdd.n4841 1560
R27864 vdd.n4831 vdd.n4822 1560
R27865 vdd.n4896 vdd.n4891 1560
R27866 vdd.n4881 vdd.n4872 1560
R27867 vdd.n4944 vdd.n4939 1560
R27868 vdd.n4929 vdd.n4920 1560
R27869 vdd.n4636 vdd.n4630 1560
R27870 vdd.n4657 vdd.n4614 1560
R27871 vdd.n4995 vdd.n4990 1560
R27872 vdd.n4980 vdd.n4971 1560
R27873 vdd.n5042 vdd.n5037 1560
R27874 vdd.n5027 vdd.n5018 1560
R27875 vdd.n5090 vdd.n5085 1560
R27876 vdd.n5075 vdd.n5066 1560
R27877 vdd.n5141 vdd.n5136 1560
R27878 vdd.n5126 vdd.n5117 1560
R27879 vdd.n5191 vdd.n5186 1560
R27880 vdd.n5176 vdd.n5167 1560
R27881 vdd.n5239 vdd.n5234 1560
R27882 vdd.n5224 vdd.n5215 1560
R27883 vdd.n5289 vdd.n5284 1560
R27884 vdd.n5274 vdd.n5265 1560
R27885 vdd.n5336 vdd.n5331 1560
R27886 vdd.n5321 vdd.n5312 1560
R27887 vdd.n5386 vdd.n5381 1560
R27888 vdd.n5371 vdd.n5362 1560
R27889 vdd.n5436 vdd.n5431 1560
R27890 vdd.n5421 vdd.n5412 1560
R27891 vdd.n5484 vdd.n5479 1560
R27892 vdd.n5469 vdd.n5460 1560
R27893 vdd.n4391 vdd.n4385 1560
R27894 vdd.n4412 vdd.n4369 1560
R27895 vdd.n5535 vdd.n5530 1560
R27896 vdd.n5520 vdd.n5511 1560
R27897 vdd.n5582 vdd.n5577 1560
R27898 vdd.n5567 vdd.n5558 1560
R27899 vdd.n5632 vdd.n5627 1560
R27900 vdd.n5617 vdd.n5608 1560
R27901 vdd.n5682 vdd.n5677 1560
R27902 vdd.n5667 vdd.n5658 1560
R27903 vdd.n5730 vdd.n5725 1560
R27904 vdd.n5715 vdd.n5706 1560
R27905 vdd.n5856 vdd.n5855 1560
R27906 vdd.n5873 vdd.n5871 1560
R27907 vdd.n5808 vdd.n5807 1560
R27908 vdd.n5825 vdd.n5823 1560
R27909 vdd.n5905 vdd.n5904 1560
R27910 vdd.n5922 vdd.n5920 1560
R27911 vdd.n5955 vdd.n5954 1560
R27912 vdd.n5972 vdd.n5970 1560
R27913 vdd.n6003 vdd.n6002 1560
R27914 vdd.n6020 vdd.n6018 1560
R27915 vdd.n4189 vdd.n4183 1560
R27916 vdd.n4210 vdd.n4170 1560
R27917 vdd.n6151 vdd.n6150 1560
R27918 vdd.n6168 vdd.n6166 1560
R27919 vdd.n6102 vdd.n6101 1560
R27920 vdd.n6119 vdd.n6117 1560
R27921 vdd.n6054 vdd.n6053 1560
R27922 vdd.n6071 vdd.n6069 1560
R27923 vdd.n6200 vdd.n6199 1560
R27924 vdd.n6217 vdd.n6215 1560
R27925 vdd.n6250 vdd.n6249 1560
R27926 vdd.n6267 vdd.n6265 1560
R27927 vdd.n6298 vdd.n6297 1560
R27928 vdd.n6315 vdd.n6313 1560
R27929 vdd.n6396 vdd.n6395 1560
R27930 vdd.n6413 vdd.n6411 1560
R27931 vdd.n6348 vdd.n6347 1560
R27932 vdd.n6365 vdd.n6363 1560
R27933 vdd.n6445 vdd.n6444 1560
R27934 vdd.n6462 vdd.n6460 1560
R27935 vdd.n6495 vdd.n6494 1560
R27936 vdd.n6512 vdd.n6510 1560
R27937 vdd.n6543 vdd.n6542 1560
R27938 vdd.n6560 vdd.n6558 1560
R27939 vdd.n3943 vdd.n3937 1560
R27940 vdd.n3964 vdd.n3924 1560
R27941 vdd.n6642 vdd.n6641 1560
R27942 vdd.n6659 vdd.n6657 1560
R27943 vdd.n6594 vdd.n6593 1560
R27944 vdd.n6611 vdd.n6609 1560
R27945 vdd.n6691 vdd.n6690 1560
R27946 vdd.n6708 vdd.n6706 1560
R27947 vdd.n6741 vdd.n6740 1560
R27948 vdd.n6758 vdd.n6756 1560
R27949 vdd.n6789 vdd.n6788 1560
R27950 vdd.n6806 vdd.n6804 1560
R27951 vdd.n701 vdd.n700 1560
R27952 vdd.n718 vdd.n716 1560
R27953 vdd.n749 vdd.n748 1560
R27954 vdd.n766 vdd.n764 1560
R27955 vdd.n851 vdd.n850 1560
R27956 vdd.n868 vdd.n866 1560
R27957 vdd.n899 vdd.n898 1560
R27958 vdd.n916 vdd.n914 1560
R27959 vdd.n947 vdd.n946 1560
R27960 vdd.n964 vdd.n962 1560
R27961 vdd.n995 vdd.n994 1560
R27962 vdd.n1012 vdd.n1010 1560
R27963 vdd.n1097 vdd.n1096 1560
R27964 vdd.n1114 vdd.n1112 1560
R27965 vdd.n2617 vdd.n2616 1560
R27966 vdd.n2634 vdd.n2632 1560
R27967 vdd.n1165 vdd.n1160 1560
R27968 vdd.n1150 vdd.n1141 1560
R27969 vdd.n1213 vdd.n1208 1560
R27970 vdd.n1198 vdd.n1189 1560
R27971 vdd.n1314 vdd.n1309 1560
R27972 vdd.n1299 vdd.n1290 1560
R27973 vdd.n1362 vdd.n1357 1560
R27974 vdd.n1347 vdd.n1338 1560
R27975 vdd.n1410 vdd.n1405 1560
R27976 vdd.n1395 vdd.n1386 1560
R27977 vdd.n1458 vdd.n1453 1560
R27978 vdd.n1443 vdd.n1434 1560
R27979 vdd.n1559 vdd.n1554 1560
R27980 vdd.n1544 vdd.n1535 1560
R27981 vdd.n672 vdd.n667 1560
R27982 vdd.n657 vdd.n648 1560
R27983 vdd.n1607 vdd.n1602 1560
R27984 vdd.n1592 vdd.n1583 1560
R27985 vdd.n1654 vdd.n1649 1560
R27986 vdd.n1639 vdd.n1630 1560
R27987 vdd.n1704 vdd.n1699 1560
R27988 vdd.n1689 vdd.n1680 1560
R27989 vdd.n1754 vdd.n1749 1560
R27990 vdd.n1739 vdd.n1730 1560
R27991 vdd.n1802 vdd.n1797 1560
R27992 vdd.n1787 vdd.n1778 1560
R27993 vdd.n1494 vdd.n1488 1560
R27994 vdd.n1515 vdd.n1472 1560
R27995 vdd.n1853 vdd.n1848 1560
R27996 vdd.n1838 vdd.n1829 1560
R27997 vdd.n1900 vdd.n1895 1560
R27998 vdd.n1885 vdd.n1876 1560
R27999 vdd.n1948 vdd.n1943 1560
R28000 vdd.n1933 vdd.n1924 1560
R28001 vdd.n1999 vdd.n1994 1560
R28002 vdd.n1984 vdd.n1975 1560
R28003 vdd.n2049 vdd.n2044 1560
R28004 vdd.n2034 vdd.n2025 1560
R28005 vdd.n2097 vdd.n2092 1560
R28006 vdd.n2082 vdd.n2073 1560
R28007 vdd.n2147 vdd.n2142 1560
R28008 vdd.n2132 vdd.n2123 1560
R28009 vdd.n2194 vdd.n2189 1560
R28010 vdd.n2179 vdd.n2170 1560
R28011 vdd.n2244 vdd.n2239 1560
R28012 vdd.n2229 vdd.n2220 1560
R28013 vdd.n2294 vdd.n2289 1560
R28014 vdd.n2279 vdd.n2270 1560
R28015 vdd.n2342 vdd.n2337 1560
R28016 vdd.n2327 vdd.n2318 1560
R28017 vdd.n1249 vdd.n1243 1560
R28018 vdd.n1270 vdd.n1227 1560
R28019 vdd.n2393 vdd.n2388 1560
R28020 vdd.n2378 vdd.n2369 1560
R28021 vdd.n2440 vdd.n2435 1560
R28022 vdd.n2425 vdd.n2416 1560
R28023 vdd.n2490 vdd.n2485 1560
R28024 vdd.n2475 vdd.n2466 1560
R28025 vdd.n2540 vdd.n2535 1560
R28026 vdd.n2525 vdd.n2516 1560
R28027 vdd.n2588 vdd.n2583 1560
R28028 vdd.n2573 vdd.n2564 1560
R28029 vdd.n2714 vdd.n2713 1560
R28030 vdd.n2731 vdd.n2729 1560
R28031 vdd.n2666 vdd.n2665 1560
R28032 vdd.n2683 vdd.n2681 1560
R28033 vdd.n2763 vdd.n2762 1560
R28034 vdd.n2780 vdd.n2778 1560
R28035 vdd.n2813 vdd.n2812 1560
R28036 vdd.n2830 vdd.n2828 1560
R28037 vdd.n2861 vdd.n2860 1560
R28038 vdd.n2878 vdd.n2876 1560
R28039 vdd.n1047 vdd.n1041 1560
R28040 vdd.n1068 vdd.n1028 1560
R28041 vdd.n3009 vdd.n3008 1560
R28042 vdd.n3026 vdd.n3024 1560
R28043 vdd.n2960 vdd.n2959 1560
R28044 vdd.n2977 vdd.n2975 1560
R28045 vdd.n2912 vdd.n2911 1560
R28046 vdd.n2929 vdd.n2927 1560
R28047 vdd.n3058 vdd.n3057 1560
R28048 vdd.n3075 vdd.n3073 1560
R28049 vdd.n3108 vdd.n3107 1560
R28050 vdd.n3125 vdd.n3123 1560
R28051 vdd.n3156 vdd.n3155 1560
R28052 vdd.n3173 vdd.n3171 1560
R28053 vdd.n3254 vdd.n3253 1560
R28054 vdd.n3271 vdd.n3269 1560
R28055 vdd.n3206 vdd.n3205 1560
R28056 vdd.n3223 vdd.n3221 1560
R28057 vdd.n3303 vdd.n3302 1560
R28058 vdd.n3320 vdd.n3318 1560
R28059 vdd.n3353 vdd.n3352 1560
R28060 vdd.n3370 vdd.n3368 1560
R28061 vdd.n3401 vdd.n3400 1560
R28062 vdd.n3418 vdd.n3416 1560
R28063 vdd.n801 vdd.n795 1560
R28064 vdd.n822 vdd.n782 1560
R28065 vdd.n3500 vdd.n3499 1560
R28066 vdd.n3517 vdd.n3515 1560
R28067 vdd.n3452 vdd.n3451 1560
R28068 vdd.n3469 vdd.n3467 1560
R28069 vdd.n3549 vdd.n3548 1560
R28070 vdd.n3566 vdd.n3564 1560
R28071 vdd.n3599 vdd.n3598 1560
R28072 vdd.n3616 vdd.n3614 1560
R28073 vdd.n3647 vdd.n3646 1560
R28074 vdd.n3664 vdd.n3662 1560
R28075 vdd.n605 vdd.n604 1560
R28076 vdd.n622 vdd.n620 1560
R28077 vdd.n3746 vdd.n3745 1560
R28078 vdd.n3763 vdd.n3761 1560
R28079 vdd.n3698 vdd.n3697 1560
R28080 vdd.n3715 vdd.n3713 1560
R28081 vdd.n6888 vdd.n6887 1560
R28082 vdd.n6905 vdd.n6903 1560
R28083 vdd.n6840 vdd.n6839 1560
R28084 vdd.n6857 vdd.n6855 1560
R28085 vdd.n10030 vdd.n10029 1560
R28086 vdd.n10047 vdd.n10045 1560
R28087 vdd.n9982 vdd.n9981 1560
R28088 vdd.n9999 vdd.n9997 1560
R28089 vdd.n10078 vdd.n10077 1560
R28090 vdd.n10095 vdd.n10093 1560
R28091 vdd.n10126 vdd.n10125 1560
R28092 vdd.n10143 vdd.n10141 1560
R28093 vdd.n10228 vdd.n10227 1560
R28094 vdd.n10245 vdd.n10243 1560
R28095 vdd.n10276 vdd.n10275 1560
R28096 vdd.n10293 vdd.n10291 1560
R28097 vdd.n10324 vdd.n10323 1560
R28098 vdd.n10341 vdd.n10339 1560
R28099 vdd.n10372 vdd.n10371 1560
R28100 vdd.n10389 vdd.n10387 1560
R28101 vdd.n10474 vdd.n10473 1560
R28102 vdd.n10491 vdd.n10489 1560
R28103 vdd.n66 vdd.n65 1560
R28104 vdd.n83 vdd.n81 1560
R28105 vdd.n18 vdd.n17 1560
R28106 vdd.n35 vdd.n33 1560
R28107 vdd.n10522 vdd.n10521 1560
R28108 vdd.n10539 vdd.n10537 1560
R28109 vdd.n10572 vdd.n10571 1560
R28110 vdd.n10589 vdd.n10587 1560
R28111 vdd.n10620 vdd.n10619 1560
R28112 vdd.n10637 vdd.n10635 1560
R28113 vdd.n10424 vdd.n10418 1560
R28114 vdd.n10445 vdd.n10405 1560
R28115 vdd.n10768 vdd.n10767 1560
R28116 vdd.n10785 vdd.n10783 1560
R28117 vdd.n10719 vdd.n10718 1560
R28118 vdd.n10736 vdd.n10734 1560
R28119 vdd.n10671 vdd.n10670 1560
R28120 vdd.n10688 vdd.n10686 1560
R28121 vdd.n10817 vdd.n10816 1560
R28122 vdd.n10834 vdd.n10832 1560
R28123 vdd.n10867 vdd.n10866 1560
R28124 vdd.n10884 vdd.n10882 1560
R28125 vdd.n10915 vdd.n10914 1560
R28126 vdd.n10932 vdd.n10930 1560
R28127 vdd.n11013 vdd.n11012 1560
R28128 vdd.n11030 vdd.n11028 1560
R28129 vdd.n10965 vdd.n10964 1560
R28130 vdd.n10982 vdd.n10980 1560
R28131 vdd.n11062 vdd.n11061 1560
R28132 vdd.n11079 vdd.n11077 1560
R28133 vdd.n11112 vdd.n11111 1560
R28134 vdd.n11129 vdd.n11127 1560
R28135 vdd.n11160 vdd.n11159 1560
R28136 vdd.n11177 vdd.n11175 1560
R28137 vdd.n10178 vdd.n10172 1560
R28138 vdd.n10199 vdd.n10159 1560
R28139 vdd.n11259 vdd.n11258 1560
R28140 vdd.n11276 vdd.n11274 1560
R28141 vdd.n11211 vdd.n11210 1560
R28142 vdd.n11228 vdd.n11226 1560
R28143 vdd.n11308 vdd.n11307 1560
R28144 vdd.n11325 vdd.n11323 1560
R28145 vdd.n11358 vdd.n11357 1560
R28146 vdd.n11375 vdd.n11373 1560
R28147 vdd.n11406 vdd.n11405 1560
R28148 vdd.n11423 vdd.n11421 1560
R28149 vdd.n11477 vdd.n11472 1560
R28150 vdd.n11462 vdd.n11453 1560
R28151 vdd.n11524 vdd.n11519 1560
R28152 vdd.n11509 vdd.n11500 1560
R28153 vdd.n11574 vdd.n11569 1560
R28154 vdd.n11559 vdd.n11550 1560
R28155 vdd.n11624 vdd.n11619 1560
R28156 vdd.n11609 vdd.n11600 1560
R28157 vdd.n11672 vdd.n11667 1560
R28158 vdd.n11657 vdd.n11648 1560
R28159 vdd.n464 vdd.n458 1560
R28160 vdd.n485 vdd.n442 1560
R28161 vdd.n11723 vdd.n11718 1560
R28162 vdd.n11708 vdd.n11699 1560
R28163 vdd.n11770 vdd.n11765 1560
R28164 vdd.n11755 vdd.n11746 1560
R28165 vdd.n11818 vdd.n11813 1560
R28166 vdd.n11803 vdd.n11794 1560
R28167 vdd.n11869 vdd.n11864 1560
R28168 vdd.n11854 vdd.n11845 1560
R28169 vdd.n11919 vdd.n11914 1560
R28170 vdd.n11904 vdd.n11895 1560
R28171 vdd.n11967 vdd.n11962 1560
R28172 vdd.n11952 vdd.n11943 1560
R28173 vdd.n12017 vdd.n12012 1560
R28174 vdd.n12002 vdd.n11993 1560
R28175 vdd.n12064 vdd.n12059 1560
R28176 vdd.n12049 vdd.n12040 1560
R28177 vdd.n12114 vdd.n12109 1560
R28178 vdd.n12099 vdd.n12090 1560
R28179 vdd.n12164 vdd.n12159 1560
R28180 vdd.n12149 vdd.n12140 1560
R28181 vdd.n12212 vdd.n12207 1560
R28182 vdd.n12197 vdd.n12188 1560
R28183 vdd.n219 vdd.n213 1560
R28184 vdd.n240 vdd.n197 1560
R28185 vdd.n12263 vdd.n12258 1560
R28186 vdd.n12248 vdd.n12239 1560
R28187 vdd.n12310 vdd.n12305 1560
R28188 vdd.n12295 vdd.n12286 1560
R28189 vdd.n12360 vdd.n12355 1560
R28190 vdd.n12345 vdd.n12336 1560
R28191 vdd.n12410 vdd.n12405 1560
R28192 vdd.n12395 vdd.n12386 1560
R28193 vdd.n12458 vdd.n12453 1560
R28194 vdd.n12443 vdd.n12434 1560
R28195 vdd.n127 vdd.n106 878.823
R28196 vdd.n127 vdd.n101 878.823
R28197 vdd.n105 vdd.n104 878.823
R28198 vdd.n104 vdd.n100 878.823
R28199 vdd.n110 vdd.n108 878.823
R28200 vdd.n121 vdd.n110 878.823
R28201 vdd.n175 vdd.n154 878.823
R28202 vdd.n175 vdd.n149 878.823
R28203 vdd.n153 vdd.n152 878.823
R28204 vdd.n152 vdd.n148 878.823
R28205 vdd.n158 vdd.n156 878.823
R28206 vdd.n169 vdd.n158 878.823
R28207 vdd.n276 vdd.n255 878.823
R28208 vdd.n276 vdd.n250 878.823
R28209 vdd.n254 vdd.n253 878.823
R28210 vdd.n253 vdd.n249 878.823
R28211 vdd.n259 vdd.n257 878.823
R28212 vdd.n270 vdd.n259 878.823
R28213 vdd.n324 vdd.n303 878.823
R28214 vdd.n324 vdd.n298 878.823
R28215 vdd.n302 vdd.n301 878.823
R28216 vdd.n301 vdd.n297 878.823
R28217 vdd.n307 vdd.n305 878.823
R28218 vdd.n318 vdd.n307 878.823
R28219 vdd.n372 vdd.n351 878.823
R28220 vdd.n372 vdd.n346 878.823
R28221 vdd.n350 vdd.n349 878.823
R28222 vdd.n349 vdd.n345 878.823
R28223 vdd.n355 vdd.n353 878.823
R28224 vdd.n366 vdd.n355 878.823
R28225 vdd.n420 vdd.n399 878.823
R28226 vdd.n420 vdd.n394 878.823
R28227 vdd.n398 vdd.n397 878.823
R28228 vdd.n397 vdd.n393 878.823
R28229 vdd.n403 vdd.n401 878.823
R28230 vdd.n414 vdd.n403 878.823
R28231 vdd.n521 vdd.n500 878.823
R28232 vdd.n521 vdd.n495 878.823
R28233 vdd.n499 vdd.n498 878.823
R28234 vdd.n498 vdd.n494 878.823
R28235 vdd.n504 vdd.n502 878.823
R28236 vdd.n515 vdd.n504 878.823
R28237 vdd.n569 vdd.n548 878.823
R28238 vdd.n569 vdd.n543 878.823
R28239 vdd.n547 vdd.n546 878.823
R28240 vdd.n546 vdd.n542 878.823
R28241 vdd.n552 vdd.n550 878.823
R28242 vdd.n563 vdd.n552 878.823
R28243 vdd.n6974 vdd.n6970 878.823
R28244 vdd.n6975 vdd.n6974 878.823
R28245 vdd.n6991 vdd.n6980 878.823
R28246 vdd.n6980 vdd.n6978 878.823
R28247 vdd.n6997 vdd.n6971 878.823
R28248 vdd.n6997 vdd.n6976 878.823
R28249 vdd.n7022 vdd.n7018 878.823
R28250 vdd.n7023 vdd.n7022 878.823
R28251 vdd.n7039 vdd.n7028 878.823
R28252 vdd.n7028 vdd.n7026 878.823
R28253 vdd.n7045 vdd.n7019 878.823
R28254 vdd.n7045 vdd.n7024 878.823
R28255 vdd.n7124 vdd.n7120 878.823
R28256 vdd.n7125 vdd.n7124 878.823
R28257 vdd.n7141 vdd.n7130 878.823
R28258 vdd.n7130 vdd.n7128 878.823
R28259 vdd.n7147 vdd.n7121 878.823
R28260 vdd.n7147 vdd.n7126 878.823
R28261 vdd.n7172 vdd.n7168 878.823
R28262 vdd.n7173 vdd.n7172 878.823
R28263 vdd.n7189 vdd.n7178 878.823
R28264 vdd.n7178 vdd.n7176 878.823
R28265 vdd.n7195 vdd.n7169 878.823
R28266 vdd.n7195 vdd.n7174 878.823
R28267 vdd.n7220 vdd.n7216 878.823
R28268 vdd.n7221 vdd.n7220 878.823
R28269 vdd.n7237 vdd.n7226 878.823
R28270 vdd.n7226 vdd.n7224 878.823
R28271 vdd.n7243 vdd.n7217 878.823
R28272 vdd.n7243 vdd.n7222 878.823
R28273 vdd.n7268 vdd.n7264 878.823
R28274 vdd.n7269 vdd.n7268 878.823
R28275 vdd.n7285 vdd.n7274 878.823
R28276 vdd.n7274 vdd.n7272 878.823
R28277 vdd.n7291 vdd.n7265 878.823
R28278 vdd.n7291 vdd.n7270 878.823
R28279 vdd.n7370 vdd.n7366 878.823
R28280 vdd.n7371 vdd.n7370 878.823
R28281 vdd.n7387 vdd.n7376 878.823
R28282 vdd.n7376 vdd.n7374 878.823
R28283 vdd.n7393 vdd.n7367 878.823
R28284 vdd.n7393 vdd.n7372 878.823
R28285 vdd.n8890 vdd.n8886 878.823
R28286 vdd.n8891 vdd.n8890 878.823
R28287 vdd.n8907 vdd.n8896 878.823
R28288 vdd.n8896 vdd.n8894 878.823
R28289 vdd.n8913 vdd.n8887 878.823
R28290 vdd.n8913 vdd.n8892 878.823
R28291 vdd.n7441 vdd.n7420 878.823
R28292 vdd.n7441 vdd.n7415 878.823
R28293 vdd.n7419 vdd.n7418 878.823
R28294 vdd.n7418 vdd.n7414 878.823
R28295 vdd.n7424 vdd.n7422 878.823
R28296 vdd.n7435 vdd.n7424 878.823
R28297 vdd.n7489 vdd.n7468 878.823
R28298 vdd.n7489 vdd.n7463 878.823
R28299 vdd.n7467 vdd.n7466 878.823
R28300 vdd.n7466 vdd.n7462 878.823
R28301 vdd.n7472 vdd.n7470 878.823
R28302 vdd.n7483 vdd.n7472 878.823
R28303 vdd.n7590 vdd.n7569 878.823
R28304 vdd.n7590 vdd.n7564 878.823
R28305 vdd.n7568 vdd.n7567 878.823
R28306 vdd.n7567 vdd.n7563 878.823
R28307 vdd.n7573 vdd.n7571 878.823
R28308 vdd.n7584 vdd.n7573 878.823
R28309 vdd.n7638 vdd.n7617 878.823
R28310 vdd.n7638 vdd.n7612 878.823
R28311 vdd.n7616 vdd.n7615 878.823
R28312 vdd.n7615 vdd.n7611 878.823
R28313 vdd.n7621 vdd.n7619 878.823
R28314 vdd.n7632 vdd.n7621 878.823
R28315 vdd.n7686 vdd.n7665 878.823
R28316 vdd.n7686 vdd.n7660 878.823
R28317 vdd.n7664 vdd.n7663 878.823
R28318 vdd.n7663 vdd.n7659 878.823
R28319 vdd.n7669 vdd.n7667 878.823
R28320 vdd.n7680 vdd.n7669 878.823
R28321 vdd.n7734 vdd.n7713 878.823
R28322 vdd.n7734 vdd.n7708 878.823
R28323 vdd.n7712 vdd.n7711 878.823
R28324 vdd.n7711 vdd.n7707 878.823
R28325 vdd.n7717 vdd.n7715 878.823
R28326 vdd.n7728 vdd.n7717 878.823
R28327 vdd.n7835 vdd.n7814 878.823
R28328 vdd.n7835 vdd.n7809 878.823
R28329 vdd.n7813 vdd.n7812 878.823
R28330 vdd.n7812 vdd.n7808 878.823
R28331 vdd.n7818 vdd.n7816 878.823
R28332 vdd.n7829 vdd.n7818 878.823
R28333 vdd.n6948 vdd.n6927 878.823
R28334 vdd.n6948 vdd.n6922 878.823
R28335 vdd.n6926 vdd.n6925 878.823
R28336 vdd.n6925 vdd.n6921 878.823
R28337 vdd.n6931 vdd.n6929 878.823
R28338 vdd.n6942 vdd.n6931 878.823
R28339 vdd.n7883 vdd.n7862 878.823
R28340 vdd.n7883 vdd.n7857 878.823
R28341 vdd.n7861 vdd.n7860 878.823
R28342 vdd.n7860 vdd.n7856 878.823
R28343 vdd.n7866 vdd.n7864 878.823
R28344 vdd.n7877 vdd.n7866 878.823
R28345 vdd.n7930 vdd.n7909 878.823
R28346 vdd.n7930 vdd.n7904 878.823
R28347 vdd.n7908 vdd.n7907 878.823
R28348 vdd.n7907 vdd.n7903 878.823
R28349 vdd.n7913 vdd.n7911 878.823
R28350 vdd.n7924 vdd.n7913 878.823
R28351 vdd.n7980 vdd.n7959 878.823
R28352 vdd.n7980 vdd.n7954 878.823
R28353 vdd.n7958 vdd.n7957 878.823
R28354 vdd.n7957 vdd.n7953 878.823
R28355 vdd.n7963 vdd.n7961 878.823
R28356 vdd.n7974 vdd.n7963 878.823
R28357 vdd.n8030 vdd.n8009 878.823
R28358 vdd.n8030 vdd.n8004 878.823
R28359 vdd.n8008 vdd.n8007 878.823
R28360 vdd.n8007 vdd.n8003 878.823
R28361 vdd.n8013 vdd.n8011 878.823
R28362 vdd.n8024 vdd.n8013 878.823
R28363 vdd.n8078 vdd.n8057 878.823
R28364 vdd.n8078 vdd.n8052 878.823
R28365 vdd.n8056 vdd.n8055 878.823
R28366 vdd.n8055 vdd.n8051 878.823
R28367 vdd.n8061 vdd.n8059 878.823
R28368 vdd.n8072 vdd.n8061 878.823
R28369 vdd.n7769 vdd.n7768 878.823
R28370 vdd.n7769 vdd.n7765 878.823
R28371 vdd.n7786 vdd.n7763 878.823
R28372 vdd.n7786 vdd.n7785 878.823
R28373 vdd.n7760 vdd.n7759 878.823
R28374 vdd.n7760 vdd.n7757 878.823
R28375 vdd.n8129 vdd.n8108 878.823
R28376 vdd.n8129 vdd.n8103 878.823
R28377 vdd.n8107 vdd.n8106 878.823
R28378 vdd.n8106 vdd.n8102 878.823
R28379 vdd.n8112 vdd.n8110 878.823
R28380 vdd.n8123 vdd.n8112 878.823
R28381 vdd.n8176 vdd.n8155 878.823
R28382 vdd.n8176 vdd.n8150 878.823
R28383 vdd.n8154 vdd.n8153 878.823
R28384 vdd.n8153 vdd.n8149 878.823
R28385 vdd.n8159 vdd.n8157 878.823
R28386 vdd.n8170 vdd.n8159 878.823
R28387 vdd.n8224 vdd.n8203 878.823
R28388 vdd.n8224 vdd.n8198 878.823
R28389 vdd.n8202 vdd.n8201 878.823
R28390 vdd.n8201 vdd.n8197 878.823
R28391 vdd.n8207 vdd.n8205 878.823
R28392 vdd.n8218 vdd.n8207 878.823
R28393 vdd.n8275 vdd.n8254 878.823
R28394 vdd.n8275 vdd.n8249 878.823
R28395 vdd.n8253 vdd.n8252 878.823
R28396 vdd.n8252 vdd.n8248 878.823
R28397 vdd.n8258 vdd.n8256 878.823
R28398 vdd.n8269 vdd.n8258 878.823
R28399 vdd.n8325 vdd.n8304 878.823
R28400 vdd.n8325 vdd.n8299 878.823
R28401 vdd.n8303 vdd.n8302 878.823
R28402 vdd.n8302 vdd.n8298 878.823
R28403 vdd.n8308 vdd.n8306 878.823
R28404 vdd.n8319 vdd.n8308 878.823
R28405 vdd.n8373 vdd.n8352 878.823
R28406 vdd.n8373 vdd.n8347 878.823
R28407 vdd.n8351 vdd.n8350 878.823
R28408 vdd.n8350 vdd.n8346 878.823
R28409 vdd.n8356 vdd.n8354 878.823
R28410 vdd.n8367 vdd.n8356 878.823
R28411 vdd.n8423 vdd.n8402 878.823
R28412 vdd.n8423 vdd.n8397 878.823
R28413 vdd.n8401 vdd.n8400 878.823
R28414 vdd.n8400 vdd.n8396 878.823
R28415 vdd.n8406 vdd.n8404 878.823
R28416 vdd.n8417 vdd.n8406 878.823
R28417 vdd.n8470 vdd.n8449 878.823
R28418 vdd.n8470 vdd.n8444 878.823
R28419 vdd.n8448 vdd.n8447 878.823
R28420 vdd.n8447 vdd.n8443 878.823
R28421 vdd.n8453 vdd.n8451 878.823
R28422 vdd.n8464 vdd.n8453 878.823
R28423 vdd.n8520 vdd.n8499 878.823
R28424 vdd.n8520 vdd.n8494 878.823
R28425 vdd.n8498 vdd.n8497 878.823
R28426 vdd.n8497 vdd.n8493 878.823
R28427 vdd.n8503 vdd.n8501 878.823
R28428 vdd.n8514 vdd.n8503 878.823
R28429 vdd.n8570 vdd.n8549 878.823
R28430 vdd.n8570 vdd.n8544 878.823
R28431 vdd.n8548 vdd.n8547 878.823
R28432 vdd.n8547 vdd.n8543 878.823
R28433 vdd.n8553 vdd.n8551 878.823
R28434 vdd.n8564 vdd.n8553 878.823
R28435 vdd.n8618 vdd.n8597 878.823
R28436 vdd.n8618 vdd.n8592 878.823
R28437 vdd.n8596 vdd.n8595 878.823
R28438 vdd.n8595 vdd.n8591 878.823
R28439 vdd.n8601 vdd.n8599 878.823
R28440 vdd.n8612 vdd.n8601 878.823
R28441 vdd.n7524 vdd.n7523 878.823
R28442 vdd.n7524 vdd.n7520 878.823
R28443 vdd.n7541 vdd.n7518 878.823
R28444 vdd.n7541 vdd.n7540 878.823
R28445 vdd.n7515 vdd.n7514 878.823
R28446 vdd.n7515 vdd.n7512 878.823
R28447 vdd.n8669 vdd.n8648 878.823
R28448 vdd.n8669 vdd.n8643 878.823
R28449 vdd.n8647 vdd.n8646 878.823
R28450 vdd.n8646 vdd.n8642 878.823
R28451 vdd.n8652 vdd.n8650 878.823
R28452 vdd.n8663 vdd.n8652 878.823
R28453 vdd.n8716 vdd.n8695 878.823
R28454 vdd.n8716 vdd.n8690 878.823
R28455 vdd.n8694 vdd.n8693 878.823
R28456 vdd.n8693 vdd.n8689 878.823
R28457 vdd.n8699 vdd.n8697 878.823
R28458 vdd.n8710 vdd.n8699 878.823
R28459 vdd.n8766 vdd.n8745 878.823
R28460 vdd.n8766 vdd.n8740 878.823
R28461 vdd.n8744 vdd.n8743 878.823
R28462 vdd.n8743 vdd.n8739 878.823
R28463 vdd.n8749 vdd.n8747 878.823
R28464 vdd.n8760 vdd.n8749 878.823
R28465 vdd.n8816 vdd.n8795 878.823
R28466 vdd.n8816 vdd.n8790 878.823
R28467 vdd.n8794 vdd.n8793 878.823
R28468 vdd.n8793 vdd.n8789 878.823
R28469 vdd.n8799 vdd.n8797 878.823
R28470 vdd.n8810 vdd.n8799 878.823
R28471 vdd.n8864 vdd.n8843 878.823
R28472 vdd.n8864 vdd.n8838 878.823
R28473 vdd.n8842 vdd.n8841 878.823
R28474 vdd.n8841 vdd.n8837 878.823
R28475 vdd.n8847 vdd.n8845 878.823
R28476 vdd.n8858 vdd.n8847 878.823
R28477 vdd.n8987 vdd.n8983 878.823
R28478 vdd.n8988 vdd.n8987 878.823
R28479 vdd.n9004 vdd.n8993 878.823
R28480 vdd.n8993 vdd.n8991 878.823
R28481 vdd.n9010 vdd.n8984 878.823
R28482 vdd.n9010 vdd.n8989 878.823
R28483 vdd.n8939 vdd.n8935 878.823
R28484 vdd.n8940 vdd.n8939 878.823
R28485 vdd.n8956 vdd.n8945 878.823
R28486 vdd.n8945 vdd.n8943 878.823
R28487 vdd.n8962 vdd.n8936 878.823
R28488 vdd.n8962 vdd.n8941 878.823
R28489 vdd.n9036 vdd.n9032 878.823
R28490 vdd.n9037 vdd.n9036 878.823
R28491 vdd.n9053 vdd.n9042 878.823
R28492 vdd.n9042 vdd.n9040 878.823
R28493 vdd.n9059 vdd.n9033 878.823
R28494 vdd.n9059 vdd.n9038 878.823
R28495 vdd.n9086 vdd.n9082 878.823
R28496 vdd.n9087 vdd.n9086 878.823
R28497 vdd.n9103 vdd.n9092 878.823
R28498 vdd.n9092 vdd.n9090 878.823
R28499 vdd.n9109 vdd.n9083 878.823
R28500 vdd.n9109 vdd.n9088 878.823
R28501 vdd.n9134 vdd.n9130 878.823
R28502 vdd.n9135 vdd.n9134 878.823
R28503 vdd.n9151 vdd.n9140 878.823
R28504 vdd.n9140 vdd.n9138 878.823
R28505 vdd.n9157 vdd.n9131 878.823
R28506 vdd.n9157 vdd.n9136 878.823
R28507 vdd.n7344 vdd.n7318 878.823
R28508 vdd.n7344 vdd.n7319 878.823
R28509 vdd.n7326 vdd.n7322 878.823
R28510 vdd.n7327 vdd.n7326 878.823
R28511 vdd.n7351 vdd.n7350 878.823
R28512 vdd.n7350 vdd.n7314 878.823
R28513 vdd.n9282 vdd.n9278 878.823
R28514 vdd.n9283 vdd.n9282 878.823
R28515 vdd.n9299 vdd.n9288 878.823
R28516 vdd.n9288 vdd.n9286 878.823
R28517 vdd.n9305 vdd.n9279 878.823
R28518 vdd.n9305 vdd.n9284 878.823
R28519 vdd.n9233 vdd.n9229 878.823
R28520 vdd.n9234 vdd.n9233 878.823
R28521 vdd.n9250 vdd.n9239 878.823
R28522 vdd.n9239 vdd.n9237 878.823
R28523 vdd.n9256 vdd.n9230 878.823
R28524 vdd.n9256 vdd.n9235 878.823
R28525 vdd.n9185 vdd.n9181 878.823
R28526 vdd.n9186 vdd.n9185 878.823
R28527 vdd.n9202 vdd.n9191 878.823
R28528 vdd.n9191 vdd.n9189 878.823
R28529 vdd.n9208 vdd.n9182 878.823
R28530 vdd.n9208 vdd.n9187 878.823
R28531 vdd.n9331 vdd.n9327 878.823
R28532 vdd.n9332 vdd.n9331 878.823
R28533 vdd.n9348 vdd.n9337 878.823
R28534 vdd.n9337 vdd.n9335 878.823
R28535 vdd.n9354 vdd.n9328 878.823
R28536 vdd.n9354 vdd.n9333 878.823
R28537 vdd.n9381 vdd.n9377 878.823
R28538 vdd.n9382 vdd.n9381 878.823
R28539 vdd.n9398 vdd.n9387 878.823
R28540 vdd.n9387 vdd.n9385 878.823
R28541 vdd.n9404 vdd.n9378 878.823
R28542 vdd.n9404 vdd.n9383 878.823
R28543 vdd.n9429 vdd.n9425 878.823
R28544 vdd.n9430 vdd.n9429 878.823
R28545 vdd.n9446 vdd.n9435 878.823
R28546 vdd.n9435 vdd.n9433 878.823
R28547 vdd.n9452 vdd.n9426 878.823
R28548 vdd.n9452 vdd.n9431 878.823
R28549 vdd.n9527 vdd.n9523 878.823
R28550 vdd.n9528 vdd.n9527 878.823
R28551 vdd.n9544 vdd.n9533 878.823
R28552 vdd.n9533 vdd.n9531 878.823
R28553 vdd.n9550 vdd.n9524 878.823
R28554 vdd.n9550 vdd.n9529 878.823
R28555 vdd.n9479 vdd.n9475 878.823
R28556 vdd.n9480 vdd.n9479 878.823
R28557 vdd.n9496 vdd.n9485 878.823
R28558 vdd.n9485 vdd.n9483 878.823
R28559 vdd.n9502 vdd.n9476 878.823
R28560 vdd.n9502 vdd.n9481 878.823
R28561 vdd.n9576 vdd.n9572 878.823
R28562 vdd.n9577 vdd.n9576 878.823
R28563 vdd.n9593 vdd.n9582 878.823
R28564 vdd.n9582 vdd.n9580 878.823
R28565 vdd.n9599 vdd.n9573 878.823
R28566 vdd.n9599 vdd.n9578 878.823
R28567 vdd.n9626 vdd.n9622 878.823
R28568 vdd.n9627 vdd.n9626 878.823
R28569 vdd.n9643 vdd.n9632 878.823
R28570 vdd.n9632 vdd.n9630 878.823
R28571 vdd.n9649 vdd.n9623 878.823
R28572 vdd.n9649 vdd.n9628 878.823
R28573 vdd.n9674 vdd.n9670 878.823
R28574 vdd.n9675 vdd.n9674 878.823
R28575 vdd.n9691 vdd.n9680 878.823
R28576 vdd.n9680 vdd.n9678 878.823
R28577 vdd.n9697 vdd.n9671 878.823
R28578 vdd.n9697 vdd.n9676 878.823
R28579 vdd.n7098 vdd.n7072 878.823
R28580 vdd.n7098 vdd.n7073 878.823
R28581 vdd.n7080 vdd.n7076 878.823
R28582 vdd.n7081 vdd.n7080 878.823
R28583 vdd.n7105 vdd.n7104 878.823
R28584 vdd.n7104 vdd.n7068 878.823
R28585 vdd.n9773 vdd.n9769 878.823
R28586 vdd.n9774 vdd.n9773 878.823
R28587 vdd.n9790 vdd.n9779 878.823
R28588 vdd.n9779 vdd.n9777 878.823
R28589 vdd.n9796 vdd.n9770 878.823
R28590 vdd.n9796 vdd.n9775 878.823
R28591 vdd.n9725 vdd.n9721 878.823
R28592 vdd.n9726 vdd.n9725 878.823
R28593 vdd.n9742 vdd.n9731 878.823
R28594 vdd.n9731 vdd.n9729 878.823
R28595 vdd.n9748 vdd.n9722 878.823
R28596 vdd.n9748 vdd.n9727 878.823
R28597 vdd.n9822 vdd.n9818 878.823
R28598 vdd.n9823 vdd.n9822 878.823
R28599 vdd.n9839 vdd.n9828 878.823
R28600 vdd.n9828 vdd.n9826 878.823
R28601 vdd.n9845 vdd.n9819 878.823
R28602 vdd.n9845 vdd.n9824 878.823
R28603 vdd.n9872 vdd.n9868 878.823
R28604 vdd.n9873 vdd.n9872 878.823
R28605 vdd.n9889 vdd.n9878 878.823
R28606 vdd.n9878 vdd.n9876 878.823
R28607 vdd.n9895 vdd.n9869 878.823
R28608 vdd.n9895 vdd.n9874 878.823
R28609 vdd.n9920 vdd.n9916 878.823
R28610 vdd.n9921 vdd.n9920 878.823
R28611 vdd.n9937 vdd.n9926 878.823
R28612 vdd.n9926 vdd.n9924 878.823
R28613 vdd.n9943 vdd.n9917 878.823
R28614 vdd.n9943 vdd.n9922 878.823
R28615 vdd.n3832 vdd.n3828 878.823
R28616 vdd.n3833 vdd.n3832 878.823
R28617 vdd.n3849 vdd.n3838 878.823
R28618 vdd.n3838 vdd.n3836 878.823
R28619 vdd.n3855 vdd.n3829 878.823
R28620 vdd.n3855 vdd.n3834 878.823
R28621 vdd.n3880 vdd.n3876 878.823
R28622 vdd.n3881 vdd.n3880 878.823
R28623 vdd.n3897 vdd.n3886 878.823
R28624 vdd.n3886 vdd.n3884 878.823
R28625 vdd.n3903 vdd.n3877 878.823
R28626 vdd.n3903 vdd.n3882 878.823
R28627 vdd.n3982 vdd.n3978 878.823
R28628 vdd.n3983 vdd.n3982 878.823
R28629 vdd.n3999 vdd.n3988 878.823
R28630 vdd.n3988 vdd.n3986 878.823
R28631 vdd.n4005 vdd.n3979 878.823
R28632 vdd.n4005 vdd.n3984 878.823
R28633 vdd.n4030 vdd.n4026 878.823
R28634 vdd.n4031 vdd.n4030 878.823
R28635 vdd.n4047 vdd.n4036 878.823
R28636 vdd.n4036 vdd.n4034 878.823
R28637 vdd.n4053 vdd.n4027 878.823
R28638 vdd.n4053 vdd.n4032 878.823
R28639 vdd.n4078 vdd.n4074 878.823
R28640 vdd.n4079 vdd.n4078 878.823
R28641 vdd.n4095 vdd.n4084 878.823
R28642 vdd.n4084 vdd.n4082 878.823
R28643 vdd.n4101 vdd.n4075 878.823
R28644 vdd.n4101 vdd.n4080 878.823
R28645 vdd.n4126 vdd.n4122 878.823
R28646 vdd.n4127 vdd.n4126 878.823
R28647 vdd.n4143 vdd.n4132 878.823
R28648 vdd.n4132 vdd.n4130 878.823
R28649 vdd.n4149 vdd.n4123 878.823
R28650 vdd.n4149 vdd.n4128 878.823
R28651 vdd.n4228 vdd.n4224 878.823
R28652 vdd.n4229 vdd.n4228 878.823
R28653 vdd.n4245 vdd.n4234 878.823
R28654 vdd.n4234 vdd.n4232 878.823
R28655 vdd.n4251 vdd.n4225 878.823
R28656 vdd.n4251 vdd.n4230 878.823
R28657 vdd.n5748 vdd.n5744 878.823
R28658 vdd.n5749 vdd.n5748 878.823
R28659 vdd.n5765 vdd.n5754 878.823
R28660 vdd.n5754 vdd.n5752 878.823
R28661 vdd.n5771 vdd.n5745 878.823
R28662 vdd.n5771 vdd.n5750 878.823
R28663 vdd.n4299 vdd.n4278 878.823
R28664 vdd.n4299 vdd.n4273 878.823
R28665 vdd.n4277 vdd.n4276 878.823
R28666 vdd.n4276 vdd.n4272 878.823
R28667 vdd.n4282 vdd.n4280 878.823
R28668 vdd.n4293 vdd.n4282 878.823
R28669 vdd.n4347 vdd.n4326 878.823
R28670 vdd.n4347 vdd.n4321 878.823
R28671 vdd.n4325 vdd.n4324 878.823
R28672 vdd.n4324 vdd.n4320 878.823
R28673 vdd.n4330 vdd.n4328 878.823
R28674 vdd.n4341 vdd.n4330 878.823
R28675 vdd.n4448 vdd.n4427 878.823
R28676 vdd.n4448 vdd.n4422 878.823
R28677 vdd.n4426 vdd.n4425 878.823
R28678 vdd.n4425 vdd.n4421 878.823
R28679 vdd.n4431 vdd.n4429 878.823
R28680 vdd.n4442 vdd.n4431 878.823
R28681 vdd.n4496 vdd.n4475 878.823
R28682 vdd.n4496 vdd.n4470 878.823
R28683 vdd.n4474 vdd.n4473 878.823
R28684 vdd.n4473 vdd.n4469 878.823
R28685 vdd.n4479 vdd.n4477 878.823
R28686 vdd.n4490 vdd.n4479 878.823
R28687 vdd.n4544 vdd.n4523 878.823
R28688 vdd.n4544 vdd.n4518 878.823
R28689 vdd.n4522 vdd.n4521 878.823
R28690 vdd.n4521 vdd.n4517 878.823
R28691 vdd.n4527 vdd.n4525 878.823
R28692 vdd.n4538 vdd.n4527 878.823
R28693 vdd.n4592 vdd.n4571 878.823
R28694 vdd.n4592 vdd.n4566 878.823
R28695 vdd.n4570 vdd.n4569 878.823
R28696 vdd.n4569 vdd.n4565 878.823
R28697 vdd.n4575 vdd.n4573 878.823
R28698 vdd.n4586 vdd.n4575 878.823
R28699 vdd.n4693 vdd.n4672 878.823
R28700 vdd.n4693 vdd.n4667 878.823
R28701 vdd.n4671 vdd.n4670 878.823
R28702 vdd.n4670 vdd.n4666 878.823
R28703 vdd.n4676 vdd.n4674 878.823
R28704 vdd.n4687 vdd.n4676 878.823
R28705 vdd.n3806 vdd.n3785 878.823
R28706 vdd.n3806 vdd.n3780 878.823
R28707 vdd.n3784 vdd.n3783 878.823
R28708 vdd.n3783 vdd.n3779 878.823
R28709 vdd.n3789 vdd.n3787 878.823
R28710 vdd.n3800 vdd.n3789 878.823
R28711 vdd.n4741 vdd.n4720 878.823
R28712 vdd.n4741 vdd.n4715 878.823
R28713 vdd.n4719 vdd.n4718 878.823
R28714 vdd.n4718 vdd.n4714 878.823
R28715 vdd.n4724 vdd.n4722 878.823
R28716 vdd.n4735 vdd.n4724 878.823
R28717 vdd.n4788 vdd.n4767 878.823
R28718 vdd.n4788 vdd.n4762 878.823
R28719 vdd.n4766 vdd.n4765 878.823
R28720 vdd.n4765 vdd.n4761 878.823
R28721 vdd.n4771 vdd.n4769 878.823
R28722 vdd.n4782 vdd.n4771 878.823
R28723 vdd.n4838 vdd.n4817 878.823
R28724 vdd.n4838 vdd.n4812 878.823
R28725 vdd.n4816 vdd.n4815 878.823
R28726 vdd.n4815 vdd.n4811 878.823
R28727 vdd.n4821 vdd.n4819 878.823
R28728 vdd.n4832 vdd.n4821 878.823
R28729 vdd.n4888 vdd.n4867 878.823
R28730 vdd.n4888 vdd.n4862 878.823
R28731 vdd.n4866 vdd.n4865 878.823
R28732 vdd.n4865 vdd.n4861 878.823
R28733 vdd.n4871 vdd.n4869 878.823
R28734 vdd.n4882 vdd.n4871 878.823
R28735 vdd.n4936 vdd.n4915 878.823
R28736 vdd.n4936 vdd.n4910 878.823
R28737 vdd.n4914 vdd.n4913 878.823
R28738 vdd.n4913 vdd.n4909 878.823
R28739 vdd.n4919 vdd.n4917 878.823
R28740 vdd.n4930 vdd.n4919 878.823
R28741 vdd.n4627 vdd.n4626 878.823
R28742 vdd.n4627 vdd.n4623 878.823
R28743 vdd.n4644 vdd.n4621 878.823
R28744 vdd.n4644 vdd.n4643 878.823
R28745 vdd.n4618 vdd.n4617 878.823
R28746 vdd.n4618 vdd.n4615 878.823
R28747 vdd.n4987 vdd.n4966 878.823
R28748 vdd.n4987 vdd.n4961 878.823
R28749 vdd.n4965 vdd.n4964 878.823
R28750 vdd.n4964 vdd.n4960 878.823
R28751 vdd.n4970 vdd.n4968 878.823
R28752 vdd.n4981 vdd.n4970 878.823
R28753 vdd.n5034 vdd.n5013 878.823
R28754 vdd.n5034 vdd.n5008 878.823
R28755 vdd.n5012 vdd.n5011 878.823
R28756 vdd.n5011 vdd.n5007 878.823
R28757 vdd.n5017 vdd.n5015 878.823
R28758 vdd.n5028 vdd.n5017 878.823
R28759 vdd.n5082 vdd.n5061 878.823
R28760 vdd.n5082 vdd.n5056 878.823
R28761 vdd.n5060 vdd.n5059 878.823
R28762 vdd.n5059 vdd.n5055 878.823
R28763 vdd.n5065 vdd.n5063 878.823
R28764 vdd.n5076 vdd.n5065 878.823
R28765 vdd.n5133 vdd.n5112 878.823
R28766 vdd.n5133 vdd.n5107 878.823
R28767 vdd.n5111 vdd.n5110 878.823
R28768 vdd.n5110 vdd.n5106 878.823
R28769 vdd.n5116 vdd.n5114 878.823
R28770 vdd.n5127 vdd.n5116 878.823
R28771 vdd.n5183 vdd.n5162 878.823
R28772 vdd.n5183 vdd.n5157 878.823
R28773 vdd.n5161 vdd.n5160 878.823
R28774 vdd.n5160 vdd.n5156 878.823
R28775 vdd.n5166 vdd.n5164 878.823
R28776 vdd.n5177 vdd.n5166 878.823
R28777 vdd.n5231 vdd.n5210 878.823
R28778 vdd.n5231 vdd.n5205 878.823
R28779 vdd.n5209 vdd.n5208 878.823
R28780 vdd.n5208 vdd.n5204 878.823
R28781 vdd.n5214 vdd.n5212 878.823
R28782 vdd.n5225 vdd.n5214 878.823
R28783 vdd.n5281 vdd.n5260 878.823
R28784 vdd.n5281 vdd.n5255 878.823
R28785 vdd.n5259 vdd.n5258 878.823
R28786 vdd.n5258 vdd.n5254 878.823
R28787 vdd.n5264 vdd.n5262 878.823
R28788 vdd.n5275 vdd.n5264 878.823
R28789 vdd.n5328 vdd.n5307 878.823
R28790 vdd.n5328 vdd.n5302 878.823
R28791 vdd.n5306 vdd.n5305 878.823
R28792 vdd.n5305 vdd.n5301 878.823
R28793 vdd.n5311 vdd.n5309 878.823
R28794 vdd.n5322 vdd.n5311 878.823
R28795 vdd.n5378 vdd.n5357 878.823
R28796 vdd.n5378 vdd.n5352 878.823
R28797 vdd.n5356 vdd.n5355 878.823
R28798 vdd.n5355 vdd.n5351 878.823
R28799 vdd.n5361 vdd.n5359 878.823
R28800 vdd.n5372 vdd.n5361 878.823
R28801 vdd.n5428 vdd.n5407 878.823
R28802 vdd.n5428 vdd.n5402 878.823
R28803 vdd.n5406 vdd.n5405 878.823
R28804 vdd.n5405 vdd.n5401 878.823
R28805 vdd.n5411 vdd.n5409 878.823
R28806 vdd.n5422 vdd.n5411 878.823
R28807 vdd.n5476 vdd.n5455 878.823
R28808 vdd.n5476 vdd.n5450 878.823
R28809 vdd.n5454 vdd.n5453 878.823
R28810 vdd.n5453 vdd.n5449 878.823
R28811 vdd.n5459 vdd.n5457 878.823
R28812 vdd.n5470 vdd.n5459 878.823
R28813 vdd.n4382 vdd.n4381 878.823
R28814 vdd.n4382 vdd.n4378 878.823
R28815 vdd.n4399 vdd.n4376 878.823
R28816 vdd.n4399 vdd.n4398 878.823
R28817 vdd.n4373 vdd.n4372 878.823
R28818 vdd.n4373 vdd.n4370 878.823
R28819 vdd.n5527 vdd.n5506 878.823
R28820 vdd.n5527 vdd.n5501 878.823
R28821 vdd.n5505 vdd.n5504 878.823
R28822 vdd.n5504 vdd.n5500 878.823
R28823 vdd.n5510 vdd.n5508 878.823
R28824 vdd.n5521 vdd.n5510 878.823
R28825 vdd.n5574 vdd.n5553 878.823
R28826 vdd.n5574 vdd.n5548 878.823
R28827 vdd.n5552 vdd.n5551 878.823
R28828 vdd.n5551 vdd.n5547 878.823
R28829 vdd.n5557 vdd.n5555 878.823
R28830 vdd.n5568 vdd.n5557 878.823
R28831 vdd.n5624 vdd.n5603 878.823
R28832 vdd.n5624 vdd.n5598 878.823
R28833 vdd.n5602 vdd.n5601 878.823
R28834 vdd.n5601 vdd.n5597 878.823
R28835 vdd.n5607 vdd.n5605 878.823
R28836 vdd.n5618 vdd.n5607 878.823
R28837 vdd.n5674 vdd.n5653 878.823
R28838 vdd.n5674 vdd.n5648 878.823
R28839 vdd.n5652 vdd.n5651 878.823
R28840 vdd.n5651 vdd.n5647 878.823
R28841 vdd.n5657 vdd.n5655 878.823
R28842 vdd.n5668 vdd.n5657 878.823
R28843 vdd.n5722 vdd.n5701 878.823
R28844 vdd.n5722 vdd.n5696 878.823
R28845 vdd.n5700 vdd.n5699 878.823
R28846 vdd.n5699 vdd.n5695 878.823
R28847 vdd.n5705 vdd.n5703 878.823
R28848 vdd.n5716 vdd.n5705 878.823
R28849 vdd.n5845 vdd.n5841 878.823
R28850 vdd.n5846 vdd.n5845 878.823
R28851 vdd.n5862 vdd.n5851 878.823
R28852 vdd.n5851 vdd.n5849 878.823
R28853 vdd.n5868 vdd.n5842 878.823
R28854 vdd.n5868 vdd.n5847 878.823
R28855 vdd.n5797 vdd.n5793 878.823
R28856 vdd.n5798 vdd.n5797 878.823
R28857 vdd.n5814 vdd.n5803 878.823
R28858 vdd.n5803 vdd.n5801 878.823
R28859 vdd.n5820 vdd.n5794 878.823
R28860 vdd.n5820 vdd.n5799 878.823
R28861 vdd.n5894 vdd.n5890 878.823
R28862 vdd.n5895 vdd.n5894 878.823
R28863 vdd.n5911 vdd.n5900 878.823
R28864 vdd.n5900 vdd.n5898 878.823
R28865 vdd.n5917 vdd.n5891 878.823
R28866 vdd.n5917 vdd.n5896 878.823
R28867 vdd.n5944 vdd.n5940 878.823
R28868 vdd.n5945 vdd.n5944 878.823
R28869 vdd.n5961 vdd.n5950 878.823
R28870 vdd.n5950 vdd.n5948 878.823
R28871 vdd.n5967 vdd.n5941 878.823
R28872 vdd.n5967 vdd.n5946 878.823
R28873 vdd.n5992 vdd.n5988 878.823
R28874 vdd.n5993 vdd.n5992 878.823
R28875 vdd.n6009 vdd.n5998 878.823
R28876 vdd.n5998 vdd.n5996 878.823
R28877 vdd.n6015 vdd.n5989 878.823
R28878 vdd.n6015 vdd.n5994 878.823
R28879 vdd.n4202 vdd.n4176 878.823
R28880 vdd.n4202 vdd.n4177 878.823
R28881 vdd.n4184 vdd.n4180 878.823
R28882 vdd.n4185 vdd.n4184 878.823
R28883 vdd.n4209 vdd.n4208 878.823
R28884 vdd.n4208 vdd.n4172 878.823
R28885 vdd.n6140 vdd.n6136 878.823
R28886 vdd.n6141 vdd.n6140 878.823
R28887 vdd.n6157 vdd.n6146 878.823
R28888 vdd.n6146 vdd.n6144 878.823
R28889 vdd.n6163 vdd.n6137 878.823
R28890 vdd.n6163 vdd.n6142 878.823
R28891 vdd.n6091 vdd.n6087 878.823
R28892 vdd.n6092 vdd.n6091 878.823
R28893 vdd.n6108 vdd.n6097 878.823
R28894 vdd.n6097 vdd.n6095 878.823
R28895 vdd.n6114 vdd.n6088 878.823
R28896 vdd.n6114 vdd.n6093 878.823
R28897 vdd.n6043 vdd.n6039 878.823
R28898 vdd.n6044 vdd.n6043 878.823
R28899 vdd.n6060 vdd.n6049 878.823
R28900 vdd.n6049 vdd.n6047 878.823
R28901 vdd.n6066 vdd.n6040 878.823
R28902 vdd.n6066 vdd.n6045 878.823
R28903 vdd.n6189 vdd.n6185 878.823
R28904 vdd.n6190 vdd.n6189 878.823
R28905 vdd.n6206 vdd.n6195 878.823
R28906 vdd.n6195 vdd.n6193 878.823
R28907 vdd.n6212 vdd.n6186 878.823
R28908 vdd.n6212 vdd.n6191 878.823
R28909 vdd.n6239 vdd.n6235 878.823
R28910 vdd.n6240 vdd.n6239 878.823
R28911 vdd.n6256 vdd.n6245 878.823
R28912 vdd.n6245 vdd.n6243 878.823
R28913 vdd.n6262 vdd.n6236 878.823
R28914 vdd.n6262 vdd.n6241 878.823
R28915 vdd.n6287 vdd.n6283 878.823
R28916 vdd.n6288 vdd.n6287 878.823
R28917 vdd.n6304 vdd.n6293 878.823
R28918 vdd.n6293 vdd.n6291 878.823
R28919 vdd.n6310 vdd.n6284 878.823
R28920 vdd.n6310 vdd.n6289 878.823
R28921 vdd.n6385 vdd.n6381 878.823
R28922 vdd.n6386 vdd.n6385 878.823
R28923 vdd.n6402 vdd.n6391 878.823
R28924 vdd.n6391 vdd.n6389 878.823
R28925 vdd.n6408 vdd.n6382 878.823
R28926 vdd.n6408 vdd.n6387 878.823
R28927 vdd.n6337 vdd.n6333 878.823
R28928 vdd.n6338 vdd.n6337 878.823
R28929 vdd.n6354 vdd.n6343 878.823
R28930 vdd.n6343 vdd.n6341 878.823
R28931 vdd.n6360 vdd.n6334 878.823
R28932 vdd.n6360 vdd.n6339 878.823
R28933 vdd.n6434 vdd.n6430 878.823
R28934 vdd.n6435 vdd.n6434 878.823
R28935 vdd.n6451 vdd.n6440 878.823
R28936 vdd.n6440 vdd.n6438 878.823
R28937 vdd.n6457 vdd.n6431 878.823
R28938 vdd.n6457 vdd.n6436 878.823
R28939 vdd.n6484 vdd.n6480 878.823
R28940 vdd.n6485 vdd.n6484 878.823
R28941 vdd.n6501 vdd.n6490 878.823
R28942 vdd.n6490 vdd.n6488 878.823
R28943 vdd.n6507 vdd.n6481 878.823
R28944 vdd.n6507 vdd.n6486 878.823
R28945 vdd.n6532 vdd.n6528 878.823
R28946 vdd.n6533 vdd.n6532 878.823
R28947 vdd.n6549 vdd.n6538 878.823
R28948 vdd.n6538 vdd.n6536 878.823
R28949 vdd.n6555 vdd.n6529 878.823
R28950 vdd.n6555 vdd.n6534 878.823
R28951 vdd.n3956 vdd.n3930 878.823
R28952 vdd.n3956 vdd.n3931 878.823
R28953 vdd.n3938 vdd.n3934 878.823
R28954 vdd.n3939 vdd.n3938 878.823
R28955 vdd.n3963 vdd.n3962 878.823
R28956 vdd.n3962 vdd.n3926 878.823
R28957 vdd.n6631 vdd.n6627 878.823
R28958 vdd.n6632 vdd.n6631 878.823
R28959 vdd.n6648 vdd.n6637 878.823
R28960 vdd.n6637 vdd.n6635 878.823
R28961 vdd.n6654 vdd.n6628 878.823
R28962 vdd.n6654 vdd.n6633 878.823
R28963 vdd.n6583 vdd.n6579 878.823
R28964 vdd.n6584 vdd.n6583 878.823
R28965 vdd.n6600 vdd.n6589 878.823
R28966 vdd.n6589 vdd.n6587 878.823
R28967 vdd.n6606 vdd.n6580 878.823
R28968 vdd.n6606 vdd.n6585 878.823
R28969 vdd.n6680 vdd.n6676 878.823
R28970 vdd.n6681 vdd.n6680 878.823
R28971 vdd.n6697 vdd.n6686 878.823
R28972 vdd.n6686 vdd.n6684 878.823
R28973 vdd.n6703 vdd.n6677 878.823
R28974 vdd.n6703 vdd.n6682 878.823
R28975 vdd.n6730 vdd.n6726 878.823
R28976 vdd.n6731 vdd.n6730 878.823
R28977 vdd.n6747 vdd.n6736 878.823
R28978 vdd.n6736 vdd.n6734 878.823
R28979 vdd.n6753 vdd.n6727 878.823
R28980 vdd.n6753 vdd.n6732 878.823
R28981 vdd.n6778 vdd.n6774 878.823
R28982 vdd.n6779 vdd.n6778 878.823
R28983 vdd.n6795 vdd.n6784 878.823
R28984 vdd.n6784 vdd.n6782 878.823
R28985 vdd.n6801 vdd.n6775 878.823
R28986 vdd.n6801 vdd.n6780 878.823
R28987 vdd.n690 vdd.n686 878.823
R28988 vdd.n691 vdd.n690 878.823
R28989 vdd.n707 vdd.n696 878.823
R28990 vdd.n696 vdd.n694 878.823
R28991 vdd.n713 vdd.n687 878.823
R28992 vdd.n713 vdd.n692 878.823
R28993 vdd.n738 vdd.n734 878.823
R28994 vdd.n739 vdd.n738 878.823
R28995 vdd.n755 vdd.n744 878.823
R28996 vdd.n744 vdd.n742 878.823
R28997 vdd.n761 vdd.n735 878.823
R28998 vdd.n761 vdd.n740 878.823
R28999 vdd.n840 vdd.n836 878.823
R29000 vdd.n841 vdd.n840 878.823
R29001 vdd.n857 vdd.n846 878.823
R29002 vdd.n846 vdd.n844 878.823
R29003 vdd.n863 vdd.n837 878.823
R29004 vdd.n863 vdd.n842 878.823
R29005 vdd.n888 vdd.n884 878.823
R29006 vdd.n889 vdd.n888 878.823
R29007 vdd.n905 vdd.n894 878.823
R29008 vdd.n894 vdd.n892 878.823
R29009 vdd.n911 vdd.n885 878.823
R29010 vdd.n911 vdd.n890 878.823
R29011 vdd.n936 vdd.n932 878.823
R29012 vdd.n937 vdd.n936 878.823
R29013 vdd.n953 vdd.n942 878.823
R29014 vdd.n942 vdd.n940 878.823
R29015 vdd.n959 vdd.n933 878.823
R29016 vdd.n959 vdd.n938 878.823
R29017 vdd.n984 vdd.n980 878.823
R29018 vdd.n985 vdd.n984 878.823
R29019 vdd.n1001 vdd.n990 878.823
R29020 vdd.n990 vdd.n988 878.823
R29021 vdd.n1007 vdd.n981 878.823
R29022 vdd.n1007 vdd.n986 878.823
R29023 vdd.n1086 vdd.n1082 878.823
R29024 vdd.n1087 vdd.n1086 878.823
R29025 vdd.n1103 vdd.n1092 878.823
R29026 vdd.n1092 vdd.n1090 878.823
R29027 vdd.n1109 vdd.n1083 878.823
R29028 vdd.n1109 vdd.n1088 878.823
R29029 vdd.n2606 vdd.n2602 878.823
R29030 vdd.n2607 vdd.n2606 878.823
R29031 vdd.n2623 vdd.n2612 878.823
R29032 vdd.n2612 vdd.n2610 878.823
R29033 vdd.n2629 vdd.n2603 878.823
R29034 vdd.n2629 vdd.n2608 878.823
R29035 vdd.n1157 vdd.n1136 878.823
R29036 vdd.n1157 vdd.n1131 878.823
R29037 vdd.n1135 vdd.n1134 878.823
R29038 vdd.n1134 vdd.n1130 878.823
R29039 vdd.n1140 vdd.n1138 878.823
R29040 vdd.n1151 vdd.n1140 878.823
R29041 vdd.n1205 vdd.n1184 878.823
R29042 vdd.n1205 vdd.n1179 878.823
R29043 vdd.n1183 vdd.n1182 878.823
R29044 vdd.n1182 vdd.n1178 878.823
R29045 vdd.n1188 vdd.n1186 878.823
R29046 vdd.n1199 vdd.n1188 878.823
R29047 vdd.n1306 vdd.n1285 878.823
R29048 vdd.n1306 vdd.n1280 878.823
R29049 vdd.n1284 vdd.n1283 878.823
R29050 vdd.n1283 vdd.n1279 878.823
R29051 vdd.n1289 vdd.n1287 878.823
R29052 vdd.n1300 vdd.n1289 878.823
R29053 vdd.n1354 vdd.n1333 878.823
R29054 vdd.n1354 vdd.n1328 878.823
R29055 vdd.n1332 vdd.n1331 878.823
R29056 vdd.n1331 vdd.n1327 878.823
R29057 vdd.n1337 vdd.n1335 878.823
R29058 vdd.n1348 vdd.n1337 878.823
R29059 vdd.n1402 vdd.n1381 878.823
R29060 vdd.n1402 vdd.n1376 878.823
R29061 vdd.n1380 vdd.n1379 878.823
R29062 vdd.n1379 vdd.n1375 878.823
R29063 vdd.n1385 vdd.n1383 878.823
R29064 vdd.n1396 vdd.n1385 878.823
R29065 vdd.n1450 vdd.n1429 878.823
R29066 vdd.n1450 vdd.n1424 878.823
R29067 vdd.n1428 vdd.n1427 878.823
R29068 vdd.n1427 vdd.n1423 878.823
R29069 vdd.n1433 vdd.n1431 878.823
R29070 vdd.n1444 vdd.n1433 878.823
R29071 vdd.n1551 vdd.n1530 878.823
R29072 vdd.n1551 vdd.n1525 878.823
R29073 vdd.n1529 vdd.n1528 878.823
R29074 vdd.n1528 vdd.n1524 878.823
R29075 vdd.n1534 vdd.n1532 878.823
R29076 vdd.n1545 vdd.n1534 878.823
R29077 vdd.n664 vdd.n643 878.823
R29078 vdd.n664 vdd.n638 878.823
R29079 vdd.n642 vdd.n641 878.823
R29080 vdd.n641 vdd.n637 878.823
R29081 vdd.n647 vdd.n645 878.823
R29082 vdd.n658 vdd.n647 878.823
R29083 vdd.n1599 vdd.n1578 878.823
R29084 vdd.n1599 vdd.n1573 878.823
R29085 vdd.n1577 vdd.n1576 878.823
R29086 vdd.n1576 vdd.n1572 878.823
R29087 vdd.n1582 vdd.n1580 878.823
R29088 vdd.n1593 vdd.n1582 878.823
R29089 vdd.n1646 vdd.n1625 878.823
R29090 vdd.n1646 vdd.n1620 878.823
R29091 vdd.n1624 vdd.n1623 878.823
R29092 vdd.n1623 vdd.n1619 878.823
R29093 vdd.n1629 vdd.n1627 878.823
R29094 vdd.n1640 vdd.n1629 878.823
R29095 vdd.n1696 vdd.n1675 878.823
R29096 vdd.n1696 vdd.n1670 878.823
R29097 vdd.n1674 vdd.n1673 878.823
R29098 vdd.n1673 vdd.n1669 878.823
R29099 vdd.n1679 vdd.n1677 878.823
R29100 vdd.n1690 vdd.n1679 878.823
R29101 vdd.n1746 vdd.n1725 878.823
R29102 vdd.n1746 vdd.n1720 878.823
R29103 vdd.n1724 vdd.n1723 878.823
R29104 vdd.n1723 vdd.n1719 878.823
R29105 vdd.n1729 vdd.n1727 878.823
R29106 vdd.n1740 vdd.n1729 878.823
R29107 vdd.n1794 vdd.n1773 878.823
R29108 vdd.n1794 vdd.n1768 878.823
R29109 vdd.n1772 vdd.n1771 878.823
R29110 vdd.n1771 vdd.n1767 878.823
R29111 vdd.n1777 vdd.n1775 878.823
R29112 vdd.n1788 vdd.n1777 878.823
R29113 vdd.n1485 vdd.n1484 878.823
R29114 vdd.n1485 vdd.n1481 878.823
R29115 vdd.n1502 vdd.n1479 878.823
R29116 vdd.n1502 vdd.n1501 878.823
R29117 vdd.n1476 vdd.n1475 878.823
R29118 vdd.n1476 vdd.n1473 878.823
R29119 vdd.n1845 vdd.n1824 878.823
R29120 vdd.n1845 vdd.n1819 878.823
R29121 vdd.n1823 vdd.n1822 878.823
R29122 vdd.n1822 vdd.n1818 878.823
R29123 vdd.n1828 vdd.n1826 878.823
R29124 vdd.n1839 vdd.n1828 878.823
R29125 vdd.n1892 vdd.n1871 878.823
R29126 vdd.n1892 vdd.n1866 878.823
R29127 vdd.n1870 vdd.n1869 878.823
R29128 vdd.n1869 vdd.n1865 878.823
R29129 vdd.n1875 vdd.n1873 878.823
R29130 vdd.n1886 vdd.n1875 878.823
R29131 vdd.n1940 vdd.n1919 878.823
R29132 vdd.n1940 vdd.n1914 878.823
R29133 vdd.n1918 vdd.n1917 878.823
R29134 vdd.n1917 vdd.n1913 878.823
R29135 vdd.n1923 vdd.n1921 878.823
R29136 vdd.n1934 vdd.n1923 878.823
R29137 vdd.n1991 vdd.n1970 878.823
R29138 vdd.n1991 vdd.n1965 878.823
R29139 vdd.n1969 vdd.n1968 878.823
R29140 vdd.n1968 vdd.n1964 878.823
R29141 vdd.n1974 vdd.n1972 878.823
R29142 vdd.n1985 vdd.n1974 878.823
R29143 vdd.n2041 vdd.n2020 878.823
R29144 vdd.n2041 vdd.n2015 878.823
R29145 vdd.n2019 vdd.n2018 878.823
R29146 vdd.n2018 vdd.n2014 878.823
R29147 vdd.n2024 vdd.n2022 878.823
R29148 vdd.n2035 vdd.n2024 878.823
R29149 vdd.n2089 vdd.n2068 878.823
R29150 vdd.n2089 vdd.n2063 878.823
R29151 vdd.n2067 vdd.n2066 878.823
R29152 vdd.n2066 vdd.n2062 878.823
R29153 vdd.n2072 vdd.n2070 878.823
R29154 vdd.n2083 vdd.n2072 878.823
R29155 vdd.n2139 vdd.n2118 878.823
R29156 vdd.n2139 vdd.n2113 878.823
R29157 vdd.n2117 vdd.n2116 878.823
R29158 vdd.n2116 vdd.n2112 878.823
R29159 vdd.n2122 vdd.n2120 878.823
R29160 vdd.n2133 vdd.n2122 878.823
R29161 vdd.n2186 vdd.n2165 878.823
R29162 vdd.n2186 vdd.n2160 878.823
R29163 vdd.n2164 vdd.n2163 878.823
R29164 vdd.n2163 vdd.n2159 878.823
R29165 vdd.n2169 vdd.n2167 878.823
R29166 vdd.n2180 vdd.n2169 878.823
R29167 vdd.n2236 vdd.n2215 878.823
R29168 vdd.n2236 vdd.n2210 878.823
R29169 vdd.n2214 vdd.n2213 878.823
R29170 vdd.n2213 vdd.n2209 878.823
R29171 vdd.n2219 vdd.n2217 878.823
R29172 vdd.n2230 vdd.n2219 878.823
R29173 vdd.n2286 vdd.n2265 878.823
R29174 vdd.n2286 vdd.n2260 878.823
R29175 vdd.n2264 vdd.n2263 878.823
R29176 vdd.n2263 vdd.n2259 878.823
R29177 vdd.n2269 vdd.n2267 878.823
R29178 vdd.n2280 vdd.n2269 878.823
R29179 vdd.n2334 vdd.n2313 878.823
R29180 vdd.n2334 vdd.n2308 878.823
R29181 vdd.n2312 vdd.n2311 878.823
R29182 vdd.n2311 vdd.n2307 878.823
R29183 vdd.n2317 vdd.n2315 878.823
R29184 vdd.n2328 vdd.n2317 878.823
R29185 vdd.n1240 vdd.n1239 878.823
R29186 vdd.n1240 vdd.n1236 878.823
R29187 vdd.n1257 vdd.n1234 878.823
R29188 vdd.n1257 vdd.n1256 878.823
R29189 vdd.n1231 vdd.n1230 878.823
R29190 vdd.n1231 vdd.n1228 878.823
R29191 vdd.n2385 vdd.n2364 878.823
R29192 vdd.n2385 vdd.n2359 878.823
R29193 vdd.n2363 vdd.n2362 878.823
R29194 vdd.n2362 vdd.n2358 878.823
R29195 vdd.n2368 vdd.n2366 878.823
R29196 vdd.n2379 vdd.n2368 878.823
R29197 vdd.n2432 vdd.n2411 878.823
R29198 vdd.n2432 vdd.n2406 878.823
R29199 vdd.n2410 vdd.n2409 878.823
R29200 vdd.n2409 vdd.n2405 878.823
R29201 vdd.n2415 vdd.n2413 878.823
R29202 vdd.n2426 vdd.n2415 878.823
R29203 vdd.n2482 vdd.n2461 878.823
R29204 vdd.n2482 vdd.n2456 878.823
R29205 vdd.n2460 vdd.n2459 878.823
R29206 vdd.n2459 vdd.n2455 878.823
R29207 vdd.n2465 vdd.n2463 878.823
R29208 vdd.n2476 vdd.n2465 878.823
R29209 vdd.n2532 vdd.n2511 878.823
R29210 vdd.n2532 vdd.n2506 878.823
R29211 vdd.n2510 vdd.n2509 878.823
R29212 vdd.n2509 vdd.n2505 878.823
R29213 vdd.n2515 vdd.n2513 878.823
R29214 vdd.n2526 vdd.n2515 878.823
R29215 vdd.n2580 vdd.n2559 878.823
R29216 vdd.n2580 vdd.n2554 878.823
R29217 vdd.n2558 vdd.n2557 878.823
R29218 vdd.n2557 vdd.n2553 878.823
R29219 vdd.n2563 vdd.n2561 878.823
R29220 vdd.n2574 vdd.n2563 878.823
R29221 vdd.n2703 vdd.n2699 878.823
R29222 vdd.n2704 vdd.n2703 878.823
R29223 vdd.n2720 vdd.n2709 878.823
R29224 vdd.n2709 vdd.n2707 878.823
R29225 vdd.n2726 vdd.n2700 878.823
R29226 vdd.n2726 vdd.n2705 878.823
R29227 vdd.n2655 vdd.n2651 878.823
R29228 vdd.n2656 vdd.n2655 878.823
R29229 vdd.n2672 vdd.n2661 878.823
R29230 vdd.n2661 vdd.n2659 878.823
R29231 vdd.n2678 vdd.n2652 878.823
R29232 vdd.n2678 vdd.n2657 878.823
R29233 vdd.n2752 vdd.n2748 878.823
R29234 vdd.n2753 vdd.n2752 878.823
R29235 vdd.n2769 vdd.n2758 878.823
R29236 vdd.n2758 vdd.n2756 878.823
R29237 vdd.n2775 vdd.n2749 878.823
R29238 vdd.n2775 vdd.n2754 878.823
R29239 vdd.n2802 vdd.n2798 878.823
R29240 vdd.n2803 vdd.n2802 878.823
R29241 vdd.n2819 vdd.n2808 878.823
R29242 vdd.n2808 vdd.n2806 878.823
R29243 vdd.n2825 vdd.n2799 878.823
R29244 vdd.n2825 vdd.n2804 878.823
R29245 vdd.n2850 vdd.n2846 878.823
R29246 vdd.n2851 vdd.n2850 878.823
R29247 vdd.n2867 vdd.n2856 878.823
R29248 vdd.n2856 vdd.n2854 878.823
R29249 vdd.n2873 vdd.n2847 878.823
R29250 vdd.n2873 vdd.n2852 878.823
R29251 vdd.n1060 vdd.n1034 878.823
R29252 vdd.n1060 vdd.n1035 878.823
R29253 vdd.n1042 vdd.n1038 878.823
R29254 vdd.n1043 vdd.n1042 878.823
R29255 vdd.n1067 vdd.n1066 878.823
R29256 vdd.n1066 vdd.n1030 878.823
R29257 vdd.n2998 vdd.n2994 878.823
R29258 vdd.n2999 vdd.n2998 878.823
R29259 vdd.n3015 vdd.n3004 878.823
R29260 vdd.n3004 vdd.n3002 878.823
R29261 vdd.n3021 vdd.n2995 878.823
R29262 vdd.n3021 vdd.n3000 878.823
R29263 vdd.n2949 vdd.n2945 878.823
R29264 vdd.n2950 vdd.n2949 878.823
R29265 vdd.n2966 vdd.n2955 878.823
R29266 vdd.n2955 vdd.n2953 878.823
R29267 vdd.n2972 vdd.n2946 878.823
R29268 vdd.n2972 vdd.n2951 878.823
R29269 vdd.n2901 vdd.n2897 878.823
R29270 vdd.n2902 vdd.n2901 878.823
R29271 vdd.n2918 vdd.n2907 878.823
R29272 vdd.n2907 vdd.n2905 878.823
R29273 vdd.n2924 vdd.n2898 878.823
R29274 vdd.n2924 vdd.n2903 878.823
R29275 vdd.n3047 vdd.n3043 878.823
R29276 vdd.n3048 vdd.n3047 878.823
R29277 vdd.n3064 vdd.n3053 878.823
R29278 vdd.n3053 vdd.n3051 878.823
R29279 vdd.n3070 vdd.n3044 878.823
R29280 vdd.n3070 vdd.n3049 878.823
R29281 vdd.n3097 vdd.n3093 878.823
R29282 vdd.n3098 vdd.n3097 878.823
R29283 vdd.n3114 vdd.n3103 878.823
R29284 vdd.n3103 vdd.n3101 878.823
R29285 vdd.n3120 vdd.n3094 878.823
R29286 vdd.n3120 vdd.n3099 878.823
R29287 vdd.n3145 vdd.n3141 878.823
R29288 vdd.n3146 vdd.n3145 878.823
R29289 vdd.n3162 vdd.n3151 878.823
R29290 vdd.n3151 vdd.n3149 878.823
R29291 vdd.n3168 vdd.n3142 878.823
R29292 vdd.n3168 vdd.n3147 878.823
R29293 vdd.n3243 vdd.n3239 878.823
R29294 vdd.n3244 vdd.n3243 878.823
R29295 vdd.n3260 vdd.n3249 878.823
R29296 vdd.n3249 vdd.n3247 878.823
R29297 vdd.n3266 vdd.n3240 878.823
R29298 vdd.n3266 vdd.n3245 878.823
R29299 vdd.n3195 vdd.n3191 878.823
R29300 vdd.n3196 vdd.n3195 878.823
R29301 vdd.n3212 vdd.n3201 878.823
R29302 vdd.n3201 vdd.n3199 878.823
R29303 vdd.n3218 vdd.n3192 878.823
R29304 vdd.n3218 vdd.n3197 878.823
R29305 vdd.n3292 vdd.n3288 878.823
R29306 vdd.n3293 vdd.n3292 878.823
R29307 vdd.n3309 vdd.n3298 878.823
R29308 vdd.n3298 vdd.n3296 878.823
R29309 vdd.n3315 vdd.n3289 878.823
R29310 vdd.n3315 vdd.n3294 878.823
R29311 vdd.n3342 vdd.n3338 878.823
R29312 vdd.n3343 vdd.n3342 878.823
R29313 vdd.n3359 vdd.n3348 878.823
R29314 vdd.n3348 vdd.n3346 878.823
R29315 vdd.n3365 vdd.n3339 878.823
R29316 vdd.n3365 vdd.n3344 878.823
R29317 vdd.n3390 vdd.n3386 878.823
R29318 vdd.n3391 vdd.n3390 878.823
R29319 vdd.n3407 vdd.n3396 878.823
R29320 vdd.n3396 vdd.n3394 878.823
R29321 vdd.n3413 vdd.n3387 878.823
R29322 vdd.n3413 vdd.n3392 878.823
R29323 vdd.n814 vdd.n788 878.823
R29324 vdd.n814 vdd.n789 878.823
R29325 vdd.n796 vdd.n792 878.823
R29326 vdd.n797 vdd.n796 878.823
R29327 vdd.n821 vdd.n820 878.823
R29328 vdd.n820 vdd.n784 878.823
R29329 vdd.n3489 vdd.n3485 878.823
R29330 vdd.n3490 vdd.n3489 878.823
R29331 vdd.n3506 vdd.n3495 878.823
R29332 vdd.n3495 vdd.n3493 878.823
R29333 vdd.n3512 vdd.n3486 878.823
R29334 vdd.n3512 vdd.n3491 878.823
R29335 vdd.n3441 vdd.n3437 878.823
R29336 vdd.n3442 vdd.n3441 878.823
R29337 vdd.n3458 vdd.n3447 878.823
R29338 vdd.n3447 vdd.n3445 878.823
R29339 vdd.n3464 vdd.n3438 878.823
R29340 vdd.n3464 vdd.n3443 878.823
R29341 vdd.n3538 vdd.n3534 878.823
R29342 vdd.n3539 vdd.n3538 878.823
R29343 vdd.n3555 vdd.n3544 878.823
R29344 vdd.n3544 vdd.n3542 878.823
R29345 vdd.n3561 vdd.n3535 878.823
R29346 vdd.n3561 vdd.n3540 878.823
R29347 vdd.n3588 vdd.n3584 878.823
R29348 vdd.n3589 vdd.n3588 878.823
R29349 vdd.n3605 vdd.n3594 878.823
R29350 vdd.n3594 vdd.n3592 878.823
R29351 vdd.n3611 vdd.n3585 878.823
R29352 vdd.n3611 vdd.n3590 878.823
R29353 vdd.n3636 vdd.n3632 878.823
R29354 vdd.n3637 vdd.n3636 878.823
R29355 vdd.n3653 vdd.n3642 878.823
R29356 vdd.n3642 vdd.n3640 878.823
R29357 vdd.n3659 vdd.n3633 878.823
R29358 vdd.n3659 vdd.n3638 878.823
R29359 vdd.n594 vdd.n590 878.823
R29360 vdd.n595 vdd.n594 878.823
R29361 vdd.n611 vdd.n600 878.823
R29362 vdd.n600 vdd.n598 878.823
R29363 vdd.n617 vdd.n591 878.823
R29364 vdd.n617 vdd.n596 878.823
R29365 vdd.n3735 vdd.n3731 878.823
R29366 vdd.n3736 vdd.n3735 878.823
R29367 vdd.n3752 vdd.n3741 878.823
R29368 vdd.n3741 vdd.n3739 878.823
R29369 vdd.n3758 vdd.n3732 878.823
R29370 vdd.n3758 vdd.n3737 878.823
R29371 vdd.n3687 vdd.n3683 878.823
R29372 vdd.n3688 vdd.n3687 878.823
R29373 vdd.n3704 vdd.n3693 878.823
R29374 vdd.n3693 vdd.n3691 878.823
R29375 vdd.n3710 vdd.n3684 878.823
R29376 vdd.n3710 vdd.n3689 878.823
R29377 vdd.n6877 vdd.n6873 878.823
R29378 vdd.n6878 vdd.n6877 878.823
R29379 vdd.n6894 vdd.n6883 878.823
R29380 vdd.n6883 vdd.n6881 878.823
R29381 vdd.n6900 vdd.n6874 878.823
R29382 vdd.n6900 vdd.n6879 878.823
R29383 vdd.n6829 vdd.n6825 878.823
R29384 vdd.n6830 vdd.n6829 878.823
R29385 vdd.n6846 vdd.n6835 878.823
R29386 vdd.n6835 vdd.n6833 878.823
R29387 vdd.n6852 vdd.n6826 878.823
R29388 vdd.n6852 vdd.n6831 878.823
R29389 vdd.n10019 vdd.n10015 878.823
R29390 vdd.n10020 vdd.n10019 878.823
R29391 vdd.n10036 vdd.n10025 878.823
R29392 vdd.n10025 vdd.n10023 878.823
R29393 vdd.n10042 vdd.n10016 878.823
R29394 vdd.n10042 vdd.n10021 878.823
R29395 vdd.n9971 vdd.n9967 878.823
R29396 vdd.n9972 vdd.n9971 878.823
R29397 vdd.n9988 vdd.n9977 878.823
R29398 vdd.n9977 vdd.n9975 878.823
R29399 vdd.n9994 vdd.n9968 878.823
R29400 vdd.n9994 vdd.n9973 878.823
R29401 vdd.n10067 vdd.n10063 878.823
R29402 vdd.n10068 vdd.n10067 878.823
R29403 vdd.n10084 vdd.n10073 878.823
R29404 vdd.n10073 vdd.n10071 878.823
R29405 vdd.n10090 vdd.n10064 878.823
R29406 vdd.n10090 vdd.n10069 878.823
R29407 vdd.n10115 vdd.n10111 878.823
R29408 vdd.n10116 vdd.n10115 878.823
R29409 vdd.n10132 vdd.n10121 878.823
R29410 vdd.n10121 vdd.n10119 878.823
R29411 vdd.n10138 vdd.n10112 878.823
R29412 vdd.n10138 vdd.n10117 878.823
R29413 vdd.n10217 vdd.n10213 878.823
R29414 vdd.n10218 vdd.n10217 878.823
R29415 vdd.n10234 vdd.n10223 878.823
R29416 vdd.n10223 vdd.n10221 878.823
R29417 vdd.n10240 vdd.n10214 878.823
R29418 vdd.n10240 vdd.n10219 878.823
R29419 vdd.n10265 vdd.n10261 878.823
R29420 vdd.n10266 vdd.n10265 878.823
R29421 vdd.n10282 vdd.n10271 878.823
R29422 vdd.n10271 vdd.n10269 878.823
R29423 vdd.n10288 vdd.n10262 878.823
R29424 vdd.n10288 vdd.n10267 878.823
R29425 vdd.n10313 vdd.n10309 878.823
R29426 vdd.n10314 vdd.n10313 878.823
R29427 vdd.n10330 vdd.n10319 878.823
R29428 vdd.n10319 vdd.n10317 878.823
R29429 vdd.n10336 vdd.n10310 878.823
R29430 vdd.n10336 vdd.n10315 878.823
R29431 vdd.n10361 vdd.n10357 878.823
R29432 vdd.n10362 vdd.n10361 878.823
R29433 vdd.n10378 vdd.n10367 878.823
R29434 vdd.n10367 vdd.n10365 878.823
R29435 vdd.n10384 vdd.n10358 878.823
R29436 vdd.n10384 vdd.n10363 878.823
R29437 vdd.n10463 vdd.n10459 878.823
R29438 vdd.n10464 vdd.n10463 878.823
R29439 vdd.n10480 vdd.n10469 878.823
R29440 vdd.n10469 vdd.n10467 878.823
R29441 vdd.n10486 vdd.n10460 878.823
R29442 vdd.n10486 vdd.n10465 878.823
R29443 vdd.n55 vdd.n51 878.823
R29444 vdd.n56 vdd.n55 878.823
R29445 vdd.n72 vdd.n61 878.823
R29446 vdd.n61 vdd.n59 878.823
R29447 vdd.n78 vdd.n52 878.823
R29448 vdd.n78 vdd.n57 878.823
R29449 vdd.n7 vdd.n3 878.823
R29450 vdd.n8 vdd.n7 878.823
R29451 vdd.n24 vdd.n13 878.823
R29452 vdd.n13 vdd.n11 878.823
R29453 vdd.n30 vdd.n4 878.823
R29454 vdd.n30 vdd.n9 878.823
R29455 vdd.n10511 vdd.n10507 878.823
R29456 vdd.n10512 vdd.n10511 878.823
R29457 vdd.n10528 vdd.n10517 878.823
R29458 vdd.n10517 vdd.n10515 878.823
R29459 vdd.n10534 vdd.n10508 878.823
R29460 vdd.n10534 vdd.n10513 878.823
R29461 vdd.n10561 vdd.n10557 878.823
R29462 vdd.n10562 vdd.n10561 878.823
R29463 vdd.n10578 vdd.n10567 878.823
R29464 vdd.n10567 vdd.n10565 878.823
R29465 vdd.n10584 vdd.n10558 878.823
R29466 vdd.n10584 vdd.n10563 878.823
R29467 vdd.n10609 vdd.n10605 878.823
R29468 vdd.n10610 vdd.n10609 878.823
R29469 vdd.n10626 vdd.n10615 878.823
R29470 vdd.n10615 vdd.n10613 878.823
R29471 vdd.n10632 vdd.n10606 878.823
R29472 vdd.n10632 vdd.n10611 878.823
R29473 vdd.n10437 vdd.n10411 878.823
R29474 vdd.n10437 vdd.n10412 878.823
R29475 vdd.n10419 vdd.n10415 878.823
R29476 vdd.n10420 vdd.n10419 878.823
R29477 vdd.n10444 vdd.n10443 878.823
R29478 vdd.n10443 vdd.n10407 878.823
R29479 vdd.n10757 vdd.n10753 878.823
R29480 vdd.n10758 vdd.n10757 878.823
R29481 vdd.n10774 vdd.n10763 878.823
R29482 vdd.n10763 vdd.n10761 878.823
R29483 vdd.n10780 vdd.n10754 878.823
R29484 vdd.n10780 vdd.n10759 878.823
R29485 vdd.n10708 vdd.n10704 878.823
R29486 vdd.n10709 vdd.n10708 878.823
R29487 vdd.n10725 vdd.n10714 878.823
R29488 vdd.n10714 vdd.n10712 878.823
R29489 vdd.n10731 vdd.n10705 878.823
R29490 vdd.n10731 vdd.n10710 878.823
R29491 vdd.n10660 vdd.n10656 878.823
R29492 vdd.n10661 vdd.n10660 878.823
R29493 vdd.n10677 vdd.n10666 878.823
R29494 vdd.n10666 vdd.n10664 878.823
R29495 vdd.n10683 vdd.n10657 878.823
R29496 vdd.n10683 vdd.n10662 878.823
R29497 vdd.n10806 vdd.n10802 878.823
R29498 vdd.n10807 vdd.n10806 878.823
R29499 vdd.n10823 vdd.n10812 878.823
R29500 vdd.n10812 vdd.n10810 878.823
R29501 vdd.n10829 vdd.n10803 878.823
R29502 vdd.n10829 vdd.n10808 878.823
R29503 vdd.n10856 vdd.n10852 878.823
R29504 vdd.n10857 vdd.n10856 878.823
R29505 vdd.n10873 vdd.n10862 878.823
R29506 vdd.n10862 vdd.n10860 878.823
R29507 vdd.n10879 vdd.n10853 878.823
R29508 vdd.n10879 vdd.n10858 878.823
R29509 vdd.n10904 vdd.n10900 878.823
R29510 vdd.n10905 vdd.n10904 878.823
R29511 vdd.n10921 vdd.n10910 878.823
R29512 vdd.n10910 vdd.n10908 878.823
R29513 vdd.n10927 vdd.n10901 878.823
R29514 vdd.n10927 vdd.n10906 878.823
R29515 vdd.n11002 vdd.n10998 878.823
R29516 vdd.n11003 vdd.n11002 878.823
R29517 vdd.n11019 vdd.n11008 878.823
R29518 vdd.n11008 vdd.n11006 878.823
R29519 vdd.n11025 vdd.n10999 878.823
R29520 vdd.n11025 vdd.n11004 878.823
R29521 vdd.n10954 vdd.n10950 878.823
R29522 vdd.n10955 vdd.n10954 878.823
R29523 vdd.n10971 vdd.n10960 878.823
R29524 vdd.n10960 vdd.n10958 878.823
R29525 vdd.n10977 vdd.n10951 878.823
R29526 vdd.n10977 vdd.n10956 878.823
R29527 vdd.n11051 vdd.n11047 878.823
R29528 vdd.n11052 vdd.n11051 878.823
R29529 vdd.n11068 vdd.n11057 878.823
R29530 vdd.n11057 vdd.n11055 878.823
R29531 vdd.n11074 vdd.n11048 878.823
R29532 vdd.n11074 vdd.n11053 878.823
R29533 vdd.n11101 vdd.n11097 878.823
R29534 vdd.n11102 vdd.n11101 878.823
R29535 vdd.n11118 vdd.n11107 878.823
R29536 vdd.n11107 vdd.n11105 878.823
R29537 vdd.n11124 vdd.n11098 878.823
R29538 vdd.n11124 vdd.n11103 878.823
R29539 vdd.n11149 vdd.n11145 878.823
R29540 vdd.n11150 vdd.n11149 878.823
R29541 vdd.n11166 vdd.n11155 878.823
R29542 vdd.n11155 vdd.n11153 878.823
R29543 vdd.n11172 vdd.n11146 878.823
R29544 vdd.n11172 vdd.n11151 878.823
R29545 vdd.n10191 vdd.n10165 878.823
R29546 vdd.n10191 vdd.n10166 878.823
R29547 vdd.n10173 vdd.n10169 878.823
R29548 vdd.n10174 vdd.n10173 878.823
R29549 vdd.n10198 vdd.n10197 878.823
R29550 vdd.n10197 vdd.n10161 878.823
R29551 vdd.n11248 vdd.n11244 878.823
R29552 vdd.n11249 vdd.n11248 878.823
R29553 vdd.n11265 vdd.n11254 878.823
R29554 vdd.n11254 vdd.n11252 878.823
R29555 vdd.n11271 vdd.n11245 878.823
R29556 vdd.n11271 vdd.n11250 878.823
R29557 vdd.n11200 vdd.n11196 878.823
R29558 vdd.n11201 vdd.n11200 878.823
R29559 vdd.n11217 vdd.n11206 878.823
R29560 vdd.n11206 vdd.n11204 878.823
R29561 vdd.n11223 vdd.n11197 878.823
R29562 vdd.n11223 vdd.n11202 878.823
R29563 vdd.n11297 vdd.n11293 878.823
R29564 vdd.n11298 vdd.n11297 878.823
R29565 vdd.n11314 vdd.n11303 878.823
R29566 vdd.n11303 vdd.n11301 878.823
R29567 vdd.n11320 vdd.n11294 878.823
R29568 vdd.n11320 vdd.n11299 878.823
R29569 vdd.n11347 vdd.n11343 878.823
R29570 vdd.n11348 vdd.n11347 878.823
R29571 vdd.n11364 vdd.n11353 878.823
R29572 vdd.n11353 vdd.n11351 878.823
R29573 vdd.n11370 vdd.n11344 878.823
R29574 vdd.n11370 vdd.n11349 878.823
R29575 vdd.n11395 vdd.n11391 878.823
R29576 vdd.n11396 vdd.n11395 878.823
R29577 vdd.n11412 vdd.n11401 878.823
R29578 vdd.n11401 vdd.n11399 878.823
R29579 vdd.n11418 vdd.n11392 878.823
R29580 vdd.n11418 vdd.n11397 878.823
R29581 vdd.n11469 vdd.n11448 878.823
R29582 vdd.n11469 vdd.n11443 878.823
R29583 vdd.n11447 vdd.n11446 878.823
R29584 vdd.n11446 vdd.n11442 878.823
R29585 vdd.n11452 vdd.n11450 878.823
R29586 vdd.n11463 vdd.n11452 878.823
R29587 vdd.n11516 vdd.n11495 878.823
R29588 vdd.n11516 vdd.n11490 878.823
R29589 vdd.n11494 vdd.n11493 878.823
R29590 vdd.n11493 vdd.n11489 878.823
R29591 vdd.n11499 vdd.n11497 878.823
R29592 vdd.n11510 vdd.n11499 878.823
R29593 vdd.n11566 vdd.n11545 878.823
R29594 vdd.n11566 vdd.n11540 878.823
R29595 vdd.n11544 vdd.n11543 878.823
R29596 vdd.n11543 vdd.n11539 878.823
R29597 vdd.n11549 vdd.n11547 878.823
R29598 vdd.n11560 vdd.n11549 878.823
R29599 vdd.n11616 vdd.n11595 878.823
R29600 vdd.n11616 vdd.n11590 878.823
R29601 vdd.n11594 vdd.n11593 878.823
R29602 vdd.n11593 vdd.n11589 878.823
R29603 vdd.n11599 vdd.n11597 878.823
R29604 vdd.n11610 vdd.n11599 878.823
R29605 vdd.n11664 vdd.n11643 878.823
R29606 vdd.n11664 vdd.n11638 878.823
R29607 vdd.n11642 vdd.n11641 878.823
R29608 vdd.n11641 vdd.n11637 878.823
R29609 vdd.n11647 vdd.n11645 878.823
R29610 vdd.n11658 vdd.n11647 878.823
R29611 vdd.n455 vdd.n454 878.823
R29612 vdd.n455 vdd.n451 878.823
R29613 vdd.n472 vdd.n449 878.823
R29614 vdd.n472 vdd.n471 878.823
R29615 vdd.n446 vdd.n445 878.823
R29616 vdd.n446 vdd.n443 878.823
R29617 vdd.n11715 vdd.n11694 878.823
R29618 vdd.n11715 vdd.n11689 878.823
R29619 vdd.n11693 vdd.n11692 878.823
R29620 vdd.n11692 vdd.n11688 878.823
R29621 vdd.n11698 vdd.n11696 878.823
R29622 vdd.n11709 vdd.n11698 878.823
R29623 vdd.n11762 vdd.n11741 878.823
R29624 vdd.n11762 vdd.n11736 878.823
R29625 vdd.n11740 vdd.n11739 878.823
R29626 vdd.n11739 vdd.n11735 878.823
R29627 vdd.n11745 vdd.n11743 878.823
R29628 vdd.n11756 vdd.n11745 878.823
R29629 vdd.n11810 vdd.n11789 878.823
R29630 vdd.n11810 vdd.n11784 878.823
R29631 vdd.n11788 vdd.n11787 878.823
R29632 vdd.n11787 vdd.n11783 878.823
R29633 vdd.n11793 vdd.n11791 878.823
R29634 vdd.n11804 vdd.n11793 878.823
R29635 vdd.n11861 vdd.n11840 878.823
R29636 vdd.n11861 vdd.n11835 878.823
R29637 vdd.n11839 vdd.n11838 878.823
R29638 vdd.n11838 vdd.n11834 878.823
R29639 vdd.n11844 vdd.n11842 878.823
R29640 vdd.n11855 vdd.n11844 878.823
R29641 vdd.n11911 vdd.n11890 878.823
R29642 vdd.n11911 vdd.n11885 878.823
R29643 vdd.n11889 vdd.n11888 878.823
R29644 vdd.n11888 vdd.n11884 878.823
R29645 vdd.n11894 vdd.n11892 878.823
R29646 vdd.n11905 vdd.n11894 878.823
R29647 vdd.n11959 vdd.n11938 878.823
R29648 vdd.n11959 vdd.n11933 878.823
R29649 vdd.n11937 vdd.n11936 878.823
R29650 vdd.n11936 vdd.n11932 878.823
R29651 vdd.n11942 vdd.n11940 878.823
R29652 vdd.n11953 vdd.n11942 878.823
R29653 vdd.n12009 vdd.n11988 878.823
R29654 vdd.n12009 vdd.n11983 878.823
R29655 vdd.n11987 vdd.n11986 878.823
R29656 vdd.n11986 vdd.n11982 878.823
R29657 vdd.n11992 vdd.n11990 878.823
R29658 vdd.n12003 vdd.n11992 878.823
R29659 vdd.n12056 vdd.n12035 878.823
R29660 vdd.n12056 vdd.n12030 878.823
R29661 vdd.n12034 vdd.n12033 878.823
R29662 vdd.n12033 vdd.n12029 878.823
R29663 vdd.n12039 vdd.n12037 878.823
R29664 vdd.n12050 vdd.n12039 878.823
R29665 vdd.n12106 vdd.n12085 878.823
R29666 vdd.n12106 vdd.n12080 878.823
R29667 vdd.n12084 vdd.n12083 878.823
R29668 vdd.n12083 vdd.n12079 878.823
R29669 vdd.n12089 vdd.n12087 878.823
R29670 vdd.n12100 vdd.n12089 878.823
R29671 vdd.n12156 vdd.n12135 878.823
R29672 vdd.n12156 vdd.n12130 878.823
R29673 vdd.n12134 vdd.n12133 878.823
R29674 vdd.n12133 vdd.n12129 878.823
R29675 vdd.n12139 vdd.n12137 878.823
R29676 vdd.n12150 vdd.n12139 878.823
R29677 vdd.n12204 vdd.n12183 878.823
R29678 vdd.n12204 vdd.n12178 878.823
R29679 vdd.n12182 vdd.n12181 878.823
R29680 vdd.n12181 vdd.n12177 878.823
R29681 vdd.n12187 vdd.n12185 878.823
R29682 vdd.n12198 vdd.n12187 878.823
R29683 vdd.n210 vdd.n209 878.823
R29684 vdd.n210 vdd.n206 878.823
R29685 vdd.n227 vdd.n204 878.823
R29686 vdd.n227 vdd.n226 878.823
R29687 vdd.n201 vdd.n200 878.823
R29688 vdd.n201 vdd.n198 878.823
R29689 vdd.n12255 vdd.n12234 878.823
R29690 vdd.n12255 vdd.n12229 878.823
R29691 vdd.n12233 vdd.n12232 878.823
R29692 vdd.n12232 vdd.n12228 878.823
R29693 vdd.n12238 vdd.n12236 878.823
R29694 vdd.n12249 vdd.n12238 878.823
R29695 vdd.n12302 vdd.n12281 878.823
R29696 vdd.n12302 vdd.n12276 878.823
R29697 vdd.n12280 vdd.n12279 878.823
R29698 vdd.n12279 vdd.n12275 878.823
R29699 vdd.n12285 vdd.n12283 878.823
R29700 vdd.n12296 vdd.n12285 878.823
R29701 vdd.n12352 vdd.n12331 878.823
R29702 vdd.n12352 vdd.n12326 878.823
R29703 vdd.n12330 vdd.n12329 878.823
R29704 vdd.n12329 vdd.n12325 878.823
R29705 vdd.n12335 vdd.n12333 878.823
R29706 vdd.n12346 vdd.n12335 878.823
R29707 vdd.n12402 vdd.n12381 878.823
R29708 vdd.n12402 vdd.n12376 878.823
R29709 vdd.n12380 vdd.n12379 878.823
R29710 vdd.n12379 vdd.n12375 878.823
R29711 vdd.n12385 vdd.n12383 878.823
R29712 vdd.n12396 vdd.n12385 878.823
R29713 vdd.n12450 vdd.n12429 878.823
R29714 vdd.n12450 vdd.n12424 878.823
R29715 vdd.n12428 vdd.n12427 878.823
R29716 vdd.n12427 vdd.n12423 878.823
R29717 vdd.n12433 vdd.n12431 878.823
R29718 vdd.n12444 vdd.n12433 878.823
R29719 vdd.n12494 vdd.n12485 681.178
R29720 vdd.n12494 vdd.n12486 681.178
R29721 vdd.n12514 vdd.n12508 681.178
R29722 vdd.n12492 vdd.n12487 681.178
R29723 vdd.n12492 vdd.n12488 681.178
R29724 vdd.n12512 vdd.n12509 681.178
R29725 vdd.n117 vdd.n108 681.178
R29726 vdd.n124 vdd.n108 681.178
R29727 vdd.n124 vdd.n105 681.178
R29728 vdd.n139 vdd.n105 681.178
R29729 vdd.n139 vdd.n106 681.178
R29730 vdd.n135 vdd.n106 681.178
R29731 vdd.n121 vdd.n120 681.178
R29732 vdd.n122 vdd.n121 681.178
R29733 vdd.n122 vdd.n100 681.178
R29734 vdd.n141 vdd.n100 681.178
R29735 vdd.n141 vdd.n101 681.178
R29736 vdd.n132 vdd.n101 681.178
R29737 vdd.n165 vdd.n156 681.178
R29738 vdd.n172 vdd.n156 681.178
R29739 vdd.n172 vdd.n153 681.178
R29740 vdd.n187 vdd.n153 681.178
R29741 vdd.n187 vdd.n154 681.178
R29742 vdd.n183 vdd.n154 681.178
R29743 vdd.n169 vdd.n168 681.178
R29744 vdd.n170 vdd.n169 681.178
R29745 vdd.n170 vdd.n148 681.178
R29746 vdd.n189 vdd.n148 681.178
R29747 vdd.n189 vdd.n149 681.178
R29748 vdd.n180 vdd.n149 681.178
R29749 vdd.n266 vdd.n257 681.178
R29750 vdd.n273 vdd.n257 681.178
R29751 vdd.n273 vdd.n254 681.178
R29752 vdd.n288 vdd.n254 681.178
R29753 vdd.n288 vdd.n255 681.178
R29754 vdd.n284 vdd.n255 681.178
R29755 vdd.n270 vdd.n269 681.178
R29756 vdd.n271 vdd.n270 681.178
R29757 vdd.n271 vdd.n249 681.178
R29758 vdd.n290 vdd.n249 681.178
R29759 vdd.n290 vdd.n250 681.178
R29760 vdd.n281 vdd.n250 681.178
R29761 vdd.n314 vdd.n305 681.178
R29762 vdd.n321 vdd.n305 681.178
R29763 vdd.n321 vdd.n302 681.178
R29764 vdd.n336 vdd.n302 681.178
R29765 vdd.n336 vdd.n303 681.178
R29766 vdd.n332 vdd.n303 681.178
R29767 vdd.n318 vdd.n317 681.178
R29768 vdd.n319 vdd.n318 681.178
R29769 vdd.n319 vdd.n297 681.178
R29770 vdd.n338 vdd.n297 681.178
R29771 vdd.n338 vdd.n298 681.178
R29772 vdd.n329 vdd.n298 681.178
R29773 vdd.n362 vdd.n353 681.178
R29774 vdd.n369 vdd.n353 681.178
R29775 vdd.n369 vdd.n350 681.178
R29776 vdd.n384 vdd.n350 681.178
R29777 vdd.n384 vdd.n351 681.178
R29778 vdd.n380 vdd.n351 681.178
R29779 vdd.n366 vdd.n365 681.178
R29780 vdd.n367 vdd.n366 681.178
R29781 vdd.n367 vdd.n345 681.178
R29782 vdd.n386 vdd.n345 681.178
R29783 vdd.n386 vdd.n346 681.178
R29784 vdd.n377 vdd.n346 681.178
R29785 vdd.n410 vdd.n401 681.178
R29786 vdd.n417 vdd.n401 681.178
R29787 vdd.n417 vdd.n398 681.178
R29788 vdd.n432 vdd.n398 681.178
R29789 vdd.n432 vdd.n399 681.178
R29790 vdd.n428 vdd.n399 681.178
R29791 vdd.n414 vdd.n413 681.178
R29792 vdd.n415 vdd.n414 681.178
R29793 vdd.n415 vdd.n393 681.178
R29794 vdd.n434 vdd.n393 681.178
R29795 vdd.n434 vdd.n394 681.178
R29796 vdd.n425 vdd.n394 681.178
R29797 vdd.n511 vdd.n502 681.178
R29798 vdd.n518 vdd.n502 681.178
R29799 vdd.n518 vdd.n499 681.178
R29800 vdd.n533 vdd.n499 681.178
R29801 vdd.n533 vdd.n500 681.178
R29802 vdd.n529 vdd.n500 681.178
R29803 vdd.n515 vdd.n514 681.178
R29804 vdd.n516 vdd.n515 681.178
R29805 vdd.n516 vdd.n494 681.178
R29806 vdd.n535 vdd.n494 681.178
R29807 vdd.n535 vdd.n495 681.178
R29808 vdd.n526 vdd.n495 681.178
R29809 vdd.n559 vdd.n550 681.178
R29810 vdd.n566 vdd.n550 681.178
R29811 vdd.n566 vdd.n547 681.178
R29812 vdd.n581 vdd.n547 681.178
R29813 vdd.n581 vdd.n548 681.178
R29814 vdd.n577 vdd.n548 681.178
R29815 vdd.n563 vdd.n562 681.178
R29816 vdd.n564 vdd.n563 681.178
R29817 vdd.n564 vdd.n542 681.178
R29818 vdd.n583 vdd.n542 681.178
R29819 vdd.n583 vdd.n543 681.178
R29820 vdd.n574 vdd.n543 681.178
R29821 vdd.n6991 vdd.n6990 681.178
R29822 vdd.n6992 vdd.n6991 681.178
R29823 vdd.n6992 vdd.n6970 681.178
R29824 vdd.n7011 vdd.n6970 681.178
R29825 vdd.n7011 vdd.n6971 681.178
R29826 vdd.n7002 vdd.n6971 681.178
R29827 vdd.n6984 vdd.n6978 681.178
R29828 vdd.n6994 vdd.n6978 681.178
R29829 vdd.n6994 vdd.n6975 681.178
R29830 vdd.n7009 vdd.n6975 681.178
R29831 vdd.n7009 vdd.n6976 681.178
R29832 vdd.n7005 vdd.n6976 681.178
R29833 vdd.n7039 vdd.n7038 681.178
R29834 vdd.n7040 vdd.n7039 681.178
R29835 vdd.n7040 vdd.n7018 681.178
R29836 vdd.n7059 vdd.n7018 681.178
R29837 vdd.n7059 vdd.n7019 681.178
R29838 vdd.n7050 vdd.n7019 681.178
R29839 vdd.n7032 vdd.n7026 681.178
R29840 vdd.n7042 vdd.n7026 681.178
R29841 vdd.n7042 vdd.n7023 681.178
R29842 vdd.n7057 vdd.n7023 681.178
R29843 vdd.n7057 vdd.n7024 681.178
R29844 vdd.n7053 vdd.n7024 681.178
R29845 vdd.n7141 vdd.n7140 681.178
R29846 vdd.n7142 vdd.n7141 681.178
R29847 vdd.n7142 vdd.n7120 681.178
R29848 vdd.n7161 vdd.n7120 681.178
R29849 vdd.n7161 vdd.n7121 681.178
R29850 vdd.n7152 vdd.n7121 681.178
R29851 vdd.n7134 vdd.n7128 681.178
R29852 vdd.n7144 vdd.n7128 681.178
R29853 vdd.n7144 vdd.n7125 681.178
R29854 vdd.n7159 vdd.n7125 681.178
R29855 vdd.n7159 vdd.n7126 681.178
R29856 vdd.n7155 vdd.n7126 681.178
R29857 vdd.n7189 vdd.n7188 681.178
R29858 vdd.n7190 vdd.n7189 681.178
R29859 vdd.n7190 vdd.n7168 681.178
R29860 vdd.n7209 vdd.n7168 681.178
R29861 vdd.n7209 vdd.n7169 681.178
R29862 vdd.n7200 vdd.n7169 681.178
R29863 vdd.n7182 vdd.n7176 681.178
R29864 vdd.n7192 vdd.n7176 681.178
R29865 vdd.n7192 vdd.n7173 681.178
R29866 vdd.n7207 vdd.n7173 681.178
R29867 vdd.n7207 vdd.n7174 681.178
R29868 vdd.n7203 vdd.n7174 681.178
R29869 vdd.n7237 vdd.n7236 681.178
R29870 vdd.n7238 vdd.n7237 681.178
R29871 vdd.n7238 vdd.n7216 681.178
R29872 vdd.n7257 vdd.n7216 681.178
R29873 vdd.n7257 vdd.n7217 681.178
R29874 vdd.n7248 vdd.n7217 681.178
R29875 vdd.n7230 vdd.n7224 681.178
R29876 vdd.n7240 vdd.n7224 681.178
R29877 vdd.n7240 vdd.n7221 681.178
R29878 vdd.n7255 vdd.n7221 681.178
R29879 vdd.n7255 vdd.n7222 681.178
R29880 vdd.n7251 vdd.n7222 681.178
R29881 vdd.n7285 vdd.n7284 681.178
R29882 vdd.n7286 vdd.n7285 681.178
R29883 vdd.n7286 vdd.n7264 681.178
R29884 vdd.n7305 vdd.n7264 681.178
R29885 vdd.n7305 vdd.n7265 681.178
R29886 vdd.n7296 vdd.n7265 681.178
R29887 vdd.n7278 vdd.n7272 681.178
R29888 vdd.n7288 vdd.n7272 681.178
R29889 vdd.n7288 vdd.n7269 681.178
R29890 vdd.n7303 vdd.n7269 681.178
R29891 vdd.n7303 vdd.n7270 681.178
R29892 vdd.n7299 vdd.n7270 681.178
R29893 vdd.n7387 vdd.n7386 681.178
R29894 vdd.n7388 vdd.n7387 681.178
R29895 vdd.n7388 vdd.n7366 681.178
R29896 vdd.n7407 vdd.n7366 681.178
R29897 vdd.n7407 vdd.n7367 681.178
R29898 vdd.n7398 vdd.n7367 681.178
R29899 vdd.n7380 vdd.n7374 681.178
R29900 vdd.n7390 vdd.n7374 681.178
R29901 vdd.n7390 vdd.n7371 681.178
R29902 vdd.n7405 vdd.n7371 681.178
R29903 vdd.n7405 vdd.n7372 681.178
R29904 vdd.n7401 vdd.n7372 681.178
R29905 vdd.n8907 vdd.n8906 681.178
R29906 vdd.n8908 vdd.n8907 681.178
R29907 vdd.n8908 vdd.n8886 681.178
R29908 vdd.n8927 vdd.n8886 681.178
R29909 vdd.n8927 vdd.n8887 681.178
R29910 vdd.n8918 vdd.n8887 681.178
R29911 vdd.n8900 vdd.n8894 681.178
R29912 vdd.n8910 vdd.n8894 681.178
R29913 vdd.n8910 vdd.n8891 681.178
R29914 vdd.n8925 vdd.n8891 681.178
R29915 vdd.n8925 vdd.n8892 681.178
R29916 vdd.n8921 vdd.n8892 681.178
R29917 vdd.n7431 vdd.n7422 681.178
R29918 vdd.n7438 vdd.n7422 681.178
R29919 vdd.n7438 vdd.n7419 681.178
R29920 vdd.n7453 vdd.n7419 681.178
R29921 vdd.n7453 vdd.n7420 681.178
R29922 vdd.n7449 vdd.n7420 681.178
R29923 vdd.n7435 vdd.n7434 681.178
R29924 vdd.n7436 vdd.n7435 681.178
R29925 vdd.n7436 vdd.n7414 681.178
R29926 vdd.n7455 vdd.n7414 681.178
R29927 vdd.n7455 vdd.n7415 681.178
R29928 vdd.n7446 vdd.n7415 681.178
R29929 vdd.n7479 vdd.n7470 681.178
R29930 vdd.n7486 vdd.n7470 681.178
R29931 vdd.n7486 vdd.n7467 681.178
R29932 vdd.n7501 vdd.n7467 681.178
R29933 vdd.n7501 vdd.n7468 681.178
R29934 vdd.n7497 vdd.n7468 681.178
R29935 vdd.n7483 vdd.n7482 681.178
R29936 vdd.n7484 vdd.n7483 681.178
R29937 vdd.n7484 vdd.n7462 681.178
R29938 vdd.n7503 vdd.n7462 681.178
R29939 vdd.n7503 vdd.n7463 681.178
R29940 vdd.n7494 vdd.n7463 681.178
R29941 vdd.n7580 vdd.n7571 681.178
R29942 vdd.n7587 vdd.n7571 681.178
R29943 vdd.n7587 vdd.n7568 681.178
R29944 vdd.n7602 vdd.n7568 681.178
R29945 vdd.n7602 vdd.n7569 681.178
R29946 vdd.n7598 vdd.n7569 681.178
R29947 vdd.n7584 vdd.n7583 681.178
R29948 vdd.n7585 vdd.n7584 681.178
R29949 vdd.n7585 vdd.n7563 681.178
R29950 vdd.n7604 vdd.n7563 681.178
R29951 vdd.n7604 vdd.n7564 681.178
R29952 vdd.n7595 vdd.n7564 681.178
R29953 vdd.n7628 vdd.n7619 681.178
R29954 vdd.n7635 vdd.n7619 681.178
R29955 vdd.n7635 vdd.n7616 681.178
R29956 vdd.n7650 vdd.n7616 681.178
R29957 vdd.n7650 vdd.n7617 681.178
R29958 vdd.n7646 vdd.n7617 681.178
R29959 vdd.n7632 vdd.n7631 681.178
R29960 vdd.n7633 vdd.n7632 681.178
R29961 vdd.n7633 vdd.n7611 681.178
R29962 vdd.n7652 vdd.n7611 681.178
R29963 vdd.n7652 vdd.n7612 681.178
R29964 vdd.n7643 vdd.n7612 681.178
R29965 vdd.n7676 vdd.n7667 681.178
R29966 vdd.n7683 vdd.n7667 681.178
R29967 vdd.n7683 vdd.n7664 681.178
R29968 vdd.n7698 vdd.n7664 681.178
R29969 vdd.n7698 vdd.n7665 681.178
R29970 vdd.n7694 vdd.n7665 681.178
R29971 vdd.n7680 vdd.n7679 681.178
R29972 vdd.n7681 vdd.n7680 681.178
R29973 vdd.n7681 vdd.n7659 681.178
R29974 vdd.n7700 vdd.n7659 681.178
R29975 vdd.n7700 vdd.n7660 681.178
R29976 vdd.n7691 vdd.n7660 681.178
R29977 vdd.n7724 vdd.n7715 681.178
R29978 vdd.n7731 vdd.n7715 681.178
R29979 vdd.n7731 vdd.n7712 681.178
R29980 vdd.n7746 vdd.n7712 681.178
R29981 vdd.n7746 vdd.n7713 681.178
R29982 vdd.n7742 vdd.n7713 681.178
R29983 vdd.n7728 vdd.n7727 681.178
R29984 vdd.n7729 vdd.n7728 681.178
R29985 vdd.n7729 vdd.n7707 681.178
R29986 vdd.n7748 vdd.n7707 681.178
R29987 vdd.n7748 vdd.n7708 681.178
R29988 vdd.n7739 vdd.n7708 681.178
R29989 vdd.n7825 vdd.n7816 681.178
R29990 vdd.n7832 vdd.n7816 681.178
R29991 vdd.n7832 vdd.n7813 681.178
R29992 vdd.n7847 vdd.n7813 681.178
R29993 vdd.n7847 vdd.n7814 681.178
R29994 vdd.n7843 vdd.n7814 681.178
R29995 vdd.n7829 vdd.n7828 681.178
R29996 vdd.n7830 vdd.n7829 681.178
R29997 vdd.n7830 vdd.n7808 681.178
R29998 vdd.n7849 vdd.n7808 681.178
R29999 vdd.n7849 vdd.n7809 681.178
R30000 vdd.n7840 vdd.n7809 681.178
R30001 vdd.n6938 vdd.n6929 681.178
R30002 vdd.n6945 vdd.n6929 681.178
R30003 vdd.n6945 vdd.n6926 681.178
R30004 vdd.n6960 vdd.n6926 681.178
R30005 vdd.n6960 vdd.n6927 681.178
R30006 vdd.n6956 vdd.n6927 681.178
R30007 vdd.n6942 vdd.n6941 681.178
R30008 vdd.n6943 vdd.n6942 681.178
R30009 vdd.n6943 vdd.n6921 681.178
R30010 vdd.n6962 vdd.n6921 681.178
R30011 vdd.n6962 vdd.n6922 681.178
R30012 vdd.n6953 vdd.n6922 681.178
R30013 vdd.n7873 vdd.n7864 681.178
R30014 vdd.n7880 vdd.n7864 681.178
R30015 vdd.n7880 vdd.n7861 681.178
R30016 vdd.n7895 vdd.n7861 681.178
R30017 vdd.n7895 vdd.n7862 681.178
R30018 vdd.n7891 vdd.n7862 681.178
R30019 vdd.n7877 vdd.n7876 681.178
R30020 vdd.n7878 vdd.n7877 681.178
R30021 vdd.n7878 vdd.n7856 681.178
R30022 vdd.n7897 vdd.n7856 681.178
R30023 vdd.n7897 vdd.n7857 681.178
R30024 vdd.n7888 vdd.n7857 681.178
R30025 vdd.n7920 vdd.n7911 681.178
R30026 vdd.n7927 vdd.n7911 681.178
R30027 vdd.n7927 vdd.n7908 681.178
R30028 vdd.n7942 vdd.n7908 681.178
R30029 vdd.n7942 vdd.n7909 681.178
R30030 vdd.n7938 vdd.n7909 681.178
R30031 vdd.n7924 vdd.n7923 681.178
R30032 vdd.n7925 vdd.n7924 681.178
R30033 vdd.n7925 vdd.n7903 681.178
R30034 vdd.n7944 vdd.n7903 681.178
R30035 vdd.n7944 vdd.n7904 681.178
R30036 vdd.n7935 vdd.n7904 681.178
R30037 vdd.n7970 vdd.n7961 681.178
R30038 vdd.n7977 vdd.n7961 681.178
R30039 vdd.n7977 vdd.n7958 681.178
R30040 vdd.n7992 vdd.n7958 681.178
R30041 vdd.n7992 vdd.n7959 681.178
R30042 vdd.n7988 vdd.n7959 681.178
R30043 vdd.n7974 vdd.n7973 681.178
R30044 vdd.n7975 vdd.n7974 681.178
R30045 vdd.n7975 vdd.n7953 681.178
R30046 vdd.n7994 vdd.n7953 681.178
R30047 vdd.n7994 vdd.n7954 681.178
R30048 vdd.n7985 vdd.n7954 681.178
R30049 vdd.n8020 vdd.n8011 681.178
R30050 vdd.n8027 vdd.n8011 681.178
R30051 vdd.n8027 vdd.n8008 681.178
R30052 vdd.n8042 vdd.n8008 681.178
R30053 vdd.n8042 vdd.n8009 681.178
R30054 vdd.n8038 vdd.n8009 681.178
R30055 vdd.n8024 vdd.n8023 681.178
R30056 vdd.n8025 vdd.n8024 681.178
R30057 vdd.n8025 vdd.n8003 681.178
R30058 vdd.n8044 vdd.n8003 681.178
R30059 vdd.n8044 vdd.n8004 681.178
R30060 vdd.n8035 vdd.n8004 681.178
R30061 vdd.n8068 vdd.n8059 681.178
R30062 vdd.n8075 vdd.n8059 681.178
R30063 vdd.n8075 vdd.n8056 681.178
R30064 vdd.n8090 vdd.n8056 681.178
R30065 vdd.n8090 vdd.n8057 681.178
R30066 vdd.n8086 vdd.n8057 681.178
R30067 vdd.n8072 vdd.n8071 681.178
R30068 vdd.n8073 vdd.n8072 681.178
R30069 vdd.n8073 vdd.n8051 681.178
R30070 vdd.n8092 vdd.n8051 681.178
R30071 vdd.n8092 vdd.n8052 681.178
R30072 vdd.n8083 vdd.n8052 681.178
R30073 vdd.n7796 vdd.n7759 681.178
R30074 vdd.n7792 vdd.n7759 681.178
R30075 vdd.n7792 vdd.n7763 681.178
R30076 vdd.n7782 vdd.n7763 681.178
R30077 vdd.n7782 vdd.n7768 681.178
R30078 vdd.n7778 vdd.n7768 681.178
R30079 vdd.n7799 vdd.n7757 681.178
R30080 vdd.n7790 vdd.n7757 681.178
R30081 vdd.n7790 vdd.n7785 681.178
R30082 vdd.n7785 vdd.n7784 681.178
R30083 vdd.n7784 vdd.n7765 681.178
R30084 vdd.n7775 vdd.n7765 681.178
R30085 vdd.n8119 vdd.n8110 681.178
R30086 vdd.n8126 vdd.n8110 681.178
R30087 vdd.n8126 vdd.n8107 681.178
R30088 vdd.n8141 vdd.n8107 681.178
R30089 vdd.n8141 vdd.n8108 681.178
R30090 vdd.n8137 vdd.n8108 681.178
R30091 vdd.n8123 vdd.n8122 681.178
R30092 vdd.n8124 vdd.n8123 681.178
R30093 vdd.n8124 vdd.n8102 681.178
R30094 vdd.n8143 vdd.n8102 681.178
R30095 vdd.n8143 vdd.n8103 681.178
R30096 vdd.n8134 vdd.n8103 681.178
R30097 vdd.n8166 vdd.n8157 681.178
R30098 vdd.n8173 vdd.n8157 681.178
R30099 vdd.n8173 vdd.n8154 681.178
R30100 vdd.n8188 vdd.n8154 681.178
R30101 vdd.n8188 vdd.n8155 681.178
R30102 vdd.n8184 vdd.n8155 681.178
R30103 vdd.n8170 vdd.n8169 681.178
R30104 vdd.n8171 vdd.n8170 681.178
R30105 vdd.n8171 vdd.n8149 681.178
R30106 vdd.n8190 vdd.n8149 681.178
R30107 vdd.n8190 vdd.n8150 681.178
R30108 vdd.n8181 vdd.n8150 681.178
R30109 vdd.n8214 vdd.n8205 681.178
R30110 vdd.n8221 vdd.n8205 681.178
R30111 vdd.n8221 vdd.n8202 681.178
R30112 vdd.n8236 vdd.n8202 681.178
R30113 vdd.n8236 vdd.n8203 681.178
R30114 vdd.n8232 vdd.n8203 681.178
R30115 vdd.n8218 vdd.n8217 681.178
R30116 vdd.n8219 vdd.n8218 681.178
R30117 vdd.n8219 vdd.n8197 681.178
R30118 vdd.n8238 vdd.n8197 681.178
R30119 vdd.n8238 vdd.n8198 681.178
R30120 vdd.n8229 vdd.n8198 681.178
R30121 vdd.n8265 vdd.n8256 681.178
R30122 vdd.n8272 vdd.n8256 681.178
R30123 vdd.n8272 vdd.n8253 681.178
R30124 vdd.n8287 vdd.n8253 681.178
R30125 vdd.n8287 vdd.n8254 681.178
R30126 vdd.n8283 vdd.n8254 681.178
R30127 vdd.n8269 vdd.n8268 681.178
R30128 vdd.n8270 vdd.n8269 681.178
R30129 vdd.n8270 vdd.n8248 681.178
R30130 vdd.n8289 vdd.n8248 681.178
R30131 vdd.n8289 vdd.n8249 681.178
R30132 vdd.n8280 vdd.n8249 681.178
R30133 vdd.n8315 vdd.n8306 681.178
R30134 vdd.n8322 vdd.n8306 681.178
R30135 vdd.n8322 vdd.n8303 681.178
R30136 vdd.n8337 vdd.n8303 681.178
R30137 vdd.n8337 vdd.n8304 681.178
R30138 vdd.n8333 vdd.n8304 681.178
R30139 vdd.n8319 vdd.n8318 681.178
R30140 vdd.n8320 vdd.n8319 681.178
R30141 vdd.n8320 vdd.n8298 681.178
R30142 vdd.n8339 vdd.n8298 681.178
R30143 vdd.n8339 vdd.n8299 681.178
R30144 vdd.n8330 vdd.n8299 681.178
R30145 vdd.n8363 vdd.n8354 681.178
R30146 vdd.n8370 vdd.n8354 681.178
R30147 vdd.n8370 vdd.n8351 681.178
R30148 vdd.n8385 vdd.n8351 681.178
R30149 vdd.n8385 vdd.n8352 681.178
R30150 vdd.n8381 vdd.n8352 681.178
R30151 vdd.n8367 vdd.n8366 681.178
R30152 vdd.n8368 vdd.n8367 681.178
R30153 vdd.n8368 vdd.n8346 681.178
R30154 vdd.n8387 vdd.n8346 681.178
R30155 vdd.n8387 vdd.n8347 681.178
R30156 vdd.n8378 vdd.n8347 681.178
R30157 vdd.n8413 vdd.n8404 681.178
R30158 vdd.n8420 vdd.n8404 681.178
R30159 vdd.n8420 vdd.n8401 681.178
R30160 vdd.n8435 vdd.n8401 681.178
R30161 vdd.n8435 vdd.n8402 681.178
R30162 vdd.n8431 vdd.n8402 681.178
R30163 vdd.n8417 vdd.n8416 681.178
R30164 vdd.n8418 vdd.n8417 681.178
R30165 vdd.n8418 vdd.n8396 681.178
R30166 vdd.n8437 vdd.n8396 681.178
R30167 vdd.n8437 vdd.n8397 681.178
R30168 vdd.n8428 vdd.n8397 681.178
R30169 vdd.n8460 vdd.n8451 681.178
R30170 vdd.n8467 vdd.n8451 681.178
R30171 vdd.n8467 vdd.n8448 681.178
R30172 vdd.n8482 vdd.n8448 681.178
R30173 vdd.n8482 vdd.n8449 681.178
R30174 vdd.n8478 vdd.n8449 681.178
R30175 vdd.n8464 vdd.n8463 681.178
R30176 vdd.n8465 vdd.n8464 681.178
R30177 vdd.n8465 vdd.n8443 681.178
R30178 vdd.n8484 vdd.n8443 681.178
R30179 vdd.n8484 vdd.n8444 681.178
R30180 vdd.n8475 vdd.n8444 681.178
R30181 vdd.n8510 vdd.n8501 681.178
R30182 vdd.n8517 vdd.n8501 681.178
R30183 vdd.n8517 vdd.n8498 681.178
R30184 vdd.n8532 vdd.n8498 681.178
R30185 vdd.n8532 vdd.n8499 681.178
R30186 vdd.n8528 vdd.n8499 681.178
R30187 vdd.n8514 vdd.n8513 681.178
R30188 vdd.n8515 vdd.n8514 681.178
R30189 vdd.n8515 vdd.n8493 681.178
R30190 vdd.n8534 vdd.n8493 681.178
R30191 vdd.n8534 vdd.n8494 681.178
R30192 vdd.n8525 vdd.n8494 681.178
R30193 vdd.n8560 vdd.n8551 681.178
R30194 vdd.n8567 vdd.n8551 681.178
R30195 vdd.n8567 vdd.n8548 681.178
R30196 vdd.n8582 vdd.n8548 681.178
R30197 vdd.n8582 vdd.n8549 681.178
R30198 vdd.n8578 vdd.n8549 681.178
R30199 vdd.n8564 vdd.n8563 681.178
R30200 vdd.n8565 vdd.n8564 681.178
R30201 vdd.n8565 vdd.n8543 681.178
R30202 vdd.n8584 vdd.n8543 681.178
R30203 vdd.n8584 vdd.n8544 681.178
R30204 vdd.n8575 vdd.n8544 681.178
R30205 vdd.n8608 vdd.n8599 681.178
R30206 vdd.n8615 vdd.n8599 681.178
R30207 vdd.n8615 vdd.n8596 681.178
R30208 vdd.n8630 vdd.n8596 681.178
R30209 vdd.n8630 vdd.n8597 681.178
R30210 vdd.n8626 vdd.n8597 681.178
R30211 vdd.n8612 vdd.n8611 681.178
R30212 vdd.n8613 vdd.n8612 681.178
R30213 vdd.n8613 vdd.n8591 681.178
R30214 vdd.n8632 vdd.n8591 681.178
R30215 vdd.n8632 vdd.n8592 681.178
R30216 vdd.n8623 vdd.n8592 681.178
R30217 vdd.n7551 vdd.n7514 681.178
R30218 vdd.n7547 vdd.n7514 681.178
R30219 vdd.n7547 vdd.n7518 681.178
R30220 vdd.n7537 vdd.n7518 681.178
R30221 vdd.n7537 vdd.n7523 681.178
R30222 vdd.n7533 vdd.n7523 681.178
R30223 vdd.n7554 vdd.n7512 681.178
R30224 vdd.n7545 vdd.n7512 681.178
R30225 vdd.n7545 vdd.n7540 681.178
R30226 vdd.n7540 vdd.n7539 681.178
R30227 vdd.n7539 vdd.n7520 681.178
R30228 vdd.n7530 vdd.n7520 681.178
R30229 vdd.n8659 vdd.n8650 681.178
R30230 vdd.n8666 vdd.n8650 681.178
R30231 vdd.n8666 vdd.n8647 681.178
R30232 vdd.n8681 vdd.n8647 681.178
R30233 vdd.n8681 vdd.n8648 681.178
R30234 vdd.n8677 vdd.n8648 681.178
R30235 vdd.n8663 vdd.n8662 681.178
R30236 vdd.n8664 vdd.n8663 681.178
R30237 vdd.n8664 vdd.n8642 681.178
R30238 vdd.n8683 vdd.n8642 681.178
R30239 vdd.n8683 vdd.n8643 681.178
R30240 vdd.n8674 vdd.n8643 681.178
R30241 vdd.n8706 vdd.n8697 681.178
R30242 vdd.n8713 vdd.n8697 681.178
R30243 vdd.n8713 vdd.n8694 681.178
R30244 vdd.n8728 vdd.n8694 681.178
R30245 vdd.n8728 vdd.n8695 681.178
R30246 vdd.n8724 vdd.n8695 681.178
R30247 vdd.n8710 vdd.n8709 681.178
R30248 vdd.n8711 vdd.n8710 681.178
R30249 vdd.n8711 vdd.n8689 681.178
R30250 vdd.n8730 vdd.n8689 681.178
R30251 vdd.n8730 vdd.n8690 681.178
R30252 vdd.n8721 vdd.n8690 681.178
R30253 vdd.n8756 vdd.n8747 681.178
R30254 vdd.n8763 vdd.n8747 681.178
R30255 vdd.n8763 vdd.n8744 681.178
R30256 vdd.n8778 vdd.n8744 681.178
R30257 vdd.n8778 vdd.n8745 681.178
R30258 vdd.n8774 vdd.n8745 681.178
R30259 vdd.n8760 vdd.n8759 681.178
R30260 vdd.n8761 vdd.n8760 681.178
R30261 vdd.n8761 vdd.n8739 681.178
R30262 vdd.n8780 vdd.n8739 681.178
R30263 vdd.n8780 vdd.n8740 681.178
R30264 vdd.n8771 vdd.n8740 681.178
R30265 vdd.n8806 vdd.n8797 681.178
R30266 vdd.n8813 vdd.n8797 681.178
R30267 vdd.n8813 vdd.n8794 681.178
R30268 vdd.n8828 vdd.n8794 681.178
R30269 vdd.n8828 vdd.n8795 681.178
R30270 vdd.n8824 vdd.n8795 681.178
R30271 vdd.n8810 vdd.n8809 681.178
R30272 vdd.n8811 vdd.n8810 681.178
R30273 vdd.n8811 vdd.n8789 681.178
R30274 vdd.n8830 vdd.n8789 681.178
R30275 vdd.n8830 vdd.n8790 681.178
R30276 vdd.n8821 vdd.n8790 681.178
R30277 vdd.n8854 vdd.n8845 681.178
R30278 vdd.n8861 vdd.n8845 681.178
R30279 vdd.n8861 vdd.n8842 681.178
R30280 vdd.n8876 vdd.n8842 681.178
R30281 vdd.n8876 vdd.n8843 681.178
R30282 vdd.n8872 vdd.n8843 681.178
R30283 vdd.n8858 vdd.n8857 681.178
R30284 vdd.n8859 vdd.n8858 681.178
R30285 vdd.n8859 vdd.n8837 681.178
R30286 vdd.n8878 vdd.n8837 681.178
R30287 vdd.n8878 vdd.n8838 681.178
R30288 vdd.n8869 vdd.n8838 681.178
R30289 vdd.n9004 vdd.n9003 681.178
R30290 vdd.n9005 vdd.n9004 681.178
R30291 vdd.n9005 vdd.n8983 681.178
R30292 vdd.n9024 vdd.n8983 681.178
R30293 vdd.n9024 vdd.n8984 681.178
R30294 vdd.n9015 vdd.n8984 681.178
R30295 vdd.n8997 vdd.n8991 681.178
R30296 vdd.n9007 vdd.n8991 681.178
R30297 vdd.n9007 vdd.n8988 681.178
R30298 vdd.n9022 vdd.n8988 681.178
R30299 vdd.n9022 vdd.n8989 681.178
R30300 vdd.n9018 vdd.n8989 681.178
R30301 vdd.n8956 vdd.n8955 681.178
R30302 vdd.n8957 vdd.n8956 681.178
R30303 vdd.n8957 vdd.n8935 681.178
R30304 vdd.n8976 vdd.n8935 681.178
R30305 vdd.n8976 vdd.n8936 681.178
R30306 vdd.n8967 vdd.n8936 681.178
R30307 vdd.n8949 vdd.n8943 681.178
R30308 vdd.n8959 vdd.n8943 681.178
R30309 vdd.n8959 vdd.n8940 681.178
R30310 vdd.n8974 vdd.n8940 681.178
R30311 vdd.n8974 vdd.n8941 681.178
R30312 vdd.n8970 vdd.n8941 681.178
R30313 vdd.n9053 vdd.n9052 681.178
R30314 vdd.n9054 vdd.n9053 681.178
R30315 vdd.n9054 vdd.n9032 681.178
R30316 vdd.n9073 vdd.n9032 681.178
R30317 vdd.n9073 vdd.n9033 681.178
R30318 vdd.n9064 vdd.n9033 681.178
R30319 vdd.n9046 vdd.n9040 681.178
R30320 vdd.n9056 vdd.n9040 681.178
R30321 vdd.n9056 vdd.n9037 681.178
R30322 vdd.n9071 vdd.n9037 681.178
R30323 vdd.n9071 vdd.n9038 681.178
R30324 vdd.n9067 vdd.n9038 681.178
R30325 vdd.n9103 vdd.n9102 681.178
R30326 vdd.n9104 vdd.n9103 681.178
R30327 vdd.n9104 vdd.n9082 681.178
R30328 vdd.n9123 vdd.n9082 681.178
R30329 vdd.n9123 vdd.n9083 681.178
R30330 vdd.n9114 vdd.n9083 681.178
R30331 vdd.n9096 vdd.n9090 681.178
R30332 vdd.n9106 vdd.n9090 681.178
R30333 vdd.n9106 vdd.n9087 681.178
R30334 vdd.n9121 vdd.n9087 681.178
R30335 vdd.n9121 vdd.n9088 681.178
R30336 vdd.n9117 vdd.n9088 681.178
R30337 vdd.n9151 vdd.n9150 681.178
R30338 vdd.n9152 vdd.n9151 681.178
R30339 vdd.n9152 vdd.n9130 681.178
R30340 vdd.n9171 vdd.n9130 681.178
R30341 vdd.n9171 vdd.n9131 681.178
R30342 vdd.n9162 vdd.n9131 681.178
R30343 vdd.n9144 vdd.n9138 681.178
R30344 vdd.n9154 vdd.n9138 681.178
R30345 vdd.n9154 vdd.n9135 681.178
R30346 vdd.n9169 vdd.n9135 681.178
R30347 vdd.n9169 vdd.n9136 681.178
R30348 vdd.n9165 vdd.n9136 681.178
R30349 vdd.n7334 vdd.n7322 681.178
R30350 vdd.n7338 vdd.n7322 681.178
R30351 vdd.n7338 vdd.n7318 681.178
R30352 vdd.n7318 vdd.n7316 681.178
R30353 vdd.n7351 vdd.n7316 681.178
R30354 vdd.n7352 vdd.n7351 681.178
R30355 vdd.n7331 vdd.n7327 681.178
R30356 vdd.n7327 vdd.n7321 681.178
R30357 vdd.n7321 vdd.n7319 681.178
R30358 vdd.n7341 vdd.n7319 681.178
R30359 vdd.n7341 vdd.n7314 681.178
R30360 vdd.n7355 vdd.n7314 681.178
R30361 vdd.n9299 vdd.n9298 681.178
R30362 vdd.n9300 vdd.n9299 681.178
R30363 vdd.n9300 vdd.n9278 681.178
R30364 vdd.n9319 vdd.n9278 681.178
R30365 vdd.n9319 vdd.n9279 681.178
R30366 vdd.n9310 vdd.n9279 681.178
R30367 vdd.n9292 vdd.n9286 681.178
R30368 vdd.n9302 vdd.n9286 681.178
R30369 vdd.n9302 vdd.n9283 681.178
R30370 vdd.n9317 vdd.n9283 681.178
R30371 vdd.n9317 vdd.n9284 681.178
R30372 vdd.n9313 vdd.n9284 681.178
R30373 vdd.n9250 vdd.n9249 681.178
R30374 vdd.n9251 vdd.n9250 681.178
R30375 vdd.n9251 vdd.n9229 681.178
R30376 vdd.n9270 vdd.n9229 681.178
R30377 vdd.n9270 vdd.n9230 681.178
R30378 vdd.n9261 vdd.n9230 681.178
R30379 vdd.n9243 vdd.n9237 681.178
R30380 vdd.n9253 vdd.n9237 681.178
R30381 vdd.n9253 vdd.n9234 681.178
R30382 vdd.n9268 vdd.n9234 681.178
R30383 vdd.n9268 vdd.n9235 681.178
R30384 vdd.n9264 vdd.n9235 681.178
R30385 vdd.n9202 vdd.n9201 681.178
R30386 vdd.n9203 vdd.n9202 681.178
R30387 vdd.n9203 vdd.n9181 681.178
R30388 vdd.n9222 vdd.n9181 681.178
R30389 vdd.n9222 vdd.n9182 681.178
R30390 vdd.n9213 vdd.n9182 681.178
R30391 vdd.n9195 vdd.n9189 681.178
R30392 vdd.n9205 vdd.n9189 681.178
R30393 vdd.n9205 vdd.n9186 681.178
R30394 vdd.n9220 vdd.n9186 681.178
R30395 vdd.n9220 vdd.n9187 681.178
R30396 vdd.n9216 vdd.n9187 681.178
R30397 vdd.n9348 vdd.n9347 681.178
R30398 vdd.n9349 vdd.n9348 681.178
R30399 vdd.n9349 vdd.n9327 681.178
R30400 vdd.n9368 vdd.n9327 681.178
R30401 vdd.n9368 vdd.n9328 681.178
R30402 vdd.n9359 vdd.n9328 681.178
R30403 vdd.n9341 vdd.n9335 681.178
R30404 vdd.n9351 vdd.n9335 681.178
R30405 vdd.n9351 vdd.n9332 681.178
R30406 vdd.n9366 vdd.n9332 681.178
R30407 vdd.n9366 vdd.n9333 681.178
R30408 vdd.n9362 vdd.n9333 681.178
R30409 vdd.n9398 vdd.n9397 681.178
R30410 vdd.n9399 vdd.n9398 681.178
R30411 vdd.n9399 vdd.n9377 681.178
R30412 vdd.n9418 vdd.n9377 681.178
R30413 vdd.n9418 vdd.n9378 681.178
R30414 vdd.n9409 vdd.n9378 681.178
R30415 vdd.n9391 vdd.n9385 681.178
R30416 vdd.n9401 vdd.n9385 681.178
R30417 vdd.n9401 vdd.n9382 681.178
R30418 vdd.n9416 vdd.n9382 681.178
R30419 vdd.n9416 vdd.n9383 681.178
R30420 vdd.n9412 vdd.n9383 681.178
R30421 vdd.n9446 vdd.n9445 681.178
R30422 vdd.n9447 vdd.n9446 681.178
R30423 vdd.n9447 vdd.n9425 681.178
R30424 vdd.n9466 vdd.n9425 681.178
R30425 vdd.n9466 vdd.n9426 681.178
R30426 vdd.n9457 vdd.n9426 681.178
R30427 vdd.n9439 vdd.n9433 681.178
R30428 vdd.n9449 vdd.n9433 681.178
R30429 vdd.n9449 vdd.n9430 681.178
R30430 vdd.n9464 vdd.n9430 681.178
R30431 vdd.n9464 vdd.n9431 681.178
R30432 vdd.n9460 vdd.n9431 681.178
R30433 vdd.n9544 vdd.n9543 681.178
R30434 vdd.n9545 vdd.n9544 681.178
R30435 vdd.n9545 vdd.n9523 681.178
R30436 vdd.n9564 vdd.n9523 681.178
R30437 vdd.n9564 vdd.n9524 681.178
R30438 vdd.n9555 vdd.n9524 681.178
R30439 vdd.n9537 vdd.n9531 681.178
R30440 vdd.n9547 vdd.n9531 681.178
R30441 vdd.n9547 vdd.n9528 681.178
R30442 vdd.n9562 vdd.n9528 681.178
R30443 vdd.n9562 vdd.n9529 681.178
R30444 vdd.n9558 vdd.n9529 681.178
R30445 vdd.n9496 vdd.n9495 681.178
R30446 vdd.n9497 vdd.n9496 681.178
R30447 vdd.n9497 vdd.n9475 681.178
R30448 vdd.n9516 vdd.n9475 681.178
R30449 vdd.n9516 vdd.n9476 681.178
R30450 vdd.n9507 vdd.n9476 681.178
R30451 vdd.n9489 vdd.n9483 681.178
R30452 vdd.n9499 vdd.n9483 681.178
R30453 vdd.n9499 vdd.n9480 681.178
R30454 vdd.n9514 vdd.n9480 681.178
R30455 vdd.n9514 vdd.n9481 681.178
R30456 vdd.n9510 vdd.n9481 681.178
R30457 vdd.n9593 vdd.n9592 681.178
R30458 vdd.n9594 vdd.n9593 681.178
R30459 vdd.n9594 vdd.n9572 681.178
R30460 vdd.n9613 vdd.n9572 681.178
R30461 vdd.n9613 vdd.n9573 681.178
R30462 vdd.n9604 vdd.n9573 681.178
R30463 vdd.n9586 vdd.n9580 681.178
R30464 vdd.n9596 vdd.n9580 681.178
R30465 vdd.n9596 vdd.n9577 681.178
R30466 vdd.n9611 vdd.n9577 681.178
R30467 vdd.n9611 vdd.n9578 681.178
R30468 vdd.n9607 vdd.n9578 681.178
R30469 vdd.n9643 vdd.n9642 681.178
R30470 vdd.n9644 vdd.n9643 681.178
R30471 vdd.n9644 vdd.n9622 681.178
R30472 vdd.n9663 vdd.n9622 681.178
R30473 vdd.n9663 vdd.n9623 681.178
R30474 vdd.n9654 vdd.n9623 681.178
R30475 vdd.n9636 vdd.n9630 681.178
R30476 vdd.n9646 vdd.n9630 681.178
R30477 vdd.n9646 vdd.n9627 681.178
R30478 vdd.n9661 vdd.n9627 681.178
R30479 vdd.n9661 vdd.n9628 681.178
R30480 vdd.n9657 vdd.n9628 681.178
R30481 vdd.n9691 vdd.n9690 681.178
R30482 vdd.n9692 vdd.n9691 681.178
R30483 vdd.n9692 vdd.n9670 681.178
R30484 vdd.n9711 vdd.n9670 681.178
R30485 vdd.n9711 vdd.n9671 681.178
R30486 vdd.n9702 vdd.n9671 681.178
R30487 vdd.n9684 vdd.n9678 681.178
R30488 vdd.n9694 vdd.n9678 681.178
R30489 vdd.n9694 vdd.n9675 681.178
R30490 vdd.n9709 vdd.n9675 681.178
R30491 vdd.n9709 vdd.n9676 681.178
R30492 vdd.n9705 vdd.n9676 681.178
R30493 vdd.n7088 vdd.n7076 681.178
R30494 vdd.n7092 vdd.n7076 681.178
R30495 vdd.n7092 vdd.n7072 681.178
R30496 vdd.n7072 vdd.n7070 681.178
R30497 vdd.n7105 vdd.n7070 681.178
R30498 vdd.n7106 vdd.n7105 681.178
R30499 vdd.n7085 vdd.n7081 681.178
R30500 vdd.n7081 vdd.n7075 681.178
R30501 vdd.n7075 vdd.n7073 681.178
R30502 vdd.n7095 vdd.n7073 681.178
R30503 vdd.n7095 vdd.n7068 681.178
R30504 vdd.n7109 vdd.n7068 681.178
R30505 vdd.n9790 vdd.n9789 681.178
R30506 vdd.n9791 vdd.n9790 681.178
R30507 vdd.n9791 vdd.n9769 681.178
R30508 vdd.n9810 vdd.n9769 681.178
R30509 vdd.n9810 vdd.n9770 681.178
R30510 vdd.n9801 vdd.n9770 681.178
R30511 vdd.n9783 vdd.n9777 681.178
R30512 vdd.n9793 vdd.n9777 681.178
R30513 vdd.n9793 vdd.n9774 681.178
R30514 vdd.n9808 vdd.n9774 681.178
R30515 vdd.n9808 vdd.n9775 681.178
R30516 vdd.n9804 vdd.n9775 681.178
R30517 vdd.n9742 vdd.n9741 681.178
R30518 vdd.n9743 vdd.n9742 681.178
R30519 vdd.n9743 vdd.n9721 681.178
R30520 vdd.n9762 vdd.n9721 681.178
R30521 vdd.n9762 vdd.n9722 681.178
R30522 vdd.n9753 vdd.n9722 681.178
R30523 vdd.n9735 vdd.n9729 681.178
R30524 vdd.n9745 vdd.n9729 681.178
R30525 vdd.n9745 vdd.n9726 681.178
R30526 vdd.n9760 vdd.n9726 681.178
R30527 vdd.n9760 vdd.n9727 681.178
R30528 vdd.n9756 vdd.n9727 681.178
R30529 vdd.n9839 vdd.n9838 681.178
R30530 vdd.n9840 vdd.n9839 681.178
R30531 vdd.n9840 vdd.n9818 681.178
R30532 vdd.n9859 vdd.n9818 681.178
R30533 vdd.n9859 vdd.n9819 681.178
R30534 vdd.n9850 vdd.n9819 681.178
R30535 vdd.n9832 vdd.n9826 681.178
R30536 vdd.n9842 vdd.n9826 681.178
R30537 vdd.n9842 vdd.n9823 681.178
R30538 vdd.n9857 vdd.n9823 681.178
R30539 vdd.n9857 vdd.n9824 681.178
R30540 vdd.n9853 vdd.n9824 681.178
R30541 vdd.n9889 vdd.n9888 681.178
R30542 vdd.n9890 vdd.n9889 681.178
R30543 vdd.n9890 vdd.n9868 681.178
R30544 vdd.n9909 vdd.n9868 681.178
R30545 vdd.n9909 vdd.n9869 681.178
R30546 vdd.n9900 vdd.n9869 681.178
R30547 vdd.n9882 vdd.n9876 681.178
R30548 vdd.n9892 vdd.n9876 681.178
R30549 vdd.n9892 vdd.n9873 681.178
R30550 vdd.n9907 vdd.n9873 681.178
R30551 vdd.n9907 vdd.n9874 681.178
R30552 vdd.n9903 vdd.n9874 681.178
R30553 vdd.n9937 vdd.n9936 681.178
R30554 vdd.n9938 vdd.n9937 681.178
R30555 vdd.n9938 vdd.n9916 681.178
R30556 vdd.n9957 vdd.n9916 681.178
R30557 vdd.n9957 vdd.n9917 681.178
R30558 vdd.n9948 vdd.n9917 681.178
R30559 vdd.n9930 vdd.n9924 681.178
R30560 vdd.n9940 vdd.n9924 681.178
R30561 vdd.n9940 vdd.n9921 681.178
R30562 vdd.n9955 vdd.n9921 681.178
R30563 vdd.n9955 vdd.n9922 681.178
R30564 vdd.n9951 vdd.n9922 681.178
R30565 vdd.n3849 vdd.n3848 681.178
R30566 vdd.n3850 vdd.n3849 681.178
R30567 vdd.n3850 vdd.n3828 681.178
R30568 vdd.n3869 vdd.n3828 681.178
R30569 vdd.n3869 vdd.n3829 681.178
R30570 vdd.n3860 vdd.n3829 681.178
R30571 vdd.n3842 vdd.n3836 681.178
R30572 vdd.n3852 vdd.n3836 681.178
R30573 vdd.n3852 vdd.n3833 681.178
R30574 vdd.n3867 vdd.n3833 681.178
R30575 vdd.n3867 vdd.n3834 681.178
R30576 vdd.n3863 vdd.n3834 681.178
R30577 vdd.n3897 vdd.n3896 681.178
R30578 vdd.n3898 vdd.n3897 681.178
R30579 vdd.n3898 vdd.n3876 681.178
R30580 vdd.n3917 vdd.n3876 681.178
R30581 vdd.n3917 vdd.n3877 681.178
R30582 vdd.n3908 vdd.n3877 681.178
R30583 vdd.n3890 vdd.n3884 681.178
R30584 vdd.n3900 vdd.n3884 681.178
R30585 vdd.n3900 vdd.n3881 681.178
R30586 vdd.n3915 vdd.n3881 681.178
R30587 vdd.n3915 vdd.n3882 681.178
R30588 vdd.n3911 vdd.n3882 681.178
R30589 vdd.n3999 vdd.n3998 681.178
R30590 vdd.n4000 vdd.n3999 681.178
R30591 vdd.n4000 vdd.n3978 681.178
R30592 vdd.n4019 vdd.n3978 681.178
R30593 vdd.n4019 vdd.n3979 681.178
R30594 vdd.n4010 vdd.n3979 681.178
R30595 vdd.n3992 vdd.n3986 681.178
R30596 vdd.n4002 vdd.n3986 681.178
R30597 vdd.n4002 vdd.n3983 681.178
R30598 vdd.n4017 vdd.n3983 681.178
R30599 vdd.n4017 vdd.n3984 681.178
R30600 vdd.n4013 vdd.n3984 681.178
R30601 vdd.n4047 vdd.n4046 681.178
R30602 vdd.n4048 vdd.n4047 681.178
R30603 vdd.n4048 vdd.n4026 681.178
R30604 vdd.n4067 vdd.n4026 681.178
R30605 vdd.n4067 vdd.n4027 681.178
R30606 vdd.n4058 vdd.n4027 681.178
R30607 vdd.n4040 vdd.n4034 681.178
R30608 vdd.n4050 vdd.n4034 681.178
R30609 vdd.n4050 vdd.n4031 681.178
R30610 vdd.n4065 vdd.n4031 681.178
R30611 vdd.n4065 vdd.n4032 681.178
R30612 vdd.n4061 vdd.n4032 681.178
R30613 vdd.n4095 vdd.n4094 681.178
R30614 vdd.n4096 vdd.n4095 681.178
R30615 vdd.n4096 vdd.n4074 681.178
R30616 vdd.n4115 vdd.n4074 681.178
R30617 vdd.n4115 vdd.n4075 681.178
R30618 vdd.n4106 vdd.n4075 681.178
R30619 vdd.n4088 vdd.n4082 681.178
R30620 vdd.n4098 vdd.n4082 681.178
R30621 vdd.n4098 vdd.n4079 681.178
R30622 vdd.n4113 vdd.n4079 681.178
R30623 vdd.n4113 vdd.n4080 681.178
R30624 vdd.n4109 vdd.n4080 681.178
R30625 vdd.n4143 vdd.n4142 681.178
R30626 vdd.n4144 vdd.n4143 681.178
R30627 vdd.n4144 vdd.n4122 681.178
R30628 vdd.n4163 vdd.n4122 681.178
R30629 vdd.n4163 vdd.n4123 681.178
R30630 vdd.n4154 vdd.n4123 681.178
R30631 vdd.n4136 vdd.n4130 681.178
R30632 vdd.n4146 vdd.n4130 681.178
R30633 vdd.n4146 vdd.n4127 681.178
R30634 vdd.n4161 vdd.n4127 681.178
R30635 vdd.n4161 vdd.n4128 681.178
R30636 vdd.n4157 vdd.n4128 681.178
R30637 vdd.n4245 vdd.n4244 681.178
R30638 vdd.n4246 vdd.n4245 681.178
R30639 vdd.n4246 vdd.n4224 681.178
R30640 vdd.n4265 vdd.n4224 681.178
R30641 vdd.n4265 vdd.n4225 681.178
R30642 vdd.n4256 vdd.n4225 681.178
R30643 vdd.n4238 vdd.n4232 681.178
R30644 vdd.n4248 vdd.n4232 681.178
R30645 vdd.n4248 vdd.n4229 681.178
R30646 vdd.n4263 vdd.n4229 681.178
R30647 vdd.n4263 vdd.n4230 681.178
R30648 vdd.n4259 vdd.n4230 681.178
R30649 vdd.n5765 vdd.n5764 681.178
R30650 vdd.n5766 vdd.n5765 681.178
R30651 vdd.n5766 vdd.n5744 681.178
R30652 vdd.n5785 vdd.n5744 681.178
R30653 vdd.n5785 vdd.n5745 681.178
R30654 vdd.n5776 vdd.n5745 681.178
R30655 vdd.n5758 vdd.n5752 681.178
R30656 vdd.n5768 vdd.n5752 681.178
R30657 vdd.n5768 vdd.n5749 681.178
R30658 vdd.n5783 vdd.n5749 681.178
R30659 vdd.n5783 vdd.n5750 681.178
R30660 vdd.n5779 vdd.n5750 681.178
R30661 vdd.n4289 vdd.n4280 681.178
R30662 vdd.n4296 vdd.n4280 681.178
R30663 vdd.n4296 vdd.n4277 681.178
R30664 vdd.n4311 vdd.n4277 681.178
R30665 vdd.n4311 vdd.n4278 681.178
R30666 vdd.n4307 vdd.n4278 681.178
R30667 vdd.n4293 vdd.n4292 681.178
R30668 vdd.n4294 vdd.n4293 681.178
R30669 vdd.n4294 vdd.n4272 681.178
R30670 vdd.n4313 vdd.n4272 681.178
R30671 vdd.n4313 vdd.n4273 681.178
R30672 vdd.n4304 vdd.n4273 681.178
R30673 vdd.n4337 vdd.n4328 681.178
R30674 vdd.n4344 vdd.n4328 681.178
R30675 vdd.n4344 vdd.n4325 681.178
R30676 vdd.n4359 vdd.n4325 681.178
R30677 vdd.n4359 vdd.n4326 681.178
R30678 vdd.n4355 vdd.n4326 681.178
R30679 vdd.n4341 vdd.n4340 681.178
R30680 vdd.n4342 vdd.n4341 681.178
R30681 vdd.n4342 vdd.n4320 681.178
R30682 vdd.n4361 vdd.n4320 681.178
R30683 vdd.n4361 vdd.n4321 681.178
R30684 vdd.n4352 vdd.n4321 681.178
R30685 vdd.n4438 vdd.n4429 681.178
R30686 vdd.n4445 vdd.n4429 681.178
R30687 vdd.n4445 vdd.n4426 681.178
R30688 vdd.n4460 vdd.n4426 681.178
R30689 vdd.n4460 vdd.n4427 681.178
R30690 vdd.n4456 vdd.n4427 681.178
R30691 vdd.n4442 vdd.n4441 681.178
R30692 vdd.n4443 vdd.n4442 681.178
R30693 vdd.n4443 vdd.n4421 681.178
R30694 vdd.n4462 vdd.n4421 681.178
R30695 vdd.n4462 vdd.n4422 681.178
R30696 vdd.n4453 vdd.n4422 681.178
R30697 vdd.n4486 vdd.n4477 681.178
R30698 vdd.n4493 vdd.n4477 681.178
R30699 vdd.n4493 vdd.n4474 681.178
R30700 vdd.n4508 vdd.n4474 681.178
R30701 vdd.n4508 vdd.n4475 681.178
R30702 vdd.n4504 vdd.n4475 681.178
R30703 vdd.n4490 vdd.n4489 681.178
R30704 vdd.n4491 vdd.n4490 681.178
R30705 vdd.n4491 vdd.n4469 681.178
R30706 vdd.n4510 vdd.n4469 681.178
R30707 vdd.n4510 vdd.n4470 681.178
R30708 vdd.n4501 vdd.n4470 681.178
R30709 vdd.n4534 vdd.n4525 681.178
R30710 vdd.n4541 vdd.n4525 681.178
R30711 vdd.n4541 vdd.n4522 681.178
R30712 vdd.n4556 vdd.n4522 681.178
R30713 vdd.n4556 vdd.n4523 681.178
R30714 vdd.n4552 vdd.n4523 681.178
R30715 vdd.n4538 vdd.n4537 681.178
R30716 vdd.n4539 vdd.n4538 681.178
R30717 vdd.n4539 vdd.n4517 681.178
R30718 vdd.n4558 vdd.n4517 681.178
R30719 vdd.n4558 vdd.n4518 681.178
R30720 vdd.n4549 vdd.n4518 681.178
R30721 vdd.n4582 vdd.n4573 681.178
R30722 vdd.n4589 vdd.n4573 681.178
R30723 vdd.n4589 vdd.n4570 681.178
R30724 vdd.n4604 vdd.n4570 681.178
R30725 vdd.n4604 vdd.n4571 681.178
R30726 vdd.n4600 vdd.n4571 681.178
R30727 vdd.n4586 vdd.n4585 681.178
R30728 vdd.n4587 vdd.n4586 681.178
R30729 vdd.n4587 vdd.n4565 681.178
R30730 vdd.n4606 vdd.n4565 681.178
R30731 vdd.n4606 vdd.n4566 681.178
R30732 vdd.n4597 vdd.n4566 681.178
R30733 vdd.n4683 vdd.n4674 681.178
R30734 vdd.n4690 vdd.n4674 681.178
R30735 vdd.n4690 vdd.n4671 681.178
R30736 vdd.n4705 vdd.n4671 681.178
R30737 vdd.n4705 vdd.n4672 681.178
R30738 vdd.n4701 vdd.n4672 681.178
R30739 vdd.n4687 vdd.n4686 681.178
R30740 vdd.n4688 vdd.n4687 681.178
R30741 vdd.n4688 vdd.n4666 681.178
R30742 vdd.n4707 vdd.n4666 681.178
R30743 vdd.n4707 vdd.n4667 681.178
R30744 vdd.n4698 vdd.n4667 681.178
R30745 vdd.n3796 vdd.n3787 681.178
R30746 vdd.n3803 vdd.n3787 681.178
R30747 vdd.n3803 vdd.n3784 681.178
R30748 vdd.n3818 vdd.n3784 681.178
R30749 vdd.n3818 vdd.n3785 681.178
R30750 vdd.n3814 vdd.n3785 681.178
R30751 vdd.n3800 vdd.n3799 681.178
R30752 vdd.n3801 vdd.n3800 681.178
R30753 vdd.n3801 vdd.n3779 681.178
R30754 vdd.n3820 vdd.n3779 681.178
R30755 vdd.n3820 vdd.n3780 681.178
R30756 vdd.n3811 vdd.n3780 681.178
R30757 vdd.n4731 vdd.n4722 681.178
R30758 vdd.n4738 vdd.n4722 681.178
R30759 vdd.n4738 vdd.n4719 681.178
R30760 vdd.n4753 vdd.n4719 681.178
R30761 vdd.n4753 vdd.n4720 681.178
R30762 vdd.n4749 vdd.n4720 681.178
R30763 vdd.n4735 vdd.n4734 681.178
R30764 vdd.n4736 vdd.n4735 681.178
R30765 vdd.n4736 vdd.n4714 681.178
R30766 vdd.n4755 vdd.n4714 681.178
R30767 vdd.n4755 vdd.n4715 681.178
R30768 vdd.n4746 vdd.n4715 681.178
R30769 vdd.n4778 vdd.n4769 681.178
R30770 vdd.n4785 vdd.n4769 681.178
R30771 vdd.n4785 vdd.n4766 681.178
R30772 vdd.n4800 vdd.n4766 681.178
R30773 vdd.n4800 vdd.n4767 681.178
R30774 vdd.n4796 vdd.n4767 681.178
R30775 vdd.n4782 vdd.n4781 681.178
R30776 vdd.n4783 vdd.n4782 681.178
R30777 vdd.n4783 vdd.n4761 681.178
R30778 vdd.n4802 vdd.n4761 681.178
R30779 vdd.n4802 vdd.n4762 681.178
R30780 vdd.n4793 vdd.n4762 681.178
R30781 vdd.n4828 vdd.n4819 681.178
R30782 vdd.n4835 vdd.n4819 681.178
R30783 vdd.n4835 vdd.n4816 681.178
R30784 vdd.n4850 vdd.n4816 681.178
R30785 vdd.n4850 vdd.n4817 681.178
R30786 vdd.n4846 vdd.n4817 681.178
R30787 vdd.n4832 vdd.n4831 681.178
R30788 vdd.n4833 vdd.n4832 681.178
R30789 vdd.n4833 vdd.n4811 681.178
R30790 vdd.n4852 vdd.n4811 681.178
R30791 vdd.n4852 vdd.n4812 681.178
R30792 vdd.n4843 vdd.n4812 681.178
R30793 vdd.n4878 vdd.n4869 681.178
R30794 vdd.n4885 vdd.n4869 681.178
R30795 vdd.n4885 vdd.n4866 681.178
R30796 vdd.n4900 vdd.n4866 681.178
R30797 vdd.n4900 vdd.n4867 681.178
R30798 vdd.n4896 vdd.n4867 681.178
R30799 vdd.n4882 vdd.n4881 681.178
R30800 vdd.n4883 vdd.n4882 681.178
R30801 vdd.n4883 vdd.n4861 681.178
R30802 vdd.n4902 vdd.n4861 681.178
R30803 vdd.n4902 vdd.n4862 681.178
R30804 vdd.n4893 vdd.n4862 681.178
R30805 vdd.n4926 vdd.n4917 681.178
R30806 vdd.n4933 vdd.n4917 681.178
R30807 vdd.n4933 vdd.n4914 681.178
R30808 vdd.n4948 vdd.n4914 681.178
R30809 vdd.n4948 vdd.n4915 681.178
R30810 vdd.n4944 vdd.n4915 681.178
R30811 vdd.n4930 vdd.n4929 681.178
R30812 vdd.n4931 vdd.n4930 681.178
R30813 vdd.n4931 vdd.n4909 681.178
R30814 vdd.n4950 vdd.n4909 681.178
R30815 vdd.n4950 vdd.n4910 681.178
R30816 vdd.n4941 vdd.n4910 681.178
R30817 vdd.n4654 vdd.n4617 681.178
R30818 vdd.n4650 vdd.n4617 681.178
R30819 vdd.n4650 vdd.n4621 681.178
R30820 vdd.n4640 vdd.n4621 681.178
R30821 vdd.n4640 vdd.n4626 681.178
R30822 vdd.n4636 vdd.n4626 681.178
R30823 vdd.n4657 vdd.n4615 681.178
R30824 vdd.n4648 vdd.n4615 681.178
R30825 vdd.n4648 vdd.n4643 681.178
R30826 vdd.n4643 vdd.n4642 681.178
R30827 vdd.n4642 vdd.n4623 681.178
R30828 vdd.n4633 vdd.n4623 681.178
R30829 vdd.n4977 vdd.n4968 681.178
R30830 vdd.n4984 vdd.n4968 681.178
R30831 vdd.n4984 vdd.n4965 681.178
R30832 vdd.n4999 vdd.n4965 681.178
R30833 vdd.n4999 vdd.n4966 681.178
R30834 vdd.n4995 vdd.n4966 681.178
R30835 vdd.n4981 vdd.n4980 681.178
R30836 vdd.n4982 vdd.n4981 681.178
R30837 vdd.n4982 vdd.n4960 681.178
R30838 vdd.n5001 vdd.n4960 681.178
R30839 vdd.n5001 vdd.n4961 681.178
R30840 vdd.n4992 vdd.n4961 681.178
R30841 vdd.n5024 vdd.n5015 681.178
R30842 vdd.n5031 vdd.n5015 681.178
R30843 vdd.n5031 vdd.n5012 681.178
R30844 vdd.n5046 vdd.n5012 681.178
R30845 vdd.n5046 vdd.n5013 681.178
R30846 vdd.n5042 vdd.n5013 681.178
R30847 vdd.n5028 vdd.n5027 681.178
R30848 vdd.n5029 vdd.n5028 681.178
R30849 vdd.n5029 vdd.n5007 681.178
R30850 vdd.n5048 vdd.n5007 681.178
R30851 vdd.n5048 vdd.n5008 681.178
R30852 vdd.n5039 vdd.n5008 681.178
R30853 vdd.n5072 vdd.n5063 681.178
R30854 vdd.n5079 vdd.n5063 681.178
R30855 vdd.n5079 vdd.n5060 681.178
R30856 vdd.n5094 vdd.n5060 681.178
R30857 vdd.n5094 vdd.n5061 681.178
R30858 vdd.n5090 vdd.n5061 681.178
R30859 vdd.n5076 vdd.n5075 681.178
R30860 vdd.n5077 vdd.n5076 681.178
R30861 vdd.n5077 vdd.n5055 681.178
R30862 vdd.n5096 vdd.n5055 681.178
R30863 vdd.n5096 vdd.n5056 681.178
R30864 vdd.n5087 vdd.n5056 681.178
R30865 vdd.n5123 vdd.n5114 681.178
R30866 vdd.n5130 vdd.n5114 681.178
R30867 vdd.n5130 vdd.n5111 681.178
R30868 vdd.n5145 vdd.n5111 681.178
R30869 vdd.n5145 vdd.n5112 681.178
R30870 vdd.n5141 vdd.n5112 681.178
R30871 vdd.n5127 vdd.n5126 681.178
R30872 vdd.n5128 vdd.n5127 681.178
R30873 vdd.n5128 vdd.n5106 681.178
R30874 vdd.n5147 vdd.n5106 681.178
R30875 vdd.n5147 vdd.n5107 681.178
R30876 vdd.n5138 vdd.n5107 681.178
R30877 vdd.n5173 vdd.n5164 681.178
R30878 vdd.n5180 vdd.n5164 681.178
R30879 vdd.n5180 vdd.n5161 681.178
R30880 vdd.n5195 vdd.n5161 681.178
R30881 vdd.n5195 vdd.n5162 681.178
R30882 vdd.n5191 vdd.n5162 681.178
R30883 vdd.n5177 vdd.n5176 681.178
R30884 vdd.n5178 vdd.n5177 681.178
R30885 vdd.n5178 vdd.n5156 681.178
R30886 vdd.n5197 vdd.n5156 681.178
R30887 vdd.n5197 vdd.n5157 681.178
R30888 vdd.n5188 vdd.n5157 681.178
R30889 vdd.n5221 vdd.n5212 681.178
R30890 vdd.n5228 vdd.n5212 681.178
R30891 vdd.n5228 vdd.n5209 681.178
R30892 vdd.n5243 vdd.n5209 681.178
R30893 vdd.n5243 vdd.n5210 681.178
R30894 vdd.n5239 vdd.n5210 681.178
R30895 vdd.n5225 vdd.n5224 681.178
R30896 vdd.n5226 vdd.n5225 681.178
R30897 vdd.n5226 vdd.n5204 681.178
R30898 vdd.n5245 vdd.n5204 681.178
R30899 vdd.n5245 vdd.n5205 681.178
R30900 vdd.n5236 vdd.n5205 681.178
R30901 vdd.n5271 vdd.n5262 681.178
R30902 vdd.n5278 vdd.n5262 681.178
R30903 vdd.n5278 vdd.n5259 681.178
R30904 vdd.n5293 vdd.n5259 681.178
R30905 vdd.n5293 vdd.n5260 681.178
R30906 vdd.n5289 vdd.n5260 681.178
R30907 vdd.n5275 vdd.n5274 681.178
R30908 vdd.n5276 vdd.n5275 681.178
R30909 vdd.n5276 vdd.n5254 681.178
R30910 vdd.n5295 vdd.n5254 681.178
R30911 vdd.n5295 vdd.n5255 681.178
R30912 vdd.n5286 vdd.n5255 681.178
R30913 vdd.n5318 vdd.n5309 681.178
R30914 vdd.n5325 vdd.n5309 681.178
R30915 vdd.n5325 vdd.n5306 681.178
R30916 vdd.n5340 vdd.n5306 681.178
R30917 vdd.n5340 vdd.n5307 681.178
R30918 vdd.n5336 vdd.n5307 681.178
R30919 vdd.n5322 vdd.n5321 681.178
R30920 vdd.n5323 vdd.n5322 681.178
R30921 vdd.n5323 vdd.n5301 681.178
R30922 vdd.n5342 vdd.n5301 681.178
R30923 vdd.n5342 vdd.n5302 681.178
R30924 vdd.n5333 vdd.n5302 681.178
R30925 vdd.n5368 vdd.n5359 681.178
R30926 vdd.n5375 vdd.n5359 681.178
R30927 vdd.n5375 vdd.n5356 681.178
R30928 vdd.n5390 vdd.n5356 681.178
R30929 vdd.n5390 vdd.n5357 681.178
R30930 vdd.n5386 vdd.n5357 681.178
R30931 vdd.n5372 vdd.n5371 681.178
R30932 vdd.n5373 vdd.n5372 681.178
R30933 vdd.n5373 vdd.n5351 681.178
R30934 vdd.n5392 vdd.n5351 681.178
R30935 vdd.n5392 vdd.n5352 681.178
R30936 vdd.n5383 vdd.n5352 681.178
R30937 vdd.n5418 vdd.n5409 681.178
R30938 vdd.n5425 vdd.n5409 681.178
R30939 vdd.n5425 vdd.n5406 681.178
R30940 vdd.n5440 vdd.n5406 681.178
R30941 vdd.n5440 vdd.n5407 681.178
R30942 vdd.n5436 vdd.n5407 681.178
R30943 vdd.n5422 vdd.n5421 681.178
R30944 vdd.n5423 vdd.n5422 681.178
R30945 vdd.n5423 vdd.n5401 681.178
R30946 vdd.n5442 vdd.n5401 681.178
R30947 vdd.n5442 vdd.n5402 681.178
R30948 vdd.n5433 vdd.n5402 681.178
R30949 vdd.n5466 vdd.n5457 681.178
R30950 vdd.n5473 vdd.n5457 681.178
R30951 vdd.n5473 vdd.n5454 681.178
R30952 vdd.n5488 vdd.n5454 681.178
R30953 vdd.n5488 vdd.n5455 681.178
R30954 vdd.n5484 vdd.n5455 681.178
R30955 vdd.n5470 vdd.n5469 681.178
R30956 vdd.n5471 vdd.n5470 681.178
R30957 vdd.n5471 vdd.n5449 681.178
R30958 vdd.n5490 vdd.n5449 681.178
R30959 vdd.n5490 vdd.n5450 681.178
R30960 vdd.n5481 vdd.n5450 681.178
R30961 vdd.n4409 vdd.n4372 681.178
R30962 vdd.n4405 vdd.n4372 681.178
R30963 vdd.n4405 vdd.n4376 681.178
R30964 vdd.n4395 vdd.n4376 681.178
R30965 vdd.n4395 vdd.n4381 681.178
R30966 vdd.n4391 vdd.n4381 681.178
R30967 vdd.n4412 vdd.n4370 681.178
R30968 vdd.n4403 vdd.n4370 681.178
R30969 vdd.n4403 vdd.n4398 681.178
R30970 vdd.n4398 vdd.n4397 681.178
R30971 vdd.n4397 vdd.n4378 681.178
R30972 vdd.n4388 vdd.n4378 681.178
R30973 vdd.n5517 vdd.n5508 681.178
R30974 vdd.n5524 vdd.n5508 681.178
R30975 vdd.n5524 vdd.n5505 681.178
R30976 vdd.n5539 vdd.n5505 681.178
R30977 vdd.n5539 vdd.n5506 681.178
R30978 vdd.n5535 vdd.n5506 681.178
R30979 vdd.n5521 vdd.n5520 681.178
R30980 vdd.n5522 vdd.n5521 681.178
R30981 vdd.n5522 vdd.n5500 681.178
R30982 vdd.n5541 vdd.n5500 681.178
R30983 vdd.n5541 vdd.n5501 681.178
R30984 vdd.n5532 vdd.n5501 681.178
R30985 vdd.n5564 vdd.n5555 681.178
R30986 vdd.n5571 vdd.n5555 681.178
R30987 vdd.n5571 vdd.n5552 681.178
R30988 vdd.n5586 vdd.n5552 681.178
R30989 vdd.n5586 vdd.n5553 681.178
R30990 vdd.n5582 vdd.n5553 681.178
R30991 vdd.n5568 vdd.n5567 681.178
R30992 vdd.n5569 vdd.n5568 681.178
R30993 vdd.n5569 vdd.n5547 681.178
R30994 vdd.n5588 vdd.n5547 681.178
R30995 vdd.n5588 vdd.n5548 681.178
R30996 vdd.n5579 vdd.n5548 681.178
R30997 vdd.n5614 vdd.n5605 681.178
R30998 vdd.n5621 vdd.n5605 681.178
R30999 vdd.n5621 vdd.n5602 681.178
R31000 vdd.n5636 vdd.n5602 681.178
R31001 vdd.n5636 vdd.n5603 681.178
R31002 vdd.n5632 vdd.n5603 681.178
R31003 vdd.n5618 vdd.n5617 681.178
R31004 vdd.n5619 vdd.n5618 681.178
R31005 vdd.n5619 vdd.n5597 681.178
R31006 vdd.n5638 vdd.n5597 681.178
R31007 vdd.n5638 vdd.n5598 681.178
R31008 vdd.n5629 vdd.n5598 681.178
R31009 vdd.n5664 vdd.n5655 681.178
R31010 vdd.n5671 vdd.n5655 681.178
R31011 vdd.n5671 vdd.n5652 681.178
R31012 vdd.n5686 vdd.n5652 681.178
R31013 vdd.n5686 vdd.n5653 681.178
R31014 vdd.n5682 vdd.n5653 681.178
R31015 vdd.n5668 vdd.n5667 681.178
R31016 vdd.n5669 vdd.n5668 681.178
R31017 vdd.n5669 vdd.n5647 681.178
R31018 vdd.n5688 vdd.n5647 681.178
R31019 vdd.n5688 vdd.n5648 681.178
R31020 vdd.n5679 vdd.n5648 681.178
R31021 vdd.n5712 vdd.n5703 681.178
R31022 vdd.n5719 vdd.n5703 681.178
R31023 vdd.n5719 vdd.n5700 681.178
R31024 vdd.n5734 vdd.n5700 681.178
R31025 vdd.n5734 vdd.n5701 681.178
R31026 vdd.n5730 vdd.n5701 681.178
R31027 vdd.n5716 vdd.n5715 681.178
R31028 vdd.n5717 vdd.n5716 681.178
R31029 vdd.n5717 vdd.n5695 681.178
R31030 vdd.n5736 vdd.n5695 681.178
R31031 vdd.n5736 vdd.n5696 681.178
R31032 vdd.n5727 vdd.n5696 681.178
R31033 vdd.n5862 vdd.n5861 681.178
R31034 vdd.n5863 vdd.n5862 681.178
R31035 vdd.n5863 vdd.n5841 681.178
R31036 vdd.n5882 vdd.n5841 681.178
R31037 vdd.n5882 vdd.n5842 681.178
R31038 vdd.n5873 vdd.n5842 681.178
R31039 vdd.n5855 vdd.n5849 681.178
R31040 vdd.n5865 vdd.n5849 681.178
R31041 vdd.n5865 vdd.n5846 681.178
R31042 vdd.n5880 vdd.n5846 681.178
R31043 vdd.n5880 vdd.n5847 681.178
R31044 vdd.n5876 vdd.n5847 681.178
R31045 vdd.n5814 vdd.n5813 681.178
R31046 vdd.n5815 vdd.n5814 681.178
R31047 vdd.n5815 vdd.n5793 681.178
R31048 vdd.n5834 vdd.n5793 681.178
R31049 vdd.n5834 vdd.n5794 681.178
R31050 vdd.n5825 vdd.n5794 681.178
R31051 vdd.n5807 vdd.n5801 681.178
R31052 vdd.n5817 vdd.n5801 681.178
R31053 vdd.n5817 vdd.n5798 681.178
R31054 vdd.n5832 vdd.n5798 681.178
R31055 vdd.n5832 vdd.n5799 681.178
R31056 vdd.n5828 vdd.n5799 681.178
R31057 vdd.n5911 vdd.n5910 681.178
R31058 vdd.n5912 vdd.n5911 681.178
R31059 vdd.n5912 vdd.n5890 681.178
R31060 vdd.n5931 vdd.n5890 681.178
R31061 vdd.n5931 vdd.n5891 681.178
R31062 vdd.n5922 vdd.n5891 681.178
R31063 vdd.n5904 vdd.n5898 681.178
R31064 vdd.n5914 vdd.n5898 681.178
R31065 vdd.n5914 vdd.n5895 681.178
R31066 vdd.n5929 vdd.n5895 681.178
R31067 vdd.n5929 vdd.n5896 681.178
R31068 vdd.n5925 vdd.n5896 681.178
R31069 vdd.n5961 vdd.n5960 681.178
R31070 vdd.n5962 vdd.n5961 681.178
R31071 vdd.n5962 vdd.n5940 681.178
R31072 vdd.n5981 vdd.n5940 681.178
R31073 vdd.n5981 vdd.n5941 681.178
R31074 vdd.n5972 vdd.n5941 681.178
R31075 vdd.n5954 vdd.n5948 681.178
R31076 vdd.n5964 vdd.n5948 681.178
R31077 vdd.n5964 vdd.n5945 681.178
R31078 vdd.n5979 vdd.n5945 681.178
R31079 vdd.n5979 vdd.n5946 681.178
R31080 vdd.n5975 vdd.n5946 681.178
R31081 vdd.n6009 vdd.n6008 681.178
R31082 vdd.n6010 vdd.n6009 681.178
R31083 vdd.n6010 vdd.n5988 681.178
R31084 vdd.n6029 vdd.n5988 681.178
R31085 vdd.n6029 vdd.n5989 681.178
R31086 vdd.n6020 vdd.n5989 681.178
R31087 vdd.n6002 vdd.n5996 681.178
R31088 vdd.n6012 vdd.n5996 681.178
R31089 vdd.n6012 vdd.n5993 681.178
R31090 vdd.n6027 vdd.n5993 681.178
R31091 vdd.n6027 vdd.n5994 681.178
R31092 vdd.n6023 vdd.n5994 681.178
R31093 vdd.n4192 vdd.n4180 681.178
R31094 vdd.n4196 vdd.n4180 681.178
R31095 vdd.n4196 vdd.n4176 681.178
R31096 vdd.n4176 vdd.n4174 681.178
R31097 vdd.n4209 vdd.n4174 681.178
R31098 vdd.n4210 vdd.n4209 681.178
R31099 vdd.n4189 vdd.n4185 681.178
R31100 vdd.n4185 vdd.n4179 681.178
R31101 vdd.n4179 vdd.n4177 681.178
R31102 vdd.n4199 vdd.n4177 681.178
R31103 vdd.n4199 vdd.n4172 681.178
R31104 vdd.n4213 vdd.n4172 681.178
R31105 vdd.n6157 vdd.n6156 681.178
R31106 vdd.n6158 vdd.n6157 681.178
R31107 vdd.n6158 vdd.n6136 681.178
R31108 vdd.n6177 vdd.n6136 681.178
R31109 vdd.n6177 vdd.n6137 681.178
R31110 vdd.n6168 vdd.n6137 681.178
R31111 vdd.n6150 vdd.n6144 681.178
R31112 vdd.n6160 vdd.n6144 681.178
R31113 vdd.n6160 vdd.n6141 681.178
R31114 vdd.n6175 vdd.n6141 681.178
R31115 vdd.n6175 vdd.n6142 681.178
R31116 vdd.n6171 vdd.n6142 681.178
R31117 vdd.n6108 vdd.n6107 681.178
R31118 vdd.n6109 vdd.n6108 681.178
R31119 vdd.n6109 vdd.n6087 681.178
R31120 vdd.n6128 vdd.n6087 681.178
R31121 vdd.n6128 vdd.n6088 681.178
R31122 vdd.n6119 vdd.n6088 681.178
R31123 vdd.n6101 vdd.n6095 681.178
R31124 vdd.n6111 vdd.n6095 681.178
R31125 vdd.n6111 vdd.n6092 681.178
R31126 vdd.n6126 vdd.n6092 681.178
R31127 vdd.n6126 vdd.n6093 681.178
R31128 vdd.n6122 vdd.n6093 681.178
R31129 vdd.n6060 vdd.n6059 681.178
R31130 vdd.n6061 vdd.n6060 681.178
R31131 vdd.n6061 vdd.n6039 681.178
R31132 vdd.n6080 vdd.n6039 681.178
R31133 vdd.n6080 vdd.n6040 681.178
R31134 vdd.n6071 vdd.n6040 681.178
R31135 vdd.n6053 vdd.n6047 681.178
R31136 vdd.n6063 vdd.n6047 681.178
R31137 vdd.n6063 vdd.n6044 681.178
R31138 vdd.n6078 vdd.n6044 681.178
R31139 vdd.n6078 vdd.n6045 681.178
R31140 vdd.n6074 vdd.n6045 681.178
R31141 vdd.n6206 vdd.n6205 681.178
R31142 vdd.n6207 vdd.n6206 681.178
R31143 vdd.n6207 vdd.n6185 681.178
R31144 vdd.n6226 vdd.n6185 681.178
R31145 vdd.n6226 vdd.n6186 681.178
R31146 vdd.n6217 vdd.n6186 681.178
R31147 vdd.n6199 vdd.n6193 681.178
R31148 vdd.n6209 vdd.n6193 681.178
R31149 vdd.n6209 vdd.n6190 681.178
R31150 vdd.n6224 vdd.n6190 681.178
R31151 vdd.n6224 vdd.n6191 681.178
R31152 vdd.n6220 vdd.n6191 681.178
R31153 vdd.n6256 vdd.n6255 681.178
R31154 vdd.n6257 vdd.n6256 681.178
R31155 vdd.n6257 vdd.n6235 681.178
R31156 vdd.n6276 vdd.n6235 681.178
R31157 vdd.n6276 vdd.n6236 681.178
R31158 vdd.n6267 vdd.n6236 681.178
R31159 vdd.n6249 vdd.n6243 681.178
R31160 vdd.n6259 vdd.n6243 681.178
R31161 vdd.n6259 vdd.n6240 681.178
R31162 vdd.n6274 vdd.n6240 681.178
R31163 vdd.n6274 vdd.n6241 681.178
R31164 vdd.n6270 vdd.n6241 681.178
R31165 vdd.n6304 vdd.n6303 681.178
R31166 vdd.n6305 vdd.n6304 681.178
R31167 vdd.n6305 vdd.n6283 681.178
R31168 vdd.n6324 vdd.n6283 681.178
R31169 vdd.n6324 vdd.n6284 681.178
R31170 vdd.n6315 vdd.n6284 681.178
R31171 vdd.n6297 vdd.n6291 681.178
R31172 vdd.n6307 vdd.n6291 681.178
R31173 vdd.n6307 vdd.n6288 681.178
R31174 vdd.n6322 vdd.n6288 681.178
R31175 vdd.n6322 vdd.n6289 681.178
R31176 vdd.n6318 vdd.n6289 681.178
R31177 vdd.n6402 vdd.n6401 681.178
R31178 vdd.n6403 vdd.n6402 681.178
R31179 vdd.n6403 vdd.n6381 681.178
R31180 vdd.n6422 vdd.n6381 681.178
R31181 vdd.n6422 vdd.n6382 681.178
R31182 vdd.n6413 vdd.n6382 681.178
R31183 vdd.n6395 vdd.n6389 681.178
R31184 vdd.n6405 vdd.n6389 681.178
R31185 vdd.n6405 vdd.n6386 681.178
R31186 vdd.n6420 vdd.n6386 681.178
R31187 vdd.n6420 vdd.n6387 681.178
R31188 vdd.n6416 vdd.n6387 681.178
R31189 vdd.n6354 vdd.n6353 681.178
R31190 vdd.n6355 vdd.n6354 681.178
R31191 vdd.n6355 vdd.n6333 681.178
R31192 vdd.n6374 vdd.n6333 681.178
R31193 vdd.n6374 vdd.n6334 681.178
R31194 vdd.n6365 vdd.n6334 681.178
R31195 vdd.n6347 vdd.n6341 681.178
R31196 vdd.n6357 vdd.n6341 681.178
R31197 vdd.n6357 vdd.n6338 681.178
R31198 vdd.n6372 vdd.n6338 681.178
R31199 vdd.n6372 vdd.n6339 681.178
R31200 vdd.n6368 vdd.n6339 681.178
R31201 vdd.n6451 vdd.n6450 681.178
R31202 vdd.n6452 vdd.n6451 681.178
R31203 vdd.n6452 vdd.n6430 681.178
R31204 vdd.n6471 vdd.n6430 681.178
R31205 vdd.n6471 vdd.n6431 681.178
R31206 vdd.n6462 vdd.n6431 681.178
R31207 vdd.n6444 vdd.n6438 681.178
R31208 vdd.n6454 vdd.n6438 681.178
R31209 vdd.n6454 vdd.n6435 681.178
R31210 vdd.n6469 vdd.n6435 681.178
R31211 vdd.n6469 vdd.n6436 681.178
R31212 vdd.n6465 vdd.n6436 681.178
R31213 vdd.n6501 vdd.n6500 681.178
R31214 vdd.n6502 vdd.n6501 681.178
R31215 vdd.n6502 vdd.n6480 681.178
R31216 vdd.n6521 vdd.n6480 681.178
R31217 vdd.n6521 vdd.n6481 681.178
R31218 vdd.n6512 vdd.n6481 681.178
R31219 vdd.n6494 vdd.n6488 681.178
R31220 vdd.n6504 vdd.n6488 681.178
R31221 vdd.n6504 vdd.n6485 681.178
R31222 vdd.n6519 vdd.n6485 681.178
R31223 vdd.n6519 vdd.n6486 681.178
R31224 vdd.n6515 vdd.n6486 681.178
R31225 vdd.n6549 vdd.n6548 681.178
R31226 vdd.n6550 vdd.n6549 681.178
R31227 vdd.n6550 vdd.n6528 681.178
R31228 vdd.n6569 vdd.n6528 681.178
R31229 vdd.n6569 vdd.n6529 681.178
R31230 vdd.n6560 vdd.n6529 681.178
R31231 vdd.n6542 vdd.n6536 681.178
R31232 vdd.n6552 vdd.n6536 681.178
R31233 vdd.n6552 vdd.n6533 681.178
R31234 vdd.n6567 vdd.n6533 681.178
R31235 vdd.n6567 vdd.n6534 681.178
R31236 vdd.n6563 vdd.n6534 681.178
R31237 vdd.n3946 vdd.n3934 681.178
R31238 vdd.n3950 vdd.n3934 681.178
R31239 vdd.n3950 vdd.n3930 681.178
R31240 vdd.n3930 vdd.n3928 681.178
R31241 vdd.n3963 vdd.n3928 681.178
R31242 vdd.n3964 vdd.n3963 681.178
R31243 vdd.n3943 vdd.n3939 681.178
R31244 vdd.n3939 vdd.n3933 681.178
R31245 vdd.n3933 vdd.n3931 681.178
R31246 vdd.n3953 vdd.n3931 681.178
R31247 vdd.n3953 vdd.n3926 681.178
R31248 vdd.n3967 vdd.n3926 681.178
R31249 vdd.n6648 vdd.n6647 681.178
R31250 vdd.n6649 vdd.n6648 681.178
R31251 vdd.n6649 vdd.n6627 681.178
R31252 vdd.n6668 vdd.n6627 681.178
R31253 vdd.n6668 vdd.n6628 681.178
R31254 vdd.n6659 vdd.n6628 681.178
R31255 vdd.n6641 vdd.n6635 681.178
R31256 vdd.n6651 vdd.n6635 681.178
R31257 vdd.n6651 vdd.n6632 681.178
R31258 vdd.n6666 vdd.n6632 681.178
R31259 vdd.n6666 vdd.n6633 681.178
R31260 vdd.n6662 vdd.n6633 681.178
R31261 vdd.n6600 vdd.n6599 681.178
R31262 vdd.n6601 vdd.n6600 681.178
R31263 vdd.n6601 vdd.n6579 681.178
R31264 vdd.n6620 vdd.n6579 681.178
R31265 vdd.n6620 vdd.n6580 681.178
R31266 vdd.n6611 vdd.n6580 681.178
R31267 vdd.n6593 vdd.n6587 681.178
R31268 vdd.n6603 vdd.n6587 681.178
R31269 vdd.n6603 vdd.n6584 681.178
R31270 vdd.n6618 vdd.n6584 681.178
R31271 vdd.n6618 vdd.n6585 681.178
R31272 vdd.n6614 vdd.n6585 681.178
R31273 vdd.n6697 vdd.n6696 681.178
R31274 vdd.n6698 vdd.n6697 681.178
R31275 vdd.n6698 vdd.n6676 681.178
R31276 vdd.n6717 vdd.n6676 681.178
R31277 vdd.n6717 vdd.n6677 681.178
R31278 vdd.n6708 vdd.n6677 681.178
R31279 vdd.n6690 vdd.n6684 681.178
R31280 vdd.n6700 vdd.n6684 681.178
R31281 vdd.n6700 vdd.n6681 681.178
R31282 vdd.n6715 vdd.n6681 681.178
R31283 vdd.n6715 vdd.n6682 681.178
R31284 vdd.n6711 vdd.n6682 681.178
R31285 vdd.n6747 vdd.n6746 681.178
R31286 vdd.n6748 vdd.n6747 681.178
R31287 vdd.n6748 vdd.n6726 681.178
R31288 vdd.n6767 vdd.n6726 681.178
R31289 vdd.n6767 vdd.n6727 681.178
R31290 vdd.n6758 vdd.n6727 681.178
R31291 vdd.n6740 vdd.n6734 681.178
R31292 vdd.n6750 vdd.n6734 681.178
R31293 vdd.n6750 vdd.n6731 681.178
R31294 vdd.n6765 vdd.n6731 681.178
R31295 vdd.n6765 vdd.n6732 681.178
R31296 vdd.n6761 vdd.n6732 681.178
R31297 vdd.n6795 vdd.n6794 681.178
R31298 vdd.n6796 vdd.n6795 681.178
R31299 vdd.n6796 vdd.n6774 681.178
R31300 vdd.n6815 vdd.n6774 681.178
R31301 vdd.n6815 vdd.n6775 681.178
R31302 vdd.n6806 vdd.n6775 681.178
R31303 vdd.n6788 vdd.n6782 681.178
R31304 vdd.n6798 vdd.n6782 681.178
R31305 vdd.n6798 vdd.n6779 681.178
R31306 vdd.n6813 vdd.n6779 681.178
R31307 vdd.n6813 vdd.n6780 681.178
R31308 vdd.n6809 vdd.n6780 681.178
R31309 vdd.n707 vdd.n706 681.178
R31310 vdd.n708 vdd.n707 681.178
R31311 vdd.n708 vdd.n686 681.178
R31312 vdd.n727 vdd.n686 681.178
R31313 vdd.n727 vdd.n687 681.178
R31314 vdd.n718 vdd.n687 681.178
R31315 vdd.n700 vdd.n694 681.178
R31316 vdd.n710 vdd.n694 681.178
R31317 vdd.n710 vdd.n691 681.178
R31318 vdd.n725 vdd.n691 681.178
R31319 vdd.n725 vdd.n692 681.178
R31320 vdd.n721 vdd.n692 681.178
R31321 vdd.n755 vdd.n754 681.178
R31322 vdd.n756 vdd.n755 681.178
R31323 vdd.n756 vdd.n734 681.178
R31324 vdd.n775 vdd.n734 681.178
R31325 vdd.n775 vdd.n735 681.178
R31326 vdd.n766 vdd.n735 681.178
R31327 vdd.n748 vdd.n742 681.178
R31328 vdd.n758 vdd.n742 681.178
R31329 vdd.n758 vdd.n739 681.178
R31330 vdd.n773 vdd.n739 681.178
R31331 vdd.n773 vdd.n740 681.178
R31332 vdd.n769 vdd.n740 681.178
R31333 vdd.n857 vdd.n856 681.178
R31334 vdd.n858 vdd.n857 681.178
R31335 vdd.n858 vdd.n836 681.178
R31336 vdd.n877 vdd.n836 681.178
R31337 vdd.n877 vdd.n837 681.178
R31338 vdd.n868 vdd.n837 681.178
R31339 vdd.n850 vdd.n844 681.178
R31340 vdd.n860 vdd.n844 681.178
R31341 vdd.n860 vdd.n841 681.178
R31342 vdd.n875 vdd.n841 681.178
R31343 vdd.n875 vdd.n842 681.178
R31344 vdd.n871 vdd.n842 681.178
R31345 vdd.n905 vdd.n904 681.178
R31346 vdd.n906 vdd.n905 681.178
R31347 vdd.n906 vdd.n884 681.178
R31348 vdd.n925 vdd.n884 681.178
R31349 vdd.n925 vdd.n885 681.178
R31350 vdd.n916 vdd.n885 681.178
R31351 vdd.n898 vdd.n892 681.178
R31352 vdd.n908 vdd.n892 681.178
R31353 vdd.n908 vdd.n889 681.178
R31354 vdd.n923 vdd.n889 681.178
R31355 vdd.n923 vdd.n890 681.178
R31356 vdd.n919 vdd.n890 681.178
R31357 vdd.n953 vdd.n952 681.178
R31358 vdd.n954 vdd.n953 681.178
R31359 vdd.n954 vdd.n932 681.178
R31360 vdd.n973 vdd.n932 681.178
R31361 vdd.n973 vdd.n933 681.178
R31362 vdd.n964 vdd.n933 681.178
R31363 vdd.n946 vdd.n940 681.178
R31364 vdd.n956 vdd.n940 681.178
R31365 vdd.n956 vdd.n937 681.178
R31366 vdd.n971 vdd.n937 681.178
R31367 vdd.n971 vdd.n938 681.178
R31368 vdd.n967 vdd.n938 681.178
R31369 vdd.n1001 vdd.n1000 681.178
R31370 vdd.n1002 vdd.n1001 681.178
R31371 vdd.n1002 vdd.n980 681.178
R31372 vdd.n1021 vdd.n980 681.178
R31373 vdd.n1021 vdd.n981 681.178
R31374 vdd.n1012 vdd.n981 681.178
R31375 vdd.n994 vdd.n988 681.178
R31376 vdd.n1004 vdd.n988 681.178
R31377 vdd.n1004 vdd.n985 681.178
R31378 vdd.n1019 vdd.n985 681.178
R31379 vdd.n1019 vdd.n986 681.178
R31380 vdd.n1015 vdd.n986 681.178
R31381 vdd.n1103 vdd.n1102 681.178
R31382 vdd.n1104 vdd.n1103 681.178
R31383 vdd.n1104 vdd.n1082 681.178
R31384 vdd.n1123 vdd.n1082 681.178
R31385 vdd.n1123 vdd.n1083 681.178
R31386 vdd.n1114 vdd.n1083 681.178
R31387 vdd.n1096 vdd.n1090 681.178
R31388 vdd.n1106 vdd.n1090 681.178
R31389 vdd.n1106 vdd.n1087 681.178
R31390 vdd.n1121 vdd.n1087 681.178
R31391 vdd.n1121 vdd.n1088 681.178
R31392 vdd.n1117 vdd.n1088 681.178
R31393 vdd.n2623 vdd.n2622 681.178
R31394 vdd.n2624 vdd.n2623 681.178
R31395 vdd.n2624 vdd.n2602 681.178
R31396 vdd.n2643 vdd.n2602 681.178
R31397 vdd.n2643 vdd.n2603 681.178
R31398 vdd.n2634 vdd.n2603 681.178
R31399 vdd.n2616 vdd.n2610 681.178
R31400 vdd.n2626 vdd.n2610 681.178
R31401 vdd.n2626 vdd.n2607 681.178
R31402 vdd.n2641 vdd.n2607 681.178
R31403 vdd.n2641 vdd.n2608 681.178
R31404 vdd.n2637 vdd.n2608 681.178
R31405 vdd.n1147 vdd.n1138 681.178
R31406 vdd.n1154 vdd.n1138 681.178
R31407 vdd.n1154 vdd.n1135 681.178
R31408 vdd.n1169 vdd.n1135 681.178
R31409 vdd.n1169 vdd.n1136 681.178
R31410 vdd.n1165 vdd.n1136 681.178
R31411 vdd.n1151 vdd.n1150 681.178
R31412 vdd.n1152 vdd.n1151 681.178
R31413 vdd.n1152 vdd.n1130 681.178
R31414 vdd.n1171 vdd.n1130 681.178
R31415 vdd.n1171 vdd.n1131 681.178
R31416 vdd.n1162 vdd.n1131 681.178
R31417 vdd.n1195 vdd.n1186 681.178
R31418 vdd.n1202 vdd.n1186 681.178
R31419 vdd.n1202 vdd.n1183 681.178
R31420 vdd.n1217 vdd.n1183 681.178
R31421 vdd.n1217 vdd.n1184 681.178
R31422 vdd.n1213 vdd.n1184 681.178
R31423 vdd.n1199 vdd.n1198 681.178
R31424 vdd.n1200 vdd.n1199 681.178
R31425 vdd.n1200 vdd.n1178 681.178
R31426 vdd.n1219 vdd.n1178 681.178
R31427 vdd.n1219 vdd.n1179 681.178
R31428 vdd.n1210 vdd.n1179 681.178
R31429 vdd.n1296 vdd.n1287 681.178
R31430 vdd.n1303 vdd.n1287 681.178
R31431 vdd.n1303 vdd.n1284 681.178
R31432 vdd.n1318 vdd.n1284 681.178
R31433 vdd.n1318 vdd.n1285 681.178
R31434 vdd.n1314 vdd.n1285 681.178
R31435 vdd.n1300 vdd.n1299 681.178
R31436 vdd.n1301 vdd.n1300 681.178
R31437 vdd.n1301 vdd.n1279 681.178
R31438 vdd.n1320 vdd.n1279 681.178
R31439 vdd.n1320 vdd.n1280 681.178
R31440 vdd.n1311 vdd.n1280 681.178
R31441 vdd.n1344 vdd.n1335 681.178
R31442 vdd.n1351 vdd.n1335 681.178
R31443 vdd.n1351 vdd.n1332 681.178
R31444 vdd.n1366 vdd.n1332 681.178
R31445 vdd.n1366 vdd.n1333 681.178
R31446 vdd.n1362 vdd.n1333 681.178
R31447 vdd.n1348 vdd.n1347 681.178
R31448 vdd.n1349 vdd.n1348 681.178
R31449 vdd.n1349 vdd.n1327 681.178
R31450 vdd.n1368 vdd.n1327 681.178
R31451 vdd.n1368 vdd.n1328 681.178
R31452 vdd.n1359 vdd.n1328 681.178
R31453 vdd.n1392 vdd.n1383 681.178
R31454 vdd.n1399 vdd.n1383 681.178
R31455 vdd.n1399 vdd.n1380 681.178
R31456 vdd.n1414 vdd.n1380 681.178
R31457 vdd.n1414 vdd.n1381 681.178
R31458 vdd.n1410 vdd.n1381 681.178
R31459 vdd.n1396 vdd.n1395 681.178
R31460 vdd.n1397 vdd.n1396 681.178
R31461 vdd.n1397 vdd.n1375 681.178
R31462 vdd.n1416 vdd.n1375 681.178
R31463 vdd.n1416 vdd.n1376 681.178
R31464 vdd.n1407 vdd.n1376 681.178
R31465 vdd.n1440 vdd.n1431 681.178
R31466 vdd.n1447 vdd.n1431 681.178
R31467 vdd.n1447 vdd.n1428 681.178
R31468 vdd.n1462 vdd.n1428 681.178
R31469 vdd.n1462 vdd.n1429 681.178
R31470 vdd.n1458 vdd.n1429 681.178
R31471 vdd.n1444 vdd.n1443 681.178
R31472 vdd.n1445 vdd.n1444 681.178
R31473 vdd.n1445 vdd.n1423 681.178
R31474 vdd.n1464 vdd.n1423 681.178
R31475 vdd.n1464 vdd.n1424 681.178
R31476 vdd.n1455 vdd.n1424 681.178
R31477 vdd.n1541 vdd.n1532 681.178
R31478 vdd.n1548 vdd.n1532 681.178
R31479 vdd.n1548 vdd.n1529 681.178
R31480 vdd.n1563 vdd.n1529 681.178
R31481 vdd.n1563 vdd.n1530 681.178
R31482 vdd.n1559 vdd.n1530 681.178
R31483 vdd.n1545 vdd.n1544 681.178
R31484 vdd.n1546 vdd.n1545 681.178
R31485 vdd.n1546 vdd.n1524 681.178
R31486 vdd.n1565 vdd.n1524 681.178
R31487 vdd.n1565 vdd.n1525 681.178
R31488 vdd.n1556 vdd.n1525 681.178
R31489 vdd.n654 vdd.n645 681.178
R31490 vdd.n661 vdd.n645 681.178
R31491 vdd.n661 vdd.n642 681.178
R31492 vdd.n676 vdd.n642 681.178
R31493 vdd.n676 vdd.n643 681.178
R31494 vdd.n672 vdd.n643 681.178
R31495 vdd.n658 vdd.n657 681.178
R31496 vdd.n659 vdd.n658 681.178
R31497 vdd.n659 vdd.n637 681.178
R31498 vdd.n678 vdd.n637 681.178
R31499 vdd.n678 vdd.n638 681.178
R31500 vdd.n669 vdd.n638 681.178
R31501 vdd.n1589 vdd.n1580 681.178
R31502 vdd.n1596 vdd.n1580 681.178
R31503 vdd.n1596 vdd.n1577 681.178
R31504 vdd.n1611 vdd.n1577 681.178
R31505 vdd.n1611 vdd.n1578 681.178
R31506 vdd.n1607 vdd.n1578 681.178
R31507 vdd.n1593 vdd.n1592 681.178
R31508 vdd.n1594 vdd.n1593 681.178
R31509 vdd.n1594 vdd.n1572 681.178
R31510 vdd.n1613 vdd.n1572 681.178
R31511 vdd.n1613 vdd.n1573 681.178
R31512 vdd.n1604 vdd.n1573 681.178
R31513 vdd.n1636 vdd.n1627 681.178
R31514 vdd.n1643 vdd.n1627 681.178
R31515 vdd.n1643 vdd.n1624 681.178
R31516 vdd.n1658 vdd.n1624 681.178
R31517 vdd.n1658 vdd.n1625 681.178
R31518 vdd.n1654 vdd.n1625 681.178
R31519 vdd.n1640 vdd.n1639 681.178
R31520 vdd.n1641 vdd.n1640 681.178
R31521 vdd.n1641 vdd.n1619 681.178
R31522 vdd.n1660 vdd.n1619 681.178
R31523 vdd.n1660 vdd.n1620 681.178
R31524 vdd.n1651 vdd.n1620 681.178
R31525 vdd.n1686 vdd.n1677 681.178
R31526 vdd.n1693 vdd.n1677 681.178
R31527 vdd.n1693 vdd.n1674 681.178
R31528 vdd.n1708 vdd.n1674 681.178
R31529 vdd.n1708 vdd.n1675 681.178
R31530 vdd.n1704 vdd.n1675 681.178
R31531 vdd.n1690 vdd.n1689 681.178
R31532 vdd.n1691 vdd.n1690 681.178
R31533 vdd.n1691 vdd.n1669 681.178
R31534 vdd.n1710 vdd.n1669 681.178
R31535 vdd.n1710 vdd.n1670 681.178
R31536 vdd.n1701 vdd.n1670 681.178
R31537 vdd.n1736 vdd.n1727 681.178
R31538 vdd.n1743 vdd.n1727 681.178
R31539 vdd.n1743 vdd.n1724 681.178
R31540 vdd.n1758 vdd.n1724 681.178
R31541 vdd.n1758 vdd.n1725 681.178
R31542 vdd.n1754 vdd.n1725 681.178
R31543 vdd.n1740 vdd.n1739 681.178
R31544 vdd.n1741 vdd.n1740 681.178
R31545 vdd.n1741 vdd.n1719 681.178
R31546 vdd.n1760 vdd.n1719 681.178
R31547 vdd.n1760 vdd.n1720 681.178
R31548 vdd.n1751 vdd.n1720 681.178
R31549 vdd.n1784 vdd.n1775 681.178
R31550 vdd.n1791 vdd.n1775 681.178
R31551 vdd.n1791 vdd.n1772 681.178
R31552 vdd.n1806 vdd.n1772 681.178
R31553 vdd.n1806 vdd.n1773 681.178
R31554 vdd.n1802 vdd.n1773 681.178
R31555 vdd.n1788 vdd.n1787 681.178
R31556 vdd.n1789 vdd.n1788 681.178
R31557 vdd.n1789 vdd.n1767 681.178
R31558 vdd.n1808 vdd.n1767 681.178
R31559 vdd.n1808 vdd.n1768 681.178
R31560 vdd.n1799 vdd.n1768 681.178
R31561 vdd.n1512 vdd.n1475 681.178
R31562 vdd.n1508 vdd.n1475 681.178
R31563 vdd.n1508 vdd.n1479 681.178
R31564 vdd.n1498 vdd.n1479 681.178
R31565 vdd.n1498 vdd.n1484 681.178
R31566 vdd.n1494 vdd.n1484 681.178
R31567 vdd.n1515 vdd.n1473 681.178
R31568 vdd.n1506 vdd.n1473 681.178
R31569 vdd.n1506 vdd.n1501 681.178
R31570 vdd.n1501 vdd.n1500 681.178
R31571 vdd.n1500 vdd.n1481 681.178
R31572 vdd.n1491 vdd.n1481 681.178
R31573 vdd.n1835 vdd.n1826 681.178
R31574 vdd.n1842 vdd.n1826 681.178
R31575 vdd.n1842 vdd.n1823 681.178
R31576 vdd.n1857 vdd.n1823 681.178
R31577 vdd.n1857 vdd.n1824 681.178
R31578 vdd.n1853 vdd.n1824 681.178
R31579 vdd.n1839 vdd.n1838 681.178
R31580 vdd.n1840 vdd.n1839 681.178
R31581 vdd.n1840 vdd.n1818 681.178
R31582 vdd.n1859 vdd.n1818 681.178
R31583 vdd.n1859 vdd.n1819 681.178
R31584 vdd.n1850 vdd.n1819 681.178
R31585 vdd.n1882 vdd.n1873 681.178
R31586 vdd.n1889 vdd.n1873 681.178
R31587 vdd.n1889 vdd.n1870 681.178
R31588 vdd.n1904 vdd.n1870 681.178
R31589 vdd.n1904 vdd.n1871 681.178
R31590 vdd.n1900 vdd.n1871 681.178
R31591 vdd.n1886 vdd.n1885 681.178
R31592 vdd.n1887 vdd.n1886 681.178
R31593 vdd.n1887 vdd.n1865 681.178
R31594 vdd.n1906 vdd.n1865 681.178
R31595 vdd.n1906 vdd.n1866 681.178
R31596 vdd.n1897 vdd.n1866 681.178
R31597 vdd.n1930 vdd.n1921 681.178
R31598 vdd.n1937 vdd.n1921 681.178
R31599 vdd.n1937 vdd.n1918 681.178
R31600 vdd.n1952 vdd.n1918 681.178
R31601 vdd.n1952 vdd.n1919 681.178
R31602 vdd.n1948 vdd.n1919 681.178
R31603 vdd.n1934 vdd.n1933 681.178
R31604 vdd.n1935 vdd.n1934 681.178
R31605 vdd.n1935 vdd.n1913 681.178
R31606 vdd.n1954 vdd.n1913 681.178
R31607 vdd.n1954 vdd.n1914 681.178
R31608 vdd.n1945 vdd.n1914 681.178
R31609 vdd.n1981 vdd.n1972 681.178
R31610 vdd.n1988 vdd.n1972 681.178
R31611 vdd.n1988 vdd.n1969 681.178
R31612 vdd.n2003 vdd.n1969 681.178
R31613 vdd.n2003 vdd.n1970 681.178
R31614 vdd.n1999 vdd.n1970 681.178
R31615 vdd.n1985 vdd.n1984 681.178
R31616 vdd.n1986 vdd.n1985 681.178
R31617 vdd.n1986 vdd.n1964 681.178
R31618 vdd.n2005 vdd.n1964 681.178
R31619 vdd.n2005 vdd.n1965 681.178
R31620 vdd.n1996 vdd.n1965 681.178
R31621 vdd.n2031 vdd.n2022 681.178
R31622 vdd.n2038 vdd.n2022 681.178
R31623 vdd.n2038 vdd.n2019 681.178
R31624 vdd.n2053 vdd.n2019 681.178
R31625 vdd.n2053 vdd.n2020 681.178
R31626 vdd.n2049 vdd.n2020 681.178
R31627 vdd.n2035 vdd.n2034 681.178
R31628 vdd.n2036 vdd.n2035 681.178
R31629 vdd.n2036 vdd.n2014 681.178
R31630 vdd.n2055 vdd.n2014 681.178
R31631 vdd.n2055 vdd.n2015 681.178
R31632 vdd.n2046 vdd.n2015 681.178
R31633 vdd.n2079 vdd.n2070 681.178
R31634 vdd.n2086 vdd.n2070 681.178
R31635 vdd.n2086 vdd.n2067 681.178
R31636 vdd.n2101 vdd.n2067 681.178
R31637 vdd.n2101 vdd.n2068 681.178
R31638 vdd.n2097 vdd.n2068 681.178
R31639 vdd.n2083 vdd.n2082 681.178
R31640 vdd.n2084 vdd.n2083 681.178
R31641 vdd.n2084 vdd.n2062 681.178
R31642 vdd.n2103 vdd.n2062 681.178
R31643 vdd.n2103 vdd.n2063 681.178
R31644 vdd.n2094 vdd.n2063 681.178
R31645 vdd.n2129 vdd.n2120 681.178
R31646 vdd.n2136 vdd.n2120 681.178
R31647 vdd.n2136 vdd.n2117 681.178
R31648 vdd.n2151 vdd.n2117 681.178
R31649 vdd.n2151 vdd.n2118 681.178
R31650 vdd.n2147 vdd.n2118 681.178
R31651 vdd.n2133 vdd.n2132 681.178
R31652 vdd.n2134 vdd.n2133 681.178
R31653 vdd.n2134 vdd.n2112 681.178
R31654 vdd.n2153 vdd.n2112 681.178
R31655 vdd.n2153 vdd.n2113 681.178
R31656 vdd.n2144 vdd.n2113 681.178
R31657 vdd.n2176 vdd.n2167 681.178
R31658 vdd.n2183 vdd.n2167 681.178
R31659 vdd.n2183 vdd.n2164 681.178
R31660 vdd.n2198 vdd.n2164 681.178
R31661 vdd.n2198 vdd.n2165 681.178
R31662 vdd.n2194 vdd.n2165 681.178
R31663 vdd.n2180 vdd.n2179 681.178
R31664 vdd.n2181 vdd.n2180 681.178
R31665 vdd.n2181 vdd.n2159 681.178
R31666 vdd.n2200 vdd.n2159 681.178
R31667 vdd.n2200 vdd.n2160 681.178
R31668 vdd.n2191 vdd.n2160 681.178
R31669 vdd.n2226 vdd.n2217 681.178
R31670 vdd.n2233 vdd.n2217 681.178
R31671 vdd.n2233 vdd.n2214 681.178
R31672 vdd.n2248 vdd.n2214 681.178
R31673 vdd.n2248 vdd.n2215 681.178
R31674 vdd.n2244 vdd.n2215 681.178
R31675 vdd.n2230 vdd.n2229 681.178
R31676 vdd.n2231 vdd.n2230 681.178
R31677 vdd.n2231 vdd.n2209 681.178
R31678 vdd.n2250 vdd.n2209 681.178
R31679 vdd.n2250 vdd.n2210 681.178
R31680 vdd.n2241 vdd.n2210 681.178
R31681 vdd.n2276 vdd.n2267 681.178
R31682 vdd.n2283 vdd.n2267 681.178
R31683 vdd.n2283 vdd.n2264 681.178
R31684 vdd.n2298 vdd.n2264 681.178
R31685 vdd.n2298 vdd.n2265 681.178
R31686 vdd.n2294 vdd.n2265 681.178
R31687 vdd.n2280 vdd.n2279 681.178
R31688 vdd.n2281 vdd.n2280 681.178
R31689 vdd.n2281 vdd.n2259 681.178
R31690 vdd.n2300 vdd.n2259 681.178
R31691 vdd.n2300 vdd.n2260 681.178
R31692 vdd.n2291 vdd.n2260 681.178
R31693 vdd.n2324 vdd.n2315 681.178
R31694 vdd.n2331 vdd.n2315 681.178
R31695 vdd.n2331 vdd.n2312 681.178
R31696 vdd.n2346 vdd.n2312 681.178
R31697 vdd.n2346 vdd.n2313 681.178
R31698 vdd.n2342 vdd.n2313 681.178
R31699 vdd.n2328 vdd.n2327 681.178
R31700 vdd.n2329 vdd.n2328 681.178
R31701 vdd.n2329 vdd.n2307 681.178
R31702 vdd.n2348 vdd.n2307 681.178
R31703 vdd.n2348 vdd.n2308 681.178
R31704 vdd.n2339 vdd.n2308 681.178
R31705 vdd.n1267 vdd.n1230 681.178
R31706 vdd.n1263 vdd.n1230 681.178
R31707 vdd.n1263 vdd.n1234 681.178
R31708 vdd.n1253 vdd.n1234 681.178
R31709 vdd.n1253 vdd.n1239 681.178
R31710 vdd.n1249 vdd.n1239 681.178
R31711 vdd.n1270 vdd.n1228 681.178
R31712 vdd.n1261 vdd.n1228 681.178
R31713 vdd.n1261 vdd.n1256 681.178
R31714 vdd.n1256 vdd.n1255 681.178
R31715 vdd.n1255 vdd.n1236 681.178
R31716 vdd.n1246 vdd.n1236 681.178
R31717 vdd.n2375 vdd.n2366 681.178
R31718 vdd.n2382 vdd.n2366 681.178
R31719 vdd.n2382 vdd.n2363 681.178
R31720 vdd.n2397 vdd.n2363 681.178
R31721 vdd.n2397 vdd.n2364 681.178
R31722 vdd.n2393 vdd.n2364 681.178
R31723 vdd.n2379 vdd.n2378 681.178
R31724 vdd.n2380 vdd.n2379 681.178
R31725 vdd.n2380 vdd.n2358 681.178
R31726 vdd.n2399 vdd.n2358 681.178
R31727 vdd.n2399 vdd.n2359 681.178
R31728 vdd.n2390 vdd.n2359 681.178
R31729 vdd.n2422 vdd.n2413 681.178
R31730 vdd.n2429 vdd.n2413 681.178
R31731 vdd.n2429 vdd.n2410 681.178
R31732 vdd.n2444 vdd.n2410 681.178
R31733 vdd.n2444 vdd.n2411 681.178
R31734 vdd.n2440 vdd.n2411 681.178
R31735 vdd.n2426 vdd.n2425 681.178
R31736 vdd.n2427 vdd.n2426 681.178
R31737 vdd.n2427 vdd.n2405 681.178
R31738 vdd.n2446 vdd.n2405 681.178
R31739 vdd.n2446 vdd.n2406 681.178
R31740 vdd.n2437 vdd.n2406 681.178
R31741 vdd.n2472 vdd.n2463 681.178
R31742 vdd.n2479 vdd.n2463 681.178
R31743 vdd.n2479 vdd.n2460 681.178
R31744 vdd.n2494 vdd.n2460 681.178
R31745 vdd.n2494 vdd.n2461 681.178
R31746 vdd.n2490 vdd.n2461 681.178
R31747 vdd.n2476 vdd.n2475 681.178
R31748 vdd.n2477 vdd.n2476 681.178
R31749 vdd.n2477 vdd.n2455 681.178
R31750 vdd.n2496 vdd.n2455 681.178
R31751 vdd.n2496 vdd.n2456 681.178
R31752 vdd.n2487 vdd.n2456 681.178
R31753 vdd.n2522 vdd.n2513 681.178
R31754 vdd.n2529 vdd.n2513 681.178
R31755 vdd.n2529 vdd.n2510 681.178
R31756 vdd.n2544 vdd.n2510 681.178
R31757 vdd.n2544 vdd.n2511 681.178
R31758 vdd.n2540 vdd.n2511 681.178
R31759 vdd.n2526 vdd.n2525 681.178
R31760 vdd.n2527 vdd.n2526 681.178
R31761 vdd.n2527 vdd.n2505 681.178
R31762 vdd.n2546 vdd.n2505 681.178
R31763 vdd.n2546 vdd.n2506 681.178
R31764 vdd.n2537 vdd.n2506 681.178
R31765 vdd.n2570 vdd.n2561 681.178
R31766 vdd.n2577 vdd.n2561 681.178
R31767 vdd.n2577 vdd.n2558 681.178
R31768 vdd.n2592 vdd.n2558 681.178
R31769 vdd.n2592 vdd.n2559 681.178
R31770 vdd.n2588 vdd.n2559 681.178
R31771 vdd.n2574 vdd.n2573 681.178
R31772 vdd.n2575 vdd.n2574 681.178
R31773 vdd.n2575 vdd.n2553 681.178
R31774 vdd.n2594 vdd.n2553 681.178
R31775 vdd.n2594 vdd.n2554 681.178
R31776 vdd.n2585 vdd.n2554 681.178
R31777 vdd.n2720 vdd.n2719 681.178
R31778 vdd.n2721 vdd.n2720 681.178
R31779 vdd.n2721 vdd.n2699 681.178
R31780 vdd.n2740 vdd.n2699 681.178
R31781 vdd.n2740 vdd.n2700 681.178
R31782 vdd.n2731 vdd.n2700 681.178
R31783 vdd.n2713 vdd.n2707 681.178
R31784 vdd.n2723 vdd.n2707 681.178
R31785 vdd.n2723 vdd.n2704 681.178
R31786 vdd.n2738 vdd.n2704 681.178
R31787 vdd.n2738 vdd.n2705 681.178
R31788 vdd.n2734 vdd.n2705 681.178
R31789 vdd.n2672 vdd.n2671 681.178
R31790 vdd.n2673 vdd.n2672 681.178
R31791 vdd.n2673 vdd.n2651 681.178
R31792 vdd.n2692 vdd.n2651 681.178
R31793 vdd.n2692 vdd.n2652 681.178
R31794 vdd.n2683 vdd.n2652 681.178
R31795 vdd.n2665 vdd.n2659 681.178
R31796 vdd.n2675 vdd.n2659 681.178
R31797 vdd.n2675 vdd.n2656 681.178
R31798 vdd.n2690 vdd.n2656 681.178
R31799 vdd.n2690 vdd.n2657 681.178
R31800 vdd.n2686 vdd.n2657 681.178
R31801 vdd.n2769 vdd.n2768 681.178
R31802 vdd.n2770 vdd.n2769 681.178
R31803 vdd.n2770 vdd.n2748 681.178
R31804 vdd.n2789 vdd.n2748 681.178
R31805 vdd.n2789 vdd.n2749 681.178
R31806 vdd.n2780 vdd.n2749 681.178
R31807 vdd.n2762 vdd.n2756 681.178
R31808 vdd.n2772 vdd.n2756 681.178
R31809 vdd.n2772 vdd.n2753 681.178
R31810 vdd.n2787 vdd.n2753 681.178
R31811 vdd.n2787 vdd.n2754 681.178
R31812 vdd.n2783 vdd.n2754 681.178
R31813 vdd.n2819 vdd.n2818 681.178
R31814 vdd.n2820 vdd.n2819 681.178
R31815 vdd.n2820 vdd.n2798 681.178
R31816 vdd.n2839 vdd.n2798 681.178
R31817 vdd.n2839 vdd.n2799 681.178
R31818 vdd.n2830 vdd.n2799 681.178
R31819 vdd.n2812 vdd.n2806 681.178
R31820 vdd.n2822 vdd.n2806 681.178
R31821 vdd.n2822 vdd.n2803 681.178
R31822 vdd.n2837 vdd.n2803 681.178
R31823 vdd.n2837 vdd.n2804 681.178
R31824 vdd.n2833 vdd.n2804 681.178
R31825 vdd.n2867 vdd.n2866 681.178
R31826 vdd.n2868 vdd.n2867 681.178
R31827 vdd.n2868 vdd.n2846 681.178
R31828 vdd.n2887 vdd.n2846 681.178
R31829 vdd.n2887 vdd.n2847 681.178
R31830 vdd.n2878 vdd.n2847 681.178
R31831 vdd.n2860 vdd.n2854 681.178
R31832 vdd.n2870 vdd.n2854 681.178
R31833 vdd.n2870 vdd.n2851 681.178
R31834 vdd.n2885 vdd.n2851 681.178
R31835 vdd.n2885 vdd.n2852 681.178
R31836 vdd.n2881 vdd.n2852 681.178
R31837 vdd.n1050 vdd.n1038 681.178
R31838 vdd.n1054 vdd.n1038 681.178
R31839 vdd.n1054 vdd.n1034 681.178
R31840 vdd.n1034 vdd.n1032 681.178
R31841 vdd.n1067 vdd.n1032 681.178
R31842 vdd.n1068 vdd.n1067 681.178
R31843 vdd.n1047 vdd.n1043 681.178
R31844 vdd.n1043 vdd.n1037 681.178
R31845 vdd.n1037 vdd.n1035 681.178
R31846 vdd.n1057 vdd.n1035 681.178
R31847 vdd.n1057 vdd.n1030 681.178
R31848 vdd.n1071 vdd.n1030 681.178
R31849 vdd.n3015 vdd.n3014 681.178
R31850 vdd.n3016 vdd.n3015 681.178
R31851 vdd.n3016 vdd.n2994 681.178
R31852 vdd.n3035 vdd.n2994 681.178
R31853 vdd.n3035 vdd.n2995 681.178
R31854 vdd.n3026 vdd.n2995 681.178
R31855 vdd.n3008 vdd.n3002 681.178
R31856 vdd.n3018 vdd.n3002 681.178
R31857 vdd.n3018 vdd.n2999 681.178
R31858 vdd.n3033 vdd.n2999 681.178
R31859 vdd.n3033 vdd.n3000 681.178
R31860 vdd.n3029 vdd.n3000 681.178
R31861 vdd.n2966 vdd.n2965 681.178
R31862 vdd.n2967 vdd.n2966 681.178
R31863 vdd.n2967 vdd.n2945 681.178
R31864 vdd.n2986 vdd.n2945 681.178
R31865 vdd.n2986 vdd.n2946 681.178
R31866 vdd.n2977 vdd.n2946 681.178
R31867 vdd.n2959 vdd.n2953 681.178
R31868 vdd.n2969 vdd.n2953 681.178
R31869 vdd.n2969 vdd.n2950 681.178
R31870 vdd.n2984 vdd.n2950 681.178
R31871 vdd.n2984 vdd.n2951 681.178
R31872 vdd.n2980 vdd.n2951 681.178
R31873 vdd.n2918 vdd.n2917 681.178
R31874 vdd.n2919 vdd.n2918 681.178
R31875 vdd.n2919 vdd.n2897 681.178
R31876 vdd.n2938 vdd.n2897 681.178
R31877 vdd.n2938 vdd.n2898 681.178
R31878 vdd.n2929 vdd.n2898 681.178
R31879 vdd.n2911 vdd.n2905 681.178
R31880 vdd.n2921 vdd.n2905 681.178
R31881 vdd.n2921 vdd.n2902 681.178
R31882 vdd.n2936 vdd.n2902 681.178
R31883 vdd.n2936 vdd.n2903 681.178
R31884 vdd.n2932 vdd.n2903 681.178
R31885 vdd.n3064 vdd.n3063 681.178
R31886 vdd.n3065 vdd.n3064 681.178
R31887 vdd.n3065 vdd.n3043 681.178
R31888 vdd.n3084 vdd.n3043 681.178
R31889 vdd.n3084 vdd.n3044 681.178
R31890 vdd.n3075 vdd.n3044 681.178
R31891 vdd.n3057 vdd.n3051 681.178
R31892 vdd.n3067 vdd.n3051 681.178
R31893 vdd.n3067 vdd.n3048 681.178
R31894 vdd.n3082 vdd.n3048 681.178
R31895 vdd.n3082 vdd.n3049 681.178
R31896 vdd.n3078 vdd.n3049 681.178
R31897 vdd.n3114 vdd.n3113 681.178
R31898 vdd.n3115 vdd.n3114 681.178
R31899 vdd.n3115 vdd.n3093 681.178
R31900 vdd.n3134 vdd.n3093 681.178
R31901 vdd.n3134 vdd.n3094 681.178
R31902 vdd.n3125 vdd.n3094 681.178
R31903 vdd.n3107 vdd.n3101 681.178
R31904 vdd.n3117 vdd.n3101 681.178
R31905 vdd.n3117 vdd.n3098 681.178
R31906 vdd.n3132 vdd.n3098 681.178
R31907 vdd.n3132 vdd.n3099 681.178
R31908 vdd.n3128 vdd.n3099 681.178
R31909 vdd.n3162 vdd.n3161 681.178
R31910 vdd.n3163 vdd.n3162 681.178
R31911 vdd.n3163 vdd.n3141 681.178
R31912 vdd.n3182 vdd.n3141 681.178
R31913 vdd.n3182 vdd.n3142 681.178
R31914 vdd.n3173 vdd.n3142 681.178
R31915 vdd.n3155 vdd.n3149 681.178
R31916 vdd.n3165 vdd.n3149 681.178
R31917 vdd.n3165 vdd.n3146 681.178
R31918 vdd.n3180 vdd.n3146 681.178
R31919 vdd.n3180 vdd.n3147 681.178
R31920 vdd.n3176 vdd.n3147 681.178
R31921 vdd.n3260 vdd.n3259 681.178
R31922 vdd.n3261 vdd.n3260 681.178
R31923 vdd.n3261 vdd.n3239 681.178
R31924 vdd.n3280 vdd.n3239 681.178
R31925 vdd.n3280 vdd.n3240 681.178
R31926 vdd.n3271 vdd.n3240 681.178
R31927 vdd.n3253 vdd.n3247 681.178
R31928 vdd.n3263 vdd.n3247 681.178
R31929 vdd.n3263 vdd.n3244 681.178
R31930 vdd.n3278 vdd.n3244 681.178
R31931 vdd.n3278 vdd.n3245 681.178
R31932 vdd.n3274 vdd.n3245 681.178
R31933 vdd.n3212 vdd.n3211 681.178
R31934 vdd.n3213 vdd.n3212 681.178
R31935 vdd.n3213 vdd.n3191 681.178
R31936 vdd.n3232 vdd.n3191 681.178
R31937 vdd.n3232 vdd.n3192 681.178
R31938 vdd.n3223 vdd.n3192 681.178
R31939 vdd.n3205 vdd.n3199 681.178
R31940 vdd.n3215 vdd.n3199 681.178
R31941 vdd.n3215 vdd.n3196 681.178
R31942 vdd.n3230 vdd.n3196 681.178
R31943 vdd.n3230 vdd.n3197 681.178
R31944 vdd.n3226 vdd.n3197 681.178
R31945 vdd.n3309 vdd.n3308 681.178
R31946 vdd.n3310 vdd.n3309 681.178
R31947 vdd.n3310 vdd.n3288 681.178
R31948 vdd.n3329 vdd.n3288 681.178
R31949 vdd.n3329 vdd.n3289 681.178
R31950 vdd.n3320 vdd.n3289 681.178
R31951 vdd.n3302 vdd.n3296 681.178
R31952 vdd.n3312 vdd.n3296 681.178
R31953 vdd.n3312 vdd.n3293 681.178
R31954 vdd.n3327 vdd.n3293 681.178
R31955 vdd.n3327 vdd.n3294 681.178
R31956 vdd.n3323 vdd.n3294 681.178
R31957 vdd.n3359 vdd.n3358 681.178
R31958 vdd.n3360 vdd.n3359 681.178
R31959 vdd.n3360 vdd.n3338 681.178
R31960 vdd.n3379 vdd.n3338 681.178
R31961 vdd.n3379 vdd.n3339 681.178
R31962 vdd.n3370 vdd.n3339 681.178
R31963 vdd.n3352 vdd.n3346 681.178
R31964 vdd.n3362 vdd.n3346 681.178
R31965 vdd.n3362 vdd.n3343 681.178
R31966 vdd.n3377 vdd.n3343 681.178
R31967 vdd.n3377 vdd.n3344 681.178
R31968 vdd.n3373 vdd.n3344 681.178
R31969 vdd.n3407 vdd.n3406 681.178
R31970 vdd.n3408 vdd.n3407 681.178
R31971 vdd.n3408 vdd.n3386 681.178
R31972 vdd.n3427 vdd.n3386 681.178
R31973 vdd.n3427 vdd.n3387 681.178
R31974 vdd.n3418 vdd.n3387 681.178
R31975 vdd.n3400 vdd.n3394 681.178
R31976 vdd.n3410 vdd.n3394 681.178
R31977 vdd.n3410 vdd.n3391 681.178
R31978 vdd.n3425 vdd.n3391 681.178
R31979 vdd.n3425 vdd.n3392 681.178
R31980 vdd.n3421 vdd.n3392 681.178
R31981 vdd.n804 vdd.n792 681.178
R31982 vdd.n808 vdd.n792 681.178
R31983 vdd.n808 vdd.n788 681.178
R31984 vdd.n788 vdd.n786 681.178
R31985 vdd.n821 vdd.n786 681.178
R31986 vdd.n822 vdd.n821 681.178
R31987 vdd.n801 vdd.n797 681.178
R31988 vdd.n797 vdd.n791 681.178
R31989 vdd.n791 vdd.n789 681.178
R31990 vdd.n811 vdd.n789 681.178
R31991 vdd.n811 vdd.n784 681.178
R31992 vdd.n825 vdd.n784 681.178
R31993 vdd.n3506 vdd.n3505 681.178
R31994 vdd.n3507 vdd.n3506 681.178
R31995 vdd.n3507 vdd.n3485 681.178
R31996 vdd.n3526 vdd.n3485 681.178
R31997 vdd.n3526 vdd.n3486 681.178
R31998 vdd.n3517 vdd.n3486 681.178
R31999 vdd.n3499 vdd.n3493 681.178
R32000 vdd.n3509 vdd.n3493 681.178
R32001 vdd.n3509 vdd.n3490 681.178
R32002 vdd.n3524 vdd.n3490 681.178
R32003 vdd.n3524 vdd.n3491 681.178
R32004 vdd.n3520 vdd.n3491 681.178
R32005 vdd.n3458 vdd.n3457 681.178
R32006 vdd.n3459 vdd.n3458 681.178
R32007 vdd.n3459 vdd.n3437 681.178
R32008 vdd.n3478 vdd.n3437 681.178
R32009 vdd.n3478 vdd.n3438 681.178
R32010 vdd.n3469 vdd.n3438 681.178
R32011 vdd.n3451 vdd.n3445 681.178
R32012 vdd.n3461 vdd.n3445 681.178
R32013 vdd.n3461 vdd.n3442 681.178
R32014 vdd.n3476 vdd.n3442 681.178
R32015 vdd.n3476 vdd.n3443 681.178
R32016 vdd.n3472 vdd.n3443 681.178
R32017 vdd.n3555 vdd.n3554 681.178
R32018 vdd.n3556 vdd.n3555 681.178
R32019 vdd.n3556 vdd.n3534 681.178
R32020 vdd.n3575 vdd.n3534 681.178
R32021 vdd.n3575 vdd.n3535 681.178
R32022 vdd.n3566 vdd.n3535 681.178
R32023 vdd.n3548 vdd.n3542 681.178
R32024 vdd.n3558 vdd.n3542 681.178
R32025 vdd.n3558 vdd.n3539 681.178
R32026 vdd.n3573 vdd.n3539 681.178
R32027 vdd.n3573 vdd.n3540 681.178
R32028 vdd.n3569 vdd.n3540 681.178
R32029 vdd.n3605 vdd.n3604 681.178
R32030 vdd.n3606 vdd.n3605 681.178
R32031 vdd.n3606 vdd.n3584 681.178
R32032 vdd.n3625 vdd.n3584 681.178
R32033 vdd.n3625 vdd.n3585 681.178
R32034 vdd.n3616 vdd.n3585 681.178
R32035 vdd.n3598 vdd.n3592 681.178
R32036 vdd.n3608 vdd.n3592 681.178
R32037 vdd.n3608 vdd.n3589 681.178
R32038 vdd.n3623 vdd.n3589 681.178
R32039 vdd.n3623 vdd.n3590 681.178
R32040 vdd.n3619 vdd.n3590 681.178
R32041 vdd.n3653 vdd.n3652 681.178
R32042 vdd.n3654 vdd.n3653 681.178
R32043 vdd.n3654 vdd.n3632 681.178
R32044 vdd.n3673 vdd.n3632 681.178
R32045 vdd.n3673 vdd.n3633 681.178
R32046 vdd.n3664 vdd.n3633 681.178
R32047 vdd.n3646 vdd.n3640 681.178
R32048 vdd.n3656 vdd.n3640 681.178
R32049 vdd.n3656 vdd.n3637 681.178
R32050 vdd.n3671 vdd.n3637 681.178
R32051 vdd.n3671 vdd.n3638 681.178
R32052 vdd.n3667 vdd.n3638 681.178
R32053 vdd.n611 vdd.n610 681.178
R32054 vdd.n612 vdd.n611 681.178
R32055 vdd.n612 vdd.n590 681.178
R32056 vdd.n631 vdd.n590 681.178
R32057 vdd.n631 vdd.n591 681.178
R32058 vdd.n622 vdd.n591 681.178
R32059 vdd.n604 vdd.n598 681.178
R32060 vdd.n614 vdd.n598 681.178
R32061 vdd.n614 vdd.n595 681.178
R32062 vdd.n629 vdd.n595 681.178
R32063 vdd.n629 vdd.n596 681.178
R32064 vdd.n625 vdd.n596 681.178
R32065 vdd.n3752 vdd.n3751 681.178
R32066 vdd.n3753 vdd.n3752 681.178
R32067 vdd.n3753 vdd.n3731 681.178
R32068 vdd.n3772 vdd.n3731 681.178
R32069 vdd.n3772 vdd.n3732 681.178
R32070 vdd.n3763 vdd.n3732 681.178
R32071 vdd.n3745 vdd.n3739 681.178
R32072 vdd.n3755 vdd.n3739 681.178
R32073 vdd.n3755 vdd.n3736 681.178
R32074 vdd.n3770 vdd.n3736 681.178
R32075 vdd.n3770 vdd.n3737 681.178
R32076 vdd.n3766 vdd.n3737 681.178
R32077 vdd.n3704 vdd.n3703 681.178
R32078 vdd.n3705 vdd.n3704 681.178
R32079 vdd.n3705 vdd.n3683 681.178
R32080 vdd.n3724 vdd.n3683 681.178
R32081 vdd.n3724 vdd.n3684 681.178
R32082 vdd.n3715 vdd.n3684 681.178
R32083 vdd.n3697 vdd.n3691 681.178
R32084 vdd.n3707 vdd.n3691 681.178
R32085 vdd.n3707 vdd.n3688 681.178
R32086 vdd.n3722 vdd.n3688 681.178
R32087 vdd.n3722 vdd.n3689 681.178
R32088 vdd.n3718 vdd.n3689 681.178
R32089 vdd.n6894 vdd.n6893 681.178
R32090 vdd.n6895 vdd.n6894 681.178
R32091 vdd.n6895 vdd.n6873 681.178
R32092 vdd.n6914 vdd.n6873 681.178
R32093 vdd.n6914 vdd.n6874 681.178
R32094 vdd.n6905 vdd.n6874 681.178
R32095 vdd.n6887 vdd.n6881 681.178
R32096 vdd.n6897 vdd.n6881 681.178
R32097 vdd.n6897 vdd.n6878 681.178
R32098 vdd.n6912 vdd.n6878 681.178
R32099 vdd.n6912 vdd.n6879 681.178
R32100 vdd.n6908 vdd.n6879 681.178
R32101 vdd.n6846 vdd.n6845 681.178
R32102 vdd.n6847 vdd.n6846 681.178
R32103 vdd.n6847 vdd.n6825 681.178
R32104 vdd.n6866 vdd.n6825 681.178
R32105 vdd.n6866 vdd.n6826 681.178
R32106 vdd.n6857 vdd.n6826 681.178
R32107 vdd.n6839 vdd.n6833 681.178
R32108 vdd.n6849 vdd.n6833 681.178
R32109 vdd.n6849 vdd.n6830 681.178
R32110 vdd.n6864 vdd.n6830 681.178
R32111 vdd.n6864 vdd.n6831 681.178
R32112 vdd.n6860 vdd.n6831 681.178
R32113 vdd.n10036 vdd.n10035 681.178
R32114 vdd.n10037 vdd.n10036 681.178
R32115 vdd.n10037 vdd.n10015 681.178
R32116 vdd.n10056 vdd.n10015 681.178
R32117 vdd.n10056 vdd.n10016 681.178
R32118 vdd.n10047 vdd.n10016 681.178
R32119 vdd.n10029 vdd.n10023 681.178
R32120 vdd.n10039 vdd.n10023 681.178
R32121 vdd.n10039 vdd.n10020 681.178
R32122 vdd.n10054 vdd.n10020 681.178
R32123 vdd.n10054 vdd.n10021 681.178
R32124 vdd.n10050 vdd.n10021 681.178
R32125 vdd.n9988 vdd.n9987 681.178
R32126 vdd.n9989 vdd.n9988 681.178
R32127 vdd.n9989 vdd.n9967 681.178
R32128 vdd.n10008 vdd.n9967 681.178
R32129 vdd.n10008 vdd.n9968 681.178
R32130 vdd.n9999 vdd.n9968 681.178
R32131 vdd.n9981 vdd.n9975 681.178
R32132 vdd.n9991 vdd.n9975 681.178
R32133 vdd.n9991 vdd.n9972 681.178
R32134 vdd.n10006 vdd.n9972 681.178
R32135 vdd.n10006 vdd.n9973 681.178
R32136 vdd.n10002 vdd.n9973 681.178
R32137 vdd.n10084 vdd.n10083 681.178
R32138 vdd.n10085 vdd.n10084 681.178
R32139 vdd.n10085 vdd.n10063 681.178
R32140 vdd.n10104 vdd.n10063 681.178
R32141 vdd.n10104 vdd.n10064 681.178
R32142 vdd.n10095 vdd.n10064 681.178
R32143 vdd.n10077 vdd.n10071 681.178
R32144 vdd.n10087 vdd.n10071 681.178
R32145 vdd.n10087 vdd.n10068 681.178
R32146 vdd.n10102 vdd.n10068 681.178
R32147 vdd.n10102 vdd.n10069 681.178
R32148 vdd.n10098 vdd.n10069 681.178
R32149 vdd.n10132 vdd.n10131 681.178
R32150 vdd.n10133 vdd.n10132 681.178
R32151 vdd.n10133 vdd.n10111 681.178
R32152 vdd.n10152 vdd.n10111 681.178
R32153 vdd.n10152 vdd.n10112 681.178
R32154 vdd.n10143 vdd.n10112 681.178
R32155 vdd.n10125 vdd.n10119 681.178
R32156 vdd.n10135 vdd.n10119 681.178
R32157 vdd.n10135 vdd.n10116 681.178
R32158 vdd.n10150 vdd.n10116 681.178
R32159 vdd.n10150 vdd.n10117 681.178
R32160 vdd.n10146 vdd.n10117 681.178
R32161 vdd.n10234 vdd.n10233 681.178
R32162 vdd.n10235 vdd.n10234 681.178
R32163 vdd.n10235 vdd.n10213 681.178
R32164 vdd.n10254 vdd.n10213 681.178
R32165 vdd.n10254 vdd.n10214 681.178
R32166 vdd.n10245 vdd.n10214 681.178
R32167 vdd.n10227 vdd.n10221 681.178
R32168 vdd.n10237 vdd.n10221 681.178
R32169 vdd.n10237 vdd.n10218 681.178
R32170 vdd.n10252 vdd.n10218 681.178
R32171 vdd.n10252 vdd.n10219 681.178
R32172 vdd.n10248 vdd.n10219 681.178
R32173 vdd.n10282 vdd.n10281 681.178
R32174 vdd.n10283 vdd.n10282 681.178
R32175 vdd.n10283 vdd.n10261 681.178
R32176 vdd.n10302 vdd.n10261 681.178
R32177 vdd.n10302 vdd.n10262 681.178
R32178 vdd.n10293 vdd.n10262 681.178
R32179 vdd.n10275 vdd.n10269 681.178
R32180 vdd.n10285 vdd.n10269 681.178
R32181 vdd.n10285 vdd.n10266 681.178
R32182 vdd.n10300 vdd.n10266 681.178
R32183 vdd.n10300 vdd.n10267 681.178
R32184 vdd.n10296 vdd.n10267 681.178
R32185 vdd.n10330 vdd.n10329 681.178
R32186 vdd.n10331 vdd.n10330 681.178
R32187 vdd.n10331 vdd.n10309 681.178
R32188 vdd.n10350 vdd.n10309 681.178
R32189 vdd.n10350 vdd.n10310 681.178
R32190 vdd.n10341 vdd.n10310 681.178
R32191 vdd.n10323 vdd.n10317 681.178
R32192 vdd.n10333 vdd.n10317 681.178
R32193 vdd.n10333 vdd.n10314 681.178
R32194 vdd.n10348 vdd.n10314 681.178
R32195 vdd.n10348 vdd.n10315 681.178
R32196 vdd.n10344 vdd.n10315 681.178
R32197 vdd.n10378 vdd.n10377 681.178
R32198 vdd.n10379 vdd.n10378 681.178
R32199 vdd.n10379 vdd.n10357 681.178
R32200 vdd.n10398 vdd.n10357 681.178
R32201 vdd.n10398 vdd.n10358 681.178
R32202 vdd.n10389 vdd.n10358 681.178
R32203 vdd.n10371 vdd.n10365 681.178
R32204 vdd.n10381 vdd.n10365 681.178
R32205 vdd.n10381 vdd.n10362 681.178
R32206 vdd.n10396 vdd.n10362 681.178
R32207 vdd.n10396 vdd.n10363 681.178
R32208 vdd.n10392 vdd.n10363 681.178
R32209 vdd.n10480 vdd.n10479 681.178
R32210 vdd.n10481 vdd.n10480 681.178
R32211 vdd.n10481 vdd.n10459 681.178
R32212 vdd.n10500 vdd.n10459 681.178
R32213 vdd.n10500 vdd.n10460 681.178
R32214 vdd.n10491 vdd.n10460 681.178
R32215 vdd.n10473 vdd.n10467 681.178
R32216 vdd.n10483 vdd.n10467 681.178
R32217 vdd.n10483 vdd.n10464 681.178
R32218 vdd.n10498 vdd.n10464 681.178
R32219 vdd.n10498 vdd.n10465 681.178
R32220 vdd.n10494 vdd.n10465 681.178
R32221 vdd.n72 vdd.n71 681.178
R32222 vdd.n73 vdd.n72 681.178
R32223 vdd.n73 vdd.n51 681.178
R32224 vdd.n92 vdd.n51 681.178
R32225 vdd.n92 vdd.n52 681.178
R32226 vdd.n83 vdd.n52 681.178
R32227 vdd.n65 vdd.n59 681.178
R32228 vdd.n75 vdd.n59 681.178
R32229 vdd.n75 vdd.n56 681.178
R32230 vdd.n90 vdd.n56 681.178
R32231 vdd.n90 vdd.n57 681.178
R32232 vdd.n86 vdd.n57 681.178
R32233 vdd.n24 vdd.n23 681.178
R32234 vdd.n25 vdd.n24 681.178
R32235 vdd.n25 vdd.n3 681.178
R32236 vdd.n44 vdd.n3 681.178
R32237 vdd.n44 vdd.n4 681.178
R32238 vdd.n35 vdd.n4 681.178
R32239 vdd.n17 vdd.n11 681.178
R32240 vdd.n27 vdd.n11 681.178
R32241 vdd.n27 vdd.n8 681.178
R32242 vdd.n42 vdd.n8 681.178
R32243 vdd.n42 vdd.n9 681.178
R32244 vdd.n38 vdd.n9 681.178
R32245 vdd.n10528 vdd.n10527 681.178
R32246 vdd.n10529 vdd.n10528 681.178
R32247 vdd.n10529 vdd.n10507 681.178
R32248 vdd.n10548 vdd.n10507 681.178
R32249 vdd.n10548 vdd.n10508 681.178
R32250 vdd.n10539 vdd.n10508 681.178
R32251 vdd.n10521 vdd.n10515 681.178
R32252 vdd.n10531 vdd.n10515 681.178
R32253 vdd.n10531 vdd.n10512 681.178
R32254 vdd.n10546 vdd.n10512 681.178
R32255 vdd.n10546 vdd.n10513 681.178
R32256 vdd.n10542 vdd.n10513 681.178
R32257 vdd.n10578 vdd.n10577 681.178
R32258 vdd.n10579 vdd.n10578 681.178
R32259 vdd.n10579 vdd.n10557 681.178
R32260 vdd.n10598 vdd.n10557 681.178
R32261 vdd.n10598 vdd.n10558 681.178
R32262 vdd.n10589 vdd.n10558 681.178
R32263 vdd.n10571 vdd.n10565 681.178
R32264 vdd.n10581 vdd.n10565 681.178
R32265 vdd.n10581 vdd.n10562 681.178
R32266 vdd.n10596 vdd.n10562 681.178
R32267 vdd.n10596 vdd.n10563 681.178
R32268 vdd.n10592 vdd.n10563 681.178
R32269 vdd.n10626 vdd.n10625 681.178
R32270 vdd.n10627 vdd.n10626 681.178
R32271 vdd.n10627 vdd.n10605 681.178
R32272 vdd.n10646 vdd.n10605 681.178
R32273 vdd.n10646 vdd.n10606 681.178
R32274 vdd.n10637 vdd.n10606 681.178
R32275 vdd.n10619 vdd.n10613 681.178
R32276 vdd.n10629 vdd.n10613 681.178
R32277 vdd.n10629 vdd.n10610 681.178
R32278 vdd.n10644 vdd.n10610 681.178
R32279 vdd.n10644 vdd.n10611 681.178
R32280 vdd.n10640 vdd.n10611 681.178
R32281 vdd.n10427 vdd.n10415 681.178
R32282 vdd.n10431 vdd.n10415 681.178
R32283 vdd.n10431 vdd.n10411 681.178
R32284 vdd.n10411 vdd.n10409 681.178
R32285 vdd.n10444 vdd.n10409 681.178
R32286 vdd.n10445 vdd.n10444 681.178
R32287 vdd.n10424 vdd.n10420 681.178
R32288 vdd.n10420 vdd.n10414 681.178
R32289 vdd.n10414 vdd.n10412 681.178
R32290 vdd.n10434 vdd.n10412 681.178
R32291 vdd.n10434 vdd.n10407 681.178
R32292 vdd.n10448 vdd.n10407 681.178
R32293 vdd.n10774 vdd.n10773 681.178
R32294 vdd.n10775 vdd.n10774 681.178
R32295 vdd.n10775 vdd.n10753 681.178
R32296 vdd.n10794 vdd.n10753 681.178
R32297 vdd.n10794 vdd.n10754 681.178
R32298 vdd.n10785 vdd.n10754 681.178
R32299 vdd.n10767 vdd.n10761 681.178
R32300 vdd.n10777 vdd.n10761 681.178
R32301 vdd.n10777 vdd.n10758 681.178
R32302 vdd.n10792 vdd.n10758 681.178
R32303 vdd.n10792 vdd.n10759 681.178
R32304 vdd.n10788 vdd.n10759 681.178
R32305 vdd.n10725 vdd.n10724 681.178
R32306 vdd.n10726 vdd.n10725 681.178
R32307 vdd.n10726 vdd.n10704 681.178
R32308 vdd.n10745 vdd.n10704 681.178
R32309 vdd.n10745 vdd.n10705 681.178
R32310 vdd.n10736 vdd.n10705 681.178
R32311 vdd.n10718 vdd.n10712 681.178
R32312 vdd.n10728 vdd.n10712 681.178
R32313 vdd.n10728 vdd.n10709 681.178
R32314 vdd.n10743 vdd.n10709 681.178
R32315 vdd.n10743 vdd.n10710 681.178
R32316 vdd.n10739 vdd.n10710 681.178
R32317 vdd.n10677 vdd.n10676 681.178
R32318 vdd.n10678 vdd.n10677 681.178
R32319 vdd.n10678 vdd.n10656 681.178
R32320 vdd.n10697 vdd.n10656 681.178
R32321 vdd.n10697 vdd.n10657 681.178
R32322 vdd.n10688 vdd.n10657 681.178
R32323 vdd.n10670 vdd.n10664 681.178
R32324 vdd.n10680 vdd.n10664 681.178
R32325 vdd.n10680 vdd.n10661 681.178
R32326 vdd.n10695 vdd.n10661 681.178
R32327 vdd.n10695 vdd.n10662 681.178
R32328 vdd.n10691 vdd.n10662 681.178
R32329 vdd.n10823 vdd.n10822 681.178
R32330 vdd.n10824 vdd.n10823 681.178
R32331 vdd.n10824 vdd.n10802 681.178
R32332 vdd.n10843 vdd.n10802 681.178
R32333 vdd.n10843 vdd.n10803 681.178
R32334 vdd.n10834 vdd.n10803 681.178
R32335 vdd.n10816 vdd.n10810 681.178
R32336 vdd.n10826 vdd.n10810 681.178
R32337 vdd.n10826 vdd.n10807 681.178
R32338 vdd.n10841 vdd.n10807 681.178
R32339 vdd.n10841 vdd.n10808 681.178
R32340 vdd.n10837 vdd.n10808 681.178
R32341 vdd.n10873 vdd.n10872 681.178
R32342 vdd.n10874 vdd.n10873 681.178
R32343 vdd.n10874 vdd.n10852 681.178
R32344 vdd.n10893 vdd.n10852 681.178
R32345 vdd.n10893 vdd.n10853 681.178
R32346 vdd.n10884 vdd.n10853 681.178
R32347 vdd.n10866 vdd.n10860 681.178
R32348 vdd.n10876 vdd.n10860 681.178
R32349 vdd.n10876 vdd.n10857 681.178
R32350 vdd.n10891 vdd.n10857 681.178
R32351 vdd.n10891 vdd.n10858 681.178
R32352 vdd.n10887 vdd.n10858 681.178
R32353 vdd.n10921 vdd.n10920 681.178
R32354 vdd.n10922 vdd.n10921 681.178
R32355 vdd.n10922 vdd.n10900 681.178
R32356 vdd.n10941 vdd.n10900 681.178
R32357 vdd.n10941 vdd.n10901 681.178
R32358 vdd.n10932 vdd.n10901 681.178
R32359 vdd.n10914 vdd.n10908 681.178
R32360 vdd.n10924 vdd.n10908 681.178
R32361 vdd.n10924 vdd.n10905 681.178
R32362 vdd.n10939 vdd.n10905 681.178
R32363 vdd.n10939 vdd.n10906 681.178
R32364 vdd.n10935 vdd.n10906 681.178
R32365 vdd.n11019 vdd.n11018 681.178
R32366 vdd.n11020 vdd.n11019 681.178
R32367 vdd.n11020 vdd.n10998 681.178
R32368 vdd.n11039 vdd.n10998 681.178
R32369 vdd.n11039 vdd.n10999 681.178
R32370 vdd.n11030 vdd.n10999 681.178
R32371 vdd.n11012 vdd.n11006 681.178
R32372 vdd.n11022 vdd.n11006 681.178
R32373 vdd.n11022 vdd.n11003 681.178
R32374 vdd.n11037 vdd.n11003 681.178
R32375 vdd.n11037 vdd.n11004 681.178
R32376 vdd.n11033 vdd.n11004 681.178
R32377 vdd.n10971 vdd.n10970 681.178
R32378 vdd.n10972 vdd.n10971 681.178
R32379 vdd.n10972 vdd.n10950 681.178
R32380 vdd.n10991 vdd.n10950 681.178
R32381 vdd.n10991 vdd.n10951 681.178
R32382 vdd.n10982 vdd.n10951 681.178
R32383 vdd.n10964 vdd.n10958 681.178
R32384 vdd.n10974 vdd.n10958 681.178
R32385 vdd.n10974 vdd.n10955 681.178
R32386 vdd.n10989 vdd.n10955 681.178
R32387 vdd.n10989 vdd.n10956 681.178
R32388 vdd.n10985 vdd.n10956 681.178
R32389 vdd.n11068 vdd.n11067 681.178
R32390 vdd.n11069 vdd.n11068 681.178
R32391 vdd.n11069 vdd.n11047 681.178
R32392 vdd.n11088 vdd.n11047 681.178
R32393 vdd.n11088 vdd.n11048 681.178
R32394 vdd.n11079 vdd.n11048 681.178
R32395 vdd.n11061 vdd.n11055 681.178
R32396 vdd.n11071 vdd.n11055 681.178
R32397 vdd.n11071 vdd.n11052 681.178
R32398 vdd.n11086 vdd.n11052 681.178
R32399 vdd.n11086 vdd.n11053 681.178
R32400 vdd.n11082 vdd.n11053 681.178
R32401 vdd.n11118 vdd.n11117 681.178
R32402 vdd.n11119 vdd.n11118 681.178
R32403 vdd.n11119 vdd.n11097 681.178
R32404 vdd.n11138 vdd.n11097 681.178
R32405 vdd.n11138 vdd.n11098 681.178
R32406 vdd.n11129 vdd.n11098 681.178
R32407 vdd.n11111 vdd.n11105 681.178
R32408 vdd.n11121 vdd.n11105 681.178
R32409 vdd.n11121 vdd.n11102 681.178
R32410 vdd.n11136 vdd.n11102 681.178
R32411 vdd.n11136 vdd.n11103 681.178
R32412 vdd.n11132 vdd.n11103 681.178
R32413 vdd.n11166 vdd.n11165 681.178
R32414 vdd.n11167 vdd.n11166 681.178
R32415 vdd.n11167 vdd.n11145 681.178
R32416 vdd.n11186 vdd.n11145 681.178
R32417 vdd.n11186 vdd.n11146 681.178
R32418 vdd.n11177 vdd.n11146 681.178
R32419 vdd.n11159 vdd.n11153 681.178
R32420 vdd.n11169 vdd.n11153 681.178
R32421 vdd.n11169 vdd.n11150 681.178
R32422 vdd.n11184 vdd.n11150 681.178
R32423 vdd.n11184 vdd.n11151 681.178
R32424 vdd.n11180 vdd.n11151 681.178
R32425 vdd.n10181 vdd.n10169 681.178
R32426 vdd.n10185 vdd.n10169 681.178
R32427 vdd.n10185 vdd.n10165 681.178
R32428 vdd.n10165 vdd.n10163 681.178
R32429 vdd.n10198 vdd.n10163 681.178
R32430 vdd.n10199 vdd.n10198 681.178
R32431 vdd.n10178 vdd.n10174 681.178
R32432 vdd.n10174 vdd.n10168 681.178
R32433 vdd.n10168 vdd.n10166 681.178
R32434 vdd.n10188 vdd.n10166 681.178
R32435 vdd.n10188 vdd.n10161 681.178
R32436 vdd.n10202 vdd.n10161 681.178
R32437 vdd.n11265 vdd.n11264 681.178
R32438 vdd.n11266 vdd.n11265 681.178
R32439 vdd.n11266 vdd.n11244 681.178
R32440 vdd.n11285 vdd.n11244 681.178
R32441 vdd.n11285 vdd.n11245 681.178
R32442 vdd.n11276 vdd.n11245 681.178
R32443 vdd.n11258 vdd.n11252 681.178
R32444 vdd.n11268 vdd.n11252 681.178
R32445 vdd.n11268 vdd.n11249 681.178
R32446 vdd.n11283 vdd.n11249 681.178
R32447 vdd.n11283 vdd.n11250 681.178
R32448 vdd.n11279 vdd.n11250 681.178
R32449 vdd.n11217 vdd.n11216 681.178
R32450 vdd.n11218 vdd.n11217 681.178
R32451 vdd.n11218 vdd.n11196 681.178
R32452 vdd.n11237 vdd.n11196 681.178
R32453 vdd.n11237 vdd.n11197 681.178
R32454 vdd.n11228 vdd.n11197 681.178
R32455 vdd.n11210 vdd.n11204 681.178
R32456 vdd.n11220 vdd.n11204 681.178
R32457 vdd.n11220 vdd.n11201 681.178
R32458 vdd.n11235 vdd.n11201 681.178
R32459 vdd.n11235 vdd.n11202 681.178
R32460 vdd.n11231 vdd.n11202 681.178
R32461 vdd.n11314 vdd.n11313 681.178
R32462 vdd.n11315 vdd.n11314 681.178
R32463 vdd.n11315 vdd.n11293 681.178
R32464 vdd.n11334 vdd.n11293 681.178
R32465 vdd.n11334 vdd.n11294 681.178
R32466 vdd.n11325 vdd.n11294 681.178
R32467 vdd.n11307 vdd.n11301 681.178
R32468 vdd.n11317 vdd.n11301 681.178
R32469 vdd.n11317 vdd.n11298 681.178
R32470 vdd.n11332 vdd.n11298 681.178
R32471 vdd.n11332 vdd.n11299 681.178
R32472 vdd.n11328 vdd.n11299 681.178
R32473 vdd.n11364 vdd.n11363 681.178
R32474 vdd.n11365 vdd.n11364 681.178
R32475 vdd.n11365 vdd.n11343 681.178
R32476 vdd.n11384 vdd.n11343 681.178
R32477 vdd.n11384 vdd.n11344 681.178
R32478 vdd.n11375 vdd.n11344 681.178
R32479 vdd.n11357 vdd.n11351 681.178
R32480 vdd.n11367 vdd.n11351 681.178
R32481 vdd.n11367 vdd.n11348 681.178
R32482 vdd.n11382 vdd.n11348 681.178
R32483 vdd.n11382 vdd.n11349 681.178
R32484 vdd.n11378 vdd.n11349 681.178
R32485 vdd.n11412 vdd.n11411 681.178
R32486 vdd.n11413 vdd.n11412 681.178
R32487 vdd.n11413 vdd.n11391 681.178
R32488 vdd.n11432 vdd.n11391 681.178
R32489 vdd.n11432 vdd.n11392 681.178
R32490 vdd.n11423 vdd.n11392 681.178
R32491 vdd.n11405 vdd.n11399 681.178
R32492 vdd.n11415 vdd.n11399 681.178
R32493 vdd.n11415 vdd.n11396 681.178
R32494 vdd.n11430 vdd.n11396 681.178
R32495 vdd.n11430 vdd.n11397 681.178
R32496 vdd.n11426 vdd.n11397 681.178
R32497 vdd.n11459 vdd.n11450 681.178
R32498 vdd.n11466 vdd.n11450 681.178
R32499 vdd.n11466 vdd.n11447 681.178
R32500 vdd.n11481 vdd.n11447 681.178
R32501 vdd.n11481 vdd.n11448 681.178
R32502 vdd.n11477 vdd.n11448 681.178
R32503 vdd.n11463 vdd.n11462 681.178
R32504 vdd.n11464 vdd.n11463 681.178
R32505 vdd.n11464 vdd.n11442 681.178
R32506 vdd.n11483 vdd.n11442 681.178
R32507 vdd.n11483 vdd.n11443 681.178
R32508 vdd.n11474 vdd.n11443 681.178
R32509 vdd.n11506 vdd.n11497 681.178
R32510 vdd.n11513 vdd.n11497 681.178
R32511 vdd.n11513 vdd.n11494 681.178
R32512 vdd.n11528 vdd.n11494 681.178
R32513 vdd.n11528 vdd.n11495 681.178
R32514 vdd.n11524 vdd.n11495 681.178
R32515 vdd.n11510 vdd.n11509 681.178
R32516 vdd.n11511 vdd.n11510 681.178
R32517 vdd.n11511 vdd.n11489 681.178
R32518 vdd.n11530 vdd.n11489 681.178
R32519 vdd.n11530 vdd.n11490 681.178
R32520 vdd.n11521 vdd.n11490 681.178
R32521 vdd.n11556 vdd.n11547 681.178
R32522 vdd.n11563 vdd.n11547 681.178
R32523 vdd.n11563 vdd.n11544 681.178
R32524 vdd.n11578 vdd.n11544 681.178
R32525 vdd.n11578 vdd.n11545 681.178
R32526 vdd.n11574 vdd.n11545 681.178
R32527 vdd.n11560 vdd.n11559 681.178
R32528 vdd.n11561 vdd.n11560 681.178
R32529 vdd.n11561 vdd.n11539 681.178
R32530 vdd.n11580 vdd.n11539 681.178
R32531 vdd.n11580 vdd.n11540 681.178
R32532 vdd.n11571 vdd.n11540 681.178
R32533 vdd.n11606 vdd.n11597 681.178
R32534 vdd.n11613 vdd.n11597 681.178
R32535 vdd.n11613 vdd.n11594 681.178
R32536 vdd.n11628 vdd.n11594 681.178
R32537 vdd.n11628 vdd.n11595 681.178
R32538 vdd.n11624 vdd.n11595 681.178
R32539 vdd.n11610 vdd.n11609 681.178
R32540 vdd.n11611 vdd.n11610 681.178
R32541 vdd.n11611 vdd.n11589 681.178
R32542 vdd.n11630 vdd.n11589 681.178
R32543 vdd.n11630 vdd.n11590 681.178
R32544 vdd.n11621 vdd.n11590 681.178
R32545 vdd.n11654 vdd.n11645 681.178
R32546 vdd.n11661 vdd.n11645 681.178
R32547 vdd.n11661 vdd.n11642 681.178
R32548 vdd.n11676 vdd.n11642 681.178
R32549 vdd.n11676 vdd.n11643 681.178
R32550 vdd.n11672 vdd.n11643 681.178
R32551 vdd.n11658 vdd.n11657 681.178
R32552 vdd.n11659 vdd.n11658 681.178
R32553 vdd.n11659 vdd.n11637 681.178
R32554 vdd.n11678 vdd.n11637 681.178
R32555 vdd.n11678 vdd.n11638 681.178
R32556 vdd.n11669 vdd.n11638 681.178
R32557 vdd.n482 vdd.n445 681.178
R32558 vdd.n478 vdd.n445 681.178
R32559 vdd.n478 vdd.n449 681.178
R32560 vdd.n468 vdd.n449 681.178
R32561 vdd.n468 vdd.n454 681.178
R32562 vdd.n464 vdd.n454 681.178
R32563 vdd.n485 vdd.n443 681.178
R32564 vdd.n476 vdd.n443 681.178
R32565 vdd.n476 vdd.n471 681.178
R32566 vdd.n471 vdd.n470 681.178
R32567 vdd.n470 vdd.n451 681.178
R32568 vdd.n461 vdd.n451 681.178
R32569 vdd.n11705 vdd.n11696 681.178
R32570 vdd.n11712 vdd.n11696 681.178
R32571 vdd.n11712 vdd.n11693 681.178
R32572 vdd.n11727 vdd.n11693 681.178
R32573 vdd.n11727 vdd.n11694 681.178
R32574 vdd.n11723 vdd.n11694 681.178
R32575 vdd.n11709 vdd.n11708 681.178
R32576 vdd.n11710 vdd.n11709 681.178
R32577 vdd.n11710 vdd.n11688 681.178
R32578 vdd.n11729 vdd.n11688 681.178
R32579 vdd.n11729 vdd.n11689 681.178
R32580 vdd.n11720 vdd.n11689 681.178
R32581 vdd.n11752 vdd.n11743 681.178
R32582 vdd.n11759 vdd.n11743 681.178
R32583 vdd.n11759 vdd.n11740 681.178
R32584 vdd.n11774 vdd.n11740 681.178
R32585 vdd.n11774 vdd.n11741 681.178
R32586 vdd.n11770 vdd.n11741 681.178
R32587 vdd.n11756 vdd.n11755 681.178
R32588 vdd.n11757 vdd.n11756 681.178
R32589 vdd.n11757 vdd.n11735 681.178
R32590 vdd.n11776 vdd.n11735 681.178
R32591 vdd.n11776 vdd.n11736 681.178
R32592 vdd.n11767 vdd.n11736 681.178
R32593 vdd.n11800 vdd.n11791 681.178
R32594 vdd.n11807 vdd.n11791 681.178
R32595 vdd.n11807 vdd.n11788 681.178
R32596 vdd.n11822 vdd.n11788 681.178
R32597 vdd.n11822 vdd.n11789 681.178
R32598 vdd.n11818 vdd.n11789 681.178
R32599 vdd.n11804 vdd.n11803 681.178
R32600 vdd.n11805 vdd.n11804 681.178
R32601 vdd.n11805 vdd.n11783 681.178
R32602 vdd.n11824 vdd.n11783 681.178
R32603 vdd.n11824 vdd.n11784 681.178
R32604 vdd.n11815 vdd.n11784 681.178
R32605 vdd.n11851 vdd.n11842 681.178
R32606 vdd.n11858 vdd.n11842 681.178
R32607 vdd.n11858 vdd.n11839 681.178
R32608 vdd.n11873 vdd.n11839 681.178
R32609 vdd.n11873 vdd.n11840 681.178
R32610 vdd.n11869 vdd.n11840 681.178
R32611 vdd.n11855 vdd.n11854 681.178
R32612 vdd.n11856 vdd.n11855 681.178
R32613 vdd.n11856 vdd.n11834 681.178
R32614 vdd.n11875 vdd.n11834 681.178
R32615 vdd.n11875 vdd.n11835 681.178
R32616 vdd.n11866 vdd.n11835 681.178
R32617 vdd.n11901 vdd.n11892 681.178
R32618 vdd.n11908 vdd.n11892 681.178
R32619 vdd.n11908 vdd.n11889 681.178
R32620 vdd.n11923 vdd.n11889 681.178
R32621 vdd.n11923 vdd.n11890 681.178
R32622 vdd.n11919 vdd.n11890 681.178
R32623 vdd.n11905 vdd.n11904 681.178
R32624 vdd.n11906 vdd.n11905 681.178
R32625 vdd.n11906 vdd.n11884 681.178
R32626 vdd.n11925 vdd.n11884 681.178
R32627 vdd.n11925 vdd.n11885 681.178
R32628 vdd.n11916 vdd.n11885 681.178
R32629 vdd.n11949 vdd.n11940 681.178
R32630 vdd.n11956 vdd.n11940 681.178
R32631 vdd.n11956 vdd.n11937 681.178
R32632 vdd.n11971 vdd.n11937 681.178
R32633 vdd.n11971 vdd.n11938 681.178
R32634 vdd.n11967 vdd.n11938 681.178
R32635 vdd.n11953 vdd.n11952 681.178
R32636 vdd.n11954 vdd.n11953 681.178
R32637 vdd.n11954 vdd.n11932 681.178
R32638 vdd.n11973 vdd.n11932 681.178
R32639 vdd.n11973 vdd.n11933 681.178
R32640 vdd.n11964 vdd.n11933 681.178
R32641 vdd.n11999 vdd.n11990 681.178
R32642 vdd.n12006 vdd.n11990 681.178
R32643 vdd.n12006 vdd.n11987 681.178
R32644 vdd.n12021 vdd.n11987 681.178
R32645 vdd.n12021 vdd.n11988 681.178
R32646 vdd.n12017 vdd.n11988 681.178
R32647 vdd.n12003 vdd.n12002 681.178
R32648 vdd.n12004 vdd.n12003 681.178
R32649 vdd.n12004 vdd.n11982 681.178
R32650 vdd.n12023 vdd.n11982 681.178
R32651 vdd.n12023 vdd.n11983 681.178
R32652 vdd.n12014 vdd.n11983 681.178
R32653 vdd.n12046 vdd.n12037 681.178
R32654 vdd.n12053 vdd.n12037 681.178
R32655 vdd.n12053 vdd.n12034 681.178
R32656 vdd.n12068 vdd.n12034 681.178
R32657 vdd.n12068 vdd.n12035 681.178
R32658 vdd.n12064 vdd.n12035 681.178
R32659 vdd.n12050 vdd.n12049 681.178
R32660 vdd.n12051 vdd.n12050 681.178
R32661 vdd.n12051 vdd.n12029 681.178
R32662 vdd.n12070 vdd.n12029 681.178
R32663 vdd.n12070 vdd.n12030 681.178
R32664 vdd.n12061 vdd.n12030 681.178
R32665 vdd.n12096 vdd.n12087 681.178
R32666 vdd.n12103 vdd.n12087 681.178
R32667 vdd.n12103 vdd.n12084 681.178
R32668 vdd.n12118 vdd.n12084 681.178
R32669 vdd.n12118 vdd.n12085 681.178
R32670 vdd.n12114 vdd.n12085 681.178
R32671 vdd.n12100 vdd.n12099 681.178
R32672 vdd.n12101 vdd.n12100 681.178
R32673 vdd.n12101 vdd.n12079 681.178
R32674 vdd.n12120 vdd.n12079 681.178
R32675 vdd.n12120 vdd.n12080 681.178
R32676 vdd.n12111 vdd.n12080 681.178
R32677 vdd.n12146 vdd.n12137 681.178
R32678 vdd.n12153 vdd.n12137 681.178
R32679 vdd.n12153 vdd.n12134 681.178
R32680 vdd.n12168 vdd.n12134 681.178
R32681 vdd.n12168 vdd.n12135 681.178
R32682 vdd.n12164 vdd.n12135 681.178
R32683 vdd.n12150 vdd.n12149 681.178
R32684 vdd.n12151 vdd.n12150 681.178
R32685 vdd.n12151 vdd.n12129 681.178
R32686 vdd.n12170 vdd.n12129 681.178
R32687 vdd.n12170 vdd.n12130 681.178
R32688 vdd.n12161 vdd.n12130 681.178
R32689 vdd.n12194 vdd.n12185 681.178
R32690 vdd.n12201 vdd.n12185 681.178
R32691 vdd.n12201 vdd.n12182 681.178
R32692 vdd.n12216 vdd.n12182 681.178
R32693 vdd.n12216 vdd.n12183 681.178
R32694 vdd.n12212 vdd.n12183 681.178
R32695 vdd.n12198 vdd.n12197 681.178
R32696 vdd.n12199 vdd.n12198 681.178
R32697 vdd.n12199 vdd.n12177 681.178
R32698 vdd.n12218 vdd.n12177 681.178
R32699 vdd.n12218 vdd.n12178 681.178
R32700 vdd.n12209 vdd.n12178 681.178
R32701 vdd.n237 vdd.n200 681.178
R32702 vdd.n233 vdd.n200 681.178
R32703 vdd.n233 vdd.n204 681.178
R32704 vdd.n223 vdd.n204 681.178
R32705 vdd.n223 vdd.n209 681.178
R32706 vdd.n219 vdd.n209 681.178
R32707 vdd.n240 vdd.n198 681.178
R32708 vdd.n231 vdd.n198 681.178
R32709 vdd.n231 vdd.n226 681.178
R32710 vdd.n226 vdd.n225 681.178
R32711 vdd.n225 vdd.n206 681.178
R32712 vdd.n216 vdd.n206 681.178
R32713 vdd.n12245 vdd.n12236 681.178
R32714 vdd.n12252 vdd.n12236 681.178
R32715 vdd.n12252 vdd.n12233 681.178
R32716 vdd.n12267 vdd.n12233 681.178
R32717 vdd.n12267 vdd.n12234 681.178
R32718 vdd.n12263 vdd.n12234 681.178
R32719 vdd.n12249 vdd.n12248 681.178
R32720 vdd.n12250 vdd.n12249 681.178
R32721 vdd.n12250 vdd.n12228 681.178
R32722 vdd.n12269 vdd.n12228 681.178
R32723 vdd.n12269 vdd.n12229 681.178
R32724 vdd.n12260 vdd.n12229 681.178
R32725 vdd.n12292 vdd.n12283 681.178
R32726 vdd.n12299 vdd.n12283 681.178
R32727 vdd.n12299 vdd.n12280 681.178
R32728 vdd.n12314 vdd.n12280 681.178
R32729 vdd.n12314 vdd.n12281 681.178
R32730 vdd.n12310 vdd.n12281 681.178
R32731 vdd.n12296 vdd.n12295 681.178
R32732 vdd.n12297 vdd.n12296 681.178
R32733 vdd.n12297 vdd.n12275 681.178
R32734 vdd.n12316 vdd.n12275 681.178
R32735 vdd.n12316 vdd.n12276 681.178
R32736 vdd.n12307 vdd.n12276 681.178
R32737 vdd.n12342 vdd.n12333 681.178
R32738 vdd.n12349 vdd.n12333 681.178
R32739 vdd.n12349 vdd.n12330 681.178
R32740 vdd.n12364 vdd.n12330 681.178
R32741 vdd.n12364 vdd.n12331 681.178
R32742 vdd.n12360 vdd.n12331 681.178
R32743 vdd.n12346 vdd.n12345 681.178
R32744 vdd.n12347 vdd.n12346 681.178
R32745 vdd.n12347 vdd.n12325 681.178
R32746 vdd.n12366 vdd.n12325 681.178
R32747 vdd.n12366 vdd.n12326 681.178
R32748 vdd.n12357 vdd.n12326 681.178
R32749 vdd.n12392 vdd.n12383 681.178
R32750 vdd.n12399 vdd.n12383 681.178
R32751 vdd.n12399 vdd.n12380 681.178
R32752 vdd.n12414 vdd.n12380 681.178
R32753 vdd.n12414 vdd.n12381 681.178
R32754 vdd.n12410 vdd.n12381 681.178
R32755 vdd.n12396 vdd.n12395 681.178
R32756 vdd.n12397 vdd.n12396 681.178
R32757 vdd.n12397 vdd.n12375 681.178
R32758 vdd.n12416 vdd.n12375 681.178
R32759 vdd.n12416 vdd.n12376 681.178
R32760 vdd.n12407 vdd.n12376 681.178
R32761 vdd.n12440 vdd.n12431 681.178
R32762 vdd.n12447 vdd.n12431 681.178
R32763 vdd.n12447 vdd.n12428 681.178
R32764 vdd.n12462 vdd.n12428 681.178
R32765 vdd.n12462 vdd.n12429 681.178
R32766 vdd.n12458 vdd.n12429 681.178
R32767 vdd.n12444 vdd.n12443 681.178
R32768 vdd.n12445 vdd.n12444 681.178
R32769 vdd.n12445 vdd.n12423 681.178
R32770 vdd.n12464 vdd.n12423 681.178
R32771 vdd.n12464 vdd.n12424 681.178
R32772 vdd.n12455 vdd.n12424 681.178
R32773 vdd.n119 vdd.n109 287.382
R32774 vdd.n123 vdd.n109 287.382
R32775 vdd.n123 vdd.n102 287.382
R32776 vdd.n140 vdd.n102 287.382
R32777 vdd.n140 vdd.n103 287.382
R32778 vdd.n134 vdd.n103 287.382
R32779 vdd.n167 vdd.n157 287.382
R32780 vdd.n171 vdd.n157 287.382
R32781 vdd.n171 vdd.n150 287.382
R32782 vdd.n188 vdd.n150 287.382
R32783 vdd.n188 vdd.n151 287.382
R32784 vdd.n182 vdd.n151 287.382
R32785 vdd.n268 vdd.n258 287.382
R32786 vdd.n272 vdd.n258 287.382
R32787 vdd.n272 vdd.n251 287.382
R32788 vdd.n289 vdd.n251 287.382
R32789 vdd.n289 vdd.n252 287.382
R32790 vdd.n283 vdd.n252 287.382
R32791 vdd.n316 vdd.n306 287.382
R32792 vdd.n320 vdd.n306 287.382
R32793 vdd.n320 vdd.n299 287.382
R32794 vdd.n337 vdd.n299 287.382
R32795 vdd.n337 vdd.n300 287.382
R32796 vdd.n331 vdd.n300 287.382
R32797 vdd.n364 vdd.n354 287.382
R32798 vdd.n368 vdd.n354 287.382
R32799 vdd.n368 vdd.n347 287.382
R32800 vdd.n385 vdd.n347 287.382
R32801 vdd.n385 vdd.n348 287.382
R32802 vdd.n379 vdd.n348 287.382
R32803 vdd.n412 vdd.n402 287.382
R32804 vdd.n416 vdd.n402 287.382
R32805 vdd.n416 vdd.n395 287.382
R32806 vdd.n433 vdd.n395 287.382
R32807 vdd.n433 vdd.n396 287.382
R32808 vdd.n427 vdd.n396 287.382
R32809 vdd.n513 vdd.n503 287.382
R32810 vdd.n517 vdd.n503 287.382
R32811 vdd.n517 vdd.n496 287.382
R32812 vdd.n534 vdd.n496 287.382
R32813 vdd.n534 vdd.n497 287.382
R32814 vdd.n528 vdd.n497 287.382
R32815 vdd.n561 vdd.n551 287.382
R32816 vdd.n565 vdd.n551 287.382
R32817 vdd.n565 vdd.n544 287.382
R32818 vdd.n582 vdd.n544 287.382
R32819 vdd.n582 vdd.n545 287.382
R32820 vdd.n576 vdd.n545 287.382
R32821 vdd.n6983 vdd.n6979 287.382
R32822 vdd.n6993 vdd.n6979 287.382
R32823 vdd.n6993 vdd.n6972 287.382
R32824 vdd.n7010 vdd.n6972 287.382
R32825 vdd.n7010 vdd.n6973 287.382
R32826 vdd.n7003 vdd.n6973 287.382
R32827 vdd.n7031 vdd.n7027 287.382
R32828 vdd.n7041 vdd.n7027 287.382
R32829 vdd.n7041 vdd.n7020 287.382
R32830 vdd.n7058 vdd.n7020 287.382
R32831 vdd.n7058 vdd.n7021 287.382
R32832 vdd.n7051 vdd.n7021 287.382
R32833 vdd.n7133 vdd.n7129 287.382
R32834 vdd.n7143 vdd.n7129 287.382
R32835 vdd.n7143 vdd.n7122 287.382
R32836 vdd.n7160 vdd.n7122 287.382
R32837 vdd.n7160 vdd.n7123 287.382
R32838 vdd.n7153 vdd.n7123 287.382
R32839 vdd.n7181 vdd.n7177 287.382
R32840 vdd.n7191 vdd.n7177 287.382
R32841 vdd.n7191 vdd.n7170 287.382
R32842 vdd.n7208 vdd.n7170 287.382
R32843 vdd.n7208 vdd.n7171 287.382
R32844 vdd.n7201 vdd.n7171 287.382
R32845 vdd.n7229 vdd.n7225 287.382
R32846 vdd.n7239 vdd.n7225 287.382
R32847 vdd.n7239 vdd.n7218 287.382
R32848 vdd.n7256 vdd.n7218 287.382
R32849 vdd.n7256 vdd.n7219 287.382
R32850 vdd.n7249 vdd.n7219 287.382
R32851 vdd.n7277 vdd.n7273 287.382
R32852 vdd.n7287 vdd.n7273 287.382
R32853 vdd.n7287 vdd.n7266 287.382
R32854 vdd.n7304 vdd.n7266 287.382
R32855 vdd.n7304 vdd.n7267 287.382
R32856 vdd.n7297 vdd.n7267 287.382
R32857 vdd.n7379 vdd.n7375 287.382
R32858 vdd.n7389 vdd.n7375 287.382
R32859 vdd.n7389 vdd.n7368 287.382
R32860 vdd.n7406 vdd.n7368 287.382
R32861 vdd.n7406 vdd.n7369 287.382
R32862 vdd.n7399 vdd.n7369 287.382
R32863 vdd.n8899 vdd.n8895 287.382
R32864 vdd.n8909 vdd.n8895 287.382
R32865 vdd.n8909 vdd.n8888 287.382
R32866 vdd.n8926 vdd.n8888 287.382
R32867 vdd.n8926 vdd.n8889 287.382
R32868 vdd.n8919 vdd.n8889 287.382
R32869 vdd.n7433 vdd.n7423 287.382
R32870 vdd.n7437 vdd.n7423 287.382
R32871 vdd.n7437 vdd.n7416 287.382
R32872 vdd.n7454 vdd.n7416 287.382
R32873 vdd.n7454 vdd.n7417 287.382
R32874 vdd.n7448 vdd.n7417 287.382
R32875 vdd.n7481 vdd.n7471 287.382
R32876 vdd.n7485 vdd.n7471 287.382
R32877 vdd.n7485 vdd.n7464 287.382
R32878 vdd.n7502 vdd.n7464 287.382
R32879 vdd.n7502 vdd.n7465 287.382
R32880 vdd.n7496 vdd.n7465 287.382
R32881 vdd.n7582 vdd.n7572 287.382
R32882 vdd.n7586 vdd.n7572 287.382
R32883 vdd.n7586 vdd.n7565 287.382
R32884 vdd.n7603 vdd.n7565 287.382
R32885 vdd.n7603 vdd.n7566 287.382
R32886 vdd.n7597 vdd.n7566 287.382
R32887 vdd.n7630 vdd.n7620 287.382
R32888 vdd.n7634 vdd.n7620 287.382
R32889 vdd.n7634 vdd.n7613 287.382
R32890 vdd.n7651 vdd.n7613 287.382
R32891 vdd.n7651 vdd.n7614 287.382
R32892 vdd.n7645 vdd.n7614 287.382
R32893 vdd.n7678 vdd.n7668 287.382
R32894 vdd.n7682 vdd.n7668 287.382
R32895 vdd.n7682 vdd.n7661 287.382
R32896 vdd.n7699 vdd.n7661 287.382
R32897 vdd.n7699 vdd.n7662 287.382
R32898 vdd.n7693 vdd.n7662 287.382
R32899 vdd.n7726 vdd.n7716 287.382
R32900 vdd.n7730 vdd.n7716 287.382
R32901 vdd.n7730 vdd.n7709 287.382
R32902 vdd.n7747 vdd.n7709 287.382
R32903 vdd.n7747 vdd.n7710 287.382
R32904 vdd.n7741 vdd.n7710 287.382
R32905 vdd.n7827 vdd.n7817 287.382
R32906 vdd.n7831 vdd.n7817 287.382
R32907 vdd.n7831 vdd.n7810 287.382
R32908 vdd.n7848 vdd.n7810 287.382
R32909 vdd.n7848 vdd.n7811 287.382
R32910 vdd.n7842 vdd.n7811 287.382
R32911 vdd.n6940 vdd.n6930 287.382
R32912 vdd.n6944 vdd.n6930 287.382
R32913 vdd.n6944 vdd.n6923 287.382
R32914 vdd.n6961 vdd.n6923 287.382
R32915 vdd.n6961 vdd.n6924 287.382
R32916 vdd.n6955 vdd.n6924 287.382
R32917 vdd.n7875 vdd.n7865 287.382
R32918 vdd.n7879 vdd.n7865 287.382
R32919 vdd.n7879 vdd.n7858 287.382
R32920 vdd.n7896 vdd.n7858 287.382
R32921 vdd.n7896 vdd.n7859 287.382
R32922 vdd.n7890 vdd.n7859 287.382
R32923 vdd.n7922 vdd.n7912 287.382
R32924 vdd.n7926 vdd.n7912 287.382
R32925 vdd.n7926 vdd.n7905 287.382
R32926 vdd.n7943 vdd.n7905 287.382
R32927 vdd.n7943 vdd.n7906 287.382
R32928 vdd.n7937 vdd.n7906 287.382
R32929 vdd.n7972 vdd.n7962 287.382
R32930 vdd.n7976 vdd.n7962 287.382
R32931 vdd.n7976 vdd.n7955 287.382
R32932 vdd.n7993 vdd.n7955 287.382
R32933 vdd.n7993 vdd.n7956 287.382
R32934 vdd.n7987 vdd.n7956 287.382
R32935 vdd.n8022 vdd.n8012 287.382
R32936 vdd.n8026 vdd.n8012 287.382
R32937 vdd.n8026 vdd.n8005 287.382
R32938 vdd.n8043 vdd.n8005 287.382
R32939 vdd.n8043 vdd.n8006 287.382
R32940 vdd.n8037 vdd.n8006 287.382
R32941 vdd.n8070 vdd.n8060 287.382
R32942 vdd.n8074 vdd.n8060 287.382
R32943 vdd.n8074 vdd.n8053 287.382
R32944 vdd.n8091 vdd.n8053 287.382
R32945 vdd.n8091 vdd.n8054 287.382
R32946 vdd.n8085 vdd.n8054 287.382
R32947 vdd.n7798 vdd.n7758 287.382
R32948 vdd.n7791 vdd.n7758 287.382
R32949 vdd.n7791 vdd.n7764 287.382
R32950 vdd.n7783 vdd.n7764 287.382
R32951 vdd.n7783 vdd.n7767 287.382
R32952 vdd.n7777 vdd.n7767 287.382
R32953 vdd.n8121 vdd.n8111 287.382
R32954 vdd.n8125 vdd.n8111 287.382
R32955 vdd.n8125 vdd.n8104 287.382
R32956 vdd.n8142 vdd.n8104 287.382
R32957 vdd.n8142 vdd.n8105 287.382
R32958 vdd.n8136 vdd.n8105 287.382
R32959 vdd.n8168 vdd.n8158 287.382
R32960 vdd.n8172 vdd.n8158 287.382
R32961 vdd.n8172 vdd.n8151 287.382
R32962 vdd.n8189 vdd.n8151 287.382
R32963 vdd.n8189 vdd.n8152 287.382
R32964 vdd.n8183 vdd.n8152 287.382
R32965 vdd.n8216 vdd.n8206 287.382
R32966 vdd.n8220 vdd.n8206 287.382
R32967 vdd.n8220 vdd.n8199 287.382
R32968 vdd.n8237 vdd.n8199 287.382
R32969 vdd.n8237 vdd.n8200 287.382
R32970 vdd.n8231 vdd.n8200 287.382
R32971 vdd.n8267 vdd.n8257 287.382
R32972 vdd.n8271 vdd.n8257 287.382
R32973 vdd.n8271 vdd.n8250 287.382
R32974 vdd.n8288 vdd.n8250 287.382
R32975 vdd.n8288 vdd.n8251 287.382
R32976 vdd.n8282 vdd.n8251 287.382
R32977 vdd.n8317 vdd.n8307 287.382
R32978 vdd.n8321 vdd.n8307 287.382
R32979 vdd.n8321 vdd.n8300 287.382
R32980 vdd.n8338 vdd.n8300 287.382
R32981 vdd.n8338 vdd.n8301 287.382
R32982 vdd.n8332 vdd.n8301 287.382
R32983 vdd.n8365 vdd.n8355 287.382
R32984 vdd.n8369 vdd.n8355 287.382
R32985 vdd.n8369 vdd.n8348 287.382
R32986 vdd.n8386 vdd.n8348 287.382
R32987 vdd.n8386 vdd.n8349 287.382
R32988 vdd.n8380 vdd.n8349 287.382
R32989 vdd.n8415 vdd.n8405 287.382
R32990 vdd.n8419 vdd.n8405 287.382
R32991 vdd.n8419 vdd.n8398 287.382
R32992 vdd.n8436 vdd.n8398 287.382
R32993 vdd.n8436 vdd.n8399 287.382
R32994 vdd.n8430 vdd.n8399 287.382
R32995 vdd.n8462 vdd.n8452 287.382
R32996 vdd.n8466 vdd.n8452 287.382
R32997 vdd.n8466 vdd.n8445 287.382
R32998 vdd.n8483 vdd.n8445 287.382
R32999 vdd.n8483 vdd.n8446 287.382
R33000 vdd.n8477 vdd.n8446 287.382
R33001 vdd.n8512 vdd.n8502 287.382
R33002 vdd.n8516 vdd.n8502 287.382
R33003 vdd.n8516 vdd.n8495 287.382
R33004 vdd.n8533 vdd.n8495 287.382
R33005 vdd.n8533 vdd.n8496 287.382
R33006 vdd.n8527 vdd.n8496 287.382
R33007 vdd.n8562 vdd.n8552 287.382
R33008 vdd.n8566 vdd.n8552 287.382
R33009 vdd.n8566 vdd.n8545 287.382
R33010 vdd.n8583 vdd.n8545 287.382
R33011 vdd.n8583 vdd.n8546 287.382
R33012 vdd.n8577 vdd.n8546 287.382
R33013 vdd.n8610 vdd.n8600 287.382
R33014 vdd.n8614 vdd.n8600 287.382
R33015 vdd.n8614 vdd.n8593 287.382
R33016 vdd.n8631 vdd.n8593 287.382
R33017 vdd.n8631 vdd.n8594 287.382
R33018 vdd.n8625 vdd.n8594 287.382
R33019 vdd.n7553 vdd.n7513 287.382
R33020 vdd.n7546 vdd.n7513 287.382
R33021 vdd.n7546 vdd.n7519 287.382
R33022 vdd.n7538 vdd.n7519 287.382
R33023 vdd.n7538 vdd.n7522 287.382
R33024 vdd.n7532 vdd.n7522 287.382
R33025 vdd.n8661 vdd.n8651 287.382
R33026 vdd.n8665 vdd.n8651 287.382
R33027 vdd.n8665 vdd.n8644 287.382
R33028 vdd.n8682 vdd.n8644 287.382
R33029 vdd.n8682 vdd.n8645 287.382
R33030 vdd.n8676 vdd.n8645 287.382
R33031 vdd.n8708 vdd.n8698 287.382
R33032 vdd.n8712 vdd.n8698 287.382
R33033 vdd.n8712 vdd.n8691 287.382
R33034 vdd.n8729 vdd.n8691 287.382
R33035 vdd.n8729 vdd.n8692 287.382
R33036 vdd.n8723 vdd.n8692 287.382
R33037 vdd.n8758 vdd.n8748 287.382
R33038 vdd.n8762 vdd.n8748 287.382
R33039 vdd.n8762 vdd.n8741 287.382
R33040 vdd.n8779 vdd.n8741 287.382
R33041 vdd.n8779 vdd.n8742 287.382
R33042 vdd.n8773 vdd.n8742 287.382
R33043 vdd.n8808 vdd.n8798 287.382
R33044 vdd.n8812 vdd.n8798 287.382
R33045 vdd.n8812 vdd.n8791 287.382
R33046 vdd.n8829 vdd.n8791 287.382
R33047 vdd.n8829 vdd.n8792 287.382
R33048 vdd.n8823 vdd.n8792 287.382
R33049 vdd.n8856 vdd.n8846 287.382
R33050 vdd.n8860 vdd.n8846 287.382
R33051 vdd.n8860 vdd.n8839 287.382
R33052 vdd.n8877 vdd.n8839 287.382
R33053 vdd.n8877 vdd.n8840 287.382
R33054 vdd.n8871 vdd.n8840 287.382
R33055 vdd.n8996 vdd.n8992 287.382
R33056 vdd.n9006 vdd.n8992 287.382
R33057 vdd.n9006 vdd.n8985 287.382
R33058 vdd.n9023 vdd.n8985 287.382
R33059 vdd.n9023 vdd.n8986 287.382
R33060 vdd.n9016 vdd.n8986 287.382
R33061 vdd.n8948 vdd.n8944 287.382
R33062 vdd.n8958 vdd.n8944 287.382
R33063 vdd.n8958 vdd.n8937 287.382
R33064 vdd.n8975 vdd.n8937 287.382
R33065 vdd.n8975 vdd.n8938 287.382
R33066 vdd.n8968 vdd.n8938 287.382
R33067 vdd.n9045 vdd.n9041 287.382
R33068 vdd.n9055 vdd.n9041 287.382
R33069 vdd.n9055 vdd.n9034 287.382
R33070 vdd.n9072 vdd.n9034 287.382
R33071 vdd.n9072 vdd.n9035 287.382
R33072 vdd.n9065 vdd.n9035 287.382
R33073 vdd.n9095 vdd.n9091 287.382
R33074 vdd.n9105 vdd.n9091 287.382
R33075 vdd.n9105 vdd.n9084 287.382
R33076 vdd.n9122 vdd.n9084 287.382
R33077 vdd.n9122 vdd.n9085 287.382
R33078 vdd.n9115 vdd.n9085 287.382
R33079 vdd.n9143 vdd.n9139 287.382
R33080 vdd.n9153 vdd.n9139 287.382
R33081 vdd.n9153 vdd.n9132 287.382
R33082 vdd.n9170 vdd.n9132 287.382
R33083 vdd.n9170 vdd.n9133 287.382
R33084 vdd.n9163 vdd.n9133 287.382
R33085 vdd.n7332 vdd.n7320 287.382
R33086 vdd.n7339 vdd.n7320 287.382
R33087 vdd.n7343 vdd.n7339 287.382
R33088 vdd.n7343 vdd.n7342 287.382
R33089 vdd.n7342 vdd.n7315 287.382
R33090 vdd.n7353 vdd.n7315 287.382
R33091 vdd.n9291 vdd.n9287 287.382
R33092 vdd.n9301 vdd.n9287 287.382
R33093 vdd.n9301 vdd.n9280 287.382
R33094 vdd.n9318 vdd.n9280 287.382
R33095 vdd.n9318 vdd.n9281 287.382
R33096 vdd.n9311 vdd.n9281 287.382
R33097 vdd.n9242 vdd.n9238 287.382
R33098 vdd.n9252 vdd.n9238 287.382
R33099 vdd.n9252 vdd.n9231 287.382
R33100 vdd.n9269 vdd.n9231 287.382
R33101 vdd.n9269 vdd.n9232 287.382
R33102 vdd.n9262 vdd.n9232 287.382
R33103 vdd.n9194 vdd.n9190 287.382
R33104 vdd.n9204 vdd.n9190 287.382
R33105 vdd.n9204 vdd.n9183 287.382
R33106 vdd.n9221 vdd.n9183 287.382
R33107 vdd.n9221 vdd.n9184 287.382
R33108 vdd.n9214 vdd.n9184 287.382
R33109 vdd.n9340 vdd.n9336 287.382
R33110 vdd.n9350 vdd.n9336 287.382
R33111 vdd.n9350 vdd.n9329 287.382
R33112 vdd.n9367 vdd.n9329 287.382
R33113 vdd.n9367 vdd.n9330 287.382
R33114 vdd.n9360 vdd.n9330 287.382
R33115 vdd.n9390 vdd.n9386 287.382
R33116 vdd.n9400 vdd.n9386 287.382
R33117 vdd.n9400 vdd.n9379 287.382
R33118 vdd.n9417 vdd.n9379 287.382
R33119 vdd.n9417 vdd.n9380 287.382
R33120 vdd.n9410 vdd.n9380 287.382
R33121 vdd.n9438 vdd.n9434 287.382
R33122 vdd.n9448 vdd.n9434 287.382
R33123 vdd.n9448 vdd.n9427 287.382
R33124 vdd.n9465 vdd.n9427 287.382
R33125 vdd.n9465 vdd.n9428 287.382
R33126 vdd.n9458 vdd.n9428 287.382
R33127 vdd.n9536 vdd.n9532 287.382
R33128 vdd.n9546 vdd.n9532 287.382
R33129 vdd.n9546 vdd.n9525 287.382
R33130 vdd.n9563 vdd.n9525 287.382
R33131 vdd.n9563 vdd.n9526 287.382
R33132 vdd.n9556 vdd.n9526 287.382
R33133 vdd.n9488 vdd.n9484 287.382
R33134 vdd.n9498 vdd.n9484 287.382
R33135 vdd.n9498 vdd.n9477 287.382
R33136 vdd.n9515 vdd.n9477 287.382
R33137 vdd.n9515 vdd.n9478 287.382
R33138 vdd.n9508 vdd.n9478 287.382
R33139 vdd.n9585 vdd.n9581 287.382
R33140 vdd.n9595 vdd.n9581 287.382
R33141 vdd.n9595 vdd.n9574 287.382
R33142 vdd.n9612 vdd.n9574 287.382
R33143 vdd.n9612 vdd.n9575 287.382
R33144 vdd.n9605 vdd.n9575 287.382
R33145 vdd.n9635 vdd.n9631 287.382
R33146 vdd.n9645 vdd.n9631 287.382
R33147 vdd.n9645 vdd.n9624 287.382
R33148 vdd.n9662 vdd.n9624 287.382
R33149 vdd.n9662 vdd.n9625 287.382
R33150 vdd.n9655 vdd.n9625 287.382
R33151 vdd.n9683 vdd.n9679 287.382
R33152 vdd.n9693 vdd.n9679 287.382
R33153 vdd.n9693 vdd.n9672 287.382
R33154 vdd.n9710 vdd.n9672 287.382
R33155 vdd.n9710 vdd.n9673 287.382
R33156 vdd.n9703 vdd.n9673 287.382
R33157 vdd.n7086 vdd.n7074 287.382
R33158 vdd.n7093 vdd.n7074 287.382
R33159 vdd.n7097 vdd.n7093 287.382
R33160 vdd.n7097 vdd.n7096 287.382
R33161 vdd.n7096 vdd.n7069 287.382
R33162 vdd.n7107 vdd.n7069 287.382
R33163 vdd.n9782 vdd.n9778 287.382
R33164 vdd.n9792 vdd.n9778 287.382
R33165 vdd.n9792 vdd.n9771 287.382
R33166 vdd.n9809 vdd.n9771 287.382
R33167 vdd.n9809 vdd.n9772 287.382
R33168 vdd.n9802 vdd.n9772 287.382
R33169 vdd.n9734 vdd.n9730 287.382
R33170 vdd.n9744 vdd.n9730 287.382
R33171 vdd.n9744 vdd.n9723 287.382
R33172 vdd.n9761 vdd.n9723 287.382
R33173 vdd.n9761 vdd.n9724 287.382
R33174 vdd.n9754 vdd.n9724 287.382
R33175 vdd.n9831 vdd.n9827 287.382
R33176 vdd.n9841 vdd.n9827 287.382
R33177 vdd.n9841 vdd.n9820 287.382
R33178 vdd.n9858 vdd.n9820 287.382
R33179 vdd.n9858 vdd.n9821 287.382
R33180 vdd.n9851 vdd.n9821 287.382
R33181 vdd.n9881 vdd.n9877 287.382
R33182 vdd.n9891 vdd.n9877 287.382
R33183 vdd.n9891 vdd.n9870 287.382
R33184 vdd.n9908 vdd.n9870 287.382
R33185 vdd.n9908 vdd.n9871 287.382
R33186 vdd.n9901 vdd.n9871 287.382
R33187 vdd.n9929 vdd.n9925 287.382
R33188 vdd.n9939 vdd.n9925 287.382
R33189 vdd.n9939 vdd.n9918 287.382
R33190 vdd.n9956 vdd.n9918 287.382
R33191 vdd.n9956 vdd.n9919 287.382
R33192 vdd.n9949 vdd.n9919 287.382
R33193 vdd.n3841 vdd.n3837 287.382
R33194 vdd.n3851 vdd.n3837 287.382
R33195 vdd.n3851 vdd.n3830 287.382
R33196 vdd.n3868 vdd.n3830 287.382
R33197 vdd.n3868 vdd.n3831 287.382
R33198 vdd.n3861 vdd.n3831 287.382
R33199 vdd.n3889 vdd.n3885 287.382
R33200 vdd.n3899 vdd.n3885 287.382
R33201 vdd.n3899 vdd.n3878 287.382
R33202 vdd.n3916 vdd.n3878 287.382
R33203 vdd.n3916 vdd.n3879 287.382
R33204 vdd.n3909 vdd.n3879 287.382
R33205 vdd.n3991 vdd.n3987 287.382
R33206 vdd.n4001 vdd.n3987 287.382
R33207 vdd.n4001 vdd.n3980 287.382
R33208 vdd.n4018 vdd.n3980 287.382
R33209 vdd.n4018 vdd.n3981 287.382
R33210 vdd.n4011 vdd.n3981 287.382
R33211 vdd.n4039 vdd.n4035 287.382
R33212 vdd.n4049 vdd.n4035 287.382
R33213 vdd.n4049 vdd.n4028 287.382
R33214 vdd.n4066 vdd.n4028 287.382
R33215 vdd.n4066 vdd.n4029 287.382
R33216 vdd.n4059 vdd.n4029 287.382
R33217 vdd.n4087 vdd.n4083 287.382
R33218 vdd.n4097 vdd.n4083 287.382
R33219 vdd.n4097 vdd.n4076 287.382
R33220 vdd.n4114 vdd.n4076 287.382
R33221 vdd.n4114 vdd.n4077 287.382
R33222 vdd.n4107 vdd.n4077 287.382
R33223 vdd.n4135 vdd.n4131 287.382
R33224 vdd.n4145 vdd.n4131 287.382
R33225 vdd.n4145 vdd.n4124 287.382
R33226 vdd.n4162 vdd.n4124 287.382
R33227 vdd.n4162 vdd.n4125 287.382
R33228 vdd.n4155 vdd.n4125 287.382
R33229 vdd.n4237 vdd.n4233 287.382
R33230 vdd.n4247 vdd.n4233 287.382
R33231 vdd.n4247 vdd.n4226 287.382
R33232 vdd.n4264 vdd.n4226 287.382
R33233 vdd.n4264 vdd.n4227 287.382
R33234 vdd.n4257 vdd.n4227 287.382
R33235 vdd.n5757 vdd.n5753 287.382
R33236 vdd.n5767 vdd.n5753 287.382
R33237 vdd.n5767 vdd.n5746 287.382
R33238 vdd.n5784 vdd.n5746 287.382
R33239 vdd.n5784 vdd.n5747 287.382
R33240 vdd.n5777 vdd.n5747 287.382
R33241 vdd.n4291 vdd.n4281 287.382
R33242 vdd.n4295 vdd.n4281 287.382
R33243 vdd.n4295 vdd.n4274 287.382
R33244 vdd.n4312 vdd.n4274 287.382
R33245 vdd.n4312 vdd.n4275 287.382
R33246 vdd.n4306 vdd.n4275 287.382
R33247 vdd.n4339 vdd.n4329 287.382
R33248 vdd.n4343 vdd.n4329 287.382
R33249 vdd.n4343 vdd.n4322 287.382
R33250 vdd.n4360 vdd.n4322 287.382
R33251 vdd.n4360 vdd.n4323 287.382
R33252 vdd.n4354 vdd.n4323 287.382
R33253 vdd.n4440 vdd.n4430 287.382
R33254 vdd.n4444 vdd.n4430 287.382
R33255 vdd.n4444 vdd.n4423 287.382
R33256 vdd.n4461 vdd.n4423 287.382
R33257 vdd.n4461 vdd.n4424 287.382
R33258 vdd.n4455 vdd.n4424 287.382
R33259 vdd.n4488 vdd.n4478 287.382
R33260 vdd.n4492 vdd.n4478 287.382
R33261 vdd.n4492 vdd.n4471 287.382
R33262 vdd.n4509 vdd.n4471 287.382
R33263 vdd.n4509 vdd.n4472 287.382
R33264 vdd.n4503 vdd.n4472 287.382
R33265 vdd.n4536 vdd.n4526 287.382
R33266 vdd.n4540 vdd.n4526 287.382
R33267 vdd.n4540 vdd.n4519 287.382
R33268 vdd.n4557 vdd.n4519 287.382
R33269 vdd.n4557 vdd.n4520 287.382
R33270 vdd.n4551 vdd.n4520 287.382
R33271 vdd.n4584 vdd.n4574 287.382
R33272 vdd.n4588 vdd.n4574 287.382
R33273 vdd.n4588 vdd.n4567 287.382
R33274 vdd.n4605 vdd.n4567 287.382
R33275 vdd.n4605 vdd.n4568 287.382
R33276 vdd.n4599 vdd.n4568 287.382
R33277 vdd.n4685 vdd.n4675 287.382
R33278 vdd.n4689 vdd.n4675 287.382
R33279 vdd.n4689 vdd.n4668 287.382
R33280 vdd.n4706 vdd.n4668 287.382
R33281 vdd.n4706 vdd.n4669 287.382
R33282 vdd.n4700 vdd.n4669 287.382
R33283 vdd.n3798 vdd.n3788 287.382
R33284 vdd.n3802 vdd.n3788 287.382
R33285 vdd.n3802 vdd.n3781 287.382
R33286 vdd.n3819 vdd.n3781 287.382
R33287 vdd.n3819 vdd.n3782 287.382
R33288 vdd.n3813 vdd.n3782 287.382
R33289 vdd.n4733 vdd.n4723 287.382
R33290 vdd.n4737 vdd.n4723 287.382
R33291 vdd.n4737 vdd.n4716 287.382
R33292 vdd.n4754 vdd.n4716 287.382
R33293 vdd.n4754 vdd.n4717 287.382
R33294 vdd.n4748 vdd.n4717 287.382
R33295 vdd.n4780 vdd.n4770 287.382
R33296 vdd.n4784 vdd.n4770 287.382
R33297 vdd.n4784 vdd.n4763 287.382
R33298 vdd.n4801 vdd.n4763 287.382
R33299 vdd.n4801 vdd.n4764 287.382
R33300 vdd.n4795 vdd.n4764 287.382
R33301 vdd.n4830 vdd.n4820 287.382
R33302 vdd.n4834 vdd.n4820 287.382
R33303 vdd.n4834 vdd.n4813 287.382
R33304 vdd.n4851 vdd.n4813 287.382
R33305 vdd.n4851 vdd.n4814 287.382
R33306 vdd.n4845 vdd.n4814 287.382
R33307 vdd.n4880 vdd.n4870 287.382
R33308 vdd.n4884 vdd.n4870 287.382
R33309 vdd.n4884 vdd.n4863 287.382
R33310 vdd.n4901 vdd.n4863 287.382
R33311 vdd.n4901 vdd.n4864 287.382
R33312 vdd.n4895 vdd.n4864 287.382
R33313 vdd.n4928 vdd.n4918 287.382
R33314 vdd.n4932 vdd.n4918 287.382
R33315 vdd.n4932 vdd.n4911 287.382
R33316 vdd.n4949 vdd.n4911 287.382
R33317 vdd.n4949 vdd.n4912 287.382
R33318 vdd.n4943 vdd.n4912 287.382
R33319 vdd.n4656 vdd.n4616 287.382
R33320 vdd.n4649 vdd.n4616 287.382
R33321 vdd.n4649 vdd.n4622 287.382
R33322 vdd.n4641 vdd.n4622 287.382
R33323 vdd.n4641 vdd.n4625 287.382
R33324 vdd.n4635 vdd.n4625 287.382
R33325 vdd.n4979 vdd.n4969 287.382
R33326 vdd.n4983 vdd.n4969 287.382
R33327 vdd.n4983 vdd.n4962 287.382
R33328 vdd.n5000 vdd.n4962 287.382
R33329 vdd.n5000 vdd.n4963 287.382
R33330 vdd.n4994 vdd.n4963 287.382
R33331 vdd.n5026 vdd.n5016 287.382
R33332 vdd.n5030 vdd.n5016 287.382
R33333 vdd.n5030 vdd.n5009 287.382
R33334 vdd.n5047 vdd.n5009 287.382
R33335 vdd.n5047 vdd.n5010 287.382
R33336 vdd.n5041 vdd.n5010 287.382
R33337 vdd.n5074 vdd.n5064 287.382
R33338 vdd.n5078 vdd.n5064 287.382
R33339 vdd.n5078 vdd.n5057 287.382
R33340 vdd.n5095 vdd.n5057 287.382
R33341 vdd.n5095 vdd.n5058 287.382
R33342 vdd.n5089 vdd.n5058 287.382
R33343 vdd.n5125 vdd.n5115 287.382
R33344 vdd.n5129 vdd.n5115 287.382
R33345 vdd.n5129 vdd.n5108 287.382
R33346 vdd.n5146 vdd.n5108 287.382
R33347 vdd.n5146 vdd.n5109 287.382
R33348 vdd.n5140 vdd.n5109 287.382
R33349 vdd.n5175 vdd.n5165 287.382
R33350 vdd.n5179 vdd.n5165 287.382
R33351 vdd.n5179 vdd.n5158 287.382
R33352 vdd.n5196 vdd.n5158 287.382
R33353 vdd.n5196 vdd.n5159 287.382
R33354 vdd.n5190 vdd.n5159 287.382
R33355 vdd.n5223 vdd.n5213 287.382
R33356 vdd.n5227 vdd.n5213 287.382
R33357 vdd.n5227 vdd.n5206 287.382
R33358 vdd.n5244 vdd.n5206 287.382
R33359 vdd.n5244 vdd.n5207 287.382
R33360 vdd.n5238 vdd.n5207 287.382
R33361 vdd.n5273 vdd.n5263 287.382
R33362 vdd.n5277 vdd.n5263 287.382
R33363 vdd.n5277 vdd.n5256 287.382
R33364 vdd.n5294 vdd.n5256 287.382
R33365 vdd.n5294 vdd.n5257 287.382
R33366 vdd.n5288 vdd.n5257 287.382
R33367 vdd.n5320 vdd.n5310 287.382
R33368 vdd.n5324 vdd.n5310 287.382
R33369 vdd.n5324 vdd.n5303 287.382
R33370 vdd.n5341 vdd.n5303 287.382
R33371 vdd.n5341 vdd.n5304 287.382
R33372 vdd.n5335 vdd.n5304 287.382
R33373 vdd.n5370 vdd.n5360 287.382
R33374 vdd.n5374 vdd.n5360 287.382
R33375 vdd.n5374 vdd.n5353 287.382
R33376 vdd.n5391 vdd.n5353 287.382
R33377 vdd.n5391 vdd.n5354 287.382
R33378 vdd.n5385 vdd.n5354 287.382
R33379 vdd.n5420 vdd.n5410 287.382
R33380 vdd.n5424 vdd.n5410 287.382
R33381 vdd.n5424 vdd.n5403 287.382
R33382 vdd.n5441 vdd.n5403 287.382
R33383 vdd.n5441 vdd.n5404 287.382
R33384 vdd.n5435 vdd.n5404 287.382
R33385 vdd.n5468 vdd.n5458 287.382
R33386 vdd.n5472 vdd.n5458 287.382
R33387 vdd.n5472 vdd.n5451 287.382
R33388 vdd.n5489 vdd.n5451 287.382
R33389 vdd.n5489 vdd.n5452 287.382
R33390 vdd.n5483 vdd.n5452 287.382
R33391 vdd.n4411 vdd.n4371 287.382
R33392 vdd.n4404 vdd.n4371 287.382
R33393 vdd.n4404 vdd.n4377 287.382
R33394 vdd.n4396 vdd.n4377 287.382
R33395 vdd.n4396 vdd.n4380 287.382
R33396 vdd.n4390 vdd.n4380 287.382
R33397 vdd.n5519 vdd.n5509 287.382
R33398 vdd.n5523 vdd.n5509 287.382
R33399 vdd.n5523 vdd.n5502 287.382
R33400 vdd.n5540 vdd.n5502 287.382
R33401 vdd.n5540 vdd.n5503 287.382
R33402 vdd.n5534 vdd.n5503 287.382
R33403 vdd.n5566 vdd.n5556 287.382
R33404 vdd.n5570 vdd.n5556 287.382
R33405 vdd.n5570 vdd.n5549 287.382
R33406 vdd.n5587 vdd.n5549 287.382
R33407 vdd.n5587 vdd.n5550 287.382
R33408 vdd.n5581 vdd.n5550 287.382
R33409 vdd.n5616 vdd.n5606 287.382
R33410 vdd.n5620 vdd.n5606 287.382
R33411 vdd.n5620 vdd.n5599 287.382
R33412 vdd.n5637 vdd.n5599 287.382
R33413 vdd.n5637 vdd.n5600 287.382
R33414 vdd.n5631 vdd.n5600 287.382
R33415 vdd.n5666 vdd.n5656 287.382
R33416 vdd.n5670 vdd.n5656 287.382
R33417 vdd.n5670 vdd.n5649 287.382
R33418 vdd.n5687 vdd.n5649 287.382
R33419 vdd.n5687 vdd.n5650 287.382
R33420 vdd.n5681 vdd.n5650 287.382
R33421 vdd.n5714 vdd.n5704 287.382
R33422 vdd.n5718 vdd.n5704 287.382
R33423 vdd.n5718 vdd.n5697 287.382
R33424 vdd.n5735 vdd.n5697 287.382
R33425 vdd.n5735 vdd.n5698 287.382
R33426 vdd.n5729 vdd.n5698 287.382
R33427 vdd.n5854 vdd.n5850 287.382
R33428 vdd.n5864 vdd.n5850 287.382
R33429 vdd.n5864 vdd.n5843 287.382
R33430 vdd.n5881 vdd.n5843 287.382
R33431 vdd.n5881 vdd.n5844 287.382
R33432 vdd.n5874 vdd.n5844 287.382
R33433 vdd.n5806 vdd.n5802 287.382
R33434 vdd.n5816 vdd.n5802 287.382
R33435 vdd.n5816 vdd.n5795 287.382
R33436 vdd.n5833 vdd.n5795 287.382
R33437 vdd.n5833 vdd.n5796 287.382
R33438 vdd.n5826 vdd.n5796 287.382
R33439 vdd.n5903 vdd.n5899 287.382
R33440 vdd.n5913 vdd.n5899 287.382
R33441 vdd.n5913 vdd.n5892 287.382
R33442 vdd.n5930 vdd.n5892 287.382
R33443 vdd.n5930 vdd.n5893 287.382
R33444 vdd.n5923 vdd.n5893 287.382
R33445 vdd.n5953 vdd.n5949 287.382
R33446 vdd.n5963 vdd.n5949 287.382
R33447 vdd.n5963 vdd.n5942 287.382
R33448 vdd.n5980 vdd.n5942 287.382
R33449 vdd.n5980 vdd.n5943 287.382
R33450 vdd.n5973 vdd.n5943 287.382
R33451 vdd.n6001 vdd.n5997 287.382
R33452 vdd.n6011 vdd.n5997 287.382
R33453 vdd.n6011 vdd.n5990 287.382
R33454 vdd.n6028 vdd.n5990 287.382
R33455 vdd.n6028 vdd.n5991 287.382
R33456 vdd.n6021 vdd.n5991 287.382
R33457 vdd.n4190 vdd.n4178 287.382
R33458 vdd.n4197 vdd.n4178 287.382
R33459 vdd.n4201 vdd.n4197 287.382
R33460 vdd.n4201 vdd.n4200 287.382
R33461 vdd.n4200 vdd.n4173 287.382
R33462 vdd.n4211 vdd.n4173 287.382
R33463 vdd.n6149 vdd.n6145 287.382
R33464 vdd.n6159 vdd.n6145 287.382
R33465 vdd.n6159 vdd.n6138 287.382
R33466 vdd.n6176 vdd.n6138 287.382
R33467 vdd.n6176 vdd.n6139 287.382
R33468 vdd.n6169 vdd.n6139 287.382
R33469 vdd.n6100 vdd.n6096 287.382
R33470 vdd.n6110 vdd.n6096 287.382
R33471 vdd.n6110 vdd.n6089 287.382
R33472 vdd.n6127 vdd.n6089 287.382
R33473 vdd.n6127 vdd.n6090 287.382
R33474 vdd.n6120 vdd.n6090 287.382
R33475 vdd.n6052 vdd.n6048 287.382
R33476 vdd.n6062 vdd.n6048 287.382
R33477 vdd.n6062 vdd.n6041 287.382
R33478 vdd.n6079 vdd.n6041 287.382
R33479 vdd.n6079 vdd.n6042 287.382
R33480 vdd.n6072 vdd.n6042 287.382
R33481 vdd.n6198 vdd.n6194 287.382
R33482 vdd.n6208 vdd.n6194 287.382
R33483 vdd.n6208 vdd.n6187 287.382
R33484 vdd.n6225 vdd.n6187 287.382
R33485 vdd.n6225 vdd.n6188 287.382
R33486 vdd.n6218 vdd.n6188 287.382
R33487 vdd.n6248 vdd.n6244 287.382
R33488 vdd.n6258 vdd.n6244 287.382
R33489 vdd.n6258 vdd.n6237 287.382
R33490 vdd.n6275 vdd.n6237 287.382
R33491 vdd.n6275 vdd.n6238 287.382
R33492 vdd.n6268 vdd.n6238 287.382
R33493 vdd.n6296 vdd.n6292 287.382
R33494 vdd.n6306 vdd.n6292 287.382
R33495 vdd.n6306 vdd.n6285 287.382
R33496 vdd.n6323 vdd.n6285 287.382
R33497 vdd.n6323 vdd.n6286 287.382
R33498 vdd.n6316 vdd.n6286 287.382
R33499 vdd.n6394 vdd.n6390 287.382
R33500 vdd.n6404 vdd.n6390 287.382
R33501 vdd.n6404 vdd.n6383 287.382
R33502 vdd.n6421 vdd.n6383 287.382
R33503 vdd.n6421 vdd.n6384 287.382
R33504 vdd.n6414 vdd.n6384 287.382
R33505 vdd.n6346 vdd.n6342 287.382
R33506 vdd.n6356 vdd.n6342 287.382
R33507 vdd.n6356 vdd.n6335 287.382
R33508 vdd.n6373 vdd.n6335 287.382
R33509 vdd.n6373 vdd.n6336 287.382
R33510 vdd.n6366 vdd.n6336 287.382
R33511 vdd.n6443 vdd.n6439 287.382
R33512 vdd.n6453 vdd.n6439 287.382
R33513 vdd.n6453 vdd.n6432 287.382
R33514 vdd.n6470 vdd.n6432 287.382
R33515 vdd.n6470 vdd.n6433 287.382
R33516 vdd.n6463 vdd.n6433 287.382
R33517 vdd.n6493 vdd.n6489 287.382
R33518 vdd.n6503 vdd.n6489 287.382
R33519 vdd.n6503 vdd.n6482 287.382
R33520 vdd.n6520 vdd.n6482 287.382
R33521 vdd.n6520 vdd.n6483 287.382
R33522 vdd.n6513 vdd.n6483 287.382
R33523 vdd.n6541 vdd.n6537 287.382
R33524 vdd.n6551 vdd.n6537 287.382
R33525 vdd.n6551 vdd.n6530 287.382
R33526 vdd.n6568 vdd.n6530 287.382
R33527 vdd.n6568 vdd.n6531 287.382
R33528 vdd.n6561 vdd.n6531 287.382
R33529 vdd.n3944 vdd.n3932 287.382
R33530 vdd.n3951 vdd.n3932 287.382
R33531 vdd.n3955 vdd.n3951 287.382
R33532 vdd.n3955 vdd.n3954 287.382
R33533 vdd.n3954 vdd.n3927 287.382
R33534 vdd.n3965 vdd.n3927 287.382
R33535 vdd.n6640 vdd.n6636 287.382
R33536 vdd.n6650 vdd.n6636 287.382
R33537 vdd.n6650 vdd.n6629 287.382
R33538 vdd.n6667 vdd.n6629 287.382
R33539 vdd.n6667 vdd.n6630 287.382
R33540 vdd.n6660 vdd.n6630 287.382
R33541 vdd.n6592 vdd.n6588 287.382
R33542 vdd.n6602 vdd.n6588 287.382
R33543 vdd.n6602 vdd.n6581 287.382
R33544 vdd.n6619 vdd.n6581 287.382
R33545 vdd.n6619 vdd.n6582 287.382
R33546 vdd.n6612 vdd.n6582 287.382
R33547 vdd.n6689 vdd.n6685 287.382
R33548 vdd.n6699 vdd.n6685 287.382
R33549 vdd.n6699 vdd.n6678 287.382
R33550 vdd.n6716 vdd.n6678 287.382
R33551 vdd.n6716 vdd.n6679 287.382
R33552 vdd.n6709 vdd.n6679 287.382
R33553 vdd.n6739 vdd.n6735 287.382
R33554 vdd.n6749 vdd.n6735 287.382
R33555 vdd.n6749 vdd.n6728 287.382
R33556 vdd.n6766 vdd.n6728 287.382
R33557 vdd.n6766 vdd.n6729 287.382
R33558 vdd.n6759 vdd.n6729 287.382
R33559 vdd.n6787 vdd.n6783 287.382
R33560 vdd.n6797 vdd.n6783 287.382
R33561 vdd.n6797 vdd.n6776 287.382
R33562 vdd.n6814 vdd.n6776 287.382
R33563 vdd.n6814 vdd.n6777 287.382
R33564 vdd.n6807 vdd.n6777 287.382
R33565 vdd.n699 vdd.n695 287.382
R33566 vdd.n709 vdd.n695 287.382
R33567 vdd.n709 vdd.n688 287.382
R33568 vdd.n726 vdd.n688 287.382
R33569 vdd.n726 vdd.n689 287.382
R33570 vdd.n719 vdd.n689 287.382
R33571 vdd.n747 vdd.n743 287.382
R33572 vdd.n757 vdd.n743 287.382
R33573 vdd.n757 vdd.n736 287.382
R33574 vdd.n774 vdd.n736 287.382
R33575 vdd.n774 vdd.n737 287.382
R33576 vdd.n767 vdd.n737 287.382
R33577 vdd.n849 vdd.n845 287.382
R33578 vdd.n859 vdd.n845 287.382
R33579 vdd.n859 vdd.n838 287.382
R33580 vdd.n876 vdd.n838 287.382
R33581 vdd.n876 vdd.n839 287.382
R33582 vdd.n869 vdd.n839 287.382
R33583 vdd.n897 vdd.n893 287.382
R33584 vdd.n907 vdd.n893 287.382
R33585 vdd.n907 vdd.n886 287.382
R33586 vdd.n924 vdd.n886 287.382
R33587 vdd.n924 vdd.n887 287.382
R33588 vdd.n917 vdd.n887 287.382
R33589 vdd.n945 vdd.n941 287.382
R33590 vdd.n955 vdd.n941 287.382
R33591 vdd.n955 vdd.n934 287.382
R33592 vdd.n972 vdd.n934 287.382
R33593 vdd.n972 vdd.n935 287.382
R33594 vdd.n965 vdd.n935 287.382
R33595 vdd.n993 vdd.n989 287.382
R33596 vdd.n1003 vdd.n989 287.382
R33597 vdd.n1003 vdd.n982 287.382
R33598 vdd.n1020 vdd.n982 287.382
R33599 vdd.n1020 vdd.n983 287.382
R33600 vdd.n1013 vdd.n983 287.382
R33601 vdd.n1095 vdd.n1091 287.382
R33602 vdd.n1105 vdd.n1091 287.382
R33603 vdd.n1105 vdd.n1084 287.382
R33604 vdd.n1122 vdd.n1084 287.382
R33605 vdd.n1122 vdd.n1085 287.382
R33606 vdd.n1115 vdd.n1085 287.382
R33607 vdd.n2615 vdd.n2611 287.382
R33608 vdd.n2625 vdd.n2611 287.382
R33609 vdd.n2625 vdd.n2604 287.382
R33610 vdd.n2642 vdd.n2604 287.382
R33611 vdd.n2642 vdd.n2605 287.382
R33612 vdd.n2635 vdd.n2605 287.382
R33613 vdd.n1149 vdd.n1139 287.382
R33614 vdd.n1153 vdd.n1139 287.382
R33615 vdd.n1153 vdd.n1132 287.382
R33616 vdd.n1170 vdd.n1132 287.382
R33617 vdd.n1170 vdd.n1133 287.382
R33618 vdd.n1164 vdd.n1133 287.382
R33619 vdd.n1197 vdd.n1187 287.382
R33620 vdd.n1201 vdd.n1187 287.382
R33621 vdd.n1201 vdd.n1180 287.382
R33622 vdd.n1218 vdd.n1180 287.382
R33623 vdd.n1218 vdd.n1181 287.382
R33624 vdd.n1212 vdd.n1181 287.382
R33625 vdd.n1298 vdd.n1288 287.382
R33626 vdd.n1302 vdd.n1288 287.382
R33627 vdd.n1302 vdd.n1281 287.382
R33628 vdd.n1319 vdd.n1281 287.382
R33629 vdd.n1319 vdd.n1282 287.382
R33630 vdd.n1313 vdd.n1282 287.382
R33631 vdd.n1346 vdd.n1336 287.382
R33632 vdd.n1350 vdd.n1336 287.382
R33633 vdd.n1350 vdd.n1329 287.382
R33634 vdd.n1367 vdd.n1329 287.382
R33635 vdd.n1367 vdd.n1330 287.382
R33636 vdd.n1361 vdd.n1330 287.382
R33637 vdd.n1394 vdd.n1384 287.382
R33638 vdd.n1398 vdd.n1384 287.382
R33639 vdd.n1398 vdd.n1377 287.382
R33640 vdd.n1415 vdd.n1377 287.382
R33641 vdd.n1415 vdd.n1378 287.382
R33642 vdd.n1409 vdd.n1378 287.382
R33643 vdd.n1442 vdd.n1432 287.382
R33644 vdd.n1446 vdd.n1432 287.382
R33645 vdd.n1446 vdd.n1425 287.382
R33646 vdd.n1463 vdd.n1425 287.382
R33647 vdd.n1463 vdd.n1426 287.382
R33648 vdd.n1457 vdd.n1426 287.382
R33649 vdd.n1543 vdd.n1533 287.382
R33650 vdd.n1547 vdd.n1533 287.382
R33651 vdd.n1547 vdd.n1526 287.382
R33652 vdd.n1564 vdd.n1526 287.382
R33653 vdd.n1564 vdd.n1527 287.382
R33654 vdd.n1558 vdd.n1527 287.382
R33655 vdd.n656 vdd.n646 287.382
R33656 vdd.n660 vdd.n646 287.382
R33657 vdd.n660 vdd.n639 287.382
R33658 vdd.n677 vdd.n639 287.382
R33659 vdd.n677 vdd.n640 287.382
R33660 vdd.n671 vdd.n640 287.382
R33661 vdd.n1591 vdd.n1581 287.382
R33662 vdd.n1595 vdd.n1581 287.382
R33663 vdd.n1595 vdd.n1574 287.382
R33664 vdd.n1612 vdd.n1574 287.382
R33665 vdd.n1612 vdd.n1575 287.382
R33666 vdd.n1606 vdd.n1575 287.382
R33667 vdd.n1638 vdd.n1628 287.382
R33668 vdd.n1642 vdd.n1628 287.382
R33669 vdd.n1642 vdd.n1621 287.382
R33670 vdd.n1659 vdd.n1621 287.382
R33671 vdd.n1659 vdd.n1622 287.382
R33672 vdd.n1653 vdd.n1622 287.382
R33673 vdd.n1688 vdd.n1678 287.382
R33674 vdd.n1692 vdd.n1678 287.382
R33675 vdd.n1692 vdd.n1671 287.382
R33676 vdd.n1709 vdd.n1671 287.382
R33677 vdd.n1709 vdd.n1672 287.382
R33678 vdd.n1703 vdd.n1672 287.382
R33679 vdd.n1738 vdd.n1728 287.382
R33680 vdd.n1742 vdd.n1728 287.382
R33681 vdd.n1742 vdd.n1721 287.382
R33682 vdd.n1759 vdd.n1721 287.382
R33683 vdd.n1759 vdd.n1722 287.382
R33684 vdd.n1753 vdd.n1722 287.382
R33685 vdd.n1786 vdd.n1776 287.382
R33686 vdd.n1790 vdd.n1776 287.382
R33687 vdd.n1790 vdd.n1769 287.382
R33688 vdd.n1807 vdd.n1769 287.382
R33689 vdd.n1807 vdd.n1770 287.382
R33690 vdd.n1801 vdd.n1770 287.382
R33691 vdd.n1514 vdd.n1474 287.382
R33692 vdd.n1507 vdd.n1474 287.382
R33693 vdd.n1507 vdd.n1480 287.382
R33694 vdd.n1499 vdd.n1480 287.382
R33695 vdd.n1499 vdd.n1483 287.382
R33696 vdd.n1493 vdd.n1483 287.382
R33697 vdd.n1837 vdd.n1827 287.382
R33698 vdd.n1841 vdd.n1827 287.382
R33699 vdd.n1841 vdd.n1820 287.382
R33700 vdd.n1858 vdd.n1820 287.382
R33701 vdd.n1858 vdd.n1821 287.382
R33702 vdd.n1852 vdd.n1821 287.382
R33703 vdd.n1884 vdd.n1874 287.382
R33704 vdd.n1888 vdd.n1874 287.382
R33705 vdd.n1888 vdd.n1867 287.382
R33706 vdd.n1905 vdd.n1867 287.382
R33707 vdd.n1905 vdd.n1868 287.382
R33708 vdd.n1899 vdd.n1868 287.382
R33709 vdd.n1932 vdd.n1922 287.382
R33710 vdd.n1936 vdd.n1922 287.382
R33711 vdd.n1936 vdd.n1915 287.382
R33712 vdd.n1953 vdd.n1915 287.382
R33713 vdd.n1953 vdd.n1916 287.382
R33714 vdd.n1947 vdd.n1916 287.382
R33715 vdd.n1983 vdd.n1973 287.382
R33716 vdd.n1987 vdd.n1973 287.382
R33717 vdd.n1987 vdd.n1966 287.382
R33718 vdd.n2004 vdd.n1966 287.382
R33719 vdd.n2004 vdd.n1967 287.382
R33720 vdd.n1998 vdd.n1967 287.382
R33721 vdd.n2033 vdd.n2023 287.382
R33722 vdd.n2037 vdd.n2023 287.382
R33723 vdd.n2037 vdd.n2016 287.382
R33724 vdd.n2054 vdd.n2016 287.382
R33725 vdd.n2054 vdd.n2017 287.382
R33726 vdd.n2048 vdd.n2017 287.382
R33727 vdd.n2081 vdd.n2071 287.382
R33728 vdd.n2085 vdd.n2071 287.382
R33729 vdd.n2085 vdd.n2064 287.382
R33730 vdd.n2102 vdd.n2064 287.382
R33731 vdd.n2102 vdd.n2065 287.382
R33732 vdd.n2096 vdd.n2065 287.382
R33733 vdd.n2131 vdd.n2121 287.382
R33734 vdd.n2135 vdd.n2121 287.382
R33735 vdd.n2135 vdd.n2114 287.382
R33736 vdd.n2152 vdd.n2114 287.382
R33737 vdd.n2152 vdd.n2115 287.382
R33738 vdd.n2146 vdd.n2115 287.382
R33739 vdd.n2178 vdd.n2168 287.382
R33740 vdd.n2182 vdd.n2168 287.382
R33741 vdd.n2182 vdd.n2161 287.382
R33742 vdd.n2199 vdd.n2161 287.382
R33743 vdd.n2199 vdd.n2162 287.382
R33744 vdd.n2193 vdd.n2162 287.382
R33745 vdd.n2228 vdd.n2218 287.382
R33746 vdd.n2232 vdd.n2218 287.382
R33747 vdd.n2232 vdd.n2211 287.382
R33748 vdd.n2249 vdd.n2211 287.382
R33749 vdd.n2249 vdd.n2212 287.382
R33750 vdd.n2243 vdd.n2212 287.382
R33751 vdd.n2278 vdd.n2268 287.382
R33752 vdd.n2282 vdd.n2268 287.382
R33753 vdd.n2282 vdd.n2261 287.382
R33754 vdd.n2299 vdd.n2261 287.382
R33755 vdd.n2299 vdd.n2262 287.382
R33756 vdd.n2293 vdd.n2262 287.382
R33757 vdd.n2326 vdd.n2316 287.382
R33758 vdd.n2330 vdd.n2316 287.382
R33759 vdd.n2330 vdd.n2309 287.382
R33760 vdd.n2347 vdd.n2309 287.382
R33761 vdd.n2347 vdd.n2310 287.382
R33762 vdd.n2341 vdd.n2310 287.382
R33763 vdd.n1269 vdd.n1229 287.382
R33764 vdd.n1262 vdd.n1229 287.382
R33765 vdd.n1262 vdd.n1235 287.382
R33766 vdd.n1254 vdd.n1235 287.382
R33767 vdd.n1254 vdd.n1238 287.382
R33768 vdd.n1248 vdd.n1238 287.382
R33769 vdd.n2377 vdd.n2367 287.382
R33770 vdd.n2381 vdd.n2367 287.382
R33771 vdd.n2381 vdd.n2360 287.382
R33772 vdd.n2398 vdd.n2360 287.382
R33773 vdd.n2398 vdd.n2361 287.382
R33774 vdd.n2392 vdd.n2361 287.382
R33775 vdd.n2424 vdd.n2414 287.382
R33776 vdd.n2428 vdd.n2414 287.382
R33777 vdd.n2428 vdd.n2407 287.382
R33778 vdd.n2445 vdd.n2407 287.382
R33779 vdd.n2445 vdd.n2408 287.382
R33780 vdd.n2439 vdd.n2408 287.382
R33781 vdd.n2474 vdd.n2464 287.382
R33782 vdd.n2478 vdd.n2464 287.382
R33783 vdd.n2478 vdd.n2457 287.382
R33784 vdd.n2495 vdd.n2457 287.382
R33785 vdd.n2495 vdd.n2458 287.382
R33786 vdd.n2489 vdd.n2458 287.382
R33787 vdd.n2524 vdd.n2514 287.382
R33788 vdd.n2528 vdd.n2514 287.382
R33789 vdd.n2528 vdd.n2507 287.382
R33790 vdd.n2545 vdd.n2507 287.382
R33791 vdd.n2545 vdd.n2508 287.382
R33792 vdd.n2539 vdd.n2508 287.382
R33793 vdd.n2572 vdd.n2562 287.382
R33794 vdd.n2576 vdd.n2562 287.382
R33795 vdd.n2576 vdd.n2555 287.382
R33796 vdd.n2593 vdd.n2555 287.382
R33797 vdd.n2593 vdd.n2556 287.382
R33798 vdd.n2587 vdd.n2556 287.382
R33799 vdd.n2712 vdd.n2708 287.382
R33800 vdd.n2722 vdd.n2708 287.382
R33801 vdd.n2722 vdd.n2701 287.382
R33802 vdd.n2739 vdd.n2701 287.382
R33803 vdd.n2739 vdd.n2702 287.382
R33804 vdd.n2732 vdd.n2702 287.382
R33805 vdd.n2664 vdd.n2660 287.382
R33806 vdd.n2674 vdd.n2660 287.382
R33807 vdd.n2674 vdd.n2653 287.382
R33808 vdd.n2691 vdd.n2653 287.382
R33809 vdd.n2691 vdd.n2654 287.382
R33810 vdd.n2684 vdd.n2654 287.382
R33811 vdd.n2761 vdd.n2757 287.382
R33812 vdd.n2771 vdd.n2757 287.382
R33813 vdd.n2771 vdd.n2750 287.382
R33814 vdd.n2788 vdd.n2750 287.382
R33815 vdd.n2788 vdd.n2751 287.382
R33816 vdd.n2781 vdd.n2751 287.382
R33817 vdd.n2811 vdd.n2807 287.382
R33818 vdd.n2821 vdd.n2807 287.382
R33819 vdd.n2821 vdd.n2800 287.382
R33820 vdd.n2838 vdd.n2800 287.382
R33821 vdd.n2838 vdd.n2801 287.382
R33822 vdd.n2831 vdd.n2801 287.382
R33823 vdd.n2859 vdd.n2855 287.382
R33824 vdd.n2869 vdd.n2855 287.382
R33825 vdd.n2869 vdd.n2848 287.382
R33826 vdd.n2886 vdd.n2848 287.382
R33827 vdd.n2886 vdd.n2849 287.382
R33828 vdd.n2879 vdd.n2849 287.382
R33829 vdd.n1048 vdd.n1036 287.382
R33830 vdd.n1055 vdd.n1036 287.382
R33831 vdd.n1059 vdd.n1055 287.382
R33832 vdd.n1059 vdd.n1058 287.382
R33833 vdd.n1058 vdd.n1031 287.382
R33834 vdd.n1069 vdd.n1031 287.382
R33835 vdd.n3007 vdd.n3003 287.382
R33836 vdd.n3017 vdd.n3003 287.382
R33837 vdd.n3017 vdd.n2996 287.382
R33838 vdd.n3034 vdd.n2996 287.382
R33839 vdd.n3034 vdd.n2997 287.382
R33840 vdd.n3027 vdd.n2997 287.382
R33841 vdd.n2958 vdd.n2954 287.382
R33842 vdd.n2968 vdd.n2954 287.382
R33843 vdd.n2968 vdd.n2947 287.382
R33844 vdd.n2985 vdd.n2947 287.382
R33845 vdd.n2985 vdd.n2948 287.382
R33846 vdd.n2978 vdd.n2948 287.382
R33847 vdd.n2910 vdd.n2906 287.382
R33848 vdd.n2920 vdd.n2906 287.382
R33849 vdd.n2920 vdd.n2899 287.382
R33850 vdd.n2937 vdd.n2899 287.382
R33851 vdd.n2937 vdd.n2900 287.382
R33852 vdd.n2930 vdd.n2900 287.382
R33853 vdd.n3056 vdd.n3052 287.382
R33854 vdd.n3066 vdd.n3052 287.382
R33855 vdd.n3066 vdd.n3045 287.382
R33856 vdd.n3083 vdd.n3045 287.382
R33857 vdd.n3083 vdd.n3046 287.382
R33858 vdd.n3076 vdd.n3046 287.382
R33859 vdd.n3106 vdd.n3102 287.382
R33860 vdd.n3116 vdd.n3102 287.382
R33861 vdd.n3116 vdd.n3095 287.382
R33862 vdd.n3133 vdd.n3095 287.382
R33863 vdd.n3133 vdd.n3096 287.382
R33864 vdd.n3126 vdd.n3096 287.382
R33865 vdd.n3154 vdd.n3150 287.382
R33866 vdd.n3164 vdd.n3150 287.382
R33867 vdd.n3164 vdd.n3143 287.382
R33868 vdd.n3181 vdd.n3143 287.382
R33869 vdd.n3181 vdd.n3144 287.382
R33870 vdd.n3174 vdd.n3144 287.382
R33871 vdd.n3252 vdd.n3248 287.382
R33872 vdd.n3262 vdd.n3248 287.382
R33873 vdd.n3262 vdd.n3241 287.382
R33874 vdd.n3279 vdd.n3241 287.382
R33875 vdd.n3279 vdd.n3242 287.382
R33876 vdd.n3272 vdd.n3242 287.382
R33877 vdd.n3204 vdd.n3200 287.382
R33878 vdd.n3214 vdd.n3200 287.382
R33879 vdd.n3214 vdd.n3193 287.382
R33880 vdd.n3231 vdd.n3193 287.382
R33881 vdd.n3231 vdd.n3194 287.382
R33882 vdd.n3224 vdd.n3194 287.382
R33883 vdd.n3301 vdd.n3297 287.382
R33884 vdd.n3311 vdd.n3297 287.382
R33885 vdd.n3311 vdd.n3290 287.382
R33886 vdd.n3328 vdd.n3290 287.382
R33887 vdd.n3328 vdd.n3291 287.382
R33888 vdd.n3321 vdd.n3291 287.382
R33889 vdd.n3351 vdd.n3347 287.382
R33890 vdd.n3361 vdd.n3347 287.382
R33891 vdd.n3361 vdd.n3340 287.382
R33892 vdd.n3378 vdd.n3340 287.382
R33893 vdd.n3378 vdd.n3341 287.382
R33894 vdd.n3371 vdd.n3341 287.382
R33895 vdd.n3399 vdd.n3395 287.382
R33896 vdd.n3409 vdd.n3395 287.382
R33897 vdd.n3409 vdd.n3388 287.382
R33898 vdd.n3426 vdd.n3388 287.382
R33899 vdd.n3426 vdd.n3389 287.382
R33900 vdd.n3419 vdd.n3389 287.382
R33901 vdd.n802 vdd.n790 287.382
R33902 vdd.n809 vdd.n790 287.382
R33903 vdd.n813 vdd.n809 287.382
R33904 vdd.n813 vdd.n812 287.382
R33905 vdd.n812 vdd.n785 287.382
R33906 vdd.n823 vdd.n785 287.382
R33907 vdd.n3498 vdd.n3494 287.382
R33908 vdd.n3508 vdd.n3494 287.382
R33909 vdd.n3508 vdd.n3487 287.382
R33910 vdd.n3525 vdd.n3487 287.382
R33911 vdd.n3525 vdd.n3488 287.382
R33912 vdd.n3518 vdd.n3488 287.382
R33913 vdd.n3450 vdd.n3446 287.382
R33914 vdd.n3460 vdd.n3446 287.382
R33915 vdd.n3460 vdd.n3439 287.382
R33916 vdd.n3477 vdd.n3439 287.382
R33917 vdd.n3477 vdd.n3440 287.382
R33918 vdd.n3470 vdd.n3440 287.382
R33919 vdd.n3547 vdd.n3543 287.382
R33920 vdd.n3557 vdd.n3543 287.382
R33921 vdd.n3557 vdd.n3536 287.382
R33922 vdd.n3574 vdd.n3536 287.382
R33923 vdd.n3574 vdd.n3537 287.382
R33924 vdd.n3567 vdd.n3537 287.382
R33925 vdd.n3597 vdd.n3593 287.382
R33926 vdd.n3607 vdd.n3593 287.382
R33927 vdd.n3607 vdd.n3586 287.382
R33928 vdd.n3624 vdd.n3586 287.382
R33929 vdd.n3624 vdd.n3587 287.382
R33930 vdd.n3617 vdd.n3587 287.382
R33931 vdd.n3645 vdd.n3641 287.382
R33932 vdd.n3655 vdd.n3641 287.382
R33933 vdd.n3655 vdd.n3634 287.382
R33934 vdd.n3672 vdd.n3634 287.382
R33935 vdd.n3672 vdd.n3635 287.382
R33936 vdd.n3665 vdd.n3635 287.382
R33937 vdd.n603 vdd.n599 287.382
R33938 vdd.n613 vdd.n599 287.382
R33939 vdd.n613 vdd.n592 287.382
R33940 vdd.n630 vdd.n592 287.382
R33941 vdd.n630 vdd.n593 287.382
R33942 vdd.n623 vdd.n593 287.382
R33943 vdd.n3744 vdd.n3740 287.382
R33944 vdd.n3754 vdd.n3740 287.382
R33945 vdd.n3754 vdd.n3733 287.382
R33946 vdd.n3771 vdd.n3733 287.382
R33947 vdd.n3771 vdd.n3734 287.382
R33948 vdd.n3764 vdd.n3734 287.382
R33949 vdd.n3696 vdd.n3692 287.382
R33950 vdd.n3706 vdd.n3692 287.382
R33951 vdd.n3706 vdd.n3685 287.382
R33952 vdd.n3723 vdd.n3685 287.382
R33953 vdd.n3723 vdd.n3686 287.382
R33954 vdd.n3716 vdd.n3686 287.382
R33955 vdd.n6886 vdd.n6882 287.382
R33956 vdd.n6896 vdd.n6882 287.382
R33957 vdd.n6896 vdd.n6875 287.382
R33958 vdd.n6913 vdd.n6875 287.382
R33959 vdd.n6913 vdd.n6876 287.382
R33960 vdd.n6906 vdd.n6876 287.382
R33961 vdd.n6838 vdd.n6834 287.382
R33962 vdd.n6848 vdd.n6834 287.382
R33963 vdd.n6848 vdd.n6827 287.382
R33964 vdd.n6865 vdd.n6827 287.382
R33965 vdd.n6865 vdd.n6828 287.382
R33966 vdd.n6858 vdd.n6828 287.382
R33967 vdd.n10028 vdd.n10024 287.382
R33968 vdd.n10038 vdd.n10024 287.382
R33969 vdd.n10038 vdd.n10017 287.382
R33970 vdd.n10055 vdd.n10017 287.382
R33971 vdd.n10055 vdd.n10018 287.382
R33972 vdd.n10048 vdd.n10018 287.382
R33973 vdd.n9980 vdd.n9976 287.382
R33974 vdd.n9990 vdd.n9976 287.382
R33975 vdd.n9990 vdd.n9969 287.382
R33976 vdd.n10007 vdd.n9969 287.382
R33977 vdd.n10007 vdd.n9970 287.382
R33978 vdd.n10000 vdd.n9970 287.382
R33979 vdd.n10076 vdd.n10072 287.382
R33980 vdd.n10086 vdd.n10072 287.382
R33981 vdd.n10086 vdd.n10065 287.382
R33982 vdd.n10103 vdd.n10065 287.382
R33983 vdd.n10103 vdd.n10066 287.382
R33984 vdd.n10096 vdd.n10066 287.382
R33985 vdd.n10124 vdd.n10120 287.382
R33986 vdd.n10134 vdd.n10120 287.382
R33987 vdd.n10134 vdd.n10113 287.382
R33988 vdd.n10151 vdd.n10113 287.382
R33989 vdd.n10151 vdd.n10114 287.382
R33990 vdd.n10144 vdd.n10114 287.382
R33991 vdd.n10226 vdd.n10222 287.382
R33992 vdd.n10236 vdd.n10222 287.382
R33993 vdd.n10236 vdd.n10215 287.382
R33994 vdd.n10253 vdd.n10215 287.382
R33995 vdd.n10253 vdd.n10216 287.382
R33996 vdd.n10246 vdd.n10216 287.382
R33997 vdd.n10274 vdd.n10270 287.382
R33998 vdd.n10284 vdd.n10270 287.382
R33999 vdd.n10284 vdd.n10263 287.382
R34000 vdd.n10301 vdd.n10263 287.382
R34001 vdd.n10301 vdd.n10264 287.382
R34002 vdd.n10294 vdd.n10264 287.382
R34003 vdd.n10322 vdd.n10318 287.382
R34004 vdd.n10332 vdd.n10318 287.382
R34005 vdd.n10332 vdd.n10311 287.382
R34006 vdd.n10349 vdd.n10311 287.382
R34007 vdd.n10349 vdd.n10312 287.382
R34008 vdd.n10342 vdd.n10312 287.382
R34009 vdd.n10370 vdd.n10366 287.382
R34010 vdd.n10380 vdd.n10366 287.382
R34011 vdd.n10380 vdd.n10359 287.382
R34012 vdd.n10397 vdd.n10359 287.382
R34013 vdd.n10397 vdd.n10360 287.382
R34014 vdd.n10390 vdd.n10360 287.382
R34015 vdd.n10472 vdd.n10468 287.382
R34016 vdd.n10482 vdd.n10468 287.382
R34017 vdd.n10482 vdd.n10461 287.382
R34018 vdd.n10499 vdd.n10461 287.382
R34019 vdd.n10499 vdd.n10462 287.382
R34020 vdd.n10492 vdd.n10462 287.382
R34021 vdd.n64 vdd.n60 287.382
R34022 vdd.n74 vdd.n60 287.382
R34023 vdd.n74 vdd.n53 287.382
R34024 vdd.n91 vdd.n53 287.382
R34025 vdd.n91 vdd.n54 287.382
R34026 vdd.n84 vdd.n54 287.382
R34027 vdd.n16 vdd.n12 287.382
R34028 vdd.n26 vdd.n12 287.382
R34029 vdd.n26 vdd.n5 287.382
R34030 vdd.n43 vdd.n5 287.382
R34031 vdd.n43 vdd.n6 287.382
R34032 vdd.n36 vdd.n6 287.382
R34033 vdd.n10520 vdd.n10516 287.382
R34034 vdd.n10530 vdd.n10516 287.382
R34035 vdd.n10530 vdd.n10509 287.382
R34036 vdd.n10547 vdd.n10509 287.382
R34037 vdd.n10547 vdd.n10510 287.382
R34038 vdd.n10540 vdd.n10510 287.382
R34039 vdd.n10570 vdd.n10566 287.382
R34040 vdd.n10580 vdd.n10566 287.382
R34041 vdd.n10580 vdd.n10559 287.382
R34042 vdd.n10597 vdd.n10559 287.382
R34043 vdd.n10597 vdd.n10560 287.382
R34044 vdd.n10590 vdd.n10560 287.382
R34045 vdd.n10618 vdd.n10614 287.382
R34046 vdd.n10628 vdd.n10614 287.382
R34047 vdd.n10628 vdd.n10607 287.382
R34048 vdd.n10645 vdd.n10607 287.382
R34049 vdd.n10645 vdd.n10608 287.382
R34050 vdd.n10638 vdd.n10608 287.382
R34051 vdd.n10425 vdd.n10413 287.382
R34052 vdd.n10432 vdd.n10413 287.382
R34053 vdd.n10436 vdd.n10432 287.382
R34054 vdd.n10436 vdd.n10435 287.382
R34055 vdd.n10435 vdd.n10408 287.382
R34056 vdd.n10446 vdd.n10408 287.382
R34057 vdd.n10766 vdd.n10762 287.382
R34058 vdd.n10776 vdd.n10762 287.382
R34059 vdd.n10776 vdd.n10755 287.382
R34060 vdd.n10793 vdd.n10755 287.382
R34061 vdd.n10793 vdd.n10756 287.382
R34062 vdd.n10786 vdd.n10756 287.382
R34063 vdd.n10717 vdd.n10713 287.382
R34064 vdd.n10727 vdd.n10713 287.382
R34065 vdd.n10727 vdd.n10706 287.382
R34066 vdd.n10744 vdd.n10706 287.382
R34067 vdd.n10744 vdd.n10707 287.382
R34068 vdd.n10737 vdd.n10707 287.382
R34069 vdd.n10669 vdd.n10665 287.382
R34070 vdd.n10679 vdd.n10665 287.382
R34071 vdd.n10679 vdd.n10658 287.382
R34072 vdd.n10696 vdd.n10658 287.382
R34073 vdd.n10696 vdd.n10659 287.382
R34074 vdd.n10689 vdd.n10659 287.382
R34075 vdd.n10815 vdd.n10811 287.382
R34076 vdd.n10825 vdd.n10811 287.382
R34077 vdd.n10825 vdd.n10804 287.382
R34078 vdd.n10842 vdd.n10804 287.382
R34079 vdd.n10842 vdd.n10805 287.382
R34080 vdd.n10835 vdd.n10805 287.382
R34081 vdd.n10865 vdd.n10861 287.382
R34082 vdd.n10875 vdd.n10861 287.382
R34083 vdd.n10875 vdd.n10854 287.382
R34084 vdd.n10892 vdd.n10854 287.382
R34085 vdd.n10892 vdd.n10855 287.382
R34086 vdd.n10885 vdd.n10855 287.382
R34087 vdd.n10913 vdd.n10909 287.382
R34088 vdd.n10923 vdd.n10909 287.382
R34089 vdd.n10923 vdd.n10902 287.382
R34090 vdd.n10940 vdd.n10902 287.382
R34091 vdd.n10940 vdd.n10903 287.382
R34092 vdd.n10933 vdd.n10903 287.382
R34093 vdd.n11011 vdd.n11007 287.382
R34094 vdd.n11021 vdd.n11007 287.382
R34095 vdd.n11021 vdd.n11000 287.382
R34096 vdd.n11038 vdd.n11000 287.382
R34097 vdd.n11038 vdd.n11001 287.382
R34098 vdd.n11031 vdd.n11001 287.382
R34099 vdd.n10963 vdd.n10959 287.382
R34100 vdd.n10973 vdd.n10959 287.382
R34101 vdd.n10973 vdd.n10952 287.382
R34102 vdd.n10990 vdd.n10952 287.382
R34103 vdd.n10990 vdd.n10953 287.382
R34104 vdd.n10983 vdd.n10953 287.382
R34105 vdd.n11060 vdd.n11056 287.382
R34106 vdd.n11070 vdd.n11056 287.382
R34107 vdd.n11070 vdd.n11049 287.382
R34108 vdd.n11087 vdd.n11049 287.382
R34109 vdd.n11087 vdd.n11050 287.382
R34110 vdd.n11080 vdd.n11050 287.382
R34111 vdd.n11110 vdd.n11106 287.382
R34112 vdd.n11120 vdd.n11106 287.382
R34113 vdd.n11120 vdd.n11099 287.382
R34114 vdd.n11137 vdd.n11099 287.382
R34115 vdd.n11137 vdd.n11100 287.382
R34116 vdd.n11130 vdd.n11100 287.382
R34117 vdd.n11158 vdd.n11154 287.382
R34118 vdd.n11168 vdd.n11154 287.382
R34119 vdd.n11168 vdd.n11147 287.382
R34120 vdd.n11185 vdd.n11147 287.382
R34121 vdd.n11185 vdd.n11148 287.382
R34122 vdd.n11178 vdd.n11148 287.382
R34123 vdd.n10179 vdd.n10167 287.382
R34124 vdd.n10186 vdd.n10167 287.382
R34125 vdd.n10190 vdd.n10186 287.382
R34126 vdd.n10190 vdd.n10189 287.382
R34127 vdd.n10189 vdd.n10162 287.382
R34128 vdd.n10200 vdd.n10162 287.382
R34129 vdd.n11257 vdd.n11253 287.382
R34130 vdd.n11267 vdd.n11253 287.382
R34131 vdd.n11267 vdd.n11246 287.382
R34132 vdd.n11284 vdd.n11246 287.382
R34133 vdd.n11284 vdd.n11247 287.382
R34134 vdd.n11277 vdd.n11247 287.382
R34135 vdd.n11209 vdd.n11205 287.382
R34136 vdd.n11219 vdd.n11205 287.382
R34137 vdd.n11219 vdd.n11198 287.382
R34138 vdd.n11236 vdd.n11198 287.382
R34139 vdd.n11236 vdd.n11199 287.382
R34140 vdd.n11229 vdd.n11199 287.382
R34141 vdd.n11306 vdd.n11302 287.382
R34142 vdd.n11316 vdd.n11302 287.382
R34143 vdd.n11316 vdd.n11295 287.382
R34144 vdd.n11333 vdd.n11295 287.382
R34145 vdd.n11333 vdd.n11296 287.382
R34146 vdd.n11326 vdd.n11296 287.382
R34147 vdd.n11356 vdd.n11352 287.382
R34148 vdd.n11366 vdd.n11352 287.382
R34149 vdd.n11366 vdd.n11345 287.382
R34150 vdd.n11383 vdd.n11345 287.382
R34151 vdd.n11383 vdd.n11346 287.382
R34152 vdd.n11376 vdd.n11346 287.382
R34153 vdd.n11404 vdd.n11400 287.382
R34154 vdd.n11414 vdd.n11400 287.382
R34155 vdd.n11414 vdd.n11393 287.382
R34156 vdd.n11431 vdd.n11393 287.382
R34157 vdd.n11431 vdd.n11394 287.382
R34158 vdd.n11424 vdd.n11394 287.382
R34159 vdd.n11461 vdd.n11451 287.382
R34160 vdd.n11465 vdd.n11451 287.382
R34161 vdd.n11465 vdd.n11444 287.382
R34162 vdd.n11482 vdd.n11444 287.382
R34163 vdd.n11482 vdd.n11445 287.382
R34164 vdd.n11476 vdd.n11445 287.382
R34165 vdd.n11508 vdd.n11498 287.382
R34166 vdd.n11512 vdd.n11498 287.382
R34167 vdd.n11512 vdd.n11491 287.382
R34168 vdd.n11529 vdd.n11491 287.382
R34169 vdd.n11529 vdd.n11492 287.382
R34170 vdd.n11523 vdd.n11492 287.382
R34171 vdd.n11558 vdd.n11548 287.382
R34172 vdd.n11562 vdd.n11548 287.382
R34173 vdd.n11562 vdd.n11541 287.382
R34174 vdd.n11579 vdd.n11541 287.382
R34175 vdd.n11579 vdd.n11542 287.382
R34176 vdd.n11573 vdd.n11542 287.382
R34177 vdd.n11608 vdd.n11598 287.382
R34178 vdd.n11612 vdd.n11598 287.382
R34179 vdd.n11612 vdd.n11591 287.382
R34180 vdd.n11629 vdd.n11591 287.382
R34181 vdd.n11629 vdd.n11592 287.382
R34182 vdd.n11623 vdd.n11592 287.382
R34183 vdd.n11656 vdd.n11646 287.382
R34184 vdd.n11660 vdd.n11646 287.382
R34185 vdd.n11660 vdd.n11639 287.382
R34186 vdd.n11677 vdd.n11639 287.382
R34187 vdd.n11677 vdd.n11640 287.382
R34188 vdd.n11671 vdd.n11640 287.382
R34189 vdd.n484 vdd.n444 287.382
R34190 vdd.n477 vdd.n444 287.382
R34191 vdd.n477 vdd.n450 287.382
R34192 vdd.n469 vdd.n450 287.382
R34193 vdd.n469 vdd.n453 287.382
R34194 vdd.n463 vdd.n453 287.382
R34195 vdd.n11707 vdd.n11697 287.382
R34196 vdd.n11711 vdd.n11697 287.382
R34197 vdd.n11711 vdd.n11690 287.382
R34198 vdd.n11728 vdd.n11690 287.382
R34199 vdd.n11728 vdd.n11691 287.382
R34200 vdd.n11722 vdd.n11691 287.382
R34201 vdd.n11754 vdd.n11744 287.382
R34202 vdd.n11758 vdd.n11744 287.382
R34203 vdd.n11758 vdd.n11737 287.382
R34204 vdd.n11775 vdd.n11737 287.382
R34205 vdd.n11775 vdd.n11738 287.382
R34206 vdd.n11769 vdd.n11738 287.382
R34207 vdd.n11802 vdd.n11792 287.382
R34208 vdd.n11806 vdd.n11792 287.382
R34209 vdd.n11806 vdd.n11785 287.382
R34210 vdd.n11823 vdd.n11785 287.382
R34211 vdd.n11823 vdd.n11786 287.382
R34212 vdd.n11817 vdd.n11786 287.382
R34213 vdd.n11853 vdd.n11843 287.382
R34214 vdd.n11857 vdd.n11843 287.382
R34215 vdd.n11857 vdd.n11836 287.382
R34216 vdd.n11874 vdd.n11836 287.382
R34217 vdd.n11874 vdd.n11837 287.382
R34218 vdd.n11868 vdd.n11837 287.382
R34219 vdd.n11903 vdd.n11893 287.382
R34220 vdd.n11907 vdd.n11893 287.382
R34221 vdd.n11907 vdd.n11886 287.382
R34222 vdd.n11924 vdd.n11886 287.382
R34223 vdd.n11924 vdd.n11887 287.382
R34224 vdd.n11918 vdd.n11887 287.382
R34225 vdd.n11951 vdd.n11941 287.382
R34226 vdd.n11955 vdd.n11941 287.382
R34227 vdd.n11955 vdd.n11934 287.382
R34228 vdd.n11972 vdd.n11934 287.382
R34229 vdd.n11972 vdd.n11935 287.382
R34230 vdd.n11966 vdd.n11935 287.382
R34231 vdd.n12001 vdd.n11991 287.382
R34232 vdd.n12005 vdd.n11991 287.382
R34233 vdd.n12005 vdd.n11984 287.382
R34234 vdd.n12022 vdd.n11984 287.382
R34235 vdd.n12022 vdd.n11985 287.382
R34236 vdd.n12016 vdd.n11985 287.382
R34237 vdd.n12048 vdd.n12038 287.382
R34238 vdd.n12052 vdd.n12038 287.382
R34239 vdd.n12052 vdd.n12031 287.382
R34240 vdd.n12069 vdd.n12031 287.382
R34241 vdd.n12069 vdd.n12032 287.382
R34242 vdd.n12063 vdd.n12032 287.382
R34243 vdd.n12098 vdd.n12088 287.382
R34244 vdd.n12102 vdd.n12088 287.382
R34245 vdd.n12102 vdd.n12081 287.382
R34246 vdd.n12119 vdd.n12081 287.382
R34247 vdd.n12119 vdd.n12082 287.382
R34248 vdd.n12113 vdd.n12082 287.382
R34249 vdd.n12148 vdd.n12138 287.382
R34250 vdd.n12152 vdd.n12138 287.382
R34251 vdd.n12152 vdd.n12131 287.382
R34252 vdd.n12169 vdd.n12131 287.382
R34253 vdd.n12169 vdd.n12132 287.382
R34254 vdd.n12163 vdd.n12132 287.382
R34255 vdd.n12196 vdd.n12186 287.382
R34256 vdd.n12200 vdd.n12186 287.382
R34257 vdd.n12200 vdd.n12179 287.382
R34258 vdd.n12217 vdd.n12179 287.382
R34259 vdd.n12217 vdd.n12180 287.382
R34260 vdd.n12211 vdd.n12180 287.382
R34261 vdd.n239 vdd.n199 287.382
R34262 vdd.n232 vdd.n199 287.382
R34263 vdd.n232 vdd.n205 287.382
R34264 vdd.n224 vdd.n205 287.382
R34265 vdd.n224 vdd.n208 287.382
R34266 vdd.n218 vdd.n208 287.382
R34267 vdd.n12247 vdd.n12237 287.382
R34268 vdd.n12251 vdd.n12237 287.382
R34269 vdd.n12251 vdd.n12230 287.382
R34270 vdd.n12268 vdd.n12230 287.382
R34271 vdd.n12268 vdd.n12231 287.382
R34272 vdd.n12262 vdd.n12231 287.382
R34273 vdd.n12294 vdd.n12284 287.382
R34274 vdd.n12298 vdd.n12284 287.382
R34275 vdd.n12298 vdd.n12277 287.382
R34276 vdd.n12315 vdd.n12277 287.382
R34277 vdd.n12315 vdd.n12278 287.382
R34278 vdd.n12309 vdd.n12278 287.382
R34279 vdd.n12344 vdd.n12334 287.382
R34280 vdd.n12348 vdd.n12334 287.382
R34281 vdd.n12348 vdd.n12327 287.382
R34282 vdd.n12365 vdd.n12327 287.382
R34283 vdd.n12365 vdd.n12328 287.382
R34284 vdd.n12359 vdd.n12328 287.382
R34285 vdd.n12394 vdd.n12384 287.382
R34286 vdd.n12398 vdd.n12384 287.382
R34287 vdd.n12398 vdd.n12377 287.382
R34288 vdd.n12415 vdd.n12377 287.382
R34289 vdd.n12415 vdd.n12378 287.382
R34290 vdd.n12409 vdd.n12378 287.382
R34291 vdd.n12442 vdd.n12432 287.382
R34292 vdd.n12446 vdd.n12432 287.382
R34293 vdd.n12446 vdd.n12425 287.382
R34294 vdd.n12463 vdd.n12425 287.382
R34295 vdd.n12463 vdd.n12426 287.382
R34296 vdd.n12457 vdd.n12426 287.382
R34297 vdd.n118 vdd.n111 242.685
R34298 vdd.n166 vdd.n159 242.685
R34299 vdd.n267 vdd.n260 242.685
R34300 vdd.n315 vdd.n308 242.685
R34301 vdd.n363 vdd.n356 242.685
R34302 vdd.n411 vdd.n404 242.685
R34303 vdd.n512 vdd.n505 242.685
R34304 vdd.n560 vdd.n553 242.685
R34305 vdd.n7432 vdd.n7425 242.685
R34306 vdd.n7480 vdd.n7473 242.685
R34307 vdd.n7581 vdd.n7574 242.685
R34308 vdd.n7629 vdd.n7622 242.685
R34309 vdd.n7677 vdd.n7670 242.685
R34310 vdd.n7725 vdd.n7718 242.685
R34311 vdd.n7826 vdd.n7819 242.685
R34312 vdd.n6939 vdd.n6932 242.685
R34313 vdd.n7874 vdd.n7867 242.685
R34314 vdd.n7921 vdd.n7914 242.685
R34315 vdd.n7971 vdd.n7964 242.685
R34316 vdd.n8021 vdd.n8014 242.685
R34317 vdd.n8069 vdd.n8062 242.685
R34318 vdd.n7797 vdd.n7756 242.685
R34319 vdd.n8120 vdd.n8113 242.685
R34320 vdd.n8167 vdd.n8160 242.685
R34321 vdd.n8215 vdd.n8208 242.685
R34322 vdd.n8266 vdd.n8259 242.685
R34323 vdd.n8316 vdd.n8309 242.685
R34324 vdd.n8364 vdd.n8357 242.685
R34325 vdd.n8414 vdd.n8407 242.685
R34326 vdd.n8461 vdd.n8454 242.685
R34327 vdd.n8511 vdd.n8504 242.685
R34328 vdd.n8561 vdd.n8554 242.685
R34329 vdd.n8609 vdd.n8602 242.685
R34330 vdd.n7552 vdd.n7511 242.685
R34331 vdd.n8660 vdd.n8653 242.685
R34332 vdd.n8707 vdd.n8700 242.685
R34333 vdd.n8757 vdd.n8750 242.685
R34334 vdd.n8807 vdd.n8800 242.685
R34335 vdd.n8855 vdd.n8848 242.685
R34336 vdd.n4290 vdd.n4283 242.685
R34337 vdd.n4338 vdd.n4331 242.685
R34338 vdd.n4439 vdd.n4432 242.685
R34339 vdd.n4487 vdd.n4480 242.685
R34340 vdd.n4535 vdd.n4528 242.685
R34341 vdd.n4583 vdd.n4576 242.685
R34342 vdd.n4684 vdd.n4677 242.685
R34343 vdd.n3797 vdd.n3790 242.685
R34344 vdd.n4732 vdd.n4725 242.685
R34345 vdd.n4779 vdd.n4772 242.685
R34346 vdd.n4829 vdd.n4822 242.685
R34347 vdd.n4879 vdd.n4872 242.685
R34348 vdd.n4927 vdd.n4920 242.685
R34349 vdd.n4655 vdd.n4614 242.685
R34350 vdd.n4978 vdd.n4971 242.685
R34351 vdd.n5025 vdd.n5018 242.685
R34352 vdd.n5073 vdd.n5066 242.685
R34353 vdd.n5124 vdd.n5117 242.685
R34354 vdd.n5174 vdd.n5167 242.685
R34355 vdd.n5222 vdd.n5215 242.685
R34356 vdd.n5272 vdd.n5265 242.685
R34357 vdd.n5319 vdd.n5312 242.685
R34358 vdd.n5369 vdd.n5362 242.685
R34359 vdd.n5419 vdd.n5412 242.685
R34360 vdd.n5467 vdd.n5460 242.685
R34361 vdd.n4410 vdd.n4369 242.685
R34362 vdd.n5518 vdd.n5511 242.685
R34363 vdd.n5565 vdd.n5558 242.685
R34364 vdd.n5615 vdd.n5608 242.685
R34365 vdd.n5665 vdd.n5658 242.685
R34366 vdd.n5713 vdd.n5706 242.685
R34367 vdd.n1148 vdd.n1141 242.685
R34368 vdd.n1196 vdd.n1189 242.685
R34369 vdd.n1297 vdd.n1290 242.685
R34370 vdd.n1345 vdd.n1338 242.685
R34371 vdd.n1393 vdd.n1386 242.685
R34372 vdd.n1441 vdd.n1434 242.685
R34373 vdd.n1542 vdd.n1535 242.685
R34374 vdd.n655 vdd.n648 242.685
R34375 vdd.n1590 vdd.n1583 242.685
R34376 vdd.n1637 vdd.n1630 242.685
R34377 vdd.n1687 vdd.n1680 242.685
R34378 vdd.n1737 vdd.n1730 242.685
R34379 vdd.n1785 vdd.n1778 242.685
R34380 vdd.n1513 vdd.n1472 242.685
R34381 vdd.n1836 vdd.n1829 242.685
R34382 vdd.n1883 vdd.n1876 242.685
R34383 vdd.n1931 vdd.n1924 242.685
R34384 vdd.n1982 vdd.n1975 242.685
R34385 vdd.n2032 vdd.n2025 242.685
R34386 vdd.n2080 vdd.n2073 242.685
R34387 vdd.n2130 vdd.n2123 242.685
R34388 vdd.n2177 vdd.n2170 242.685
R34389 vdd.n2227 vdd.n2220 242.685
R34390 vdd.n2277 vdd.n2270 242.685
R34391 vdd.n2325 vdd.n2318 242.685
R34392 vdd.n1268 vdd.n1227 242.685
R34393 vdd.n2376 vdd.n2369 242.685
R34394 vdd.n2423 vdd.n2416 242.685
R34395 vdd.n2473 vdd.n2466 242.685
R34396 vdd.n2523 vdd.n2516 242.685
R34397 vdd.n2571 vdd.n2564 242.685
R34398 vdd.n11460 vdd.n11453 242.685
R34399 vdd.n11507 vdd.n11500 242.685
R34400 vdd.n11557 vdd.n11550 242.685
R34401 vdd.n11607 vdd.n11600 242.685
R34402 vdd.n11655 vdd.n11648 242.685
R34403 vdd.n483 vdd.n442 242.685
R34404 vdd.n11706 vdd.n11699 242.685
R34405 vdd.n11753 vdd.n11746 242.685
R34406 vdd.n11801 vdd.n11794 242.685
R34407 vdd.n11852 vdd.n11845 242.685
R34408 vdd.n11902 vdd.n11895 242.685
R34409 vdd.n11950 vdd.n11943 242.685
R34410 vdd.n12000 vdd.n11993 242.685
R34411 vdd.n12047 vdd.n12040 242.685
R34412 vdd.n12097 vdd.n12090 242.685
R34413 vdd.n12147 vdd.n12140 242.685
R34414 vdd.n12195 vdd.n12188 242.685
R34415 vdd.n238 vdd.n197 242.685
R34416 vdd.n12246 vdd.n12239 242.685
R34417 vdd.n12293 vdd.n12286 242.685
R34418 vdd.n12343 vdd.n12336 242.685
R34419 vdd.n12393 vdd.n12386 242.685
R34420 vdd.n12441 vdd.n12434 242.685
R34421 vdd.n133 vdd.n130 242.684
R34422 vdd.n181 vdd.n178 242.684
R34423 vdd.n282 vdd.n279 242.684
R34424 vdd.n330 vdd.n327 242.684
R34425 vdd.n378 vdd.n375 242.684
R34426 vdd.n426 vdd.n423 242.684
R34427 vdd.n527 vdd.n524 242.684
R34428 vdd.n575 vdd.n572 242.684
R34429 vdd.n6985 vdd.n6981 242.684
R34430 vdd.n7004 vdd.n7000 242.684
R34431 vdd.n7033 vdd.n7029 242.684
R34432 vdd.n7052 vdd.n7048 242.684
R34433 vdd.n7135 vdd.n7131 242.684
R34434 vdd.n7154 vdd.n7150 242.684
R34435 vdd.n7183 vdd.n7179 242.684
R34436 vdd.n7202 vdd.n7198 242.684
R34437 vdd.n7231 vdd.n7227 242.684
R34438 vdd.n7250 vdd.n7246 242.684
R34439 vdd.n7279 vdd.n7275 242.684
R34440 vdd.n7298 vdd.n7294 242.684
R34441 vdd.n7381 vdd.n7377 242.684
R34442 vdd.n7400 vdd.n7396 242.684
R34443 vdd.n8901 vdd.n8897 242.684
R34444 vdd.n8920 vdd.n8916 242.684
R34445 vdd.n7447 vdd.n7444 242.684
R34446 vdd.n7495 vdd.n7492 242.684
R34447 vdd.n7596 vdd.n7593 242.684
R34448 vdd.n7644 vdd.n7641 242.684
R34449 vdd.n7692 vdd.n7689 242.684
R34450 vdd.n7740 vdd.n7737 242.684
R34451 vdd.n7841 vdd.n7838 242.684
R34452 vdd.n6954 vdd.n6951 242.684
R34453 vdd.n7889 vdd.n7886 242.684
R34454 vdd.n7936 vdd.n7933 242.684
R34455 vdd.n7986 vdd.n7983 242.684
R34456 vdd.n8036 vdd.n8033 242.684
R34457 vdd.n8084 vdd.n8081 242.684
R34458 vdd.n7776 vdd.n7772 242.684
R34459 vdd.n8135 vdd.n8132 242.684
R34460 vdd.n8182 vdd.n8179 242.684
R34461 vdd.n8230 vdd.n8227 242.684
R34462 vdd.n8281 vdd.n8278 242.684
R34463 vdd.n8331 vdd.n8328 242.684
R34464 vdd.n8379 vdd.n8376 242.684
R34465 vdd.n8429 vdd.n8426 242.684
R34466 vdd.n8476 vdd.n8473 242.684
R34467 vdd.n8526 vdd.n8523 242.684
R34468 vdd.n8576 vdd.n8573 242.684
R34469 vdd.n8624 vdd.n8621 242.684
R34470 vdd.n7531 vdd.n7527 242.684
R34471 vdd.n8675 vdd.n8672 242.684
R34472 vdd.n8722 vdd.n8719 242.684
R34473 vdd.n8772 vdd.n8769 242.684
R34474 vdd.n8822 vdd.n8819 242.684
R34475 vdd.n8870 vdd.n8867 242.684
R34476 vdd.n8998 vdd.n8994 242.684
R34477 vdd.n9017 vdd.n9013 242.684
R34478 vdd.n8950 vdd.n8946 242.684
R34479 vdd.n8969 vdd.n8965 242.684
R34480 vdd.n9047 vdd.n9043 242.684
R34481 vdd.n9066 vdd.n9062 242.684
R34482 vdd.n9097 vdd.n9093 242.684
R34483 vdd.n9116 vdd.n9112 242.684
R34484 vdd.n9145 vdd.n9141 242.684
R34485 vdd.n9164 vdd.n9160 242.684
R34486 vdd.n7333 vdd.n7325 242.684
R34487 vdd.n7354 vdd.n7312 242.684
R34488 vdd.n9293 vdd.n9289 242.684
R34489 vdd.n9312 vdd.n9308 242.684
R34490 vdd.n9244 vdd.n9240 242.684
R34491 vdd.n9263 vdd.n9259 242.684
R34492 vdd.n9196 vdd.n9192 242.684
R34493 vdd.n9215 vdd.n9211 242.684
R34494 vdd.n9342 vdd.n9338 242.684
R34495 vdd.n9361 vdd.n9357 242.684
R34496 vdd.n9392 vdd.n9388 242.684
R34497 vdd.n9411 vdd.n9407 242.684
R34498 vdd.n9440 vdd.n9436 242.684
R34499 vdd.n9459 vdd.n9455 242.684
R34500 vdd.n9538 vdd.n9534 242.684
R34501 vdd.n9557 vdd.n9553 242.684
R34502 vdd.n9490 vdd.n9486 242.684
R34503 vdd.n9509 vdd.n9505 242.684
R34504 vdd.n9587 vdd.n9583 242.684
R34505 vdd.n9606 vdd.n9602 242.684
R34506 vdd.n9637 vdd.n9633 242.684
R34507 vdd.n9656 vdd.n9652 242.684
R34508 vdd.n9685 vdd.n9681 242.684
R34509 vdd.n9704 vdd.n9700 242.684
R34510 vdd.n7087 vdd.n7079 242.684
R34511 vdd.n7108 vdd.n7066 242.684
R34512 vdd.n9784 vdd.n9780 242.684
R34513 vdd.n9803 vdd.n9799 242.684
R34514 vdd.n9736 vdd.n9732 242.684
R34515 vdd.n9755 vdd.n9751 242.684
R34516 vdd.n9833 vdd.n9829 242.684
R34517 vdd.n9852 vdd.n9848 242.684
R34518 vdd.n9883 vdd.n9879 242.684
R34519 vdd.n9902 vdd.n9898 242.684
R34520 vdd.n9931 vdd.n9927 242.684
R34521 vdd.n9950 vdd.n9946 242.684
R34522 vdd.n3843 vdd.n3839 242.684
R34523 vdd.n3862 vdd.n3858 242.684
R34524 vdd.n3891 vdd.n3887 242.684
R34525 vdd.n3910 vdd.n3906 242.684
R34526 vdd.n3993 vdd.n3989 242.684
R34527 vdd.n4012 vdd.n4008 242.684
R34528 vdd.n4041 vdd.n4037 242.684
R34529 vdd.n4060 vdd.n4056 242.684
R34530 vdd.n4089 vdd.n4085 242.684
R34531 vdd.n4108 vdd.n4104 242.684
R34532 vdd.n4137 vdd.n4133 242.684
R34533 vdd.n4156 vdd.n4152 242.684
R34534 vdd.n4239 vdd.n4235 242.684
R34535 vdd.n4258 vdd.n4254 242.684
R34536 vdd.n5759 vdd.n5755 242.684
R34537 vdd.n5778 vdd.n5774 242.684
R34538 vdd.n4305 vdd.n4302 242.684
R34539 vdd.n4353 vdd.n4350 242.684
R34540 vdd.n4454 vdd.n4451 242.684
R34541 vdd.n4502 vdd.n4499 242.684
R34542 vdd.n4550 vdd.n4547 242.684
R34543 vdd.n4598 vdd.n4595 242.684
R34544 vdd.n4699 vdd.n4696 242.684
R34545 vdd.n3812 vdd.n3809 242.684
R34546 vdd.n4747 vdd.n4744 242.684
R34547 vdd.n4794 vdd.n4791 242.684
R34548 vdd.n4844 vdd.n4841 242.684
R34549 vdd.n4894 vdd.n4891 242.684
R34550 vdd.n4942 vdd.n4939 242.684
R34551 vdd.n4634 vdd.n4630 242.684
R34552 vdd.n4993 vdd.n4990 242.684
R34553 vdd.n5040 vdd.n5037 242.684
R34554 vdd.n5088 vdd.n5085 242.684
R34555 vdd.n5139 vdd.n5136 242.684
R34556 vdd.n5189 vdd.n5186 242.684
R34557 vdd.n5237 vdd.n5234 242.684
R34558 vdd.n5287 vdd.n5284 242.684
R34559 vdd.n5334 vdd.n5331 242.684
R34560 vdd.n5384 vdd.n5381 242.684
R34561 vdd.n5434 vdd.n5431 242.684
R34562 vdd.n5482 vdd.n5479 242.684
R34563 vdd.n4389 vdd.n4385 242.684
R34564 vdd.n5533 vdd.n5530 242.684
R34565 vdd.n5580 vdd.n5577 242.684
R34566 vdd.n5630 vdd.n5627 242.684
R34567 vdd.n5680 vdd.n5677 242.684
R34568 vdd.n5728 vdd.n5725 242.684
R34569 vdd.n5856 vdd.n5852 242.684
R34570 vdd.n5875 vdd.n5871 242.684
R34571 vdd.n5808 vdd.n5804 242.684
R34572 vdd.n5827 vdd.n5823 242.684
R34573 vdd.n5905 vdd.n5901 242.684
R34574 vdd.n5924 vdd.n5920 242.684
R34575 vdd.n5955 vdd.n5951 242.684
R34576 vdd.n5974 vdd.n5970 242.684
R34577 vdd.n6003 vdd.n5999 242.684
R34578 vdd.n6022 vdd.n6018 242.684
R34579 vdd.n4191 vdd.n4183 242.684
R34580 vdd.n4212 vdd.n4170 242.684
R34581 vdd.n6151 vdd.n6147 242.684
R34582 vdd.n6170 vdd.n6166 242.684
R34583 vdd.n6102 vdd.n6098 242.684
R34584 vdd.n6121 vdd.n6117 242.684
R34585 vdd.n6054 vdd.n6050 242.684
R34586 vdd.n6073 vdd.n6069 242.684
R34587 vdd.n6200 vdd.n6196 242.684
R34588 vdd.n6219 vdd.n6215 242.684
R34589 vdd.n6250 vdd.n6246 242.684
R34590 vdd.n6269 vdd.n6265 242.684
R34591 vdd.n6298 vdd.n6294 242.684
R34592 vdd.n6317 vdd.n6313 242.684
R34593 vdd.n6396 vdd.n6392 242.684
R34594 vdd.n6415 vdd.n6411 242.684
R34595 vdd.n6348 vdd.n6344 242.684
R34596 vdd.n6367 vdd.n6363 242.684
R34597 vdd.n6445 vdd.n6441 242.684
R34598 vdd.n6464 vdd.n6460 242.684
R34599 vdd.n6495 vdd.n6491 242.684
R34600 vdd.n6514 vdd.n6510 242.684
R34601 vdd.n6543 vdd.n6539 242.684
R34602 vdd.n6562 vdd.n6558 242.684
R34603 vdd.n3945 vdd.n3937 242.684
R34604 vdd.n3966 vdd.n3924 242.684
R34605 vdd.n6642 vdd.n6638 242.684
R34606 vdd.n6661 vdd.n6657 242.684
R34607 vdd.n6594 vdd.n6590 242.684
R34608 vdd.n6613 vdd.n6609 242.684
R34609 vdd.n6691 vdd.n6687 242.684
R34610 vdd.n6710 vdd.n6706 242.684
R34611 vdd.n6741 vdd.n6737 242.684
R34612 vdd.n6760 vdd.n6756 242.684
R34613 vdd.n6789 vdd.n6785 242.684
R34614 vdd.n6808 vdd.n6804 242.684
R34615 vdd.n701 vdd.n697 242.684
R34616 vdd.n720 vdd.n716 242.684
R34617 vdd.n749 vdd.n745 242.684
R34618 vdd.n768 vdd.n764 242.684
R34619 vdd.n851 vdd.n847 242.684
R34620 vdd.n870 vdd.n866 242.684
R34621 vdd.n899 vdd.n895 242.684
R34622 vdd.n918 vdd.n914 242.684
R34623 vdd.n947 vdd.n943 242.684
R34624 vdd.n966 vdd.n962 242.684
R34625 vdd.n995 vdd.n991 242.684
R34626 vdd.n1014 vdd.n1010 242.684
R34627 vdd.n1097 vdd.n1093 242.684
R34628 vdd.n1116 vdd.n1112 242.684
R34629 vdd.n2617 vdd.n2613 242.684
R34630 vdd.n2636 vdd.n2632 242.684
R34631 vdd.n1163 vdd.n1160 242.684
R34632 vdd.n1211 vdd.n1208 242.684
R34633 vdd.n1312 vdd.n1309 242.684
R34634 vdd.n1360 vdd.n1357 242.684
R34635 vdd.n1408 vdd.n1405 242.684
R34636 vdd.n1456 vdd.n1453 242.684
R34637 vdd.n1557 vdd.n1554 242.684
R34638 vdd.n670 vdd.n667 242.684
R34639 vdd.n1605 vdd.n1602 242.684
R34640 vdd.n1652 vdd.n1649 242.684
R34641 vdd.n1702 vdd.n1699 242.684
R34642 vdd.n1752 vdd.n1749 242.684
R34643 vdd.n1800 vdd.n1797 242.684
R34644 vdd.n1492 vdd.n1488 242.684
R34645 vdd.n1851 vdd.n1848 242.684
R34646 vdd.n1898 vdd.n1895 242.684
R34647 vdd.n1946 vdd.n1943 242.684
R34648 vdd.n1997 vdd.n1994 242.684
R34649 vdd.n2047 vdd.n2044 242.684
R34650 vdd.n2095 vdd.n2092 242.684
R34651 vdd.n2145 vdd.n2142 242.684
R34652 vdd.n2192 vdd.n2189 242.684
R34653 vdd.n2242 vdd.n2239 242.684
R34654 vdd.n2292 vdd.n2289 242.684
R34655 vdd.n2340 vdd.n2337 242.684
R34656 vdd.n1247 vdd.n1243 242.684
R34657 vdd.n2391 vdd.n2388 242.684
R34658 vdd.n2438 vdd.n2435 242.684
R34659 vdd.n2488 vdd.n2485 242.684
R34660 vdd.n2538 vdd.n2535 242.684
R34661 vdd.n2586 vdd.n2583 242.684
R34662 vdd.n2714 vdd.n2710 242.684
R34663 vdd.n2733 vdd.n2729 242.684
R34664 vdd.n2666 vdd.n2662 242.684
R34665 vdd.n2685 vdd.n2681 242.684
R34666 vdd.n2763 vdd.n2759 242.684
R34667 vdd.n2782 vdd.n2778 242.684
R34668 vdd.n2813 vdd.n2809 242.684
R34669 vdd.n2832 vdd.n2828 242.684
R34670 vdd.n2861 vdd.n2857 242.684
R34671 vdd.n2880 vdd.n2876 242.684
R34672 vdd.n1049 vdd.n1041 242.684
R34673 vdd.n1070 vdd.n1028 242.684
R34674 vdd.n3009 vdd.n3005 242.684
R34675 vdd.n3028 vdd.n3024 242.684
R34676 vdd.n2960 vdd.n2956 242.684
R34677 vdd.n2979 vdd.n2975 242.684
R34678 vdd.n2912 vdd.n2908 242.684
R34679 vdd.n2931 vdd.n2927 242.684
R34680 vdd.n3058 vdd.n3054 242.684
R34681 vdd.n3077 vdd.n3073 242.684
R34682 vdd.n3108 vdd.n3104 242.684
R34683 vdd.n3127 vdd.n3123 242.684
R34684 vdd.n3156 vdd.n3152 242.684
R34685 vdd.n3175 vdd.n3171 242.684
R34686 vdd.n3254 vdd.n3250 242.684
R34687 vdd.n3273 vdd.n3269 242.684
R34688 vdd.n3206 vdd.n3202 242.684
R34689 vdd.n3225 vdd.n3221 242.684
R34690 vdd.n3303 vdd.n3299 242.684
R34691 vdd.n3322 vdd.n3318 242.684
R34692 vdd.n3353 vdd.n3349 242.684
R34693 vdd.n3372 vdd.n3368 242.684
R34694 vdd.n3401 vdd.n3397 242.684
R34695 vdd.n3420 vdd.n3416 242.684
R34696 vdd.n803 vdd.n795 242.684
R34697 vdd.n824 vdd.n782 242.684
R34698 vdd.n3500 vdd.n3496 242.684
R34699 vdd.n3519 vdd.n3515 242.684
R34700 vdd.n3452 vdd.n3448 242.684
R34701 vdd.n3471 vdd.n3467 242.684
R34702 vdd.n3549 vdd.n3545 242.684
R34703 vdd.n3568 vdd.n3564 242.684
R34704 vdd.n3599 vdd.n3595 242.684
R34705 vdd.n3618 vdd.n3614 242.684
R34706 vdd.n3647 vdd.n3643 242.684
R34707 vdd.n3666 vdd.n3662 242.684
R34708 vdd.n605 vdd.n601 242.684
R34709 vdd.n624 vdd.n620 242.684
R34710 vdd.n3746 vdd.n3742 242.684
R34711 vdd.n3765 vdd.n3761 242.684
R34712 vdd.n3698 vdd.n3694 242.684
R34713 vdd.n3717 vdd.n3713 242.684
R34714 vdd.n6888 vdd.n6884 242.684
R34715 vdd.n6907 vdd.n6903 242.684
R34716 vdd.n6840 vdd.n6836 242.684
R34717 vdd.n6859 vdd.n6855 242.684
R34718 vdd.n10030 vdd.n10026 242.684
R34719 vdd.n10049 vdd.n10045 242.684
R34720 vdd.n9982 vdd.n9978 242.684
R34721 vdd.n10001 vdd.n9997 242.684
R34722 vdd.n10078 vdd.n10074 242.684
R34723 vdd.n10097 vdd.n10093 242.684
R34724 vdd.n10126 vdd.n10122 242.684
R34725 vdd.n10145 vdd.n10141 242.684
R34726 vdd.n10228 vdd.n10224 242.684
R34727 vdd.n10247 vdd.n10243 242.684
R34728 vdd.n10276 vdd.n10272 242.684
R34729 vdd.n10295 vdd.n10291 242.684
R34730 vdd.n10324 vdd.n10320 242.684
R34731 vdd.n10343 vdd.n10339 242.684
R34732 vdd.n10372 vdd.n10368 242.684
R34733 vdd.n10391 vdd.n10387 242.684
R34734 vdd.n10474 vdd.n10470 242.684
R34735 vdd.n10493 vdd.n10489 242.684
R34736 vdd.n66 vdd.n62 242.684
R34737 vdd.n85 vdd.n81 242.684
R34738 vdd.n18 vdd.n14 242.684
R34739 vdd.n37 vdd.n33 242.684
R34740 vdd.n10522 vdd.n10518 242.684
R34741 vdd.n10541 vdd.n10537 242.684
R34742 vdd.n10572 vdd.n10568 242.684
R34743 vdd.n10591 vdd.n10587 242.684
R34744 vdd.n10620 vdd.n10616 242.684
R34745 vdd.n10639 vdd.n10635 242.684
R34746 vdd.n10426 vdd.n10418 242.684
R34747 vdd.n10447 vdd.n10405 242.684
R34748 vdd.n10768 vdd.n10764 242.684
R34749 vdd.n10787 vdd.n10783 242.684
R34750 vdd.n10719 vdd.n10715 242.684
R34751 vdd.n10738 vdd.n10734 242.684
R34752 vdd.n10671 vdd.n10667 242.684
R34753 vdd.n10690 vdd.n10686 242.684
R34754 vdd.n10817 vdd.n10813 242.684
R34755 vdd.n10836 vdd.n10832 242.684
R34756 vdd.n10867 vdd.n10863 242.684
R34757 vdd.n10886 vdd.n10882 242.684
R34758 vdd.n10915 vdd.n10911 242.684
R34759 vdd.n10934 vdd.n10930 242.684
R34760 vdd.n11013 vdd.n11009 242.684
R34761 vdd.n11032 vdd.n11028 242.684
R34762 vdd.n10965 vdd.n10961 242.684
R34763 vdd.n10984 vdd.n10980 242.684
R34764 vdd.n11062 vdd.n11058 242.684
R34765 vdd.n11081 vdd.n11077 242.684
R34766 vdd.n11112 vdd.n11108 242.684
R34767 vdd.n11131 vdd.n11127 242.684
R34768 vdd.n11160 vdd.n11156 242.684
R34769 vdd.n11179 vdd.n11175 242.684
R34770 vdd.n10180 vdd.n10172 242.684
R34771 vdd.n10201 vdd.n10159 242.684
R34772 vdd.n11259 vdd.n11255 242.684
R34773 vdd.n11278 vdd.n11274 242.684
R34774 vdd.n11211 vdd.n11207 242.684
R34775 vdd.n11230 vdd.n11226 242.684
R34776 vdd.n11308 vdd.n11304 242.684
R34777 vdd.n11327 vdd.n11323 242.684
R34778 vdd.n11358 vdd.n11354 242.684
R34779 vdd.n11377 vdd.n11373 242.684
R34780 vdd.n11406 vdd.n11402 242.684
R34781 vdd.n11425 vdd.n11421 242.684
R34782 vdd.n11475 vdd.n11472 242.684
R34783 vdd.n11522 vdd.n11519 242.684
R34784 vdd.n11572 vdd.n11569 242.684
R34785 vdd.n11622 vdd.n11619 242.684
R34786 vdd.n11670 vdd.n11667 242.684
R34787 vdd.n462 vdd.n458 242.684
R34788 vdd.n11721 vdd.n11718 242.684
R34789 vdd.n11768 vdd.n11765 242.684
R34790 vdd.n11816 vdd.n11813 242.684
R34791 vdd.n11867 vdd.n11864 242.684
R34792 vdd.n11917 vdd.n11914 242.684
R34793 vdd.n11965 vdd.n11962 242.684
R34794 vdd.n12015 vdd.n12012 242.684
R34795 vdd.n12062 vdd.n12059 242.684
R34796 vdd.n12112 vdd.n12109 242.684
R34797 vdd.n12162 vdd.n12159 242.684
R34798 vdd.n12210 vdd.n12207 242.684
R34799 vdd.n217 vdd.n213 242.684
R34800 vdd.n12261 vdd.n12258 242.684
R34801 vdd.n12308 vdd.n12305 242.684
R34802 vdd.n12358 vdd.n12355 242.684
R34803 vdd.n12408 vdd.n12405 242.684
R34804 vdd.n12456 vdd.n12453 242.684
R34805 vdd.n12507 vdd.n12498 93.7417
R34806 vdd.n12516 vdd.n12472 93.7417
R34807 vdd.n12484 vdd.n12475 93.7417
R34808 vdd.n137 vdd.n128 93.7417
R34809 vdd.n128 vdd.n99 93.7417
R34810 vdd.n126 vdd.n97 93.7417
R34811 vdd.n143 vdd.n97 93.7417
R34812 vdd.n112 vdd.n107 93.7417
R34813 vdd.n113 vdd.n112 93.7417
R34814 vdd.n185 vdd.n176 93.7417
R34815 vdd.n176 vdd.n147 93.7417
R34816 vdd.n174 vdd.n145 93.7417
R34817 vdd.n191 vdd.n145 93.7417
R34818 vdd.n160 vdd.n155 93.7417
R34819 vdd.n161 vdd.n160 93.7417
R34820 vdd.n286 vdd.n277 93.7417
R34821 vdd.n277 vdd.n248 93.7417
R34822 vdd.n275 vdd.n246 93.7417
R34823 vdd.n292 vdd.n246 93.7417
R34824 vdd.n261 vdd.n256 93.7417
R34825 vdd.n262 vdd.n261 93.7417
R34826 vdd.n334 vdd.n325 93.7417
R34827 vdd.n325 vdd.n296 93.7417
R34828 vdd.n323 vdd.n294 93.7417
R34829 vdd.n340 vdd.n294 93.7417
R34830 vdd.n309 vdd.n304 93.7417
R34831 vdd.n310 vdd.n309 93.7417
R34832 vdd.n382 vdd.n373 93.7417
R34833 vdd.n373 vdd.n344 93.7417
R34834 vdd.n371 vdd.n342 93.7417
R34835 vdd.n388 vdd.n342 93.7417
R34836 vdd.n357 vdd.n352 93.7417
R34837 vdd.n358 vdd.n357 93.7417
R34838 vdd.n430 vdd.n421 93.7417
R34839 vdd.n421 vdd.n392 93.7417
R34840 vdd.n419 vdd.n390 93.7417
R34841 vdd.n436 vdd.n390 93.7417
R34842 vdd.n405 vdd.n400 93.7417
R34843 vdd.n406 vdd.n405 93.7417
R34844 vdd.n531 vdd.n522 93.7417
R34845 vdd.n522 vdd.n493 93.7417
R34846 vdd.n520 vdd.n491 93.7417
R34847 vdd.n537 vdd.n491 93.7417
R34848 vdd.n506 vdd.n501 93.7417
R34849 vdd.n507 vdd.n506 93.7417
R34850 vdd.n579 vdd.n570 93.7417
R34851 vdd.n570 vdd.n541 93.7417
R34852 vdd.n568 vdd.n539 93.7417
R34853 vdd.n585 vdd.n539 93.7417
R34854 vdd.n554 vdd.n549 93.7417
R34855 vdd.n555 vdd.n554 93.7417
R34856 vdd.n6998 vdd.n6969 93.7417
R34857 vdd.n7007 vdd.n6998 93.7417
R34858 vdd.n7013 vdd.n6967 93.7417
R34859 vdd.n6996 vdd.n6967 93.7417
R34860 vdd.n6988 vdd.n6987 93.7417
R34861 vdd.n6987 vdd.n6977 93.7417
R34862 vdd.n7046 vdd.n7017 93.7417
R34863 vdd.n7055 vdd.n7046 93.7417
R34864 vdd.n7061 vdd.n7015 93.7417
R34865 vdd.n7044 vdd.n7015 93.7417
R34866 vdd.n7036 vdd.n7035 93.7417
R34867 vdd.n7035 vdd.n7025 93.7417
R34868 vdd.n7148 vdd.n7119 93.7417
R34869 vdd.n7157 vdd.n7148 93.7417
R34870 vdd.n7163 vdd.n7117 93.7417
R34871 vdd.n7146 vdd.n7117 93.7417
R34872 vdd.n7138 vdd.n7137 93.7417
R34873 vdd.n7137 vdd.n7127 93.7417
R34874 vdd.n7196 vdd.n7167 93.7417
R34875 vdd.n7205 vdd.n7196 93.7417
R34876 vdd.n7211 vdd.n7165 93.7417
R34877 vdd.n7194 vdd.n7165 93.7417
R34878 vdd.n7186 vdd.n7185 93.7417
R34879 vdd.n7185 vdd.n7175 93.7417
R34880 vdd.n7244 vdd.n7215 93.7417
R34881 vdd.n7253 vdd.n7244 93.7417
R34882 vdd.n7259 vdd.n7213 93.7417
R34883 vdd.n7242 vdd.n7213 93.7417
R34884 vdd.n7234 vdd.n7233 93.7417
R34885 vdd.n7233 vdd.n7223 93.7417
R34886 vdd.n7292 vdd.n7263 93.7417
R34887 vdd.n7301 vdd.n7292 93.7417
R34888 vdd.n7307 vdd.n7261 93.7417
R34889 vdd.n7290 vdd.n7261 93.7417
R34890 vdd.n7282 vdd.n7281 93.7417
R34891 vdd.n7281 vdd.n7271 93.7417
R34892 vdd.n7394 vdd.n7365 93.7417
R34893 vdd.n7403 vdd.n7394 93.7417
R34894 vdd.n7409 vdd.n7363 93.7417
R34895 vdd.n7392 vdd.n7363 93.7417
R34896 vdd.n7384 vdd.n7383 93.7417
R34897 vdd.n7383 vdd.n7373 93.7417
R34898 vdd.n8914 vdd.n8885 93.7417
R34899 vdd.n8923 vdd.n8914 93.7417
R34900 vdd.n8929 vdd.n8883 93.7417
R34901 vdd.n8912 vdd.n8883 93.7417
R34902 vdd.n8904 vdd.n8903 93.7417
R34903 vdd.n8903 vdd.n8893 93.7417
R34904 vdd.n7451 vdd.n7442 93.7417
R34905 vdd.n7442 vdd.n7413 93.7417
R34906 vdd.n7440 vdd.n7411 93.7417
R34907 vdd.n7457 vdd.n7411 93.7417
R34908 vdd.n7426 vdd.n7421 93.7417
R34909 vdd.n7427 vdd.n7426 93.7417
R34910 vdd.n7499 vdd.n7490 93.7417
R34911 vdd.n7490 vdd.n7461 93.7417
R34912 vdd.n7488 vdd.n7459 93.7417
R34913 vdd.n7505 vdd.n7459 93.7417
R34914 vdd.n7474 vdd.n7469 93.7417
R34915 vdd.n7475 vdd.n7474 93.7417
R34916 vdd.n7600 vdd.n7591 93.7417
R34917 vdd.n7591 vdd.n7562 93.7417
R34918 vdd.n7589 vdd.n7560 93.7417
R34919 vdd.n7606 vdd.n7560 93.7417
R34920 vdd.n7575 vdd.n7570 93.7417
R34921 vdd.n7576 vdd.n7575 93.7417
R34922 vdd.n7648 vdd.n7639 93.7417
R34923 vdd.n7639 vdd.n7610 93.7417
R34924 vdd.n7637 vdd.n7608 93.7417
R34925 vdd.n7654 vdd.n7608 93.7417
R34926 vdd.n7623 vdd.n7618 93.7417
R34927 vdd.n7624 vdd.n7623 93.7417
R34928 vdd.n7696 vdd.n7687 93.7417
R34929 vdd.n7687 vdd.n7658 93.7417
R34930 vdd.n7685 vdd.n7656 93.7417
R34931 vdd.n7702 vdd.n7656 93.7417
R34932 vdd.n7671 vdd.n7666 93.7417
R34933 vdd.n7672 vdd.n7671 93.7417
R34934 vdd.n7744 vdd.n7735 93.7417
R34935 vdd.n7735 vdd.n7706 93.7417
R34936 vdd.n7733 vdd.n7704 93.7417
R34937 vdd.n7750 vdd.n7704 93.7417
R34938 vdd.n7719 vdd.n7714 93.7417
R34939 vdd.n7720 vdd.n7719 93.7417
R34940 vdd.n7845 vdd.n7836 93.7417
R34941 vdd.n7836 vdd.n7807 93.7417
R34942 vdd.n7834 vdd.n7805 93.7417
R34943 vdd.n7851 vdd.n7805 93.7417
R34944 vdd.n7820 vdd.n7815 93.7417
R34945 vdd.n7821 vdd.n7820 93.7417
R34946 vdd.n6958 vdd.n6949 93.7417
R34947 vdd.n6949 vdd.n6920 93.7417
R34948 vdd.n6947 vdd.n6918 93.7417
R34949 vdd.n6964 vdd.n6918 93.7417
R34950 vdd.n6933 vdd.n6928 93.7417
R34951 vdd.n6934 vdd.n6933 93.7417
R34952 vdd.n7893 vdd.n7884 93.7417
R34953 vdd.n7884 vdd.n7855 93.7417
R34954 vdd.n7882 vdd.n7853 93.7417
R34955 vdd.n7899 vdd.n7853 93.7417
R34956 vdd.n7868 vdd.n7863 93.7417
R34957 vdd.n7869 vdd.n7868 93.7417
R34958 vdd.n7940 vdd.n7931 93.7417
R34959 vdd.n7931 vdd.n7902 93.7417
R34960 vdd.n7929 vdd.n7900 93.7417
R34961 vdd.n7946 vdd.n7900 93.7417
R34962 vdd.n7915 vdd.n7910 93.7417
R34963 vdd.n7916 vdd.n7915 93.7417
R34964 vdd.n7990 vdd.n7981 93.7417
R34965 vdd.n7981 vdd.n7952 93.7417
R34966 vdd.n7979 vdd.n7950 93.7417
R34967 vdd.n7996 vdd.n7950 93.7417
R34968 vdd.n7965 vdd.n7960 93.7417
R34969 vdd.n7966 vdd.n7965 93.7417
R34970 vdd.n8040 vdd.n8031 93.7417
R34971 vdd.n8031 vdd.n8002 93.7417
R34972 vdd.n8029 vdd.n8000 93.7417
R34973 vdd.n8046 vdd.n8000 93.7417
R34974 vdd.n8015 vdd.n8010 93.7417
R34975 vdd.n8016 vdd.n8015 93.7417
R34976 vdd.n8088 vdd.n8079 93.7417
R34977 vdd.n8079 vdd.n8050 93.7417
R34978 vdd.n8077 vdd.n8048 93.7417
R34979 vdd.n8094 vdd.n8048 93.7417
R34980 vdd.n8063 vdd.n8058 93.7417
R34981 vdd.n8064 vdd.n8063 93.7417
R34982 vdd.n7780 vdd.n7770 93.7417
R34983 vdd.n7773 vdd.n7770 93.7417
R34984 vdd.n7787 vdd.n7762 93.7417
R34985 vdd.n7788 vdd.n7787 93.7417
R34986 vdd.n7794 vdd.n7761 93.7417
R34987 vdd.n7761 vdd.n7755 93.7417
R34988 vdd.n8139 vdd.n8130 93.7417
R34989 vdd.n8130 vdd.n8101 93.7417
R34990 vdd.n8128 vdd.n8099 93.7417
R34991 vdd.n8145 vdd.n8099 93.7417
R34992 vdd.n8114 vdd.n8109 93.7417
R34993 vdd.n8115 vdd.n8114 93.7417
R34994 vdd.n8186 vdd.n8177 93.7417
R34995 vdd.n8177 vdd.n8148 93.7417
R34996 vdd.n8175 vdd.n8146 93.7417
R34997 vdd.n8192 vdd.n8146 93.7417
R34998 vdd.n8161 vdd.n8156 93.7417
R34999 vdd.n8162 vdd.n8161 93.7417
R35000 vdd.n8234 vdd.n8225 93.7417
R35001 vdd.n8225 vdd.n8196 93.7417
R35002 vdd.n8223 vdd.n8194 93.7417
R35003 vdd.n8240 vdd.n8194 93.7417
R35004 vdd.n8209 vdd.n8204 93.7417
R35005 vdd.n8210 vdd.n8209 93.7417
R35006 vdd.n8285 vdd.n8276 93.7417
R35007 vdd.n8276 vdd.n8247 93.7417
R35008 vdd.n8274 vdd.n8245 93.7417
R35009 vdd.n8291 vdd.n8245 93.7417
R35010 vdd.n8260 vdd.n8255 93.7417
R35011 vdd.n8261 vdd.n8260 93.7417
R35012 vdd.n8335 vdd.n8326 93.7417
R35013 vdd.n8326 vdd.n8297 93.7417
R35014 vdd.n8324 vdd.n8295 93.7417
R35015 vdd.n8341 vdd.n8295 93.7417
R35016 vdd.n8310 vdd.n8305 93.7417
R35017 vdd.n8311 vdd.n8310 93.7417
R35018 vdd.n8383 vdd.n8374 93.7417
R35019 vdd.n8374 vdd.n8345 93.7417
R35020 vdd.n8372 vdd.n8343 93.7417
R35021 vdd.n8389 vdd.n8343 93.7417
R35022 vdd.n8358 vdd.n8353 93.7417
R35023 vdd.n8359 vdd.n8358 93.7417
R35024 vdd.n8433 vdd.n8424 93.7417
R35025 vdd.n8424 vdd.n8395 93.7417
R35026 vdd.n8422 vdd.n8393 93.7417
R35027 vdd.n8439 vdd.n8393 93.7417
R35028 vdd.n8408 vdd.n8403 93.7417
R35029 vdd.n8409 vdd.n8408 93.7417
R35030 vdd.n8480 vdd.n8471 93.7417
R35031 vdd.n8471 vdd.n8442 93.7417
R35032 vdd.n8469 vdd.n8440 93.7417
R35033 vdd.n8486 vdd.n8440 93.7417
R35034 vdd.n8455 vdd.n8450 93.7417
R35035 vdd.n8456 vdd.n8455 93.7417
R35036 vdd.n8530 vdd.n8521 93.7417
R35037 vdd.n8521 vdd.n8492 93.7417
R35038 vdd.n8519 vdd.n8490 93.7417
R35039 vdd.n8536 vdd.n8490 93.7417
R35040 vdd.n8505 vdd.n8500 93.7417
R35041 vdd.n8506 vdd.n8505 93.7417
R35042 vdd.n8580 vdd.n8571 93.7417
R35043 vdd.n8571 vdd.n8542 93.7417
R35044 vdd.n8569 vdd.n8540 93.7417
R35045 vdd.n8586 vdd.n8540 93.7417
R35046 vdd.n8555 vdd.n8550 93.7417
R35047 vdd.n8556 vdd.n8555 93.7417
R35048 vdd.n8628 vdd.n8619 93.7417
R35049 vdd.n8619 vdd.n8590 93.7417
R35050 vdd.n8617 vdd.n8588 93.7417
R35051 vdd.n8634 vdd.n8588 93.7417
R35052 vdd.n8603 vdd.n8598 93.7417
R35053 vdd.n8604 vdd.n8603 93.7417
R35054 vdd.n7535 vdd.n7525 93.7417
R35055 vdd.n7528 vdd.n7525 93.7417
R35056 vdd.n7542 vdd.n7517 93.7417
R35057 vdd.n7543 vdd.n7542 93.7417
R35058 vdd.n7549 vdd.n7516 93.7417
R35059 vdd.n7516 vdd.n7510 93.7417
R35060 vdd.n8679 vdd.n8670 93.7417
R35061 vdd.n8670 vdd.n8641 93.7417
R35062 vdd.n8668 vdd.n8639 93.7417
R35063 vdd.n8685 vdd.n8639 93.7417
R35064 vdd.n8654 vdd.n8649 93.7417
R35065 vdd.n8655 vdd.n8654 93.7417
R35066 vdd.n8726 vdd.n8717 93.7417
R35067 vdd.n8717 vdd.n8688 93.7417
R35068 vdd.n8715 vdd.n8686 93.7417
R35069 vdd.n8732 vdd.n8686 93.7417
R35070 vdd.n8701 vdd.n8696 93.7417
R35071 vdd.n8702 vdd.n8701 93.7417
R35072 vdd.n8776 vdd.n8767 93.7417
R35073 vdd.n8767 vdd.n8738 93.7417
R35074 vdd.n8765 vdd.n8736 93.7417
R35075 vdd.n8782 vdd.n8736 93.7417
R35076 vdd.n8751 vdd.n8746 93.7417
R35077 vdd.n8752 vdd.n8751 93.7417
R35078 vdd.n8826 vdd.n8817 93.7417
R35079 vdd.n8817 vdd.n8788 93.7417
R35080 vdd.n8815 vdd.n8786 93.7417
R35081 vdd.n8832 vdd.n8786 93.7417
R35082 vdd.n8801 vdd.n8796 93.7417
R35083 vdd.n8802 vdd.n8801 93.7417
R35084 vdd.n8874 vdd.n8865 93.7417
R35085 vdd.n8865 vdd.n8836 93.7417
R35086 vdd.n8863 vdd.n8834 93.7417
R35087 vdd.n8880 vdd.n8834 93.7417
R35088 vdd.n8849 vdd.n8844 93.7417
R35089 vdd.n8850 vdd.n8849 93.7417
R35090 vdd.n9011 vdd.n8982 93.7417
R35091 vdd.n9020 vdd.n9011 93.7417
R35092 vdd.n9026 vdd.n8980 93.7417
R35093 vdd.n9009 vdd.n8980 93.7417
R35094 vdd.n9001 vdd.n9000 93.7417
R35095 vdd.n9000 vdd.n8990 93.7417
R35096 vdd.n8963 vdd.n8934 93.7417
R35097 vdd.n8972 vdd.n8963 93.7417
R35098 vdd.n8978 vdd.n8932 93.7417
R35099 vdd.n8961 vdd.n8932 93.7417
R35100 vdd.n8953 vdd.n8952 93.7417
R35101 vdd.n8952 vdd.n8942 93.7417
R35102 vdd.n9060 vdd.n9031 93.7417
R35103 vdd.n9069 vdd.n9060 93.7417
R35104 vdd.n9075 vdd.n9029 93.7417
R35105 vdd.n9058 vdd.n9029 93.7417
R35106 vdd.n9050 vdd.n9049 93.7417
R35107 vdd.n9049 vdd.n9039 93.7417
R35108 vdd.n9110 vdd.n9081 93.7417
R35109 vdd.n9119 vdd.n9110 93.7417
R35110 vdd.n9125 vdd.n9079 93.7417
R35111 vdd.n9108 vdd.n9079 93.7417
R35112 vdd.n9100 vdd.n9099 93.7417
R35113 vdd.n9099 vdd.n9089 93.7417
R35114 vdd.n9158 vdd.n9129 93.7417
R35115 vdd.n9167 vdd.n9158 93.7417
R35116 vdd.n9173 vdd.n9127 93.7417
R35117 vdd.n9156 vdd.n9127 93.7417
R35118 vdd.n9148 vdd.n9147 93.7417
R35119 vdd.n9147 vdd.n9137 93.7417
R35120 vdd.n7349 vdd.n7348 93.7417
R35121 vdd.n7349 vdd.n7313 93.7417
R35122 vdd.n7346 vdd.n7345 93.7417
R35123 vdd.n7345 vdd.n7317 93.7417
R35124 vdd.n7336 vdd.n7323 93.7417
R35125 vdd.n7329 vdd.n7323 93.7417
R35126 vdd.n9306 vdd.n9277 93.7417
R35127 vdd.n9315 vdd.n9306 93.7417
R35128 vdd.n9321 vdd.n9275 93.7417
R35129 vdd.n9304 vdd.n9275 93.7417
R35130 vdd.n9296 vdd.n9295 93.7417
R35131 vdd.n9295 vdd.n9285 93.7417
R35132 vdd.n9257 vdd.n9228 93.7417
R35133 vdd.n9266 vdd.n9257 93.7417
R35134 vdd.n9272 vdd.n9226 93.7417
R35135 vdd.n9255 vdd.n9226 93.7417
R35136 vdd.n9247 vdd.n9246 93.7417
R35137 vdd.n9246 vdd.n9236 93.7417
R35138 vdd.n9209 vdd.n9180 93.7417
R35139 vdd.n9218 vdd.n9209 93.7417
R35140 vdd.n9224 vdd.n9178 93.7417
R35141 vdd.n9207 vdd.n9178 93.7417
R35142 vdd.n9199 vdd.n9198 93.7417
R35143 vdd.n9198 vdd.n9188 93.7417
R35144 vdd.n9355 vdd.n9326 93.7417
R35145 vdd.n9364 vdd.n9355 93.7417
R35146 vdd.n9370 vdd.n9324 93.7417
R35147 vdd.n9353 vdd.n9324 93.7417
R35148 vdd.n9345 vdd.n9344 93.7417
R35149 vdd.n9344 vdd.n9334 93.7417
R35150 vdd.n9405 vdd.n9376 93.7417
R35151 vdd.n9414 vdd.n9405 93.7417
R35152 vdd.n9420 vdd.n9374 93.7417
R35153 vdd.n9403 vdd.n9374 93.7417
R35154 vdd.n9395 vdd.n9394 93.7417
R35155 vdd.n9394 vdd.n9384 93.7417
R35156 vdd.n9453 vdd.n9424 93.7417
R35157 vdd.n9462 vdd.n9453 93.7417
R35158 vdd.n9468 vdd.n9422 93.7417
R35159 vdd.n9451 vdd.n9422 93.7417
R35160 vdd.n9443 vdd.n9442 93.7417
R35161 vdd.n9442 vdd.n9432 93.7417
R35162 vdd.n9551 vdd.n9522 93.7417
R35163 vdd.n9560 vdd.n9551 93.7417
R35164 vdd.n9566 vdd.n9520 93.7417
R35165 vdd.n9549 vdd.n9520 93.7417
R35166 vdd.n9541 vdd.n9540 93.7417
R35167 vdd.n9540 vdd.n9530 93.7417
R35168 vdd.n9503 vdd.n9474 93.7417
R35169 vdd.n9512 vdd.n9503 93.7417
R35170 vdd.n9518 vdd.n9472 93.7417
R35171 vdd.n9501 vdd.n9472 93.7417
R35172 vdd.n9493 vdd.n9492 93.7417
R35173 vdd.n9492 vdd.n9482 93.7417
R35174 vdd.n9600 vdd.n9571 93.7417
R35175 vdd.n9609 vdd.n9600 93.7417
R35176 vdd.n9615 vdd.n9569 93.7417
R35177 vdd.n9598 vdd.n9569 93.7417
R35178 vdd.n9590 vdd.n9589 93.7417
R35179 vdd.n9589 vdd.n9579 93.7417
R35180 vdd.n9650 vdd.n9621 93.7417
R35181 vdd.n9659 vdd.n9650 93.7417
R35182 vdd.n9665 vdd.n9619 93.7417
R35183 vdd.n9648 vdd.n9619 93.7417
R35184 vdd.n9640 vdd.n9639 93.7417
R35185 vdd.n9639 vdd.n9629 93.7417
R35186 vdd.n9698 vdd.n9669 93.7417
R35187 vdd.n9707 vdd.n9698 93.7417
R35188 vdd.n9713 vdd.n9667 93.7417
R35189 vdd.n9696 vdd.n9667 93.7417
R35190 vdd.n9688 vdd.n9687 93.7417
R35191 vdd.n9687 vdd.n9677 93.7417
R35192 vdd.n7103 vdd.n7102 93.7417
R35193 vdd.n7103 vdd.n7067 93.7417
R35194 vdd.n7100 vdd.n7099 93.7417
R35195 vdd.n7099 vdd.n7071 93.7417
R35196 vdd.n7090 vdd.n7077 93.7417
R35197 vdd.n7083 vdd.n7077 93.7417
R35198 vdd.n9797 vdd.n9768 93.7417
R35199 vdd.n9806 vdd.n9797 93.7417
R35200 vdd.n9812 vdd.n9766 93.7417
R35201 vdd.n9795 vdd.n9766 93.7417
R35202 vdd.n9787 vdd.n9786 93.7417
R35203 vdd.n9786 vdd.n9776 93.7417
R35204 vdd.n9749 vdd.n9720 93.7417
R35205 vdd.n9758 vdd.n9749 93.7417
R35206 vdd.n9764 vdd.n9718 93.7417
R35207 vdd.n9747 vdd.n9718 93.7417
R35208 vdd.n9739 vdd.n9738 93.7417
R35209 vdd.n9738 vdd.n9728 93.7417
R35210 vdd.n9846 vdd.n9817 93.7417
R35211 vdd.n9855 vdd.n9846 93.7417
R35212 vdd.n9861 vdd.n9815 93.7417
R35213 vdd.n9844 vdd.n9815 93.7417
R35214 vdd.n9836 vdd.n9835 93.7417
R35215 vdd.n9835 vdd.n9825 93.7417
R35216 vdd.n9896 vdd.n9867 93.7417
R35217 vdd.n9905 vdd.n9896 93.7417
R35218 vdd.n9911 vdd.n9865 93.7417
R35219 vdd.n9894 vdd.n9865 93.7417
R35220 vdd.n9886 vdd.n9885 93.7417
R35221 vdd.n9885 vdd.n9875 93.7417
R35222 vdd.n9944 vdd.n9915 93.7417
R35223 vdd.n9953 vdd.n9944 93.7417
R35224 vdd.n9959 vdd.n9913 93.7417
R35225 vdd.n9942 vdd.n9913 93.7417
R35226 vdd.n9934 vdd.n9933 93.7417
R35227 vdd.n9933 vdd.n9923 93.7417
R35228 vdd.n3856 vdd.n3827 93.7417
R35229 vdd.n3865 vdd.n3856 93.7417
R35230 vdd.n3871 vdd.n3825 93.7417
R35231 vdd.n3854 vdd.n3825 93.7417
R35232 vdd.n3846 vdd.n3845 93.7417
R35233 vdd.n3845 vdd.n3835 93.7417
R35234 vdd.n3904 vdd.n3875 93.7417
R35235 vdd.n3913 vdd.n3904 93.7417
R35236 vdd.n3919 vdd.n3873 93.7417
R35237 vdd.n3902 vdd.n3873 93.7417
R35238 vdd.n3894 vdd.n3893 93.7417
R35239 vdd.n3893 vdd.n3883 93.7417
R35240 vdd.n4006 vdd.n3977 93.7417
R35241 vdd.n4015 vdd.n4006 93.7417
R35242 vdd.n4021 vdd.n3975 93.7417
R35243 vdd.n4004 vdd.n3975 93.7417
R35244 vdd.n3996 vdd.n3995 93.7417
R35245 vdd.n3995 vdd.n3985 93.7417
R35246 vdd.n4054 vdd.n4025 93.7417
R35247 vdd.n4063 vdd.n4054 93.7417
R35248 vdd.n4069 vdd.n4023 93.7417
R35249 vdd.n4052 vdd.n4023 93.7417
R35250 vdd.n4044 vdd.n4043 93.7417
R35251 vdd.n4043 vdd.n4033 93.7417
R35252 vdd.n4102 vdd.n4073 93.7417
R35253 vdd.n4111 vdd.n4102 93.7417
R35254 vdd.n4117 vdd.n4071 93.7417
R35255 vdd.n4100 vdd.n4071 93.7417
R35256 vdd.n4092 vdd.n4091 93.7417
R35257 vdd.n4091 vdd.n4081 93.7417
R35258 vdd.n4150 vdd.n4121 93.7417
R35259 vdd.n4159 vdd.n4150 93.7417
R35260 vdd.n4165 vdd.n4119 93.7417
R35261 vdd.n4148 vdd.n4119 93.7417
R35262 vdd.n4140 vdd.n4139 93.7417
R35263 vdd.n4139 vdd.n4129 93.7417
R35264 vdd.n4252 vdd.n4223 93.7417
R35265 vdd.n4261 vdd.n4252 93.7417
R35266 vdd.n4267 vdd.n4221 93.7417
R35267 vdd.n4250 vdd.n4221 93.7417
R35268 vdd.n4242 vdd.n4241 93.7417
R35269 vdd.n4241 vdd.n4231 93.7417
R35270 vdd.n5772 vdd.n5743 93.7417
R35271 vdd.n5781 vdd.n5772 93.7417
R35272 vdd.n5787 vdd.n5741 93.7417
R35273 vdd.n5770 vdd.n5741 93.7417
R35274 vdd.n5762 vdd.n5761 93.7417
R35275 vdd.n5761 vdd.n5751 93.7417
R35276 vdd.n4309 vdd.n4300 93.7417
R35277 vdd.n4300 vdd.n4271 93.7417
R35278 vdd.n4298 vdd.n4269 93.7417
R35279 vdd.n4315 vdd.n4269 93.7417
R35280 vdd.n4284 vdd.n4279 93.7417
R35281 vdd.n4285 vdd.n4284 93.7417
R35282 vdd.n4357 vdd.n4348 93.7417
R35283 vdd.n4348 vdd.n4319 93.7417
R35284 vdd.n4346 vdd.n4317 93.7417
R35285 vdd.n4363 vdd.n4317 93.7417
R35286 vdd.n4332 vdd.n4327 93.7417
R35287 vdd.n4333 vdd.n4332 93.7417
R35288 vdd.n4458 vdd.n4449 93.7417
R35289 vdd.n4449 vdd.n4420 93.7417
R35290 vdd.n4447 vdd.n4418 93.7417
R35291 vdd.n4464 vdd.n4418 93.7417
R35292 vdd.n4433 vdd.n4428 93.7417
R35293 vdd.n4434 vdd.n4433 93.7417
R35294 vdd.n4506 vdd.n4497 93.7417
R35295 vdd.n4497 vdd.n4468 93.7417
R35296 vdd.n4495 vdd.n4466 93.7417
R35297 vdd.n4512 vdd.n4466 93.7417
R35298 vdd.n4481 vdd.n4476 93.7417
R35299 vdd.n4482 vdd.n4481 93.7417
R35300 vdd.n4554 vdd.n4545 93.7417
R35301 vdd.n4545 vdd.n4516 93.7417
R35302 vdd.n4543 vdd.n4514 93.7417
R35303 vdd.n4560 vdd.n4514 93.7417
R35304 vdd.n4529 vdd.n4524 93.7417
R35305 vdd.n4530 vdd.n4529 93.7417
R35306 vdd.n4602 vdd.n4593 93.7417
R35307 vdd.n4593 vdd.n4564 93.7417
R35308 vdd.n4591 vdd.n4562 93.7417
R35309 vdd.n4608 vdd.n4562 93.7417
R35310 vdd.n4577 vdd.n4572 93.7417
R35311 vdd.n4578 vdd.n4577 93.7417
R35312 vdd.n4703 vdd.n4694 93.7417
R35313 vdd.n4694 vdd.n4665 93.7417
R35314 vdd.n4692 vdd.n4663 93.7417
R35315 vdd.n4709 vdd.n4663 93.7417
R35316 vdd.n4678 vdd.n4673 93.7417
R35317 vdd.n4679 vdd.n4678 93.7417
R35318 vdd.n3816 vdd.n3807 93.7417
R35319 vdd.n3807 vdd.n3778 93.7417
R35320 vdd.n3805 vdd.n3776 93.7417
R35321 vdd.n3822 vdd.n3776 93.7417
R35322 vdd.n3791 vdd.n3786 93.7417
R35323 vdd.n3792 vdd.n3791 93.7417
R35324 vdd.n4751 vdd.n4742 93.7417
R35325 vdd.n4742 vdd.n4713 93.7417
R35326 vdd.n4740 vdd.n4711 93.7417
R35327 vdd.n4757 vdd.n4711 93.7417
R35328 vdd.n4726 vdd.n4721 93.7417
R35329 vdd.n4727 vdd.n4726 93.7417
R35330 vdd.n4798 vdd.n4789 93.7417
R35331 vdd.n4789 vdd.n4760 93.7417
R35332 vdd.n4787 vdd.n4758 93.7417
R35333 vdd.n4804 vdd.n4758 93.7417
R35334 vdd.n4773 vdd.n4768 93.7417
R35335 vdd.n4774 vdd.n4773 93.7417
R35336 vdd.n4848 vdd.n4839 93.7417
R35337 vdd.n4839 vdd.n4810 93.7417
R35338 vdd.n4837 vdd.n4808 93.7417
R35339 vdd.n4854 vdd.n4808 93.7417
R35340 vdd.n4823 vdd.n4818 93.7417
R35341 vdd.n4824 vdd.n4823 93.7417
R35342 vdd.n4898 vdd.n4889 93.7417
R35343 vdd.n4889 vdd.n4860 93.7417
R35344 vdd.n4887 vdd.n4858 93.7417
R35345 vdd.n4904 vdd.n4858 93.7417
R35346 vdd.n4873 vdd.n4868 93.7417
R35347 vdd.n4874 vdd.n4873 93.7417
R35348 vdd.n4946 vdd.n4937 93.7417
R35349 vdd.n4937 vdd.n4908 93.7417
R35350 vdd.n4935 vdd.n4906 93.7417
R35351 vdd.n4952 vdd.n4906 93.7417
R35352 vdd.n4921 vdd.n4916 93.7417
R35353 vdd.n4922 vdd.n4921 93.7417
R35354 vdd.n4638 vdd.n4628 93.7417
R35355 vdd.n4631 vdd.n4628 93.7417
R35356 vdd.n4645 vdd.n4620 93.7417
R35357 vdd.n4646 vdd.n4645 93.7417
R35358 vdd.n4652 vdd.n4619 93.7417
R35359 vdd.n4619 vdd.n4613 93.7417
R35360 vdd.n4997 vdd.n4988 93.7417
R35361 vdd.n4988 vdd.n4959 93.7417
R35362 vdd.n4986 vdd.n4957 93.7417
R35363 vdd.n5003 vdd.n4957 93.7417
R35364 vdd.n4972 vdd.n4967 93.7417
R35365 vdd.n4973 vdd.n4972 93.7417
R35366 vdd.n5044 vdd.n5035 93.7417
R35367 vdd.n5035 vdd.n5006 93.7417
R35368 vdd.n5033 vdd.n5004 93.7417
R35369 vdd.n5050 vdd.n5004 93.7417
R35370 vdd.n5019 vdd.n5014 93.7417
R35371 vdd.n5020 vdd.n5019 93.7417
R35372 vdd.n5092 vdd.n5083 93.7417
R35373 vdd.n5083 vdd.n5054 93.7417
R35374 vdd.n5081 vdd.n5052 93.7417
R35375 vdd.n5098 vdd.n5052 93.7417
R35376 vdd.n5067 vdd.n5062 93.7417
R35377 vdd.n5068 vdd.n5067 93.7417
R35378 vdd.n5143 vdd.n5134 93.7417
R35379 vdd.n5134 vdd.n5105 93.7417
R35380 vdd.n5132 vdd.n5103 93.7417
R35381 vdd.n5149 vdd.n5103 93.7417
R35382 vdd.n5118 vdd.n5113 93.7417
R35383 vdd.n5119 vdd.n5118 93.7417
R35384 vdd.n5193 vdd.n5184 93.7417
R35385 vdd.n5184 vdd.n5155 93.7417
R35386 vdd.n5182 vdd.n5153 93.7417
R35387 vdd.n5199 vdd.n5153 93.7417
R35388 vdd.n5168 vdd.n5163 93.7417
R35389 vdd.n5169 vdd.n5168 93.7417
R35390 vdd.n5241 vdd.n5232 93.7417
R35391 vdd.n5232 vdd.n5203 93.7417
R35392 vdd.n5230 vdd.n5201 93.7417
R35393 vdd.n5247 vdd.n5201 93.7417
R35394 vdd.n5216 vdd.n5211 93.7417
R35395 vdd.n5217 vdd.n5216 93.7417
R35396 vdd.n5291 vdd.n5282 93.7417
R35397 vdd.n5282 vdd.n5253 93.7417
R35398 vdd.n5280 vdd.n5251 93.7417
R35399 vdd.n5297 vdd.n5251 93.7417
R35400 vdd.n5266 vdd.n5261 93.7417
R35401 vdd.n5267 vdd.n5266 93.7417
R35402 vdd.n5338 vdd.n5329 93.7417
R35403 vdd.n5329 vdd.n5300 93.7417
R35404 vdd.n5327 vdd.n5298 93.7417
R35405 vdd.n5344 vdd.n5298 93.7417
R35406 vdd.n5313 vdd.n5308 93.7417
R35407 vdd.n5314 vdd.n5313 93.7417
R35408 vdd.n5388 vdd.n5379 93.7417
R35409 vdd.n5379 vdd.n5350 93.7417
R35410 vdd.n5377 vdd.n5348 93.7417
R35411 vdd.n5394 vdd.n5348 93.7417
R35412 vdd.n5363 vdd.n5358 93.7417
R35413 vdd.n5364 vdd.n5363 93.7417
R35414 vdd.n5438 vdd.n5429 93.7417
R35415 vdd.n5429 vdd.n5400 93.7417
R35416 vdd.n5427 vdd.n5398 93.7417
R35417 vdd.n5444 vdd.n5398 93.7417
R35418 vdd.n5413 vdd.n5408 93.7417
R35419 vdd.n5414 vdd.n5413 93.7417
R35420 vdd.n5486 vdd.n5477 93.7417
R35421 vdd.n5477 vdd.n5448 93.7417
R35422 vdd.n5475 vdd.n5446 93.7417
R35423 vdd.n5492 vdd.n5446 93.7417
R35424 vdd.n5461 vdd.n5456 93.7417
R35425 vdd.n5462 vdd.n5461 93.7417
R35426 vdd.n4393 vdd.n4383 93.7417
R35427 vdd.n4386 vdd.n4383 93.7417
R35428 vdd.n4400 vdd.n4375 93.7417
R35429 vdd.n4401 vdd.n4400 93.7417
R35430 vdd.n4407 vdd.n4374 93.7417
R35431 vdd.n4374 vdd.n4368 93.7417
R35432 vdd.n5537 vdd.n5528 93.7417
R35433 vdd.n5528 vdd.n5499 93.7417
R35434 vdd.n5526 vdd.n5497 93.7417
R35435 vdd.n5543 vdd.n5497 93.7417
R35436 vdd.n5512 vdd.n5507 93.7417
R35437 vdd.n5513 vdd.n5512 93.7417
R35438 vdd.n5584 vdd.n5575 93.7417
R35439 vdd.n5575 vdd.n5546 93.7417
R35440 vdd.n5573 vdd.n5544 93.7417
R35441 vdd.n5590 vdd.n5544 93.7417
R35442 vdd.n5559 vdd.n5554 93.7417
R35443 vdd.n5560 vdd.n5559 93.7417
R35444 vdd.n5634 vdd.n5625 93.7417
R35445 vdd.n5625 vdd.n5596 93.7417
R35446 vdd.n5623 vdd.n5594 93.7417
R35447 vdd.n5640 vdd.n5594 93.7417
R35448 vdd.n5609 vdd.n5604 93.7417
R35449 vdd.n5610 vdd.n5609 93.7417
R35450 vdd.n5684 vdd.n5675 93.7417
R35451 vdd.n5675 vdd.n5646 93.7417
R35452 vdd.n5673 vdd.n5644 93.7417
R35453 vdd.n5690 vdd.n5644 93.7417
R35454 vdd.n5659 vdd.n5654 93.7417
R35455 vdd.n5660 vdd.n5659 93.7417
R35456 vdd.n5732 vdd.n5723 93.7417
R35457 vdd.n5723 vdd.n5694 93.7417
R35458 vdd.n5721 vdd.n5692 93.7417
R35459 vdd.n5738 vdd.n5692 93.7417
R35460 vdd.n5707 vdd.n5702 93.7417
R35461 vdd.n5708 vdd.n5707 93.7417
R35462 vdd.n5869 vdd.n5840 93.7417
R35463 vdd.n5878 vdd.n5869 93.7417
R35464 vdd.n5884 vdd.n5838 93.7417
R35465 vdd.n5867 vdd.n5838 93.7417
R35466 vdd.n5859 vdd.n5858 93.7417
R35467 vdd.n5858 vdd.n5848 93.7417
R35468 vdd.n5821 vdd.n5792 93.7417
R35469 vdd.n5830 vdd.n5821 93.7417
R35470 vdd.n5836 vdd.n5790 93.7417
R35471 vdd.n5819 vdd.n5790 93.7417
R35472 vdd.n5811 vdd.n5810 93.7417
R35473 vdd.n5810 vdd.n5800 93.7417
R35474 vdd.n5918 vdd.n5889 93.7417
R35475 vdd.n5927 vdd.n5918 93.7417
R35476 vdd.n5933 vdd.n5887 93.7417
R35477 vdd.n5916 vdd.n5887 93.7417
R35478 vdd.n5908 vdd.n5907 93.7417
R35479 vdd.n5907 vdd.n5897 93.7417
R35480 vdd.n5968 vdd.n5939 93.7417
R35481 vdd.n5977 vdd.n5968 93.7417
R35482 vdd.n5983 vdd.n5937 93.7417
R35483 vdd.n5966 vdd.n5937 93.7417
R35484 vdd.n5958 vdd.n5957 93.7417
R35485 vdd.n5957 vdd.n5947 93.7417
R35486 vdd.n6016 vdd.n5987 93.7417
R35487 vdd.n6025 vdd.n6016 93.7417
R35488 vdd.n6031 vdd.n5985 93.7417
R35489 vdd.n6014 vdd.n5985 93.7417
R35490 vdd.n6006 vdd.n6005 93.7417
R35491 vdd.n6005 vdd.n5995 93.7417
R35492 vdd.n4207 vdd.n4206 93.7417
R35493 vdd.n4207 vdd.n4171 93.7417
R35494 vdd.n4204 vdd.n4203 93.7417
R35495 vdd.n4203 vdd.n4175 93.7417
R35496 vdd.n4194 vdd.n4181 93.7417
R35497 vdd.n4187 vdd.n4181 93.7417
R35498 vdd.n6164 vdd.n6135 93.7417
R35499 vdd.n6173 vdd.n6164 93.7417
R35500 vdd.n6179 vdd.n6133 93.7417
R35501 vdd.n6162 vdd.n6133 93.7417
R35502 vdd.n6154 vdd.n6153 93.7417
R35503 vdd.n6153 vdd.n6143 93.7417
R35504 vdd.n6115 vdd.n6086 93.7417
R35505 vdd.n6124 vdd.n6115 93.7417
R35506 vdd.n6130 vdd.n6084 93.7417
R35507 vdd.n6113 vdd.n6084 93.7417
R35508 vdd.n6105 vdd.n6104 93.7417
R35509 vdd.n6104 vdd.n6094 93.7417
R35510 vdd.n6067 vdd.n6038 93.7417
R35511 vdd.n6076 vdd.n6067 93.7417
R35512 vdd.n6082 vdd.n6036 93.7417
R35513 vdd.n6065 vdd.n6036 93.7417
R35514 vdd.n6057 vdd.n6056 93.7417
R35515 vdd.n6056 vdd.n6046 93.7417
R35516 vdd.n6213 vdd.n6184 93.7417
R35517 vdd.n6222 vdd.n6213 93.7417
R35518 vdd.n6228 vdd.n6182 93.7417
R35519 vdd.n6211 vdd.n6182 93.7417
R35520 vdd.n6203 vdd.n6202 93.7417
R35521 vdd.n6202 vdd.n6192 93.7417
R35522 vdd.n6263 vdd.n6234 93.7417
R35523 vdd.n6272 vdd.n6263 93.7417
R35524 vdd.n6278 vdd.n6232 93.7417
R35525 vdd.n6261 vdd.n6232 93.7417
R35526 vdd.n6253 vdd.n6252 93.7417
R35527 vdd.n6252 vdd.n6242 93.7417
R35528 vdd.n6311 vdd.n6282 93.7417
R35529 vdd.n6320 vdd.n6311 93.7417
R35530 vdd.n6326 vdd.n6280 93.7417
R35531 vdd.n6309 vdd.n6280 93.7417
R35532 vdd.n6301 vdd.n6300 93.7417
R35533 vdd.n6300 vdd.n6290 93.7417
R35534 vdd.n6409 vdd.n6380 93.7417
R35535 vdd.n6418 vdd.n6409 93.7417
R35536 vdd.n6424 vdd.n6378 93.7417
R35537 vdd.n6407 vdd.n6378 93.7417
R35538 vdd.n6399 vdd.n6398 93.7417
R35539 vdd.n6398 vdd.n6388 93.7417
R35540 vdd.n6361 vdd.n6332 93.7417
R35541 vdd.n6370 vdd.n6361 93.7417
R35542 vdd.n6376 vdd.n6330 93.7417
R35543 vdd.n6359 vdd.n6330 93.7417
R35544 vdd.n6351 vdd.n6350 93.7417
R35545 vdd.n6350 vdd.n6340 93.7417
R35546 vdd.n6458 vdd.n6429 93.7417
R35547 vdd.n6467 vdd.n6458 93.7417
R35548 vdd.n6473 vdd.n6427 93.7417
R35549 vdd.n6456 vdd.n6427 93.7417
R35550 vdd.n6448 vdd.n6447 93.7417
R35551 vdd.n6447 vdd.n6437 93.7417
R35552 vdd.n6508 vdd.n6479 93.7417
R35553 vdd.n6517 vdd.n6508 93.7417
R35554 vdd.n6523 vdd.n6477 93.7417
R35555 vdd.n6506 vdd.n6477 93.7417
R35556 vdd.n6498 vdd.n6497 93.7417
R35557 vdd.n6497 vdd.n6487 93.7417
R35558 vdd.n6556 vdd.n6527 93.7417
R35559 vdd.n6565 vdd.n6556 93.7417
R35560 vdd.n6571 vdd.n6525 93.7417
R35561 vdd.n6554 vdd.n6525 93.7417
R35562 vdd.n6546 vdd.n6545 93.7417
R35563 vdd.n6545 vdd.n6535 93.7417
R35564 vdd.n3961 vdd.n3960 93.7417
R35565 vdd.n3961 vdd.n3925 93.7417
R35566 vdd.n3958 vdd.n3957 93.7417
R35567 vdd.n3957 vdd.n3929 93.7417
R35568 vdd.n3948 vdd.n3935 93.7417
R35569 vdd.n3941 vdd.n3935 93.7417
R35570 vdd.n6655 vdd.n6626 93.7417
R35571 vdd.n6664 vdd.n6655 93.7417
R35572 vdd.n6670 vdd.n6624 93.7417
R35573 vdd.n6653 vdd.n6624 93.7417
R35574 vdd.n6645 vdd.n6644 93.7417
R35575 vdd.n6644 vdd.n6634 93.7417
R35576 vdd.n6607 vdd.n6578 93.7417
R35577 vdd.n6616 vdd.n6607 93.7417
R35578 vdd.n6622 vdd.n6576 93.7417
R35579 vdd.n6605 vdd.n6576 93.7417
R35580 vdd.n6597 vdd.n6596 93.7417
R35581 vdd.n6596 vdd.n6586 93.7417
R35582 vdd.n6704 vdd.n6675 93.7417
R35583 vdd.n6713 vdd.n6704 93.7417
R35584 vdd.n6719 vdd.n6673 93.7417
R35585 vdd.n6702 vdd.n6673 93.7417
R35586 vdd.n6694 vdd.n6693 93.7417
R35587 vdd.n6693 vdd.n6683 93.7417
R35588 vdd.n6754 vdd.n6725 93.7417
R35589 vdd.n6763 vdd.n6754 93.7417
R35590 vdd.n6769 vdd.n6723 93.7417
R35591 vdd.n6752 vdd.n6723 93.7417
R35592 vdd.n6744 vdd.n6743 93.7417
R35593 vdd.n6743 vdd.n6733 93.7417
R35594 vdd.n6802 vdd.n6773 93.7417
R35595 vdd.n6811 vdd.n6802 93.7417
R35596 vdd.n6817 vdd.n6771 93.7417
R35597 vdd.n6800 vdd.n6771 93.7417
R35598 vdd.n6792 vdd.n6791 93.7417
R35599 vdd.n6791 vdd.n6781 93.7417
R35600 vdd.n714 vdd.n685 93.7417
R35601 vdd.n723 vdd.n714 93.7417
R35602 vdd.n729 vdd.n683 93.7417
R35603 vdd.n712 vdd.n683 93.7417
R35604 vdd.n704 vdd.n703 93.7417
R35605 vdd.n703 vdd.n693 93.7417
R35606 vdd.n762 vdd.n733 93.7417
R35607 vdd.n771 vdd.n762 93.7417
R35608 vdd.n777 vdd.n731 93.7417
R35609 vdd.n760 vdd.n731 93.7417
R35610 vdd.n752 vdd.n751 93.7417
R35611 vdd.n751 vdd.n741 93.7417
R35612 vdd.n864 vdd.n835 93.7417
R35613 vdd.n873 vdd.n864 93.7417
R35614 vdd.n879 vdd.n833 93.7417
R35615 vdd.n862 vdd.n833 93.7417
R35616 vdd.n854 vdd.n853 93.7417
R35617 vdd.n853 vdd.n843 93.7417
R35618 vdd.n912 vdd.n883 93.7417
R35619 vdd.n921 vdd.n912 93.7417
R35620 vdd.n927 vdd.n881 93.7417
R35621 vdd.n910 vdd.n881 93.7417
R35622 vdd.n902 vdd.n901 93.7417
R35623 vdd.n901 vdd.n891 93.7417
R35624 vdd.n960 vdd.n931 93.7417
R35625 vdd.n969 vdd.n960 93.7417
R35626 vdd.n975 vdd.n929 93.7417
R35627 vdd.n958 vdd.n929 93.7417
R35628 vdd.n950 vdd.n949 93.7417
R35629 vdd.n949 vdd.n939 93.7417
R35630 vdd.n1008 vdd.n979 93.7417
R35631 vdd.n1017 vdd.n1008 93.7417
R35632 vdd.n1023 vdd.n977 93.7417
R35633 vdd.n1006 vdd.n977 93.7417
R35634 vdd.n998 vdd.n997 93.7417
R35635 vdd.n997 vdd.n987 93.7417
R35636 vdd.n1110 vdd.n1081 93.7417
R35637 vdd.n1119 vdd.n1110 93.7417
R35638 vdd.n1125 vdd.n1079 93.7417
R35639 vdd.n1108 vdd.n1079 93.7417
R35640 vdd.n1100 vdd.n1099 93.7417
R35641 vdd.n1099 vdd.n1089 93.7417
R35642 vdd.n2630 vdd.n2601 93.7417
R35643 vdd.n2639 vdd.n2630 93.7417
R35644 vdd.n2645 vdd.n2599 93.7417
R35645 vdd.n2628 vdd.n2599 93.7417
R35646 vdd.n2620 vdd.n2619 93.7417
R35647 vdd.n2619 vdd.n2609 93.7417
R35648 vdd.n1167 vdd.n1158 93.7417
R35649 vdd.n1158 vdd.n1129 93.7417
R35650 vdd.n1156 vdd.n1127 93.7417
R35651 vdd.n1173 vdd.n1127 93.7417
R35652 vdd.n1142 vdd.n1137 93.7417
R35653 vdd.n1143 vdd.n1142 93.7417
R35654 vdd.n1215 vdd.n1206 93.7417
R35655 vdd.n1206 vdd.n1177 93.7417
R35656 vdd.n1204 vdd.n1175 93.7417
R35657 vdd.n1221 vdd.n1175 93.7417
R35658 vdd.n1190 vdd.n1185 93.7417
R35659 vdd.n1191 vdd.n1190 93.7417
R35660 vdd.n1316 vdd.n1307 93.7417
R35661 vdd.n1307 vdd.n1278 93.7417
R35662 vdd.n1305 vdd.n1276 93.7417
R35663 vdd.n1322 vdd.n1276 93.7417
R35664 vdd.n1291 vdd.n1286 93.7417
R35665 vdd.n1292 vdd.n1291 93.7417
R35666 vdd.n1364 vdd.n1355 93.7417
R35667 vdd.n1355 vdd.n1326 93.7417
R35668 vdd.n1353 vdd.n1324 93.7417
R35669 vdd.n1370 vdd.n1324 93.7417
R35670 vdd.n1339 vdd.n1334 93.7417
R35671 vdd.n1340 vdd.n1339 93.7417
R35672 vdd.n1412 vdd.n1403 93.7417
R35673 vdd.n1403 vdd.n1374 93.7417
R35674 vdd.n1401 vdd.n1372 93.7417
R35675 vdd.n1418 vdd.n1372 93.7417
R35676 vdd.n1387 vdd.n1382 93.7417
R35677 vdd.n1388 vdd.n1387 93.7417
R35678 vdd.n1460 vdd.n1451 93.7417
R35679 vdd.n1451 vdd.n1422 93.7417
R35680 vdd.n1449 vdd.n1420 93.7417
R35681 vdd.n1466 vdd.n1420 93.7417
R35682 vdd.n1435 vdd.n1430 93.7417
R35683 vdd.n1436 vdd.n1435 93.7417
R35684 vdd.n1561 vdd.n1552 93.7417
R35685 vdd.n1552 vdd.n1523 93.7417
R35686 vdd.n1550 vdd.n1521 93.7417
R35687 vdd.n1567 vdd.n1521 93.7417
R35688 vdd.n1536 vdd.n1531 93.7417
R35689 vdd.n1537 vdd.n1536 93.7417
R35690 vdd.n674 vdd.n665 93.7417
R35691 vdd.n665 vdd.n636 93.7417
R35692 vdd.n663 vdd.n634 93.7417
R35693 vdd.n680 vdd.n634 93.7417
R35694 vdd.n649 vdd.n644 93.7417
R35695 vdd.n650 vdd.n649 93.7417
R35696 vdd.n1609 vdd.n1600 93.7417
R35697 vdd.n1600 vdd.n1571 93.7417
R35698 vdd.n1598 vdd.n1569 93.7417
R35699 vdd.n1615 vdd.n1569 93.7417
R35700 vdd.n1584 vdd.n1579 93.7417
R35701 vdd.n1585 vdd.n1584 93.7417
R35702 vdd.n1656 vdd.n1647 93.7417
R35703 vdd.n1647 vdd.n1618 93.7417
R35704 vdd.n1645 vdd.n1616 93.7417
R35705 vdd.n1662 vdd.n1616 93.7417
R35706 vdd.n1631 vdd.n1626 93.7417
R35707 vdd.n1632 vdd.n1631 93.7417
R35708 vdd.n1706 vdd.n1697 93.7417
R35709 vdd.n1697 vdd.n1668 93.7417
R35710 vdd.n1695 vdd.n1666 93.7417
R35711 vdd.n1712 vdd.n1666 93.7417
R35712 vdd.n1681 vdd.n1676 93.7417
R35713 vdd.n1682 vdd.n1681 93.7417
R35714 vdd.n1756 vdd.n1747 93.7417
R35715 vdd.n1747 vdd.n1718 93.7417
R35716 vdd.n1745 vdd.n1716 93.7417
R35717 vdd.n1762 vdd.n1716 93.7417
R35718 vdd.n1731 vdd.n1726 93.7417
R35719 vdd.n1732 vdd.n1731 93.7417
R35720 vdd.n1804 vdd.n1795 93.7417
R35721 vdd.n1795 vdd.n1766 93.7417
R35722 vdd.n1793 vdd.n1764 93.7417
R35723 vdd.n1810 vdd.n1764 93.7417
R35724 vdd.n1779 vdd.n1774 93.7417
R35725 vdd.n1780 vdd.n1779 93.7417
R35726 vdd.n1496 vdd.n1486 93.7417
R35727 vdd.n1489 vdd.n1486 93.7417
R35728 vdd.n1503 vdd.n1478 93.7417
R35729 vdd.n1504 vdd.n1503 93.7417
R35730 vdd.n1510 vdd.n1477 93.7417
R35731 vdd.n1477 vdd.n1471 93.7417
R35732 vdd.n1855 vdd.n1846 93.7417
R35733 vdd.n1846 vdd.n1817 93.7417
R35734 vdd.n1844 vdd.n1815 93.7417
R35735 vdd.n1861 vdd.n1815 93.7417
R35736 vdd.n1830 vdd.n1825 93.7417
R35737 vdd.n1831 vdd.n1830 93.7417
R35738 vdd.n1902 vdd.n1893 93.7417
R35739 vdd.n1893 vdd.n1864 93.7417
R35740 vdd.n1891 vdd.n1862 93.7417
R35741 vdd.n1908 vdd.n1862 93.7417
R35742 vdd.n1877 vdd.n1872 93.7417
R35743 vdd.n1878 vdd.n1877 93.7417
R35744 vdd.n1950 vdd.n1941 93.7417
R35745 vdd.n1941 vdd.n1912 93.7417
R35746 vdd.n1939 vdd.n1910 93.7417
R35747 vdd.n1956 vdd.n1910 93.7417
R35748 vdd.n1925 vdd.n1920 93.7417
R35749 vdd.n1926 vdd.n1925 93.7417
R35750 vdd.n2001 vdd.n1992 93.7417
R35751 vdd.n1992 vdd.n1963 93.7417
R35752 vdd.n1990 vdd.n1961 93.7417
R35753 vdd.n2007 vdd.n1961 93.7417
R35754 vdd.n1976 vdd.n1971 93.7417
R35755 vdd.n1977 vdd.n1976 93.7417
R35756 vdd.n2051 vdd.n2042 93.7417
R35757 vdd.n2042 vdd.n2013 93.7417
R35758 vdd.n2040 vdd.n2011 93.7417
R35759 vdd.n2057 vdd.n2011 93.7417
R35760 vdd.n2026 vdd.n2021 93.7417
R35761 vdd.n2027 vdd.n2026 93.7417
R35762 vdd.n2099 vdd.n2090 93.7417
R35763 vdd.n2090 vdd.n2061 93.7417
R35764 vdd.n2088 vdd.n2059 93.7417
R35765 vdd.n2105 vdd.n2059 93.7417
R35766 vdd.n2074 vdd.n2069 93.7417
R35767 vdd.n2075 vdd.n2074 93.7417
R35768 vdd.n2149 vdd.n2140 93.7417
R35769 vdd.n2140 vdd.n2111 93.7417
R35770 vdd.n2138 vdd.n2109 93.7417
R35771 vdd.n2155 vdd.n2109 93.7417
R35772 vdd.n2124 vdd.n2119 93.7417
R35773 vdd.n2125 vdd.n2124 93.7417
R35774 vdd.n2196 vdd.n2187 93.7417
R35775 vdd.n2187 vdd.n2158 93.7417
R35776 vdd.n2185 vdd.n2156 93.7417
R35777 vdd.n2202 vdd.n2156 93.7417
R35778 vdd.n2171 vdd.n2166 93.7417
R35779 vdd.n2172 vdd.n2171 93.7417
R35780 vdd.n2246 vdd.n2237 93.7417
R35781 vdd.n2237 vdd.n2208 93.7417
R35782 vdd.n2235 vdd.n2206 93.7417
R35783 vdd.n2252 vdd.n2206 93.7417
R35784 vdd.n2221 vdd.n2216 93.7417
R35785 vdd.n2222 vdd.n2221 93.7417
R35786 vdd.n2296 vdd.n2287 93.7417
R35787 vdd.n2287 vdd.n2258 93.7417
R35788 vdd.n2285 vdd.n2256 93.7417
R35789 vdd.n2302 vdd.n2256 93.7417
R35790 vdd.n2271 vdd.n2266 93.7417
R35791 vdd.n2272 vdd.n2271 93.7417
R35792 vdd.n2344 vdd.n2335 93.7417
R35793 vdd.n2335 vdd.n2306 93.7417
R35794 vdd.n2333 vdd.n2304 93.7417
R35795 vdd.n2350 vdd.n2304 93.7417
R35796 vdd.n2319 vdd.n2314 93.7417
R35797 vdd.n2320 vdd.n2319 93.7417
R35798 vdd.n1251 vdd.n1241 93.7417
R35799 vdd.n1244 vdd.n1241 93.7417
R35800 vdd.n1258 vdd.n1233 93.7417
R35801 vdd.n1259 vdd.n1258 93.7417
R35802 vdd.n1265 vdd.n1232 93.7417
R35803 vdd.n1232 vdd.n1226 93.7417
R35804 vdd.n2395 vdd.n2386 93.7417
R35805 vdd.n2386 vdd.n2357 93.7417
R35806 vdd.n2384 vdd.n2355 93.7417
R35807 vdd.n2401 vdd.n2355 93.7417
R35808 vdd.n2370 vdd.n2365 93.7417
R35809 vdd.n2371 vdd.n2370 93.7417
R35810 vdd.n2442 vdd.n2433 93.7417
R35811 vdd.n2433 vdd.n2404 93.7417
R35812 vdd.n2431 vdd.n2402 93.7417
R35813 vdd.n2448 vdd.n2402 93.7417
R35814 vdd.n2417 vdd.n2412 93.7417
R35815 vdd.n2418 vdd.n2417 93.7417
R35816 vdd.n2492 vdd.n2483 93.7417
R35817 vdd.n2483 vdd.n2454 93.7417
R35818 vdd.n2481 vdd.n2452 93.7417
R35819 vdd.n2498 vdd.n2452 93.7417
R35820 vdd.n2467 vdd.n2462 93.7417
R35821 vdd.n2468 vdd.n2467 93.7417
R35822 vdd.n2542 vdd.n2533 93.7417
R35823 vdd.n2533 vdd.n2504 93.7417
R35824 vdd.n2531 vdd.n2502 93.7417
R35825 vdd.n2548 vdd.n2502 93.7417
R35826 vdd.n2517 vdd.n2512 93.7417
R35827 vdd.n2518 vdd.n2517 93.7417
R35828 vdd.n2590 vdd.n2581 93.7417
R35829 vdd.n2581 vdd.n2552 93.7417
R35830 vdd.n2579 vdd.n2550 93.7417
R35831 vdd.n2596 vdd.n2550 93.7417
R35832 vdd.n2565 vdd.n2560 93.7417
R35833 vdd.n2566 vdd.n2565 93.7417
R35834 vdd.n2727 vdd.n2698 93.7417
R35835 vdd.n2736 vdd.n2727 93.7417
R35836 vdd.n2742 vdd.n2696 93.7417
R35837 vdd.n2725 vdd.n2696 93.7417
R35838 vdd.n2717 vdd.n2716 93.7417
R35839 vdd.n2716 vdd.n2706 93.7417
R35840 vdd.n2679 vdd.n2650 93.7417
R35841 vdd.n2688 vdd.n2679 93.7417
R35842 vdd.n2694 vdd.n2648 93.7417
R35843 vdd.n2677 vdd.n2648 93.7417
R35844 vdd.n2669 vdd.n2668 93.7417
R35845 vdd.n2668 vdd.n2658 93.7417
R35846 vdd.n2776 vdd.n2747 93.7417
R35847 vdd.n2785 vdd.n2776 93.7417
R35848 vdd.n2791 vdd.n2745 93.7417
R35849 vdd.n2774 vdd.n2745 93.7417
R35850 vdd.n2766 vdd.n2765 93.7417
R35851 vdd.n2765 vdd.n2755 93.7417
R35852 vdd.n2826 vdd.n2797 93.7417
R35853 vdd.n2835 vdd.n2826 93.7417
R35854 vdd.n2841 vdd.n2795 93.7417
R35855 vdd.n2824 vdd.n2795 93.7417
R35856 vdd.n2816 vdd.n2815 93.7417
R35857 vdd.n2815 vdd.n2805 93.7417
R35858 vdd.n2874 vdd.n2845 93.7417
R35859 vdd.n2883 vdd.n2874 93.7417
R35860 vdd.n2889 vdd.n2843 93.7417
R35861 vdd.n2872 vdd.n2843 93.7417
R35862 vdd.n2864 vdd.n2863 93.7417
R35863 vdd.n2863 vdd.n2853 93.7417
R35864 vdd.n1065 vdd.n1064 93.7417
R35865 vdd.n1065 vdd.n1029 93.7417
R35866 vdd.n1062 vdd.n1061 93.7417
R35867 vdd.n1061 vdd.n1033 93.7417
R35868 vdd.n1052 vdd.n1039 93.7417
R35869 vdd.n1045 vdd.n1039 93.7417
R35870 vdd.n3022 vdd.n2993 93.7417
R35871 vdd.n3031 vdd.n3022 93.7417
R35872 vdd.n3037 vdd.n2991 93.7417
R35873 vdd.n3020 vdd.n2991 93.7417
R35874 vdd.n3012 vdd.n3011 93.7417
R35875 vdd.n3011 vdd.n3001 93.7417
R35876 vdd.n2973 vdd.n2944 93.7417
R35877 vdd.n2982 vdd.n2973 93.7417
R35878 vdd.n2988 vdd.n2942 93.7417
R35879 vdd.n2971 vdd.n2942 93.7417
R35880 vdd.n2963 vdd.n2962 93.7417
R35881 vdd.n2962 vdd.n2952 93.7417
R35882 vdd.n2925 vdd.n2896 93.7417
R35883 vdd.n2934 vdd.n2925 93.7417
R35884 vdd.n2940 vdd.n2894 93.7417
R35885 vdd.n2923 vdd.n2894 93.7417
R35886 vdd.n2915 vdd.n2914 93.7417
R35887 vdd.n2914 vdd.n2904 93.7417
R35888 vdd.n3071 vdd.n3042 93.7417
R35889 vdd.n3080 vdd.n3071 93.7417
R35890 vdd.n3086 vdd.n3040 93.7417
R35891 vdd.n3069 vdd.n3040 93.7417
R35892 vdd.n3061 vdd.n3060 93.7417
R35893 vdd.n3060 vdd.n3050 93.7417
R35894 vdd.n3121 vdd.n3092 93.7417
R35895 vdd.n3130 vdd.n3121 93.7417
R35896 vdd.n3136 vdd.n3090 93.7417
R35897 vdd.n3119 vdd.n3090 93.7417
R35898 vdd.n3111 vdd.n3110 93.7417
R35899 vdd.n3110 vdd.n3100 93.7417
R35900 vdd.n3169 vdd.n3140 93.7417
R35901 vdd.n3178 vdd.n3169 93.7417
R35902 vdd.n3184 vdd.n3138 93.7417
R35903 vdd.n3167 vdd.n3138 93.7417
R35904 vdd.n3159 vdd.n3158 93.7417
R35905 vdd.n3158 vdd.n3148 93.7417
R35906 vdd.n3267 vdd.n3238 93.7417
R35907 vdd.n3276 vdd.n3267 93.7417
R35908 vdd.n3282 vdd.n3236 93.7417
R35909 vdd.n3265 vdd.n3236 93.7417
R35910 vdd.n3257 vdd.n3256 93.7417
R35911 vdd.n3256 vdd.n3246 93.7417
R35912 vdd.n3219 vdd.n3190 93.7417
R35913 vdd.n3228 vdd.n3219 93.7417
R35914 vdd.n3234 vdd.n3188 93.7417
R35915 vdd.n3217 vdd.n3188 93.7417
R35916 vdd.n3209 vdd.n3208 93.7417
R35917 vdd.n3208 vdd.n3198 93.7417
R35918 vdd.n3316 vdd.n3287 93.7417
R35919 vdd.n3325 vdd.n3316 93.7417
R35920 vdd.n3331 vdd.n3285 93.7417
R35921 vdd.n3314 vdd.n3285 93.7417
R35922 vdd.n3306 vdd.n3305 93.7417
R35923 vdd.n3305 vdd.n3295 93.7417
R35924 vdd.n3366 vdd.n3337 93.7417
R35925 vdd.n3375 vdd.n3366 93.7417
R35926 vdd.n3381 vdd.n3335 93.7417
R35927 vdd.n3364 vdd.n3335 93.7417
R35928 vdd.n3356 vdd.n3355 93.7417
R35929 vdd.n3355 vdd.n3345 93.7417
R35930 vdd.n3414 vdd.n3385 93.7417
R35931 vdd.n3423 vdd.n3414 93.7417
R35932 vdd.n3429 vdd.n3383 93.7417
R35933 vdd.n3412 vdd.n3383 93.7417
R35934 vdd.n3404 vdd.n3403 93.7417
R35935 vdd.n3403 vdd.n3393 93.7417
R35936 vdd.n819 vdd.n818 93.7417
R35937 vdd.n819 vdd.n783 93.7417
R35938 vdd.n816 vdd.n815 93.7417
R35939 vdd.n815 vdd.n787 93.7417
R35940 vdd.n806 vdd.n793 93.7417
R35941 vdd.n799 vdd.n793 93.7417
R35942 vdd.n3513 vdd.n3484 93.7417
R35943 vdd.n3522 vdd.n3513 93.7417
R35944 vdd.n3528 vdd.n3482 93.7417
R35945 vdd.n3511 vdd.n3482 93.7417
R35946 vdd.n3503 vdd.n3502 93.7417
R35947 vdd.n3502 vdd.n3492 93.7417
R35948 vdd.n3465 vdd.n3436 93.7417
R35949 vdd.n3474 vdd.n3465 93.7417
R35950 vdd.n3480 vdd.n3434 93.7417
R35951 vdd.n3463 vdd.n3434 93.7417
R35952 vdd.n3455 vdd.n3454 93.7417
R35953 vdd.n3454 vdd.n3444 93.7417
R35954 vdd.n3562 vdd.n3533 93.7417
R35955 vdd.n3571 vdd.n3562 93.7417
R35956 vdd.n3577 vdd.n3531 93.7417
R35957 vdd.n3560 vdd.n3531 93.7417
R35958 vdd.n3552 vdd.n3551 93.7417
R35959 vdd.n3551 vdd.n3541 93.7417
R35960 vdd.n3612 vdd.n3583 93.7417
R35961 vdd.n3621 vdd.n3612 93.7417
R35962 vdd.n3627 vdd.n3581 93.7417
R35963 vdd.n3610 vdd.n3581 93.7417
R35964 vdd.n3602 vdd.n3601 93.7417
R35965 vdd.n3601 vdd.n3591 93.7417
R35966 vdd.n3660 vdd.n3631 93.7417
R35967 vdd.n3669 vdd.n3660 93.7417
R35968 vdd.n3675 vdd.n3629 93.7417
R35969 vdd.n3658 vdd.n3629 93.7417
R35970 vdd.n3650 vdd.n3649 93.7417
R35971 vdd.n3649 vdd.n3639 93.7417
R35972 vdd.n618 vdd.n589 93.7417
R35973 vdd.n627 vdd.n618 93.7417
R35974 vdd.n633 vdd.n587 93.7417
R35975 vdd.n616 vdd.n587 93.7417
R35976 vdd.n608 vdd.n607 93.7417
R35977 vdd.n607 vdd.n597 93.7417
R35978 vdd.n3759 vdd.n3730 93.7417
R35979 vdd.n3768 vdd.n3759 93.7417
R35980 vdd.n3774 vdd.n3728 93.7417
R35981 vdd.n3757 vdd.n3728 93.7417
R35982 vdd.n3749 vdd.n3748 93.7417
R35983 vdd.n3748 vdd.n3738 93.7417
R35984 vdd.n3711 vdd.n3682 93.7417
R35985 vdd.n3720 vdd.n3711 93.7417
R35986 vdd.n3726 vdd.n3680 93.7417
R35987 vdd.n3709 vdd.n3680 93.7417
R35988 vdd.n3701 vdd.n3700 93.7417
R35989 vdd.n3700 vdd.n3690 93.7417
R35990 vdd.n6901 vdd.n6872 93.7417
R35991 vdd.n6910 vdd.n6901 93.7417
R35992 vdd.n6916 vdd.n6870 93.7417
R35993 vdd.n6899 vdd.n6870 93.7417
R35994 vdd.n6891 vdd.n6890 93.7417
R35995 vdd.n6890 vdd.n6880 93.7417
R35996 vdd.n6853 vdd.n6824 93.7417
R35997 vdd.n6862 vdd.n6853 93.7417
R35998 vdd.n6868 vdd.n6822 93.7417
R35999 vdd.n6851 vdd.n6822 93.7417
R36000 vdd.n6843 vdd.n6842 93.7417
R36001 vdd.n6842 vdd.n6832 93.7417
R36002 vdd.n10043 vdd.n10014 93.7417
R36003 vdd.n10052 vdd.n10043 93.7417
R36004 vdd.n10058 vdd.n10012 93.7417
R36005 vdd.n10041 vdd.n10012 93.7417
R36006 vdd.n10033 vdd.n10032 93.7417
R36007 vdd.n10032 vdd.n10022 93.7417
R36008 vdd.n9995 vdd.n9966 93.7417
R36009 vdd.n10004 vdd.n9995 93.7417
R36010 vdd.n10010 vdd.n9964 93.7417
R36011 vdd.n9993 vdd.n9964 93.7417
R36012 vdd.n9985 vdd.n9984 93.7417
R36013 vdd.n9984 vdd.n9974 93.7417
R36014 vdd.n10091 vdd.n10062 93.7417
R36015 vdd.n10100 vdd.n10091 93.7417
R36016 vdd.n10106 vdd.n10060 93.7417
R36017 vdd.n10089 vdd.n10060 93.7417
R36018 vdd.n10081 vdd.n10080 93.7417
R36019 vdd.n10080 vdd.n10070 93.7417
R36020 vdd.n10139 vdd.n10110 93.7417
R36021 vdd.n10148 vdd.n10139 93.7417
R36022 vdd.n10154 vdd.n10108 93.7417
R36023 vdd.n10137 vdd.n10108 93.7417
R36024 vdd.n10129 vdd.n10128 93.7417
R36025 vdd.n10128 vdd.n10118 93.7417
R36026 vdd.n10241 vdd.n10212 93.7417
R36027 vdd.n10250 vdd.n10241 93.7417
R36028 vdd.n10256 vdd.n10210 93.7417
R36029 vdd.n10239 vdd.n10210 93.7417
R36030 vdd.n10231 vdd.n10230 93.7417
R36031 vdd.n10230 vdd.n10220 93.7417
R36032 vdd.n10289 vdd.n10260 93.7417
R36033 vdd.n10298 vdd.n10289 93.7417
R36034 vdd.n10304 vdd.n10258 93.7417
R36035 vdd.n10287 vdd.n10258 93.7417
R36036 vdd.n10279 vdd.n10278 93.7417
R36037 vdd.n10278 vdd.n10268 93.7417
R36038 vdd.n10337 vdd.n10308 93.7417
R36039 vdd.n10346 vdd.n10337 93.7417
R36040 vdd.n10352 vdd.n10306 93.7417
R36041 vdd.n10335 vdd.n10306 93.7417
R36042 vdd.n10327 vdd.n10326 93.7417
R36043 vdd.n10326 vdd.n10316 93.7417
R36044 vdd.n10385 vdd.n10356 93.7417
R36045 vdd.n10394 vdd.n10385 93.7417
R36046 vdd.n10400 vdd.n10354 93.7417
R36047 vdd.n10383 vdd.n10354 93.7417
R36048 vdd.n10375 vdd.n10374 93.7417
R36049 vdd.n10374 vdd.n10364 93.7417
R36050 vdd.n10487 vdd.n10458 93.7417
R36051 vdd.n10496 vdd.n10487 93.7417
R36052 vdd.n10502 vdd.n10456 93.7417
R36053 vdd.n10485 vdd.n10456 93.7417
R36054 vdd.n10477 vdd.n10476 93.7417
R36055 vdd.n10476 vdd.n10466 93.7417
R36056 vdd.n79 vdd.n50 93.7417
R36057 vdd.n88 vdd.n79 93.7417
R36058 vdd.n94 vdd.n48 93.7417
R36059 vdd.n77 vdd.n48 93.7417
R36060 vdd.n69 vdd.n68 93.7417
R36061 vdd.n68 vdd.n58 93.7417
R36062 vdd.n31 vdd.n2 93.7417
R36063 vdd.n40 vdd.n31 93.7417
R36064 vdd.n46 vdd.n0 93.7417
R36065 vdd.n29 vdd.n0 93.7417
R36066 vdd.n21 vdd.n20 93.7417
R36067 vdd.n20 vdd.n10 93.7417
R36068 vdd.n10535 vdd.n10506 93.7417
R36069 vdd.n10544 vdd.n10535 93.7417
R36070 vdd.n10550 vdd.n10504 93.7417
R36071 vdd.n10533 vdd.n10504 93.7417
R36072 vdd.n10525 vdd.n10524 93.7417
R36073 vdd.n10524 vdd.n10514 93.7417
R36074 vdd.n10585 vdd.n10556 93.7417
R36075 vdd.n10594 vdd.n10585 93.7417
R36076 vdd.n10600 vdd.n10554 93.7417
R36077 vdd.n10583 vdd.n10554 93.7417
R36078 vdd.n10575 vdd.n10574 93.7417
R36079 vdd.n10574 vdd.n10564 93.7417
R36080 vdd.n10633 vdd.n10604 93.7417
R36081 vdd.n10642 vdd.n10633 93.7417
R36082 vdd.n10648 vdd.n10602 93.7417
R36083 vdd.n10631 vdd.n10602 93.7417
R36084 vdd.n10623 vdd.n10622 93.7417
R36085 vdd.n10622 vdd.n10612 93.7417
R36086 vdd.n10442 vdd.n10441 93.7417
R36087 vdd.n10442 vdd.n10406 93.7417
R36088 vdd.n10439 vdd.n10438 93.7417
R36089 vdd.n10438 vdd.n10410 93.7417
R36090 vdd.n10429 vdd.n10416 93.7417
R36091 vdd.n10422 vdd.n10416 93.7417
R36092 vdd.n10781 vdd.n10752 93.7417
R36093 vdd.n10790 vdd.n10781 93.7417
R36094 vdd.n10796 vdd.n10750 93.7417
R36095 vdd.n10779 vdd.n10750 93.7417
R36096 vdd.n10771 vdd.n10770 93.7417
R36097 vdd.n10770 vdd.n10760 93.7417
R36098 vdd.n10732 vdd.n10703 93.7417
R36099 vdd.n10741 vdd.n10732 93.7417
R36100 vdd.n10747 vdd.n10701 93.7417
R36101 vdd.n10730 vdd.n10701 93.7417
R36102 vdd.n10722 vdd.n10721 93.7417
R36103 vdd.n10721 vdd.n10711 93.7417
R36104 vdd.n10684 vdd.n10655 93.7417
R36105 vdd.n10693 vdd.n10684 93.7417
R36106 vdd.n10699 vdd.n10653 93.7417
R36107 vdd.n10682 vdd.n10653 93.7417
R36108 vdd.n10674 vdd.n10673 93.7417
R36109 vdd.n10673 vdd.n10663 93.7417
R36110 vdd.n10830 vdd.n10801 93.7417
R36111 vdd.n10839 vdd.n10830 93.7417
R36112 vdd.n10845 vdd.n10799 93.7417
R36113 vdd.n10828 vdd.n10799 93.7417
R36114 vdd.n10820 vdd.n10819 93.7417
R36115 vdd.n10819 vdd.n10809 93.7417
R36116 vdd.n10880 vdd.n10851 93.7417
R36117 vdd.n10889 vdd.n10880 93.7417
R36118 vdd.n10895 vdd.n10849 93.7417
R36119 vdd.n10878 vdd.n10849 93.7417
R36120 vdd.n10870 vdd.n10869 93.7417
R36121 vdd.n10869 vdd.n10859 93.7417
R36122 vdd.n10928 vdd.n10899 93.7417
R36123 vdd.n10937 vdd.n10928 93.7417
R36124 vdd.n10943 vdd.n10897 93.7417
R36125 vdd.n10926 vdd.n10897 93.7417
R36126 vdd.n10918 vdd.n10917 93.7417
R36127 vdd.n10917 vdd.n10907 93.7417
R36128 vdd.n11026 vdd.n10997 93.7417
R36129 vdd.n11035 vdd.n11026 93.7417
R36130 vdd.n11041 vdd.n10995 93.7417
R36131 vdd.n11024 vdd.n10995 93.7417
R36132 vdd.n11016 vdd.n11015 93.7417
R36133 vdd.n11015 vdd.n11005 93.7417
R36134 vdd.n10978 vdd.n10949 93.7417
R36135 vdd.n10987 vdd.n10978 93.7417
R36136 vdd.n10993 vdd.n10947 93.7417
R36137 vdd.n10976 vdd.n10947 93.7417
R36138 vdd.n10968 vdd.n10967 93.7417
R36139 vdd.n10967 vdd.n10957 93.7417
R36140 vdd.n11075 vdd.n11046 93.7417
R36141 vdd.n11084 vdd.n11075 93.7417
R36142 vdd.n11090 vdd.n11044 93.7417
R36143 vdd.n11073 vdd.n11044 93.7417
R36144 vdd.n11065 vdd.n11064 93.7417
R36145 vdd.n11064 vdd.n11054 93.7417
R36146 vdd.n11125 vdd.n11096 93.7417
R36147 vdd.n11134 vdd.n11125 93.7417
R36148 vdd.n11140 vdd.n11094 93.7417
R36149 vdd.n11123 vdd.n11094 93.7417
R36150 vdd.n11115 vdd.n11114 93.7417
R36151 vdd.n11114 vdd.n11104 93.7417
R36152 vdd.n11173 vdd.n11144 93.7417
R36153 vdd.n11182 vdd.n11173 93.7417
R36154 vdd.n11188 vdd.n11142 93.7417
R36155 vdd.n11171 vdd.n11142 93.7417
R36156 vdd.n11163 vdd.n11162 93.7417
R36157 vdd.n11162 vdd.n11152 93.7417
R36158 vdd.n10196 vdd.n10195 93.7417
R36159 vdd.n10196 vdd.n10160 93.7417
R36160 vdd.n10193 vdd.n10192 93.7417
R36161 vdd.n10192 vdd.n10164 93.7417
R36162 vdd.n10183 vdd.n10170 93.7417
R36163 vdd.n10176 vdd.n10170 93.7417
R36164 vdd.n11272 vdd.n11243 93.7417
R36165 vdd.n11281 vdd.n11272 93.7417
R36166 vdd.n11287 vdd.n11241 93.7417
R36167 vdd.n11270 vdd.n11241 93.7417
R36168 vdd.n11262 vdd.n11261 93.7417
R36169 vdd.n11261 vdd.n11251 93.7417
R36170 vdd.n11224 vdd.n11195 93.7417
R36171 vdd.n11233 vdd.n11224 93.7417
R36172 vdd.n11239 vdd.n11193 93.7417
R36173 vdd.n11222 vdd.n11193 93.7417
R36174 vdd.n11214 vdd.n11213 93.7417
R36175 vdd.n11213 vdd.n11203 93.7417
R36176 vdd.n11321 vdd.n11292 93.7417
R36177 vdd.n11330 vdd.n11321 93.7417
R36178 vdd.n11336 vdd.n11290 93.7417
R36179 vdd.n11319 vdd.n11290 93.7417
R36180 vdd.n11311 vdd.n11310 93.7417
R36181 vdd.n11310 vdd.n11300 93.7417
R36182 vdd.n11371 vdd.n11342 93.7417
R36183 vdd.n11380 vdd.n11371 93.7417
R36184 vdd.n11386 vdd.n11340 93.7417
R36185 vdd.n11369 vdd.n11340 93.7417
R36186 vdd.n11361 vdd.n11360 93.7417
R36187 vdd.n11360 vdd.n11350 93.7417
R36188 vdd.n11419 vdd.n11390 93.7417
R36189 vdd.n11428 vdd.n11419 93.7417
R36190 vdd.n11434 vdd.n11388 93.7417
R36191 vdd.n11417 vdd.n11388 93.7417
R36192 vdd.n11409 vdd.n11408 93.7417
R36193 vdd.n11408 vdd.n11398 93.7417
R36194 vdd.n11479 vdd.n11470 93.7417
R36195 vdd.n11470 vdd.n11441 93.7417
R36196 vdd.n11468 vdd.n11439 93.7417
R36197 vdd.n11485 vdd.n11439 93.7417
R36198 vdd.n11454 vdd.n11449 93.7417
R36199 vdd.n11455 vdd.n11454 93.7417
R36200 vdd.n11526 vdd.n11517 93.7417
R36201 vdd.n11517 vdd.n11488 93.7417
R36202 vdd.n11515 vdd.n11486 93.7417
R36203 vdd.n11532 vdd.n11486 93.7417
R36204 vdd.n11501 vdd.n11496 93.7417
R36205 vdd.n11502 vdd.n11501 93.7417
R36206 vdd.n11576 vdd.n11567 93.7417
R36207 vdd.n11567 vdd.n11538 93.7417
R36208 vdd.n11565 vdd.n11536 93.7417
R36209 vdd.n11582 vdd.n11536 93.7417
R36210 vdd.n11551 vdd.n11546 93.7417
R36211 vdd.n11552 vdd.n11551 93.7417
R36212 vdd.n11626 vdd.n11617 93.7417
R36213 vdd.n11617 vdd.n11588 93.7417
R36214 vdd.n11615 vdd.n11586 93.7417
R36215 vdd.n11632 vdd.n11586 93.7417
R36216 vdd.n11601 vdd.n11596 93.7417
R36217 vdd.n11602 vdd.n11601 93.7417
R36218 vdd.n11674 vdd.n11665 93.7417
R36219 vdd.n11665 vdd.n11636 93.7417
R36220 vdd.n11663 vdd.n11634 93.7417
R36221 vdd.n11680 vdd.n11634 93.7417
R36222 vdd.n11649 vdd.n11644 93.7417
R36223 vdd.n11650 vdd.n11649 93.7417
R36224 vdd.n466 vdd.n456 93.7417
R36225 vdd.n459 vdd.n456 93.7417
R36226 vdd.n473 vdd.n448 93.7417
R36227 vdd.n474 vdd.n473 93.7417
R36228 vdd.n480 vdd.n447 93.7417
R36229 vdd.n447 vdd.n441 93.7417
R36230 vdd.n11725 vdd.n11716 93.7417
R36231 vdd.n11716 vdd.n11687 93.7417
R36232 vdd.n11714 vdd.n11685 93.7417
R36233 vdd.n11731 vdd.n11685 93.7417
R36234 vdd.n11700 vdd.n11695 93.7417
R36235 vdd.n11701 vdd.n11700 93.7417
R36236 vdd.n11772 vdd.n11763 93.7417
R36237 vdd.n11763 vdd.n11734 93.7417
R36238 vdd.n11761 vdd.n11732 93.7417
R36239 vdd.n11778 vdd.n11732 93.7417
R36240 vdd.n11747 vdd.n11742 93.7417
R36241 vdd.n11748 vdd.n11747 93.7417
R36242 vdd.n11820 vdd.n11811 93.7417
R36243 vdd.n11811 vdd.n11782 93.7417
R36244 vdd.n11809 vdd.n11780 93.7417
R36245 vdd.n11826 vdd.n11780 93.7417
R36246 vdd.n11795 vdd.n11790 93.7417
R36247 vdd.n11796 vdd.n11795 93.7417
R36248 vdd.n11871 vdd.n11862 93.7417
R36249 vdd.n11862 vdd.n11833 93.7417
R36250 vdd.n11860 vdd.n11831 93.7417
R36251 vdd.n11877 vdd.n11831 93.7417
R36252 vdd.n11846 vdd.n11841 93.7417
R36253 vdd.n11847 vdd.n11846 93.7417
R36254 vdd.n11921 vdd.n11912 93.7417
R36255 vdd.n11912 vdd.n11883 93.7417
R36256 vdd.n11910 vdd.n11881 93.7417
R36257 vdd.n11927 vdd.n11881 93.7417
R36258 vdd.n11896 vdd.n11891 93.7417
R36259 vdd.n11897 vdd.n11896 93.7417
R36260 vdd.n11969 vdd.n11960 93.7417
R36261 vdd.n11960 vdd.n11931 93.7417
R36262 vdd.n11958 vdd.n11929 93.7417
R36263 vdd.n11975 vdd.n11929 93.7417
R36264 vdd.n11944 vdd.n11939 93.7417
R36265 vdd.n11945 vdd.n11944 93.7417
R36266 vdd.n12019 vdd.n12010 93.7417
R36267 vdd.n12010 vdd.n11981 93.7417
R36268 vdd.n12008 vdd.n11979 93.7417
R36269 vdd.n12025 vdd.n11979 93.7417
R36270 vdd.n11994 vdd.n11989 93.7417
R36271 vdd.n11995 vdd.n11994 93.7417
R36272 vdd.n12066 vdd.n12057 93.7417
R36273 vdd.n12057 vdd.n12028 93.7417
R36274 vdd.n12055 vdd.n12026 93.7417
R36275 vdd.n12072 vdd.n12026 93.7417
R36276 vdd.n12041 vdd.n12036 93.7417
R36277 vdd.n12042 vdd.n12041 93.7417
R36278 vdd.n12116 vdd.n12107 93.7417
R36279 vdd.n12107 vdd.n12078 93.7417
R36280 vdd.n12105 vdd.n12076 93.7417
R36281 vdd.n12122 vdd.n12076 93.7417
R36282 vdd.n12091 vdd.n12086 93.7417
R36283 vdd.n12092 vdd.n12091 93.7417
R36284 vdd.n12166 vdd.n12157 93.7417
R36285 vdd.n12157 vdd.n12128 93.7417
R36286 vdd.n12155 vdd.n12126 93.7417
R36287 vdd.n12172 vdd.n12126 93.7417
R36288 vdd.n12141 vdd.n12136 93.7417
R36289 vdd.n12142 vdd.n12141 93.7417
R36290 vdd.n12214 vdd.n12205 93.7417
R36291 vdd.n12205 vdd.n12176 93.7417
R36292 vdd.n12203 vdd.n12174 93.7417
R36293 vdd.n12220 vdd.n12174 93.7417
R36294 vdd.n12189 vdd.n12184 93.7417
R36295 vdd.n12190 vdd.n12189 93.7417
R36296 vdd.n221 vdd.n211 93.7417
R36297 vdd.n214 vdd.n211 93.7417
R36298 vdd.n228 vdd.n203 93.7417
R36299 vdd.n229 vdd.n228 93.7417
R36300 vdd.n235 vdd.n202 93.7417
R36301 vdd.n202 vdd.n196 93.7417
R36302 vdd.n12265 vdd.n12256 93.7417
R36303 vdd.n12256 vdd.n12227 93.7417
R36304 vdd.n12254 vdd.n12225 93.7417
R36305 vdd.n12271 vdd.n12225 93.7417
R36306 vdd.n12240 vdd.n12235 93.7417
R36307 vdd.n12241 vdd.n12240 93.7417
R36308 vdd.n12312 vdd.n12303 93.7417
R36309 vdd.n12303 vdd.n12274 93.7417
R36310 vdd.n12301 vdd.n12272 93.7417
R36311 vdd.n12318 vdd.n12272 93.7417
R36312 vdd.n12287 vdd.n12282 93.7417
R36313 vdd.n12288 vdd.n12287 93.7417
R36314 vdd.n12362 vdd.n12353 93.7417
R36315 vdd.n12353 vdd.n12324 93.7417
R36316 vdd.n12351 vdd.n12322 93.7417
R36317 vdd.n12368 vdd.n12322 93.7417
R36318 vdd.n12337 vdd.n12332 93.7417
R36319 vdd.n12338 vdd.n12337 93.7417
R36320 vdd.n12412 vdd.n12403 93.7417
R36321 vdd.n12403 vdd.n12374 93.7417
R36322 vdd.n12401 vdd.n12372 93.7417
R36323 vdd.n12418 vdd.n12372 93.7417
R36324 vdd.n12387 vdd.n12382 93.7417
R36325 vdd.n12388 vdd.n12387 93.7417
R36326 vdd.n12460 vdd.n12451 93.7417
R36327 vdd.n12451 vdd.n12422 93.7417
R36328 vdd.n12449 vdd.n12420 93.7417
R36329 vdd.n12466 vdd.n12420 93.7417
R36330 vdd.n12435 vdd.n12430 93.7417
R36331 vdd.n12436 vdd.n12435 93.7417
R36332 vdd.n116 vdd.n115 84.1148
R36333 vdd.n136 vdd.n129 84.1148
R36334 vdd.n164 vdd.n163 84.1148
R36335 vdd.n184 vdd.n177 84.1148
R36336 vdd.n265 vdd.n264 84.1148
R36337 vdd.n285 vdd.n278 84.1148
R36338 vdd.n313 vdd.n312 84.1148
R36339 vdd.n333 vdd.n326 84.1148
R36340 vdd.n361 vdd.n360 84.1148
R36341 vdd.n381 vdd.n374 84.1148
R36342 vdd.n409 vdd.n408 84.1148
R36343 vdd.n429 vdd.n422 84.1148
R36344 vdd.n510 vdd.n509 84.1148
R36345 vdd.n530 vdd.n523 84.1148
R36346 vdd.n558 vdd.n557 84.1148
R36347 vdd.n578 vdd.n571 84.1148
R36348 vdd.n7006 vdd.n6999 84.1148
R36349 vdd.n6986 vdd.n6982 84.1148
R36350 vdd.n7054 vdd.n7047 84.1148
R36351 vdd.n7034 vdd.n7030 84.1148
R36352 vdd.n7156 vdd.n7149 84.1148
R36353 vdd.n7136 vdd.n7132 84.1148
R36354 vdd.n7204 vdd.n7197 84.1148
R36355 vdd.n7184 vdd.n7180 84.1148
R36356 vdd.n7252 vdd.n7245 84.1148
R36357 vdd.n7232 vdd.n7228 84.1148
R36358 vdd.n7300 vdd.n7293 84.1148
R36359 vdd.n7280 vdd.n7276 84.1148
R36360 vdd.n7402 vdd.n7395 84.1148
R36361 vdd.n7382 vdd.n7378 84.1148
R36362 vdd.n8922 vdd.n8915 84.1148
R36363 vdd.n8902 vdd.n8898 84.1148
R36364 vdd.n7430 vdd.n7429 84.1148
R36365 vdd.n7450 vdd.n7443 84.1148
R36366 vdd.n7478 vdd.n7477 84.1148
R36367 vdd.n7498 vdd.n7491 84.1148
R36368 vdd.n7579 vdd.n7578 84.1148
R36369 vdd.n7599 vdd.n7592 84.1148
R36370 vdd.n7627 vdd.n7626 84.1148
R36371 vdd.n7647 vdd.n7640 84.1148
R36372 vdd.n7675 vdd.n7674 84.1148
R36373 vdd.n7695 vdd.n7688 84.1148
R36374 vdd.n7723 vdd.n7722 84.1148
R36375 vdd.n7743 vdd.n7736 84.1148
R36376 vdd.n7824 vdd.n7823 84.1148
R36377 vdd.n7844 vdd.n7837 84.1148
R36378 vdd.n6937 vdd.n6936 84.1148
R36379 vdd.n6957 vdd.n6950 84.1148
R36380 vdd.n7872 vdd.n7871 84.1148
R36381 vdd.n7892 vdd.n7885 84.1148
R36382 vdd.n7919 vdd.n7918 84.1148
R36383 vdd.n7939 vdd.n7932 84.1148
R36384 vdd.n7969 vdd.n7968 84.1148
R36385 vdd.n7989 vdd.n7982 84.1148
R36386 vdd.n8019 vdd.n8018 84.1148
R36387 vdd.n8039 vdd.n8032 84.1148
R36388 vdd.n8067 vdd.n8066 84.1148
R36389 vdd.n8087 vdd.n8080 84.1148
R36390 vdd.n7795 vdd.n7754 84.1148
R36391 vdd.n7779 vdd.n7771 84.1148
R36392 vdd.n8118 vdd.n8117 84.1148
R36393 vdd.n8138 vdd.n8131 84.1148
R36394 vdd.n8165 vdd.n8164 84.1148
R36395 vdd.n8185 vdd.n8178 84.1148
R36396 vdd.n8213 vdd.n8212 84.1148
R36397 vdd.n8233 vdd.n8226 84.1148
R36398 vdd.n8264 vdd.n8263 84.1148
R36399 vdd.n8284 vdd.n8277 84.1148
R36400 vdd.n8314 vdd.n8313 84.1148
R36401 vdd.n8334 vdd.n8327 84.1148
R36402 vdd.n8362 vdd.n8361 84.1148
R36403 vdd.n8382 vdd.n8375 84.1148
R36404 vdd.n8412 vdd.n8411 84.1148
R36405 vdd.n8432 vdd.n8425 84.1148
R36406 vdd.n8459 vdd.n8458 84.1148
R36407 vdd.n8479 vdd.n8472 84.1148
R36408 vdd.n8509 vdd.n8508 84.1148
R36409 vdd.n8529 vdd.n8522 84.1148
R36410 vdd.n8559 vdd.n8558 84.1148
R36411 vdd.n8579 vdd.n8572 84.1148
R36412 vdd.n8607 vdd.n8606 84.1148
R36413 vdd.n8627 vdd.n8620 84.1148
R36414 vdd.n7550 vdd.n7509 84.1148
R36415 vdd.n7534 vdd.n7526 84.1148
R36416 vdd.n8658 vdd.n8657 84.1148
R36417 vdd.n8678 vdd.n8671 84.1148
R36418 vdd.n8705 vdd.n8704 84.1148
R36419 vdd.n8725 vdd.n8718 84.1148
R36420 vdd.n8755 vdd.n8754 84.1148
R36421 vdd.n8775 vdd.n8768 84.1148
R36422 vdd.n8805 vdd.n8804 84.1148
R36423 vdd.n8825 vdd.n8818 84.1148
R36424 vdd.n8853 vdd.n8852 84.1148
R36425 vdd.n8873 vdd.n8866 84.1148
R36426 vdd.n9019 vdd.n9012 84.1148
R36427 vdd.n8999 vdd.n8995 84.1148
R36428 vdd.n8971 vdd.n8964 84.1148
R36429 vdd.n8951 vdd.n8947 84.1148
R36430 vdd.n9068 vdd.n9061 84.1148
R36431 vdd.n9048 vdd.n9044 84.1148
R36432 vdd.n9118 vdd.n9111 84.1148
R36433 vdd.n9098 vdd.n9094 84.1148
R36434 vdd.n9166 vdd.n9159 84.1148
R36435 vdd.n9146 vdd.n9142 84.1148
R36436 vdd.n7357 vdd.n7356 84.1148
R36437 vdd.n7330 vdd.n7324 84.1148
R36438 vdd.n9314 vdd.n9307 84.1148
R36439 vdd.n9294 vdd.n9290 84.1148
R36440 vdd.n9265 vdd.n9258 84.1148
R36441 vdd.n9245 vdd.n9241 84.1148
R36442 vdd.n9217 vdd.n9210 84.1148
R36443 vdd.n9197 vdd.n9193 84.1148
R36444 vdd.n9363 vdd.n9356 84.1148
R36445 vdd.n9343 vdd.n9339 84.1148
R36446 vdd.n9413 vdd.n9406 84.1148
R36447 vdd.n9393 vdd.n9389 84.1148
R36448 vdd.n9461 vdd.n9454 84.1148
R36449 vdd.n9441 vdd.n9437 84.1148
R36450 vdd.n9559 vdd.n9552 84.1148
R36451 vdd.n9539 vdd.n9535 84.1148
R36452 vdd.n9511 vdd.n9504 84.1148
R36453 vdd.n9491 vdd.n9487 84.1148
R36454 vdd.n9608 vdd.n9601 84.1148
R36455 vdd.n9588 vdd.n9584 84.1148
R36456 vdd.n9658 vdd.n9651 84.1148
R36457 vdd.n9638 vdd.n9634 84.1148
R36458 vdd.n9706 vdd.n9699 84.1148
R36459 vdd.n9686 vdd.n9682 84.1148
R36460 vdd.n7111 vdd.n7110 84.1148
R36461 vdd.n7084 vdd.n7078 84.1148
R36462 vdd.n9805 vdd.n9798 84.1148
R36463 vdd.n9785 vdd.n9781 84.1148
R36464 vdd.n9757 vdd.n9750 84.1148
R36465 vdd.n9737 vdd.n9733 84.1148
R36466 vdd.n9854 vdd.n9847 84.1148
R36467 vdd.n9834 vdd.n9830 84.1148
R36468 vdd.n9904 vdd.n9897 84.1148
R36469 vdd.n9884 vdd.n9880 84.1148
R36470 vdd.n9952 vdd.n9945 84.1148
R36471 vdd.n9932 vdd.n9928 84.1148
R36472 vdd.n3864 vdd.n3857 84.1148
R36473 vdd.n3844 vdd.n3840 84.1148
R36474 vdd.n3912 vdd.n3905 84.1148
R36475 vdd.n3892 vdd.n3888 84.1148
R36476 vdd.n4014 vdd.n4007 84.1148
R36477 vdd.n3994 vdd.n3990 84.1148
R36478 vdd.n4062 vdd.n4055 84.1148
R36479 vdd.n4042 vdd.n4038 84.1148
R36480 vdd.n4110 vdd.n4103 84.1148
R36481 vdd.n4090 vdd.n4086 84.1148
R36482 vdd.n4158 vdd.n4151 84.1148
R36483 vdd.n4138 vdd.n4134 84.1148
R36484 vdd.n4260 vdd.n4253 84.1148
R36485 vdd.n4240 vdd.n4236 84.1148
R36486 vdd.n5780 vdd.n5773 84.1148
R36487 vdd.n5760 vdd.n5756 84.1148
R36488 vdd.n4288 vdd.n4287 84.1148
R36489 vdd.n4308 vdd.n4301 84.1148
R36490 vdd.n4336 vdd.n4335 84.1148
R36491 vdd.n4356 vdd.n4349 84.1148
R36492 vdd.n4437 vdd.n4436 84.1148
R36493 vdd.n4457 vdd.n4450 84.1148
R36494 vdd.n4485 vdd.n4484 84.1148
R36495 vdd.n4505 vdd.n4498 84.1148
R36496 vdd.n4533 vdd.n4532 84.1148
R36497 vdd.n4553 vdd.n4546 84.1148
R36498 vdd.n4581 vdd.n4580 84.1148
R36499 vdd.n4601 vdd.n4594 84.1148
R36500 vdd.n4682 vdd.n4681 84.1148
R36501 vdd.n4702 vdd.n4695 84.1148
R36502 vdd.n3795 vdd.n3794 84.1148
R36503 vdd.n3815 vdd.n3808 84.1148
R36504 vdd.n4730 vdd.n4729 84.1148
R36505 vdd.n4750 vdd.n4743 84.1148
R36506 vdd.n4777 vdd.n4776 84.1148
R36507 vdd.n4797 vdd.n4790 84.1148
R36508 vdd.n4827 vdd.n4826 84.1148
R36509 vdd.n4847 vdd.n4840 84.1148
R36510 vdd.n4877 vdd.n4876 84.1148
R36511 vdd.n4897 vdd.n4890 84.1148
R36512 vdd.n4925 vdd.n4924 84.1148
R36513 vdd.n4945 vdd.n4938 84.1148
R36514 vdd.n4653 vdd.n4612 84.1148
R36515 vdd.n4637 vdd.n4629 84.1148
R36516 vdd.n4976 vdd.n4975 84.1148
R36517 vdd.n4996 vdd.n4989 84.1148
R36518 vdd.n5023 vdd.n5022 84.1148
R36519 vdd.n5043 vdd.n5036 84.1148
R36520 vdd.n5071 vdd.n5070 84.1148
R36521 vdd.n5091 vdd.n5084 84.1148
R36522 vdd.n5122 vdd.n5121 84.1148
R36523 vdd.n5142 vdd.n5135 84.1148
R36524 vdd.n5172 vdd.n5171 84.1148
R36525 vdd.n5192 vdd.n5185 84.1148
R36526 vdd.n5220 vdd.n5219 84.1148
R36527 vdd.n5240 vdd.n5233 84.1148
R36528 vdd.n5270 vdd.n5269 84.1148
R36529 vdd.n5290 vdd.n5283 84.1148
R36530 vdd.n5317 vdd.n5316 84.1148
R36531 vdd.n5337 vdd.n5330 84.1148
R36532 vdd.n5367 vdd.n5366 84.1148
R36533 vdd.n5387 vdd.n5380 84.1148
R36534 vdd.n5417 vdd.n5416 84.1148
R36535 vdd.n5437 vdd.n5430 84.1148
R36536 vdd.n5465 vdd.n5464 84.1148
R36537 vdd.n5485 vdd.n5478 84.1148
R36538 vdd.n4408 vdd.n4367 84.1148
R36539 vdd.n4392 vdd.n4384 84.1148
R36540 vdd.n5516 vdd.n5515 84.1148
R36541 vdd.n5536 vdd.n5529 84.1148
R36542 vdd.n5563 vdd.n5562 84.1148
R36543 vdd.n5583 vdd.n5576 84.1148
R36544 vdd.n5613 vdd.n5612 84.1148
R36545 vdd.n5633 vdd.n5626 84.1148
R36546 vdd.n5663 vdd.n5662 84.1148
R36547 vdd.n5683 vdd.n5676 84.1148
R36548 vdd.n5711 vdd.n5710 84.1148
R36549 vdd.n5731 vdd.n5724 84.1148
R36550 vdd.n5877 vdd.n5870 84.1148
R36551 vdd.n5857 vdd.n5853 84.1148
R36552 vdd.n5829 vdd.n5822 84.1148
R36553 vdd.n5809 vdd.n5805 84.1148
R36554 vdd.n5926 vdd.n5919 84.1148
R36555 vdd.n5906 vdd.n5902 84.1148
R36556 vdd.n5976 vdd.n5969 84.1148
R36557 vdd.n5956 vdd.n5952 84.1148
R36558 vdd.n6024 vdd.n6017 84.1148
R36559 vdd.n6004 vdd.n6000 84.1148
R36560 vdd.n4215 vdd.n4214 84.1148
R36561 vdd.n4188 vdd.n4182 84.1148
R36562 vdd.n6172 vdd.n6165 84.1148
R36563 vdd.n6152 vdd.n6148 84.1148
R36564 vdd.n6123 vdd.n6116 84.1148
R36565 vdd.n6103 vdd.n6099 84.1148
R36566 vdd.n6075 vdd.n6068 84.1148
R36567 vdd.n6055 vdd.n6051 84.1148
R36568 vdd.n6221 vdd.n6214 84.1148
R36569 vdd.n6201 vdd.n6197 84.1148
R36570 vdd.n6271 vdd.n6264 84.1148
R36571 vdd.n6251 vdd.n6247 84.1148
R36572 vdd.n6319 vdd.n6312 84.1148
R36573 vdd.n6299 vdd.n6295 84.1148
R36574 vdd.n6417 vdd.n6410 84.1148
R36575 vdd.n6397 vdd.n6393 84.1148
R36576 vdd.n6369 vdd.n6362 84.1148
R36577 vdd.n6349 vdd.n6345 84.1148
R36578 vdd.n6466 vdd.n6459 84.1148
R36579 vdd.n6446 vdd.n6442 84.1148
R36580 vdd.n6516 vdd.n6509 84.1148
R36581 vdd.n6496 vdd.n6492 84.1148
R36582 vdd.n6564 vdd.n6557 84.1148
R36583 vdd.n6544 vdd.n6540 84.1148
R36584 vdd.n3969 vdd.n3968 84.1148
R36585 vdd.n3942 vdd.n3936 84.1148
R36586 vdd.n6663 vdd.n6656 84.1148
R36587 vdd.n6643 vdd.n6639 84.1148
R36588 vdd.n6615 vdd.n6608 84.1148
R36589 vdd.n6595 vdd.n6591 84.1148
R36590 vdd.n6712 vdd.n6705 84.1148
R36591 vdd.n6692 vdd.n6688 84.1148
R36592 vdd.n6762 vdd.n6755 84.1148
R36593 vdd.n6742 vdd.n6738 84.1148
R36594 vdd.n6810 vdd.n6803 84.1148
R36595 vdd.n6790 vdd.n6786 84.1148
R36596 vdd.n722 vdd.n715 84.1148
R36597 vdd.n702 vdd.n698 84.1148
R36598 vdd.n770 vdd.n763 84.1148
R36599 vdd.n750 vdd.n746 84.1148
R36600 vdd.n872 vdd.n865 84.1148
R36601 vdd.n852 vdd.n848 84.1148
R36602 vdd.n920 vdd.n913 84.1148
R36603 vdd.n900 vdd.n896 84.1148
R36604 vdd.n968 vdd.n961 84.1148
R36605 vdd.n948 vdd.n944 84.1148
R36606 vdd.n1016 vdd.n1009 84.1148
R36607 vdd.n996 vdd.n992 84.1148
R36608 vdd.n1118 vdd.n1111 84.1148
R36609 vdd.n1098 vdd.n1094 84.1148
R36610 vdd.n2638 vdd.n2631 84.1148
R36611 vdd.n2618 vdd.n2614 84.1148
R36612 vdd.n1146 vdd.n1145 84.1148
R36613 vdd.n1166 vdd.n1159 84.1148
R36614 vdd.n1194 vdd.n1193 84.1148
R36615 vdd.n1214 vdd.n1207 84.1148
R36616 vdd.n1295 vdd.n1294 84.1148
R36617 vdd.n1315 vdd.n1308 84.1148
R36618 vdd.n1343 vdd.n1342 84.1148
R36619 vdd.n1363 vdd.n1356 84.1148
R36620 vdd.n1391 vdd.n1390 84.1148
R36621 vdd.n1411 vdd.n1404 84.1148
R36622 vdd.n1439 vdd.n1438 84.1148
R36623 vdd.n1459 vdd.n1452 84.1148
R36624 vdd.n1540 vdd.n1539 84.1148
R36625 vdd.n1560 vdd.n1553 84.1148
R36626 vdd.n653 vdd.n652 84.1148
R36627 vdd.n673 vdd.n666 84.1148
R36628 vdd.n1588 vdd.n1587 84.1148
R36629 vdd.n1608 vdd.n1601 84.1148
R36630 vdd.n1635 vdd.n1634 84.1148
R36631 vdd.n1655 vdd.n1648 84.1148
R36632 vdd.n1685 vdd.n1684 84.1148
R36633 vdd.n1705 vdd.n1698 84.1148
R36634 vdd.n1735 vdd.n1734 84.1148
R36635 vdd.n1755 vdd.n1748 84.1148
R36636 vdd.n1783 vdd.n1782 84.1148
R36637 vdd.n1803 vdd.n1796 84.1148
R36638 vdd.n1511 vdd.n1470 84.1148
R36639 vdd.n1495 vdd.n1487 84.1148
R36640 vdd.n1834 vdd.n1833 84.1148
R36641 vdd.n1854 vdd.n1847 84.1148
R36642 vdd.n1881 vdd.n1880 84.1148
R36643 vdd.n1901 vdd.n1894 84.1148
R36644 vdd.n1929 vdd.n1928 84.1148
R36645 vdd.n1949 vdd.n1942 84.1148
R36646 vdd.n1980 vdd.n1979 84.1148
R36647 vdd.n2000 vdd.n1993 84.1148
R36648 vdd.n2030 vdd.n2029 84.1148
R36649 vdd.n2050 vdd.n2043 84.1148
R36650 vdd.n2078 vdd.n2077 84.1148
R36651 vdd.n2098 vdd.n2091 84.1148
R36652 vdd.n2128 vdd.n2127 84.1148
R36653 vdd.n2148 vdd.n2141 84.1148
R36654 vdd.n2175 vdd.n2174 84.1148
R36655 vdd.n2195 vdd.n2188 84.1148
R36656 vdd.n2225 vdd.n2224 84.1148
R36657 vdd.n2245 vdd.n2238 84.1148
R36658 vdd.n2275 vdd.n2274 84.1148
R36659 vdd.n2295 vdd.n2288 84.1148
R36660 vdd.n2323 vdd.n2322 84.1148
R36661 vdd.n2343 vdd.n2336 84.1148
R36662 vdd.n1266 vdd.n1225 84.1148
R36663 vdd.n1250 vdd.n1242 84.1148
R36664 vdd.n2374 vdd.n2373 84.1148
R36665 vdd.n2394 vdd.n2387 84.1148
R36666 vdd.n2421 vdd.n2420 84.1148
R36667 vdd.n2441 vdd.n2434 84.1148
R36668 vdd.n2471 vdd.n2470 84.1148
R36669 vdd.n2491 vdd.n2484 84.1148
R36670 vdd.n2521 vdd.n2520 84.1148
R36671 vdd.n2541 vdd.n2534 84.1148
R36672 vdd.n2569 vdd.n2568 84.1148
R36673 vdd.n2589 vdd.n2582 84.1148
R36674 vdd.n2735 vdd.n2728 84.1148
R36675 vdd.n2715 vdd.n2711 84.1148
R36676 vdd.n2687 vdd.n2680 84.1148
R36677 vdd.n2667 vdd.n2663 84.1148
R36678 vdd.n2784 vdd.n2777 84.1148
R36679 vdd.n2764 vdd.n2760 84.1148
R36680 vdd.n2834 vdd.n2827 84.1148
R36681 vdd.n2814 vdd.n2810 84.1148
R36682 vdd.n2882 vdd.n2875 84.1148
R36683 vdd.n2862 vdd.n2858 84.1148
R36684 vdd.n1073 vdd.n1072 84.1148
R36685 vdd.n1046 vdd.n1040 84.1148
R36686 vdd.n3030 vdd.n3023 84.1148
R36687 vdd.n3010 vdd.n3006 84.1148
R36688 vdd.n2981 vdd.n2974 84.1148
R36689 vdd.n2961 vdd.n2957 84.1148
R36690 vdd.n2933 vdd.n2926 84.1148
R36691 vdd.n2913 vdd.n2909 84.1148
R36692 vdd.n3079 vdd.n3072 84.1148
R36693 vdd.n3059 vdd.n3055 84.1148
R36694 vdd.n3129 vdd.n3122 84.1148
R36695 vdd.n3109 vdd.n3105 84.1148
R36696 vdd.n3177 vdd.n3170 84.1148
R36697 vdd.n3157 vdd.n3153 84.1148
R36698 vdd.n3275 vdd.n3268 84.1148
R36699 vdd.n3255 vdd.n3251 84.1148
R36700 vdd.n3227 vdd.n3220 84.1148
R36701 vdd.n3207 vdd.n3203 84.1148
R36702 vdd.n3324 vdd.n3317 84.1148
R36703 vdd.n3304 vdd.n3300 84.1148
R36704 vdd.n3374 vdd.n3367 84.1148
R36705 vdd.n3354 vdd.n3350 84.1148
R36706 vdd.n3422 vdd.n3415 84.1148
R36707 vdd.n3402 vdd.n3398 84.1148
R36708 vdd.n827 vdd.n826 84.1148
R36709 vdd.n800 vdd.n794 84.1148
R36710 vdd.n3521 vdd.n3514 84.1148
R36711 vdd.n3501 vdd.n3497 84.1148
R36712 vdd.n3473 vdd.n3466 84.1148
R36713 vdd.n3453 vdd.n3449 84.1148
R36714 vdd.n3570 vdd.n3563 84.1148
R36715 vdd.n3550 vdd.n3546 84.1148
R36716 vdd.n3620 vdd.n3613 84.1148
R36717 vdd.n3600 vdd.n3596 84.1148
R36718 vdd.n3668 vdd.n3661 84.1148
R36719 vdd.n3648 vdd.n3644 84.1148
R36720 vdd.n626 vdd.n619 84.1148
R36721 vdd.n606 vdd.n602 84.1148
R36722 vdd.n3767 vdd.n3760 84.1148
R36723 vdd.n3747 vdd.n3743 84.1148
R36724 vdd.n3719 vdd.n3712 84.1148
R36725 vdd.n3699 vdd.n3695 84.1148
R36726 vdd.n6909 vdd.n6902 84.1148
R36727 vdd.n6889 vdd.n6885 84.1148
R36728 vdd.n6861 vdd.n6854 84.1148
R36729 vdd.n6841 vdd.n6837 84.1148
R36730 vdd.n10051 vdd.n10044 84.1148
R36731 vdd.n10031 vdd.n10027 84.1148
R36732 vdd.n10003 vdd.n9996 84.1148
R36733 vdd.n9983 vdd.n9979 84.1148
R36734 vdd.n10099 vdd.n10092 84.1148
R36735 vdd.n10079 vdd.n10075 84.1148
R36736 vdd.n10147 vdd.n10140 84.1148
R36737 vdd.n10127 vdd.n10123 84.1148
R36738 vdd.n10249 vdd.n10242 84.1148
R36739 vdd.n10229 vdd.n10225 84.1148
R36740 vdd.n10297 vdd.n10290 84.1148
R36741 vdd.n10277 vdd.n10273 84.1148
R36742 vdd.n10345 vdd.n10338 84.1148
R36743 vdd.n10325 vdd.n10321 84.1148
R36744 vdd.n10393 vdd.n10386 84.1148
R36745 vdd.n10373 vdd.n10369 84.1148
R36746 vdd.n10495 vdd.n10488 84.1148
R36747 vdd.n10475 vdd.n10471 84.1148
R36748 vdd.n87 vdd.n80 84.1148
R36749 vdd.n67 vdd.n63 84.1148
R36750 vdd.n39 vdd.n32 84.1148
R36751 vdd.n19 vdd.n15 84.1148
R36752 vdd.n10543 vdd.n10536 84.1148
R36753 vdd.n10523 vdd.n10519 84.1148
R36754 vdd.n10593 vdd.n10586 84.1148
R36755 vdd.n10573 vdd.n10569 84.1148
R36756 vdd.n10641 vdd.n10634 84.1148
R36757 vdd.n10621 vdd.n10617 84.1148
R36758 vdd.n10450 vdd.n10449 84.1148
R36759 vdd.n10423 vdd.n10417 84.1148
R36760 vdd.n10789 vdd.n10782 84.1148
R36761 vdd.n10769 vdd.n10765 84.1148
R36762 vdd.n10740 vdd.n10733 84.1148
R36763 vdd.n10720 vdd.n10716 84.1148
R36764 vdd.n10692 vdd.n10685 84.1148
R36765 vdd.n10672 vdd.n10668 84.1148
R36766 vdd.n10838 vdd.n10831 84.1148
R36767 vdd.n10818 vdd.n10814 84.1148
R36768 vdd.n10888 vdd.n10881 84.1148
R36769 vdd.n10868 vdd.n10864 84.1148
R36770 vdd.n10936 vdd.n10929 84.1148
R36771 vdd.n10916 vdd.n10912 84.1148
R36772 vdd.n11034 vdd.n11027 84.1148
R36773 vdd.n11014 vdd.n11010 84.1148
R36774 vdd.n10986 vdd.n10979 84.1148
R36775 vdd.n10966 vdd.n10962 84.1148
R36776 vdd.n11083 vdd.n11076 84.1148
R36777 vdd.n11063 vdd.n11059 84.1148
R36778 vdd.n11133 vdd.n11126 84.1148
R36779 vdd.n11113 vdd.n11109 84.1148
R36780 vdd.n11181 vdd.n11174 84.1148
R36781 vdd.n11161 vdd.n11157 84.1148
R36782 vdd.n10204 vdd.n10203 84.1148
R36783 vdd.n10177 vdd.n10171 84.1148
R36784 vdd.n11280 vdd.n11273 84.1148
R36785 vdd.n11260 vdd.n11256 84.1148
R36786 vdd.n11232 vdd.n11225 84.1148
R36787 vdd.n11212 vdd.n11208 84.1148
R36788 vdd.n11329 vdd.n11322 84.1148
R36789 vdd.n11309 vdd.n11305 84.1148
R36790 vdd.n11379 vdd.n11372 84.1148
R36791 vdd.n11359 vdd.n11355 84.1148
R36792 vdd.n11427 vdd.n11420 84.1148
R36793 vdd.n11407 vdd.n11403 84.1148
R36794 vdd.n11458 vdd.n11457 84.1148
R36795 vdd.n11478 vdd.n11471 84.1148
R36796 vdd.n11505 vdd.n11504 84.1148
R36797 vdd.n11525 vdd.n11518 84.1148
R36798 vdd.n11555 vdd.n11554 84.1148
R36799 vdd.n11575 vdd.n11568 84.1148
R36800 vdd.n11605 vdd.n11604 84.1148
R36801 vdd.n11625 vdd.n11618 84.1148
R36802 vdd.n11653 vdd.n11652 84.1148
R36803 vdd.n11673 vdd.n11666 84.1148
R36804 vdd.n481 vdd.n440 84.1148
R36805 vdd.n465 vdd.n457 84.1148
R36806 vdd.n11704 vdd.n11703 84.1148
R36807 vdd.n11724 vdd.n11717 84.1148
R36808 vdd.n11751 vdd.n11750 84.1148
R36809 vdd.n11771 vdd.n11764 84.1148
R36810 vdd.n11799 vdd.n11798 84.1148
R36811 vdd.n11819 vdd.n11812 84.1148
R36812 vdd.n11850 vdd.n11849 84.1148
R36813 vdd.n11870 vdd.n11863 84.1148
R36814 vdd.n11900 vdd.n11899 84.1148
R36815 vdd.n11920 vdd.n11913 84.1148
R36816 vdd.n11948 vdd.n11947 84.1148
R36817 vdd.n11968 vdd.n11961 84.1148
R36818 vdd.n11998 vdd.n11997 84.1148
R36819 vdd.n12018 vdd.n12011 84.1148
R36820 vdd.n12045 vdd.n12044 84.1148
R36821 vdd.n12065 vdd.n12058 84.1148
R36822 vdd.n12095 vdd.n12094 84.1148
R36823 vdd.n12115 vdd.n12108 84.1148
R36824 vdd.n12145 vdd.n12144 84.1148
R36825 vdd.n12165 vdd.n12158 84.1148
R36826 vdd.n12193 vdd.n12192 84.1148
R36827 vdd.n12213 vdd.n12206 84.1148
R36828 vdd.n236 vdd.n195 84.1148
R36829 vdd.n220 vdd.n212 84.1148
R36830 vdd.n12244 vdd.n12243 84.1148
R36831 vdd.n12264 vdd.n12257 84.1148
R36832 vdd.n12291 vdd.n12290 84.1148
R36833 vdd.n12311 vdd.n12304 84.1148
R36834 vdd.n12341 vdd.n12340 84.1148
R36835 vdd.n12361 vdd.n12354 84.1148
R36836 vdd.n12391 vdd.n12390 84.1148
R36837 vdd.n12411 vdd.n12404 84.1148
R36838 vdd.n12439 vdd.n12438 84.1148
R36839 vdd.n12459 vdd.n12452 84.1148
R36840 vdd.n12506 vdd.n12500 63.3004
R36841 vdd.n12483 vdd.n12477 63.3004
R36842 vdd.n115 vdd.n114 63.3004
R36843 vdd.n131 vdd.n129 63.3004
R36844 vdd.n163 vdd.n162 63.3004
R36845 vdd.n179 vdd.n177 63.3004
R36846 vdd.n264 vdd.n263 63.3004
R36847 vdd.n280 vdd.n278 63.3004
R36848 vdd.n312 vdd.n311 63.3004
R36849 vdd.n328 vdd.n326 63.3004
R36850 vdd.n360 vdd.n359 63.3004
R36851 vdd.n376 vdd.n374 63.3004
R36852 vdd.n408 vdd.n407 63.3004
R36853 vdd.n424 vdd.n422 63.3004
R36854 vdd.n509 vdd.n508 63.3004
R36855 vdd.n525 vdd.n523 63.3004
R36856 vdd.n557 vdd.n556 63.3004
R36857 vdd.n573 vdd.n571 63.3004
R36858 vdd.n7001 vdd.n6999 63.3004
R36859 vdd.n6989 vdd.n6986 63.3004
R36860 vdd.n7049 vdd.n7047 63.3004
R36861 vdd.n7037 vdd.n7034 63.3004
R36862 vdd.n7151 vdd.n7149 63.3004
R36863 vdd.n7139 vdd.n7136 63.3004
R36864 vdd.n7199 vdd.n7197 63.3004
R36865 vdd.n7187 vdd.n7184 63.3004
R36866 vdd.n7247 vdd.n7245 63.3004
R36867 vdd.n7235 vdd.n7232 63.3004
R36868 vdd.n7295 vdd.n7293 63.3004
R36869 vdd.n7283 vdd.n7280 63.3004
R36870 vdd.n7397 vdd.n7395 63.3004
R36871 vdd.n7385 vdd.n7382 63.3004
R36872 vdd.n8917 vdd.n8915 63.3004
R36873 vdd.n8905 vdd.n8902 63.3004
R36874 vdd.n7429 vdd.n7428 63.3004
R36875 vdd.n7445 vdd.n7443 63.3004
R36876 vdd.n7477 vdd.n7476 63.3004
R36877 vdd.n7493 vdd.n7491 63.3004
R36878 vdd.n7578 vdd.n7577 63.3004
R36879 vdd.n7594 vdd.n7592 63.3004
R36880 vdd.n7626 vdd.n7625 63.3004
R36881 vdd.n7642 vdd.n7640 63.3004
R36882 vdd.n7674 vdd.n7673 63.3004
R36883 vdd.n7690 vdd.n7688 63.3004
R36884 vdd.n7722 vdd.n7721 63.3004
R36885 vdd.n7738 vdd.n7736 63.3004
R36886 vdd.n7823 vdd.n7822 63.3004
R36887 vdd.n7839 vdd.n7837 63.3004
R36888 vdd.n6936 vdd.n6935 63.3004
R36889 vdd.n6952 vdd.n6950 63.3004
R36890 vdd.n7871 vdd.n7870 63.3004
R36891 vdd.n7887 vdd.n7885 63.3004
R36892 vdd.n7918 vdd.n7917 63.3004
R36893 vdd.n7934 vdd.n7932 63.3004
R36894 vdd.n7968 vdd.n7967 63.3004
R36895 vdd.n7984 vdd.n7982 63.3004
R36896 vdd.n8018 vdd.n8017 63.3004
R36897 vdd.n8034 vdd.n8032 63.3004
R36898 vdd.n8066 vdd.n8065 63.3004
R36899 vdd.n8082 vdd.n8080 63.3004
R36900 vdd.n7774 vdd.n7771 63.3004
R36901 vdd.n8117 vdd.n8116 63.3004
R36902 vdd.n8133 vdd.n8131 63.3004
R36903 vdd.n8164 vdd.n8163 63.3004
R36904 vdd.n8180 vdd.n8178 63.3004
R36905 vdd.n8212 vdd.n8211 63.3004
R36906 vdd.n8228 vdd.n8226 63.3004
R36907 vdd.n8263 vdd.n8262 63.3004
R36908 vdd.n8279 vdd.n8277 63.3004
R36909 vdd.n8313 vdd.n8312 63.3004
R36910 vdd.n8329 vdd.n8327 63.3004
R36911 vdd.n8361 vdd.n8360 63.3004
R36912 vdd.n8377 vdd.n8375 63.3004
R36913 vdd.n8411 vdd.n8410 63.3004
R36914 vdd.n8427 vdd.n8425 63.3004
R36915 vdd.n8458 vdd.n8457 63.3004
R36916 vdd.n8474 vdd.n8472 63.3004
R36917 vdd.n8508 vdd.n8507 63.3004
R36918 vdd.n8524 vdd.n8522 63.3004
R36919 vdd.n8558 vdd.n8557 63.3004
R36920 vdd.n8574 vdd.n8572 63.3004
R36921 vdd.n8606 vdd.n8605 63.3004
R36922 vdd.n8622 vdd.n8620 63.3004
R36923 vdd.n7529 vdd.n7526 63.3004
R36924 vdd.n8657 vdd.n8656 63.3004
R36925 vdd.n8673 vdd.n8671 63.3004
R36926 vdd.n8704 vdd.n8703 63.3004
R36927 vdd.n8720 vdd.n8718 63.3004
R36928 vdd.n8754 vdd.n8753 63.3004
R36929 vdd.n8770 vdd.n8768 63.3004
R36930 vdd.n8804 vdd.n8803 63.3004
R36931 vdd.n8820 vdd.n8818 63.3004
R36932 vdd.n8852 vdd.n8851 63.3004
R36933 vdd.n8868 vdd.n8866 63.3004
R36934 vdd.n9014 vdd.n9012 63.3004
R36935 vdd.n9002 vdd.n8999 63.3004
R36936 vdd.n8966 vdd.n8964 63.3004
R36937 vdd.n8954 vdd.n8951 63.3004
R36938 vdd.n9063 vdd.n9061 63.3004
R36939 vdd.n9051 vdd.n9048 63.3004
R36940 vdd.n9113 vdd.n9111 63.3004
R36941 vdd.n9101 vdd.n9098 63.3004
R36942 vdd.n9161 vdd.n9159 63.3004
R36943 vdd.n9149 vdd.n9146 63.3004
R36944 vdd.n7335 vdd.n7324 63.3004
R36945 vdd.n9309 vdd.n9307 63.3004
R36946 vdd.n9297 vdd.n9294 63.3004
R36947 vdd.n9260 vdd.n9258 63.3004
R36948 vdd.n9248 vdd.n9245 63.3004
R36949 vdd.n9212 vdd.n9210 63.3004
R36950 vdd.n9200 vdd.n9197 63.3004
R36951 vdd.n9358 vdd.n9356 63.3004
R36952 vdd.n9346 vdd.n9343 63.3004
R36953 vdd.n9408 vdd.n9406 63.3004
R36954 vdd.n9396 vdd.n9393 63.3004
R36955 vdd.n9456 vdd.n9454 63.3004
R36956 vdd.n9444 vdd.n9441 63.3004
R36957 vdd.n9554 vdd.n9552 63.3004
R36958 vdd.n9542 vdd.n9539 63.3004
R36959 vdd.n9506 vdd.n9504 63.3004
R36960 vdd.n9494 vdd.n9491 63.3004
R36961 vdd.n9603 vdd.n9601 63.3004
R36962 vdd.n9591 vdd.n9588 63.3004
R36963 vdd.n9653 vdd.n9651 63.3004
R36964 vdd.n9641 vdd.n9638 63.3004
R36965 vdd.n9701 vdd.n9699 63.3004
R36966 vdd.n9689 vdd.n9686 63.3004
R36967 vdd.n7089 vdd.n7078 63.3004
R36968 vdd.n9800 vdd.n9798 63.3004
R36969 vdd.n9788 vdd.n9785 63.3004
R36970 vdd.n9752 vdd.n9750 63.3004
R36971 vdd.n9740 vdd.n9737 63.3004
R36972 vdd.n9849 vdd.n9847 63.3004
R36973 vdd.n9837 vdd.n9834 63.3004
R36974 vdd.n9899 vdd.n9897 63.3004
R36975 vdd.n9887 vdd.n9884 63.3004
R36976 vdd.n9947 vdd.n9945 63.3004
R36977 vdd.n9935 vdd.n9932 63.3004
R36978 vdd.n3859 vdd.n3857 63.3004
R36979 vdd.n3847 vdd.n3844 63.3004
R36980 vdd.n3907 vdd.n3905 63.3004
R36981 vdd.n3895 vdd.n3892 63.3004
R36982 vdd.n4009 vdd.n4007 63.3004
R36983 vdd.n3997 vdd.n3994 63.3004
R36984 vdd.n4057 vdd.n4055 63.3004
R36985 vdd.n4045 vdd.n4042 63.3004
R36986 vdd.n4105 vdd.n4103 63.3004
R36987 vdd.n4093 vdd.n4090 63.3004
R36988 vdd.n4153 vdd.n4151 63.3004
R36989 vdd.n4141 vdd.n4138 63.3004
R36990 vdd.n4255 vdd.n4253 63.3004
R36991 vdd.n4243 vdd.n4240 63.3004
R36992 vdd.n5775 vdd.n5773 63.3004
R36993 vdd.n5763 vdd.n5760 63.3004
R36994 vdd.n4287 vdd.n4286 63.3004
R36995 vdd.n4303 vdd.n4301 63.3004
R36996 vdd.n4335 vdd.n4334 63.3004
R36997 vdd.n4351 vdd.n4349 63.3004
R36998 vdd.n4436 vdd.n4435 63.3004
R36999 vdd.n4452 vdd.n4450 63.3004
R37000 vdd.n4484 vdd.n4483 63.3004
R37001 vdd.n4500 vdd.n4498 63.3004
R37002 vdd.n4532 vdd.n4531 63.3004
R37003 vdd.n4548 vdd.n4546 63.3004
R37004 vdd.n4580 vdd.n4579 63.3004
R37005 vdd.n4596 vdd.n4594 63.3004
R37006 vdd.n4681 vdd.n4680 63.3004
R37007 vdd.n4697 vdd.n4695 63.3004
R37008 vdd.n3794 vdd.n3793 63.3004
R37009 vdd.n3810 vdd.n3808 63.3004
R37010 vdd.n4729 vdd.n4728 63.3004
R37011 vdd.n4745 vdd.n4743 63.3004
R37012 vdd.n4776 vdd.n4775 63.3004
R37013 vdd.n4792 vdd.n4790 63.3004
R37014 vdd.n4826 vdd.n4825 63.3004
R37015 vdd.n4842 vdd.n4840 63.3004
R37016 vdd.n4876 vdd.n4875 63.3004
R37017 vdd.n4892 vdd.n4890 63.3004
R37018 vdd.n4924 vdd.n4923 63.3004
R37019 vdd.n4940 vdd.n4938 63.3004
R37020 vdd.n4632 vdd.n4629 63.3004
R37021 vdd.n4975 vdd.n4974 63.3004
R37022 vdd.n4991 vdd.n4989 63.3004
R37023 vdd.n5022 vdd.n5021 63.3004
R37024 vdd.n5038 vdd.n5036 63.3004
R37025 vdd.n5070 vdd.n5069 63.3004
R37026 vdd.n5086 vdd.n5084 63.3004
R37027 vdd.n5121 vdd.n5120 63.3004
R37028 vdd.n5137 vdd.n5135 63.3004
R37029 vdd.n5171 vdd.n5170 63.3004
R37030 vdd.n5187 vdd.n5185 63.3004
R37031 vdd.n5219 vdd.n5218 63.3004
R37032 vdd.n5235 vdd.n5233 63.3004
R37033 vdd.n5269 vdd.n5268 63.3004
R37034 vdd.n5285 vdd.n5283 63.3004
R37035 vdd.n5316 vdd.n5315 63.3004
R37036 vdd.n5332 vdd.n5330 63.3004
R37037 vdd.n5366 vdd.n5365 63.3004
R37038 vdd.n5382 vdd.n5380 63.3004
R37039 vdd.n5416 vdd.n5415 63.3004
R37040 vdd.n5432 vdd.n5430 63.3004
R37041 vdd.n5464 vdd.n5463 63.3004
R37042 vdd.n5480 vdd.n5478 63.3004
R37043 vdd.n4387 vdd.n4384 63.3004
R37044 vdd.n5515 vdd.n5514 63.3004
R37045 vdd.n5531 vdd.n5529 63.3004
R37046 vdd.n5562 vdd.n5561 63.3004
R37047 vdd.n5578 vdd.n5576 63.3004
R37048 vdd.n5612 vdd.n5611 63.3004
R37049 vdd.n5628 vdd.n5626 63.3004
R37050 vdd.n5662 vdd.n5661 63.3004
R37051 vdd.n5678 vdd.n5676 63.3004
R37052 vdd.n5710 vdd.n5709 63.3004
R37053 vdd.n5726 vdd.n5724 63.3004
R37054 vdd.n5872 vdd.n5870 63.3004
R37055 vdd.n5860 vdd.n5857 63.3004
R37056 vdd.n5824 vdd.n5822 63.3004
R37057 vdd.n5812 vdd.n5809 63.3004
R37058 vdd.n5921 vdd.n5919 63.3004
R37059 vdd.n5909 vdd.n5906 63.3004
R37060 vdd.n5971 vdd.n5969 63.3004
R37061 vdd.n5959 vdd.n5956 63.3004
R37062 vdd.n6019 vdd.n6017 63.3004
R37063 vdd.n6007 vdd.n6004 63.3004
R37064 vdd.n4193 vdd.n4182 63.3004
R37065 vdd.n6167 vdd.n6165 63.3004
R37066 vdd.n6155 vdd.n6152 63.3004
R37067 vdd.n6118 vdd.n6116 63.3004
R37068 vdd.n6106 vdd.n6103 63.3004
R37069 vdd.n6070 vdd.n6068 63.3004
R37070 vdd.n6058 vdd.n6055 63.3004
R37071 vdd.n6216 vdd.n6214 63.3004
R37072 vdd.n6204 vdd.n6201 63.3004
R37073 vdd.n6266 vdd.n6264 63.3004
R37074 vdd.n6254 vdd.n6251 63.3004
R37075 vdd.n6314 vdd.n6312 63.3004
R37076 vdd.n6302 vdd.n6299 63.3004
R37077 vdd.n6412 vdd.n6410 63.3004
R37078 vdd.n6400 vdd.n6397 63.3004
R37079 vdd.n6364 vdd.n6362 63.3004
R37080 vdd.n6352 vdd.n6349 63.3004
R37081 vdd.n6461 vdd.n6459 63.3004
R37082 vdd.n6449 vdd.n6446 63.3004
R37083 vdd.n6511 vdd.n6509 63.3004
R37084 vdd.n6499 vdd.n6496 63.3004
R37085 vdd.n6559 vdd.n6557 63.3004
R37086 vdd.n6547 vdd.n6544 63.3004
R37087 vdd.n3947 vdd.n3936 63.3004
R37088 vdd.n6658 vdd.n6656 63.3004
R37089 vdd.n6646 vdd.n6643 63.3004
R37090 vdd.n6610 vdd.n6608 63.3004
R37091 vdd.n6598 vdd.n6595 63.3004
R37092 vdd.n6707 vdd.n6705 63.3004
R37093 vdd.n6695 vdd.n6692 63.3004
R37094 vdd.n6757 vdd.n6755 63.3004
R37095 vdd.n6745 vdd.n6742 63.3004
R37096 vdd.n6805 vdd.n6803 63.3004
R37097 vdd.n6793 vdd.n6790 63.3004
R37098 vdd.n717 vdd.n715 63.3004
R37099 vdd.n705 vdd.n702 63.3004
R37100 vdd.n765 vdd.n763 63.3004
R37101 vdd.n753 vdd.n750 63.3004
R37102 vdd.n867 vdd.n865 63.3004
R37103 vdd.n855 vdd.n852 63.3004
R37104 vdd.n915 vdd.n913 63.3004
R37105 vdd.n903 vdd.n900 63.3004
R37106 vdd.n963 vdd.n961 63.3004
R37107 vdd.n951 vdd.n948 63.3004
R37108 vdd.n1011 vdd.n1009 63.3004
R37109 vdd.n999 vdd.n996 63.3004
R37110 vdd.n1113 vdd.n1111 63.3004
R37111 vdd.n1101 vdd.n1098 63.3004
R37112 vdd.n2633 vdd.n2631 63.3004
R37113 vdd.n2621 vdd.n2618 63.3004
R37114 vdd.n1145 vdd.n1144 63.3004
R37115 vdd.n1161 vdd.n1159 63.3004
R37116 vdd.n1193 vdd.n1192 63.3004
R37117 vdd.n1209 vdd.n1207 63.3004
R37118 vdd.n1294 vdd.n1293 63.3004
R37119 vdd.n1310 vdd.n1308 63.3004
R37120 vdd.n1342 vdd.n1341 63.3004
R37121 vdd.n1358 vdd.n1356 63.3004
R37122 vdd.n1390 vdd.n1389 63.3004
R37123 vdd.n1406 vdd.n1404 63.3004
R37124 vdd.n1438 vdd.n1437 63.3004
R37125 vdd.n1454 vdd.n1452 63.3004
R37126 vdd.n1539 vdd.n1538 63.3004
R37127 vdd.n1555 vdd.n1553 63.3004
R37128 vdd.n652 vdd.n651 63.3004
R37129 vdd.n668 vdd.n666 63.3004
R37130 vdd.n1587 vdd.n1586 63.3004
R37131 vdd.n1603 vdd.n1601 63.3004
R37132 vdd.n1634 vdd.n1633 63.3004
R37133 vdd.n1650 vdd.n1648 63.3004
R37134 vdd.n1684 vdd.n1683 63.3004
R37135 vdd.n1700 vdd.n1698 63.3004
R37136 vdd.n1734 vdd.n1733 63.3004
R37137 vdd.n1750 vdd.n1748 63.3004
R37138 vdd.n1782 vdd.n1781 63.3004
R37139 vdd.n1798 vdd.n1796 63.3004
R37140 vdd.n1490 vdd.n1487 63.3004
R37141 vdd.n1833 vdd.n1832 63.3004
R37142 vdd.n1849 vdd.n1847 63.3004
R37143 vdd.n1880 vdd.n1879 63.3004
R37144 vdd.n1896 vdd.n1894 63.3004
R37145 vdd.n1928 vdd.n1927 63.3004
R37146 vdd.n1944 vdd.n1942 63.3004
R37147 vdd.n1979 vdd.n1978 63.3004
R37148 vdd.n1995 vdd.n1993 63.3004
R37149 vdd.n2029 vdd.n2028 63.3004
R37150 vdd.n2045 vdd.n2043 63.3004
R37151 vdd.n2077 vdd.n2076 63.3004
R37152 vdd.n2093 vdd.n2091 63.3004
R37153 vdd.n2127 vdd.n2126 63.3004
R37154 vdd.n2143 vdd.n2141 63.3004
R37155 vdd.n2174 vdd.n2173 63.3004
R37156 vdd.n2190 vdd.n2188 63.3004
R37157 vdd.n2224 vdd.n2223 63.3004
R37158 vdd.n2240 vdd.n2238 63.3004
R37159 vdd.n2274 vdd.n2273 63.3004
R37160 vdd.n2290 vdd.n2288 63.3004
R37161 vdd.n2322 vdd.n2321 63.3004
R37162 vdd.n2338 vdd.n2336 63.3004
R37163 vdd.n1245 vdd.n1242 63.3004
R37164 vdd.n2373 vdd.n2372 63.3004
R37165 vdd.n2389 vdd.n2387 63.3004
R37166 vdd.n2420 vdd.n2419 63.3004
R37167 vdd.n2436 vdd.n2434 63.3004
R37168 vdd.n2470 vdd.n2469 63.3004
R37169 vdd.n2486 vdd.n2484 63.3004
R37170 vdd.n2520 vdd.n2519 63.3004
R37171 vdd.n2536 vdd.n2534 63.3004
R37172 vdd.n2568 vdd.n2567 63.3004
R37173 vdd.n2584 vdd.n2582 63.3004
R37174 vdd.n2730 vdd.n2728 63.3004
R37175 vdd.n2718 vdd.n2715 63.3004
R37176 vdd.n2682 vdd.n2680 63.3004
R37177 vdd.n2670 vdd.n2667 63.3004
R37178 vdd.n2779 vdd.n2777 63.3004
R37179 vdd.n2767 vdd.n2764 63.3004
R37180 vdd.n2829 vdd.n2827 63.3004
R37181 vdd.n2817 vdd.n2814 63.3004
R37182 vdd.n2877 vdd.n2875 63.3004
R37183 vdd.n2865 vdd.n2862 63.3004
R37184 vdd.n1051 vdd.n1040 63.3004
R37185 vdd.n3025 vdd.n3023 63.3004
R37186 vdd.n3013 vdd.n3010 63.3004
R37187 vdd.n2976 vdd.n2974 63.3004
R37188 vdd.n2964 vdd.n2961 63.3004
R37189 vdd.n2928 vdd.n2926 63.3004
R37190 vdd.n2916 vdd.n2913 63.3004
R37191 vdd.n3074 vdd.n3072 63.3004
R37192 vdd.n3062 vdd.n3059 63.3004
R37193 vdd.n3124 vdd.n3122 63.3004
R37194 vdd.n3112 vdd.n3109 63.3004
R37195 vdd.n3172 vdd.n3170 63.3004
R37196 vdd.n3160 vdd.n3157 63.3004
R37197 vdd.n3270 vdd.n3268 63.3004
R37198 vdd.n3258 vdd.n3255 63.3004
R37199 vdd.n3222 vdd.n3220 63.3004
R37200 vdd.n3210 vdd.n3207 63.3004
R37201 vdd.n3319 vdd.n3317 63.3004
R37202 vdd.n3307 vdd.n3304 63.3004
R37203 vdd.n3369 vdd.n3367 63.3004
R37204 vdd.n3357 vdd.n3354 63.3004
R37205 vdd.n3417 vdd.n3415 63.3004
R37206 vdd.n3405 vdd.n3402 63.3004
R37207 vdd.n805 vdd.n794 63.3004
R37208 vdd.n3516 vdd.n3514 63.3004
R37209 vdd.n3504 vdd.n3501 63.3004
R37210 vdd.n3468 vdd.n3466 63.3004
R37211 vdd.n3456 vdd.n3453 63.3004
R37212 vdd.n3565 vdd.n3563 63.3004
R37213 vdd.n3553 vdd.n3550 63.3004
R37214 vdd.n3615 vdd.n3613 63.3004
R37215 vdd.n3603 vdd.n3600 63.3004
R37216 vdd.n3663 vdd.n3661 63.3004
R37217 vdd.n3651 vdd.n3648 63.3004
R37218 vdd.n621 vdd.n619 63.3004
R37219 vdd.n609 vdd.n606 63.3004
R37220 vdd.n3762 vdd.n3760 63.3004
R37221 vdd.n3750 vdd.n3747 63.3004
R37222 vdd.n3714 vdd.n3712 63.3004
R37223 vdd.n3702 vdd.n3699 63.3004
R37224 vdd.n6904 vdd.n6902 63.3004
R37225 vdd.n6892 vdd.n6889 63.3004
R37226 vdd.n6856 vdd.n6854 63.3004
R37227 vdd.n6844 vdd.n6841 63.3004
R37228 vdd.n10046 vdd.n10044 63.3004
R37229 vdd.n10034 vdd.n10031 63.3004
R37230 vdd.n9998 vdd.n9996 63.3004
R37231 vdd.n9986 vdd.n9983 63.3004
R37232 vdd.n10094 vdd.n10092 63.3004
R37233 vdd.n10082 vdd.n10079 63.3004
R37234 vdd.n10142 vdd.n10140 63.3004
R37235 vdd.n10130 vdd.n10127 63.3004
R37236 vdd.n10244 vdd.n10242 63.3004
R37237 vdd.n10232 vdd.n10229 63.3004
R37238 vdd.n10292 vdd.n10290 63.3004
R37239 vdd.n10280 vdd.n10277 63.3004
R37240 vdd.n10340 vdd.n10338 63.3004
R37241 vdd.n10328 vdd.n10325 63.3004
R37242 vdd.n10388 vdd.n10386 63.3004
R37243 vdd.n10376 vdd.n10373 63.3004
R37244 vdd.n10490 vdd.n10488 63.3004
R37245 vdd.n10478 vdd.n10475 63.3004
R37246 vdd.n82 vdd.n80 63.3004
R37247 vdd.n70 vdd.n67 63.3004
R37248 vdd.n34 vdd.n32 63.3004
R37249 vdd.n22 vdd.n19 63.3004
R37250 vdd.n10538 vdd.n10536 63.3004
R37251 vdd.n10526 vdd.n10523 63.3004
R37252 vdd.n10588 vdd.n10586 63.3004
R37253 vdd.n10576 vdd.n10573 63.3004
R37254 vdd.n10636 vdd.n10634 63.3004
R37255 vdd.n10624 vdd.n10621 63.3004
R37256 vdd.n10428 vdd.n10417 63.3004
R37257 vdd.n10784 vdd.n10782 63.3004
R37258 vdd.n10772 vdd.n10769 63.3004
R37259 vdd.n10735 vdd.n10733 63.3004
R37260 vdd.n10723 vdd.n10720 63.3004
R37261 vdd.n10687 vdd.n10685 63.3004
R37262 vdd.n10675 vdd.n10672 63.3004
R37263 vdd.n10833 vdd.n10831 63.3004
R37264 vdd.n10821 vdd.n10818 63.3004
R37265 vdd.n10883 vdd.n10881 63.3004
R37266 vdd.n10871 vdd.n10868 63.3004
R37267 vdd.n10931 vdd.n10929 63.3004
R37268 vdd.n10919 vdd.n10916 63.3004
R37269 vdd.n11029 vdd.n11027 63.3004
R37270 vdd.n11017 vdd.n11014 63.3004
R37271 vdd.n10981 vdd.n10979 63.3004
R37272 vdd.n10969 vdd.n10966 63.3004
R37273 vdd.n11078 vdd.n11076 63.3004
R37274 vdd.n11066 vdd.n11063 63.3004
R37275 vdd.n11128 vdd.n11126 63.3004
R37276 vdd.n11116 vdd.n11113 63.3004
R37277 vdd.n11176 vdd.n11174 63.3004
R37278 vdd.n11164 vdd.n11161 63.3004
R37279 vdd.n10182 vdd.n10171 63.3004
R37280 vdd.n11275 vdd.n11273 63.3004
R37281 vdd.n11263 vdd.n11260 63.3004
R37282 vdd.n11227 vdd.n11225 63.3004
R37283 vdd.n11215 vdd.n11212 63.3004
R37284 vdd.n11324 vdd.n11322 63.3004
R37285 vdd.n11312 vdd.n11309 63.3004
R37286 vdd.n11374 vdd.n11372 63.3004
R37287 vdd.n11362 vdd.n11359 63.3004
R37288 vdd.n11422 vdd.n11420 63.3004
R37289 vdd.n11410 vdd.n11407 63.3004
R37290 vdd.n11457 vdd.n11456 63.3004
R37291 vdd.n11473 vdd.n11471 63.3004
R37292 vdd.n11504 vdd.n11503 63.3004
R37293 vdd.n11520 vdd.n11518 63.3004
R37294 vdd.n11554 vdd.n11553 63.3004
R37295 vdd.n11570 vdd.n11568 63.3004
R37296 vdd.n11604 vdd.n11603 63.3004
R37297 vdd.n11620 vdd.n11618 63.3004
R37298 vdd.n11652 vdd.n11651 63.3004
R37299 vdd.n11668 vdd.n11666 63.3004
R37300 vdd.n460 vdd.n457 63.3004
R37301 vdd.n11703 vdd.n11702 63.3004
R37302 vdd.n11719 vdd.n11717 63.3004
R37303 vdd.n11750 vdd.n11749 63.3004
R37304 vdd.n11766 vdd.n11764 63.3004
R37305 vdd.n11798 vdd.n11797 63.3004
R37306 vdd.n11814 vdd.n11812 63.3004
R37307 vdd.n11849 vdd.n11848 63.3004
R37308 vdd.n11865 vdd.n11863 63.3004
R37309 vdd.n11899 vdd.n11898 63.3004
R37310 vdd.n11915 vdd.n11913 63.3004
R37311 vdd.n11947 vdd.n11946 63.3004
R37312 vdd.n11963 vdd.n11961 63.3004
R37313 vdd.n11997 vdd.n11996 63.3004
R37314 vdd.n12013 vdd.n12011 63.3004
R37315 vdd.n12044 vdd.n12043 63.3004
R37316 vdd.n12060 vdd.n12058 63.3004
R37317 vdd.n12094 vdd.n12093 63.3004
R37318 vdd.n12110 vdd.n12108 63.3004
R37319 vdd.n12144 vdd.n12143 63.3004
R37320 vdd.n12160 vdd.n12158 63.3004
R37321 vdd.n12192 vdd.n12191 63.3004
R37322 vdd.n12208 vdd.n12206 63.3004
R37323 vdd.n215 vdd.n212 63.3004
R37324 vdd.n12243 vdd.n12242 63.3004
R37325 vdd.n12259 vdd.n12257 63.3004
R37326 vdd.n12290 vdd.n12289 63.3004
R37327 vdd.n12306 vdd.n12304 63.3004
R37328 vdd.n12340 vdd.n12339 63.3004
R37329 vdd.n12356 vdd.n12354 63.3004
R37330 vdd.n12390 vdd.n12389 63.3004
R37331 vdd.n12406 vdd.n12404 63.3004
R37332 vdd.n12438 vdd.n12437 63.3004
R37333 vdd.n12454 vdd.n12452 63.3004
R37334 vdd.n7801 vdd.n7754 50.8372
R37335 vdd.n7556 vdd.n7509 50.8372
R37336 vdd.n7358 vdd.n7357 50.8372
R37337 vdd.n7112 vdd.n7111 50.8372
R37338 vdd.n4659 vdd.n4612 50.8372
R37339 vdd.n4414 vdd.n4367 50.8372
R37340 vdd.n4216 vdd.n4215 50.8372
R37341 vdd.n3970 vdd.n3969 50.8372
R37342 vdd.n1517 vdd.n1470 50.8372
R37343 vdd.n1272 vdd.n1225 50.8372
R37344 vdd.n1074 vdd.n1073 50.8372
R37345 vdd.n828 vdd.n827 50.8372
R37346 vdd.n10451 vdd.n10450 50.8372
R37347 vdd.n10205 vdd.n10204 50.8372
R37348 vdd.n487 vdd.n440 50.8372
R37349 vdd.n242 vdd.n195 50.8372
R37350 vdd.n12491 vdd.n12489 35.2919
R37351 vdd.n12491 vdd.n12490 35.2919
R37352 vdd.n12511 vdd.n12510 35.2919
R37353 vdd.n116 vdd.n107 35.2919
R37354 vdd.n125 vdd.n107 35.2919
R37355 vdd.n126 vdd.n125 35.2919
R37356 vdd.n138 vdd.n126 35.2919
R37357 vdd.n138 vdd.n137 35.2919
R37358 vdd.n137 vdd.n136 35.2919
R37359 vdd.n164 vdd.n155 35.2919
R37360 vdd.n173 vdd.n155 35.2919
R37361 vdd.n174 vdd.n173 35.2919
R37362 vdd.n186 vdd.n174 35.2919
R37363 vdd.n186 vdd.n185 35.2919
R37364 vdd.n185 vdd.n184 35.2919
R37365 vdd.n265 vdd.n256 35.2919
R37366 vdd.n274 vdd.n256 35.2919
R37367 vdd.n275 vdd.n274 35.2919
R37368 vdd.n287 vdd.n275 35.2919
R37369 vdd.n287 vdd.n286 35.2919
R37370 vdd.n286 vdd.n285 35.2919
R37371 vdd.n313 vdd.n304 35.2919
R37372 vdd.n322 vdd.n304 35.2919
R37373 vdd.n323 vdd.n322 35.2919
R37374 vdd.n335 vdd.n323 35.2919
R37375 vdd.n335 vdd.n334 35.2919
R37376 vdd.n334 vdd.n333 35.2919
R37377 vdd.n361 vdd.n352 35.2919
R37378 vdd.n370 vdd.n352 35.2919
R37379 vdd.n371 vdd.n370 35.2919
R37380 vdd.n383 vdd.n371 35.2919
R37381 vdd.n383 vdd.n382 35.2919
R37382 vdd.n382 vdd.n381 35.2919
R37383 vdd.n409 vdd.n400 35.2919
R37384 vdd.n418 vdd.n400 35.2919
R37385 vdd.n419 vdd.n418 35.2919
R37386 vdd.n431 vdd.n419 35.2919
R37387 vdd.n431 vdd.n430 35.2919
R37388 vdd.n430 vdd.n429 35.2919
R37389 vdd.n510 vdd.n501 35.2919
R37390 vdd.n519 vdd.n501 35.2919
R37391 vdd.n520 vdd.n519 35.2919
R37392 vdd.n532 vdd.n520 35.2919
R37393 vdd.n532 vdd.n531 35.2919
R37394 vdd.n531 vdd.n530 35.2919
R37395 vdd.n558 vdd.n549 35.2919
R37396 vdd.n567 vdd.n549 35.2919
R37397 vdd.n568 vdd.n567 35.2919
R37398 vdd.n580 vdd.n568 35.2919
R37399 vdd.n580 vdd.n579 35.2919
R37400 vdd.n579 vdd.n578 35.2919
R37401 vdd.n6982 vdd.n6977 35.2919
R37402 vdd.n6995 vdd.n6977 35.2919
R37403 vdd.n6996 vdd.n6995 35.2919
R37404 vdd.n7008 vdd.n6996 35.2919
R37405 vdd.n7008 vdd.n7007 35.2919
R37406 vdd.n7007 vdd.n7006 35.2919
R37407 vdd.n7030 vdd.n7025 35.2919
R37408 vdd.n7043 vdd.n7025 35.2919
R37409 vdd.n7044 vdd.n7043 35.2919
R37410 vdd.n7056 vdd.n7044 35.2919
R37411 vdd.n7056 vdd.n7055 35.2919
R37412 vdd.n7055 vdd.n7054 35.2919
R37413 vdd.n7132 vdd.n7127 35.2919
R37414 vdd.n7145 vdd.n7127 35.2919
R37415 vdd.n7146 vdd.n7145 35.2919
R37416 vdd.n7158 vdd.n7146 35.2919
R37417 vdd.n7158 vdd.n7157 35.2919
R37418 vdd.n7157 vdd.n7156 35.2919
R37419 vdd.n7180 vdd.n7175 35.2919
R37420 vdd.n7193 vdd.n7175 35.2919
R37421 vdd.n7194 vdd.n7193 35.2919
R37422 vdd.n7206 vdd.n7194 35.2919
R37423 vdd.n7206 vdd.n7205 35.2919
R37424 vdd.n7205 vdd.n7204 35.2919
R37425 vdd.n7228 vdd.n7223 35.2919
R37426 vdd.n7241 vdd.n7223 35.2919
R37427 vdd.n7242 vdd.n7241 35.2919
R37428 vdd.n7254 vdd.n7242 35.2919
R37429 vdd.n7254 vdd.n7253 35.2919
R37430 vdd.n7253 vdd.n7252 35.2919
R37431 vdd.n7276 vdd.n7271 35.2919
R37432 vdd.n7289 vdd.n7271 35.2919
R37433 vdd.n7290 vdd.n7289 35.2919
R37434 vdd.n7302 vdd.n7290 35.2919
R37435 vdd.n7302 vdd.n7301 35.2919
R37436 vdd.n7301 vdd.n7300 35.2919
R37437 vdd.n7378 vdd.n7373 35.2919
R37438 vdd.n7391 vdd.n7373 35.2919
R37439 vdd.n7392 vdd.n7391 35.2919
R37440 vdd.n7404 vdd.n7392 35.2919
R37441 vdd.n7404 vdd.n7403 35.2919
R37442 vdd.n7403 vdd.n7402 35.2919
R37443 vdd.n8898 vdd.n8893 35.2919
R37444 vdd.n8911 vdd.n8893 35.2919
R37445 vdd.n8912 vdd.n8911 35.2919
R37446 vdd.n8924 vdd.n8912 35.2919
R37447 vdd.n8924 vdd.n8923 35.2919
R37448 vdd.n8923 vdd.n8922 35.2919
R37449 vdd.n7430 vdd.n7421 35.2919
R37450 vdd.n7439 vdd.n7421 35.2919
R37451 vdd.n7440 vdd.n7439 35.2919
R37452 vdd.n7452 vdd.n7440 35.2919
R37453 vdd.n7452 vdd.n7451 35.2919
R37454 vdd.n7451 vdd.n7450 35.2919
R37455 vdd.n7478 vdd.n7469 35.2919
R37456 vdd.n7487 vdd.n7469 35.2919
R37457 vdd.n7488 vdd.n7487 35.2919
R37458 vdd.n7500 vdd.n7488 35.2919
R37459 vdd.n7500 vdd.n7499 35.2919
R37460 vdd.n7499 vdd.n7498 35.2919
R37461 vdd.n7579 vdd.n7570 35.2919
R37462 vdd.n7588 vdd.n7570 35.2919
R37463 vdd.n7589 vdd.n7588 35.2919
R37464 vdd.n7601 vdd.n7589 35.2919
R37465 vdd.n7601 vdd.n7600 35.2919
R37466 vdd.n7600 vdd.n7599 35.2919
R37467 vdd.n7627 vdd.n7618 35.2919
R37468 vdd.n7636 vdd.n7618 35.2919
R37469 vdd.n7637 vdd.n7636 35.2919
R37470 vdd.n7649 vdd.n7637 35.2919
R37471 vdd.n7649 vdd.n7648 35.2919
R37472 vdd.n7648 vdd.n7647 35.2919
R37473 vdd.n7675 vdd.n7666 35.2919
R37474 vdd.n7684 vdd.n7666 35.2919
R37475 vdd.n7685 vdd.n7684 35.2919
R37476 vdd.n7697 vdd.n7685 35.2919
R37477 vdd.n7697 vdd.n7696 35.2919
R37478 vdd.n7696 vdd.n7695 35.2919
R37479 vdd.n7723 vdd.n7714 35.2919
R37480 vdd.n7732 vdd.n7714 35.2919
R37481 vdd.n7733 vdd.n7732 35.2919
R37482 vdd.n7745 vdd.n7733 35.2919
R37483 vdd.n7745 vdd.n7744 35.2919
R37484 vdd.n7744 vdd.n7743 35.2919
R37485 vdd.n7824 vdd.n7815 35.2919
R37486 vdd.n7833 vdd.n7815 35.2919
R37487 vdd.n7834 vdd.n7833 35.2919
R37488 vdd.n7846 vdd.n7834 35.2919
R37489 vdd.n7846 vdd.n7845 35.2919
R37490 vdd.n7845 vdd.n7844 35.2919
R37491 vdd.n6937 vdd.n6928 35.2919
R37492 vdd.n6946 vdd.n6928 35.2919
R37493 vdd.n6947 vdd.n6946 35.2919
R37494 vdd.n6959 vdd.n6947 35.2919
R37495 vdd.n6959 vdd.n6958 35.2919
R37496 vdd.n6958 vdd.n6957 35.2919
R37497 vdd.n7872 vdd.n7863 35.2919
R37498 vdd.n7881 vdd.n7863 35.2919
R37499 vdd.n7882 vdd.n7881 35.2919
R37500 vdd.n7894 vdd.n7882 35.2919
R37501 vdd.n7894 vdd.n7893 35.2919
R37502 vdd.n7893 vdd.n7892 35.2919
R37503 vdd.n7919 vdd.n7910 35.2919
R37504 vdd.n7928 vdd.n7910 35.2919
R37505 vdd.n7929 vdd.n7928 35.2919
R37506 vdd.n7941 vdd.n7929 35.2919
R37507 vdd.n7941 vdd.n7940 35.2919
R37508 vdd.n7940 vdd.n7939 35.2919
R37509 vdd.n7969 vdd.n7960 35.2919
R37510 vdd.n7978 vdd.n7960 35.2919
R37511 vdd.n7979 vdd.n7978 35.2919
R37512 vdd.n7991 vdd.n7979 35.2919
R37513 vdd.n7991 vdd.n7990 35.2919
R37514 vdd.n7990 vdd.n7989 35.2919
R37515 vdd.n8019 vdd.n8010 35.2919
R37516 vdd.n8028 vdd.n8010 35.2919
R37517 vdd.n8029 vdd.n8028 35.2919
R37518 vdd.n8041 vdd.n8029 35.2919
R37519 vdd.n8041 vdd.n8040 35.2919
R37520 vdd.n8040 vdd.n8039 35.2919
R37521 vdd.n8067 vdd.n8058 35.2919
R37522 vdd.n8076 vdd.n8058 35.2919
R37523 vdd.n8077 vdd.n8076 35.2919
R37524 vdd.n8089 vdd.n8077 35.2919
R37525 vdd.n8089 vdd.n8088 35.2919
R37526 vdd.n8088 vdd.n8087 35.2919
R37527 vdd.n7795 vdd.n7794 35.2919
R37528 vdd.n7794 vdd.n7793 35.2919
R37529 vdd.n7793 vdd.n7762 35.2919
R37530 vdd.n7781 vdd.n7762 35.2919
R37531 vdd.n7781 vdd.n7780 35.2919
R37532 vdd.n7780 vdd.n7779 35.2919
R37533 vdd.n8118 vdd.n8109 35.2919
R37534 vdd.n8127 vdd.n8109 35.2919
R37535 vdd.n8128 vdd.n8127 35.2919
R37536 vdd.n8140 vdd.n8128 35.2919
R37537 vdd.n8140 vdd.n8139 35.2919
R37538 vdd.n8139 vdd.n8138 35.2919
R37539 vdd.n8165 vdd.n8156 35.2919
R37540 vdd.n8174 vdd.n8156 35.2919
R37541 vdd.n8175 vdd.n8174 35.2919
R37542 vdd.n8187 vdd.n8175 35.2919
R37543 vdd.n8187 vdd.n8186 35.2919
R37544 vdd.n8186 vdd.n8185 35.2919
R37545 vdd.n8213 vdd.n8204 35.2919
R37546 vdd.n8222 vdd.n8204 35.2919
R37547 vdd.n8223 vdd.n8222 35.2919
R37548 vdd.n8235 vdd.n8223 35.2919
R37549 vdd.n8235 vdd.n8234 35.2919
R37550 vdd.n8234 vdd.n8233 35.2919
R37551 vdd.n8264 vdd.n8255 35.2919
R37552 vdd.n8273 vdd.n8255 35.2919
R37553 vdd.n8274 vdd.n8273 35.2919
R37554 vdd.n8286 vdd.n8274 35.2919
R37555 vdd.n8286 vdd.n8285 35.2919
R37556 vdd.n8285 vdd.n8284 35.2919
R37557 vdd.n8314 vdd.n8305 35.2919
R37558 vdd.n8323 vdd.n8305 35.2919
R37559 vdd.n8324 vdd.n8323 35.2919
R37560 vdd.n8336 vdd.n8324 35.2919
R37561 vdd.n8336 vdd.n8335 35.2919
R37562 vdd.n8335 vdd.n8334 35.2919
R37563 vdd.n8362 vdd.n8353 35.2919
R37564 vdd.n8371 vdd.n8353 35.2919
R37565 vdd.n8372 vdd.n8371 35.2919
R37566 vdd.n8384 vdd.n8372 35.2919
R37567 vdd.n8384 vdd.n8383 35.2919
R37568 vdd.n8383 vdd.n8382 35.2919
R37569 vdd.n8412 vdd.n8403 35.2919
R37570 vdd.n8421 vdd.n8403 35.2919
R37571 vdd.n8422 vdd.n8421 35.2919
R37572 vdd.n8434 vdd.n8422 35.2919
R37573 vdd.n8434 vdd.n8433 35.2919
R37574 vdd.n8433 vdd.n8432 35.2919
R37575 vdd.n8459 vdd.n8450 35.2919
R37576 vdd.n8468 vdd.n8450 35.2919
R37577 vdd.n8469 vdd.n8468 35.2919
R37578 vdd.n8481 vdd.n8469 35.2919
R37579 vdd.n8481 vdd.n8480 35.2919
R37580 vdd.n8480 vdd.n8479 35.2919
R37581 vdd.n8509 vdd.n8500 35.2919
R37582 vdd.n8518 vdd.n8500 35.2919
R37583 vdd.n8519 vdd.n8518 35.2919
R37584 vdd.n8531 vdd.n8519 35.2919
R37585 vdd.n8531 vdd.n8530 35.2919
R37586 vdd.n8530 vdd.n8529 35.2919
R37587 vdd.n8559 vdd.n8550 35.2919
R37588 vdd.n8568 vdd.n8550 35.2919
R37589 vdd.n8569 vdd.n8568 35.2919
R37590 vdd.n8581 vdd.n8569 35.2919
R37591 vdd.n8581 vdd.n8580 35.2919
R37592 vdd.n8580 vdd.n8579 35.2919
R37593 vdd.n8607 vdd.n8598 35.2919
R37594 vdd.n8616 vdd.n8598 35.2919
R37595 vdd.n8617 vdd.n8616 35.2919
R37596 vdd.n8629 vdd.n8617 35.2919
R37597 vdd.n8629 vdd.n8628 35.2919
R37598 vdd.n8628 vdd.n8627 35.2919
R37599 vdd.n7550 vdd.n7549 35.2919
R37600 vdd.n7549 vdd.n7548 35.2919
R37601 vdd.n7548 vdd.n7517 35.2919
R37602 vdd.n7536 vdd.n7517 35.2919
R37603 vdd.n7536 vdd.n7535 35.2919
R37604 vdd.n7535 vdd.n7534 35.2919
R37605 vdd.n8658 vdd.n8649 35.2919
R37606 vdd.n8667 vdd.n8649 35.2919
R37607 vdd.n8668 vdd.n8667 35.2919
R37608 vdd.n8680 vdd.n8668 35.2919
R37609 vdd.n8680 vdd.n8679 35.2919
R37610 vdd.n8679 vdd.n8678 35.2919
R37611 vdd.n8705 vdd.n8696 35.2919
R37612 vdd.n8714 vdd.n8696 35.2919
R37613 vdd.n8715 vdd.n8714 35.2919
R37614 vdd.n8727 vdd.n8715 35.2919
R37615 vdd.n8727 vdd.n8726 35.2919
R37616 vdd.n8726 vdd.n8725 35.2919
R37617 vdd.n8755 vdd.n8746 35.2919
R37618 vdd.n8764 vdd.n8746 35.2919
R37619 vdd.n8765 vdd.n8764 35.2919
R37620 vdd.n8777 vdd.n8765 35.2919
R37621 vdd.n8777 vdd.n8776 35.2919
R37622 vdd.n8776 vdd.n8775 35.2919
R37623 vdd.n8805 vdd.n8796 35.2919
R37624 vdd.n8814 vdd.n8796 35.2919
R37625 vdd.n8815 vdd.n8814 35.2919
R37626 vdd.n8827 vdd.n8815 35.2919
R37627 vdd.n8827 vdd.n8826 35.2919
R37628 vdd.n8826 vdd.n8825 35.2919
R37629 vdd.n8853 vdd.n8844 35.2919
R37630 vdd.n8862 vdd.n8844 35.2919
R37631 vdd.n8863 vdd.n8862 35.2919
R37632 vdd.n8875 vdd.n8863 35.2919
R37633 vdd.n8875 vdd.n8874 35.2919
R37634 vdd.n8874 vdd.n8873 35.2919
R37635 vdd.n8995 vdd.n8990 35.2919
R37636 vdd.n9008 vdd.n8990 35.2919
R37637 vdd.n9009 vdd.n9008 35.2919
R37638 vdd.n9021 vdd.n9009 35.2919
R37639 vdd.n9021 vdd.n9020 35.2919
R37640 vdd.n9020 vdd.n9019 35.2919
R37641 vdd.n8947 vdd.n8942 35.2919
R37642 vdd.n8960 vdd.n8942 35.2919
R37643 vdd.n8961 vdd.n8960 35.2919
R37644 vdd.n8973 vdd.n8961 35.2919
R37645 vdd.n8973 vdd.n8972 35.2919
R37646 vdd.n8972 vdd.n8971 35.2919
R37647 vdd.n9044 vdd.n9039 35.2919
R37648 vdd.n9057 vdd.n9039 35.2919
R37649 vdd.n9058 vdd.n9057 35.2919
R37650 vdd.n9070 vdd.n9058 35.2919
R37651 vdd.n9070 vdd.n9069 35.2919
R37652 vdd.n9069 vdd.n9068 35.2919
R37653 vdd.n9094 vdd.n9089 35.2919
R37654 vdd.n9107 vdd.n9089 35.2919
R37655 vdd.n9108 vdd.n9107 35.2919
R37656 vdd.n9120 vdd.n9108 35.2919
R37657 vdd.n9120 vdd.n9119 35.2919
R37658 vdd.n9119 vdd.n9118 35.2919
R37659 vdd.n9142 vdd.n9137 35.2919
R37660 vdd.n9155 vdd.n9137 35.2919
R37661 vdd.n9156 vdd.n9155 35.2919
R37662 vdd.n9168 vdd.n9156 35.2919
R37663 vdd.n9168 vdd.n9167 35.2919
R37664 vdd.n9167 vdd.n9166 35.2919
R37665 vdd.n7330 vdd.n7329 35.2919
R37666 vdd.n7329 vdd.n7328 35.2919
R37667 vdd.n7328 vdd.n7317 35.2919
R37668 vdd.n7340 vdd.n7317 35.2919
R37669 vdd.n7340 vdd.n7313 35.2919
R37670 vdd.n7356 vdd.n7313 35.2919
R37671 vdd.n9290 vdd.n9285 35.2919
R37672 vdd.n9303 vdd.n9285 35.2919
R37673 vdd.n9304 vdd.n9303 35.2919
R37674 vdd.n9316 vdd.n9304 35.2919
R37675 vdd.n9316 vdd.n9315 35.2919
R37676 vdd.n9315 vdd.n9314 35.2919
R37677 vdd.n9241 vdd.n9236 35.2919
R37678 vdd.n9254 vdd.n9236 35.2919
R37679 vdd.n9255 vdd.n9254 35.2919
R37680 vdd.n9267 vdd.n9255 35.2919
R37681 vdd.n9267 vdd.n9266 35.2919
R37682 vdd.n9266 vdd.n9265 35.2919
R37683 vdd.n9193 vdd.n9188 35.2919
R37684 vdd.n9206 vdd.n9188 35.2919
R37685 vdd.n9207 vdd.n9206 35.2919
R37686 vdd.n9219 vdd.n9207 35.2919
R37687 vdd.n9219 vdd.n9218 35.2919
R37688 vdd.n9218 vdd.n9217 35.2919
R37689 vdd.n9339 vdd.n9334 35.2919
R37690 vdd.n9352 vdd.n9334 35.2919
R37691 vdd.n9353 vdd.n9352 35.2919
R37692 vdd.n9365 vdd.n9353 35.2919
R37693 vdd.n9365 vdd.n9364 35.2919
R37694 vdd.n9364 vdd.n9363 35.2919
R37695 vdd.n9389 vdd.n9384 35.2919
R37696 vdd.n9402 vdd.n9384 35.2919
R37697 vdd.n9403 vdd.n9402 35.2919
R37698 vdd.n9415 vdd.n9403 35.2919
R37699 vdd.n9415 vdd.n9414 35.2919
R37700 vdd.n9414 vdd.n9413 35.2919
R37701 vdd.n9437 vdd.n9432 35.2919
R37702 vdd.n9450 vdd.n9432 35.2919
R37703 vdd.n9451 vdd.n9450 35.2919
R37704 vdd.n9463 vdd.n9451 35.2919
R37705 vdd.n9463 vdd.n9462 35.2919
R37706 vdd.n9462 vdd.n9461 35.2919
R37707 vdd.n9535 vdd.n9530 35.2919
R37708 vdd.n9548 vdd.n9530 35.2919
R37709 vdd.n9549 vdd.n9548 35.2919
R37710 vdd.n9561 vdd.n9549 35.2919
R37711 vdd.n9561 vdd.n9560 35.2919
R37712 vdd.n9560 vdd.n9559 35.2919
R37713 vdd.n9487 vdd.n9482 35.2919
R37714 vdd.n9500 vdd.n9482 35.2919
R37715 vdd.n9501 vdd.n9500 35.2919
R37716 vdd.n9513 vdd.n9501 35.2919
R37717 vdd.n9513 vdd.n9512 35.2919
R37718 vdd.n9512 vdd.n9511 35.2919
R37719 vdd.n9584 vdd.n9579 35.2919
R37720 vdd.n9597 vdd.n9579 35.2919
R37721 vdd.n9598 vdd.n9597 35.2919
R37722 vdd.n9610 vdd.n9598 35.2919
R37723 vdd.n9610 vdd.n9609 35.2919
R37724 vdd.n9609 vdd.n9608 35.2919
R37725 vdd.n9634 vdd.n9629 35.2919
R37726 vdd.n9647 vdd.n9629 35.2919
R37727 vdd.n9648 vdd.n9647 35.2919
R37728 vdd.n9660 vdd.n9648 35.2919
R37729 vdd.n9660 vdd.n9659 35.2919
R37730 vdd.n9659 vdd.n9658 35.2919
R37731 vdd.n9682 vdd.n9677 35.2919
R37732 vdd.n9695 vdd.n9677 35.2919
R37733 vdd.n9696 vdd.n9695 35.2919
R37734 vdd.n9708 vdd.n9696 35.2919
R37735 vdd.n9708 vdd.n9707 35.2919
R37736 vdd.n9707 vdd.n9706 35.2919
R37737 vdd.n7084 vdd.n7083 35.2919
R37738 vdd.n7083 vdd.n7082 35.2919
R37739 vdd.n7082 vdd.n7071 35.2919
R37740 vdd.n7094 vdd.n7071 35.2919
R37741 vdd.n7094 vdd.n7067 35.2919
R37742 vdd.n7110 vdd.n7067 35.2919
R37743 vdd.n9781 vdd.n9776 35.2919
R37744 vdd.n9794 vdd.n9776 35.2919
R37745 vdd.n9795 vdd.n9794 35.2919
R37746 vdd.n9807 vdd.n9795 35.2919
R37747 vdd.n9807 vdd.n9806 35.2919
R37748 vdd.n9806 vdd.n9805 35.2919
R37749 vdd.n9733 vdd.n9728 35.2919
R37750 vdd.n9746 vdd.n9728 35.2919
R37751 vdd.n9747 vdd.n9746 35.2919
R37752 vdd.n9759 vdd.n9747 35.2919
R37753 vdd.n9759 vdd.n9758 35.2919
R37754 vdd.n9758 vdd.n9757 35.2919
R37755 vdd.n9830 vdd.n9825 35.2919
R37756 vdd.n9843 vdd.n9825 35.2919
R37757 vdd.n9844 vdd.n9843 35.2919
R37758 vdd.n9856 vdd.n9844 35.2919
R37759 vdd.n9856 vdd.n9855 35.2919
R37760 vdd.n9855 vdd.n9854 35.2919
R37761 vdd.n9880 vdd.n9875 35.2919
R37762 vdd.n9893 vdd.n9875 35.2919
R37763 vdd.n9894 vdd.n9893 35.2919
R37764 vdd.n9906 vdd.n9894 35.2919
R37765 vdd.n9906 vdd.n9905 35.2919
R37766 vdd.n9905 vdd.n9904 35.2919
R37767 vdd.n9928 vdd.n9923 35.2919
R37768 vdd.n9941 vdd.n9923 35.2919
R37769 vdd.n9942 vdd.n9941 35.2919
R37770 vdd.n9954 vdd.n9942 35.2919
R37771 vdd.n9954 vdd.n9953 35.2919
R37772 vdd.n9953 vdd.n9952 35.2919
R37773 vdd.n3840 vdd.n3835 35.2919
R37774 vdd.n3853 vdd.n3835 35.2919
R37775 vdd.n3854 vdd.n3853 35.2919
R37776 vdd.n3866 vdd.n3854 35.2919
R37777 vdd.n3866 vdd.n3865 35.2919
R37778 vdd.n3865 vdd.n3864 35.2919
R37779 vdd.n3888 vdd.n3883 35.2919
R37780 vdd.n3901 vdd.n3883 35.2919
R37781 vdd.n3902 vdd.n3901 35.2919
R37782 vdd.n3914 vdd.n3902 35.2919
R37783 vdd.n3914 vdd.n3913 35.2919
R37784 vdd.n3913 vdd.n3912 35.2919
R37785 vdd.n3990 vdd.n3985 35.2919
R37786 vdd.n4003 vdd.n3985 35.2919
R37787 vdd.n4004 vdd.n4003 35.2919
R37788 vdd.n4016 vdd.n4004 35.2919
R37789 vdd.n4016 vdd.n4015 35.2919
R37790 vdd.n4015 vdd.n4014 35.2919
R37791 vdd.n4038 vdd.n4033 35.2919
R37792 vdd.n4051 vdd.n4033 35.2919
R37793 vdd.n4052 vdd.n4051 35.2919
R37794 vdd.n4064 vdd.n4052 35.2919
R37795 vdd.n4064 vdd.n4063 35.2919
R37796 vdd.n4063 vdd.n4062 35.2919
R37797 vdd.n4086 vdd.n4081 35.2919
R37798 vdd.n4099 vdd.n4081 35.2919
R37799 vdd.n4100 vdd.n4099 35.2919
R37800 vdd.n4112 vdd.n4100 35.2919
R37801 vdd.n4112 vdd.n4111 35.2919
R37802 vdd.n4111 vdd.n4110 35.2919
R37803 vdd.n4134 vdd.n4129 35.2919
R37804 vdd.n4147 vdd.n4129 35.2919
R37805 vdd.n4148 vdd.n4147 35.2919
R37806 vdd.n4160 vdd.n4148 35.2919
R37807 vdd.n4160 vdd.n4159 35.2919
R37808 vdd.n4159 vdd.n4158 35.2919
R37809 vdd.n4236 vdd.n4231 35.2919
R37810 vdd.n4249 vdd.n4231 35.2919
R37811 vdd.n4250 vdd.n4249 35.2919
R37812 vdd.n4262 vdd.n4250 35.2919
R37813 vdd.n4262 vdd.n4261 35.2919
R37814 vdd.n4261 vdd.n4260 35.2919
R37815 vdd.n5756 vdd.n5751 35.2919
R37816 vdd.n5769 vdd.n5751 35.2919
R37817 vdd.n5770 vdd.n5769 35.2919
R37818 vdd.n5782 vdd.n5770 35.2919
R37819 vdd.n5782 vdd.n5781 35.2919
R37820 vdd.n5781 vdd.n5780 35.2919
R37821 vdd.n4288 vdd.n4279 35.2919
R37822 vdd.n4297 vdd.n4279 35.2919
R37823 vdd.n4298 vdd.n4297 35.2919
R37824 vdd.n4310 vdd.n4298 35.2919
R37825 vdd.n4310 vdd.n4309 35.2919
R37826 vdd.n4309 vdd.n4308 35.2919
R37827 vdd.n4336 vdd.n4327 35.2919
R37828 vdd.n4345 vdd.n4327 35.2919
R37829 vdd.n4346 vdd.n4345 35.2919
R37830 vdd.n4358 vdd.n4346 35.2919
R37831 vdd.n4358 vdd.n4357 35.2919
R37832 vdd.n4357 vdd.n4356 35.2919
R37833 vdd.n4437 vdd.n4428 35.2919
R37834 vdd.n4446 vdd.n4428 35.2919
R37835 vdd.n4447 vdd.n4446 35.2919
R37836 vdd.n4459 vdd.n4447 35.2919
R37837 vdd.n4459 vdd.n4458 35.2919
R37838 vdd.n4458 vdd.n4457 35.2919
R37839 vdd.n4485 vdd.n4476 35.2919
R37840 vdd.n4494 vdd.n4476 35.2919
R37841 vdd.n4495 vdd.n4494 35.2919
R37842 vdd.n4507 vdd.n4495 35.2919
R37843 vdd.n4507 vdd.n4506 35.2919
R37844 vdd.n4506 vdd.n4505 35.2919
R37845 vdd.n4533 vdd.n4524 35.2919
R37846 vdd.n4542 vdd.n4524 35.2919
R37847 vdd.n4543 vdd.n4542 35.2919
R37848 vdd.n4555 vdd.n4543 35.2919
R37849 vdd.n4555 vdd.n4554 35.2919
R37850 vdd.n4554 vdd.n4553 35.2919
R37851 vdd.n4581 vdd.n4572 35.2919
R37852 vdd.n4590 vdd.n4572 35.2919
R37853 vdd.n4591 vdd.n4590 35.2919
R37854 vdd.n4603 vdd.n4591 35.2919
R37855 vdd.n4603 vdd.n4602 35.2919
R37856 vdd.n4602 vdd.n4601 35.2919
R37857 vdd.n4682 vdd.n4673 35.2919
R37858 vdd.n4691 vdd.n4673 35.2919
R37859 vdd.n4692 vdd.n4691 35.2919
R37860 vdd.n4704 vdd.n4692 35.2919
R37861 vdd.n4704 vdd.n4703 35.2919
R37862 vdd.n4703 vdd.n4702 35.2919
R37863 vdd.n3795 vdd.n3786 35.2919
R37864 vdd.n3804 vdd.n3786 35.2919
R37865 vdd.n3805 vdd.n3804 35.2919
R37866 vdd.n3817 vdd.n3805 35.2919
R37867 vdd.n3817 vdd.n3816 35.2919
R37868 vdd.n3816 vdd.n3815 35.2919
R37869 vdd.n4730 vdd.n4721 35.2919
R37870 vdd.n4739 vdd.n4721 35.2919
R37871 vdd.n4740 vdd.n4739 35.2919
R37872 vdd.n4752 vdd.n4740 35.2919
R37873 vdd.n4752 vdd.n4751 35.2919
R37874 vdd.n4751 vdd.n4750 35.2919
R37875 vdd.n4777 vdd.n4768 35.2919
R37876 vdd.n4786 vdd.n4768 35.2919
R37877 vdd.n4787 vdd.n4786 35.2919
R37878 vdd.n4799 vdd.n4787 35.2919
R37879 vdd.n4799 vdd.n4798 35.2919
R37880 vdd.n4798 vdd.n4797 35.2919
R37881 vdd.n4827 vdd.n4818 35.2919
R37882 vdd.n4836 vdd.n4818 35.2919
R37883 vdd.n4837 vdd.n4836 35.2919
R37884 vdd.n4849 vdd.n4837 35.2919
R37885 vdd.n4849 vdd.n4848 35.2919
R37886 vdd.n4848 vdd.n4847 35.2919
R37887 vdd.n4877 vdd.n4868 35.2919
R37888 vdd.n4886 vdd.n4868 35.2919
R37889 vdd.n4887 vdd.n4886 35.2919
R37890 vdd.n4899 vdd.n4887 35.2919
R37891 vdd.n4899 vdd.n4898 35.2919
R37892 vdd.n4898 vdd.n4897 35.2919
R37893 vdd.n4925 vdd.n4916 35.2919
R37894 vdd.n4934 vdd.n4916 35.2919
R37895 vdd.n4935 vdd.n4934 35.2919
R37896 vdd.n4947 vdd.n4935 35.2919
R37897 vdd.n4947 vdd.n4946 35.2919
R37898 vdd.n4946 vdd.n4945 35.2919
R37899 vdd.n4653 vdd.n4652 35.2919
R37900 vdd.n4652 vdd.n4651 35.2919
R37901 vdd.n4651 vdd.n4620 35.2919
R37902 vdd.n4639 vdd.n4620 35.2919
R37903 vdd.n4639 vdd.n4638 35.2919
R37904 vdd.n4638 vdd.n4637 35.2919
R37905 vdd.n4976 vdd.n4967 35.2919
R37906 vdd.n4985 vdd.n4967 35.2919
R37907 vdd.n4986 vdd.n4985 35.2919
R37908 vdd.n4998 vdd.n4986 35.2919
R37909 vdd.n4998 vdd.n4997 35.2919
R37910 vdd.n4997 vdd.n4996 35.2919
R37911 vdd.n5023 vdd.n5014 35.2919
R37912 vdd.n5032 vdd.n5014 35.2919
R37913 vdd.n5033 vdd.n5032 35.2919
R37914 vdd.n5045 vdd.n5033 35.2919
R37915 vdd.n5045 vdd.n5044 35.2919
R37916 vdd.n5044 vdd.n5043 35.2919
R37917 vdd.n5071 vdd.n5062 35.2919
R37918 vdd.n5080 vdd.n5062 35.2919
R37919 vdd.n5081 vdd.n5080 35.2919
R37920 vdd.n5093 vdd.n5081 35.2919
R37921 vdd.n5093 vdd.n5092 35.2919
R37922 vdd.n5092 vdd.n5091 35.2919
R37923 vdd.n5122 vdd.n5113 35.2919
R37924 vdd.n5131 vdd.n5113 35.2919
R37925 vdd.n5132 vdd.n5131 35.2919
R37926 vdd.n5144 vdd.n5132 35.2919
R37927 vdd.n5144 vdd.n5143 35.2919
R37928 vdd.n5143 vdd.n5142 35.2919
R37929 vdd.n5172 vdd.n5163 35.2919
R37930 vdd.n5181 vdd.n5163 35.2919
R37931 vdd.n5182 vdd.n5181 35.2919
R37932 vdd.n5194 vdd.n5182 35.2919
R37933 vdd.n5194 vdd.n5193 35.2919
R37934 vdd.n5193 vdd.n5192 35.2919
R37935 vdd.n5220 vdd.n5211 35.2919
R37936 vdd.n5229 vdd.n5211 35.2919
R37937 vdd.n5230 vdd.n5229 35.2919
R37938 vdd.n5242 vdd.n5230 35.2919
R37939 vdd.n5242 vdd.n5241 35.2919
R37940 vdd.n5241 vdd.n5240 35.2919
R37941 vdd.n5270 vdd.n5261 35.2919
R37942 vdd.n5279 vdd.n5261 35.2919
R37943 vdd.n5280 vdd.n5279 35.2919
R37944 vdd.n5292 vdd.n5280 35.2919
R37945 vdd.n5292 vdd.n5291 35.2919
R37946 vdd.n5291 vdd.n5290 35.2919
R37947 vdd.n5317 vdd.n5308 35.2919
R37948 vdd.n5326 vdd.n5308 35.2919
R37949 vdd.n5327 vdd.n5326 35.2919
R37950 vdd.n5339 vdd.n5327 35.2919
R37951 vdd.n5339 vdd.n5338 35.2919
R37952 vdd.n5338 vdd.n5337 35.2919
R37953 vdd.n5367 vdd.n5358 35.2919
R37954 vdd.n5376 vdd.n5358 35.2919
R37955 vdd.n5377 vdd.n5376 35.2919
R37956 vdd.n5389 vdd.n5377 35.2919
R37957 vdd.n5389 vdd.n5388 35.2919
R37958 vdd.n5388 vdd.n5387 35.2919
R37959 vdd.n5417 vdd.n5408 35.2919
R37960 vdd.n5426 vdd.n5408 35.2919
R37961 vdd.n5427 vdd.n5426 35.2919
R37962 vdd.n5439 vdd.n5427 35.2919
R37963 vdd.n5439 vdd.n5438 35.2919
R37964 vdd.n5438 vdd.n5437 35.2919
R37965 vdd.n5465 vdd.n5456 35.2919
R37966 vdd.n5474 vdd.n5456 35.2919
R37967 vdd.n5475 vdd.n5474 35.2919
R37968 vdd.n5487 vdd.n5475 35.2919
R37969 vdd.n5487 vdd.n5486 35.2919
R37970 vdd.n5486 vdd.n5485 35.2919
R37971 vdd.n4408 vdd.n4407 35.2919
R37972 vdd.n4407 vdd.n4406 35.2919
R37973 vdd.n4406 vdd.n4375 35.2919
R37974 vdd.n4394 vdd.n4375 35.2919
R37975 vdd.n4394 vdd.n4393 35.2919
R37976 vdd.n4393 vdd.n4392 35.2919
R37977 vdd.n5516 vdd.n5507 35.2919
R37978 vdd.n5525 vdd.n5507 35.2919
R37979 vdd.n5526 vdd.n5525 35.2919
R37980 vdd.n5538 vdd.n5526 35.2919
R37981 vdd.n5538 vdd.n5537 35.2919
R37982 vdd.n5537 vdd.n5536 35.2919
R37983 vdd.n5563 vdd.n5554 35.2919
R37984 vdd.n5572 vdd.n5554 35.2919
R37985 vdd.n5573 vdd.n5572 35.2919
R37986 vdd.n5585 vdd.n5573 35.2919
R37987 vdd.n5585 vdd.n5584 35.2919
R37988 vdd.n5584 vdd.n5583 35.2919
R37989 vdd.n5613 vdd.n5604 35.2919
R37990 vdd.n5622 vdd.n5604 35.2919
R37991 vdd.n5623 vdd.n5622 35.2919
R37992 vdd.n5635 vdd.n5623 35.2919
R37993 vdd.n5635 vdd.n5634 35.2919
R37994 vdd.n5634 vdd.n5633 35.2919
R37995 vdd.n5663 vdd.n5654 35.2919
R37996 vdd.n5672 vdd.n5654 35.2919
R37997 vdd.n5673 vdd.n5672 35.2919
R37998 vdd.n5685 vdd.n5673 35.2919
R37999 vdd.n5685 vdd.n5684 35.2919
R38000 vdd.n5684 vdd.n5683 35.2919
R38001 vdd.n5711 vdd.n5702 35.2919
R38002 vdd.n5720 vdd.n5702 35.2919
R38003 vdd.n5721 vdd.n5720 35.2919
R38004 vdd.n5733 vdd.n5721 35.2919
R38005 vdd.n5733 vdd.n5732 35.2919
R38006 vdd.n5732 vdd.n5731 35.2919
R38007 vdd.n5853 vdd.n5848 35.2919
R38008 vdd.n5866 vdd.n5848 35.2919
R38009 vdd.n5867 vdd.n5866 35.2919
R38010 vdd.n5879 vdd.n5867 35.2919
R38011 vdd.n5879 vdd.n5878 35.2919
R38012 vdd.n5878 vdd.n5877 35.2919
R38013 vdd.n5805 vdd.n5800 35.2919
R38014 vdd.n5818 vdd.n5800 35.2919
R38015 vdd.n5819 vdd.n5818 35.2919
R38016 vdd.n5831 vdd.n5819 35.2919
R38017 vdd.n5831 vdd.n5830 35.2919
R38018 vdd.n5830 vdd.n5829 35.2919
R38019 vdd.n5902 vdd.n5897 35.2919
R38020 vdd.n5915 vdd.n5897 35.2919
R38021 vdd.n5916 vdd.n5915 35.2919
R38022 vdd.n5928 vdd.n5916 35.2919
R38023 vdd.n5928 vdd.n5927 35.2919
R38024 vdd.n5927 vdd.n5926 35.2919
R38025 vdd.n5952 vdd.n5947 35.2919
R38026 vdd.n5965 vdd.n5947 35.2919
R38027 vdd.n5966 vdd.n5965 35.2919
R38028 vdd.n5978 vdd.n5966 35.2919
R38029 vdd.n5978 vdd.n5977 35.2919
R38030 vdd.n5977 vdd.n5976 35.2919
R38031 vdd.n6000 vdd.n5995 35.2919
R38032 vdd.n6013 vdd.n5995 35.2919
R38033 vdd.n6014 vdd.n6013 35.2919
R38034 vdd.n6026 vdd.n6014 35.2919
R38035 vdd.n6026 vdd.n6025 35.2919
R38036 vdd.n6025 vdd.n6024 35.2919
R38037 vdd.n4188 vdd.n4187 35.2919
R38038 vdd.n4187 vdd.n4186 35.2919
R38039 vdd.n4186 vdd.n4175 35.2919
R38040 vdd.n4198 vdd.n4175 35.2919
R38041 vdd.n4198 vdd.n4171 35.2919
R38042 vdd.n4214 vdd.n4171 35.2919
R38043 vdd.n6148 vdd.n6143 35.2919
R38044 vdd.n6161 vdd.n6143 35.2919
R38045 vdd.n6162 vdd.n6161 35.2919
R38046 vdd.n6174 vdd.n6162 35.2919
R38047 vdd.n6174 vdd.n6173 35.2919
R38048 vdd.n6173 vdd.n6172 35.2919
R38049 vdd.n6099 vdd.n6094 35.2919
R38050 vdd.n6112 vdd.n6094 35.2919
R38051 vdd.n6113 vdd.n6112 35.2919
R38052 vdd.n6125 vdd.n6113 35.2919
R38053 vdd.n6125 vdd.n6124 35.2919
R38054 vdd.n6124 vdd.n6123 35.2919
R38055 vdd.n6051 vdd.n6046 35.2919
R38056 vdd.n6064 vdd.n6046 35.2919
R38057 vdd.n6065 vdd.n6064 35.2919
R38058 vdd.n6077 vdd.n6065 35.2919
R38059 vdd.n6077 vdd.n6076 35.2919
R38060 vdd.n6076 vdd.n6075 35.2919
R38061 vdd.n6197 vdd.n6192 35.2919
R38062 vdd.n6210 vdd.n6192 35.2919
R38063 vdd.n6211 vdd.n6210 35.2919
R38064 vdd.n6223 vdd.n6211 35.2919
R38065 vdd.n6223 vdd.n6222 35.2919
R38066 vdd.n6222 vdd.n6221 35.2919
R38067 vdd.n6247 vdd.n6242 35.2919
R38068 vdd.n6260 vdd.n6242 35.2919
R38069 vdd.n6261 vdd.n6260 35.2919
R38070 vdd.n6273 vdd.n6261 35.2919
R38071 vdd.n6273 vdd.n6272 35.2919
R38072 vdd.n6272 vdd.n6271 35.2919
R38073 vdd.n6295 vdd.n6290 35.2919
R38074 vdd.n6308 vdd.n6290 35.2919
R38075 vdd.n6309 vdd.n6308 35.2919
R38076 vdd.n6321 vdd.n6309 35.2919
R38077 vdd.n6321 vdd.n6320 35.2919
R38078 vdd.n6320 vdd.n6319 35.2919
R38079 vdd.n6393 vdd.n6388 35.2919
R38080 vdd.n6406 vdd.n6388 35.2919
R38081 vdd.n6407 vdd.n6406 35.2919
R38082 vdd.n6419 vdd.n6407 35.2919
R38083 vdd.n6419 vdd.n6418 35.2919
R38084 vdd.n6418 vdd.n6417 35.2919
R38085 vdd.n6345 vdd.n6340 35.2919
R38086 vdd.n6358 vdd.n6340 35.2919
R38087 vdd.n6359 vdd.n6358 35.2919
R38088 vdd.n6371 vdd.n6359 35.2919
R38089 vdd.n6371 vdd.n6370 35.2919
R38090 vdd.n6370 vdd.n6369 35.2919
R38091 vdd.n6442 vdd.n6437 35.2919
R38092 vdd.n6455 vdd.n6437 35.2919
R38093 vdd.n6456 vdd.n6455 35.2919
R38094 vdd.n6468 vdd.n6456 35.2919
R38095 vdd.n6468 vdd.n6467 35.2919
R38096 vdd.n6467 vdd.n6466 35.2919
R38097 vdd.n6492 vdd.n6487 35.2919
R38098 vdd.n6505 vdd.n6487 35.2919
R38099 vdd.n6506 vdd.n6505 35.2919
R38100 vdd.n6518 vdd.n6506 35.2919
R38101 vdd.n6518 vdd.n6517 35.2919
R38102 vdd.n6517 vdd.n6516 35.2919
R38103 vdd.n6540 vdd.n6535 35.2919
R38104 vdd.n6553 vdd.n6535 35.2919
R38105 vdd.n6554 vdd.n6553 35.2919
R38106 vdd.n6566 vdd.n6554 35.2919
R38107 vdd.n6566 vdd.n6565 35.2919
R38108 vdd.n6565 vdd.n6564 35.2919
R38109 vdd.n3942 vdd.n3941 35.2919
R38110 vdd.n3941 vdd.n3940 35.2919
R38111 vdd.n3940 vdd.n3929 35.2919
R38112 vdd.n3952 vdd.n3929 35.2919
R38113 vdd.n3952 vdd.n3925 35.2919
R38114 vdd.n3968 vdd.n3925 35.2919
R38115 vdd.n6639 vdd.n6634 35.2919
R38116 vdd.n6652 vdd.n6634 35.2919
R38117 vdd.n6653 vdd.n6652 35.2919
R38118 vdd.n6665 vdd.n6653 35.2919
R38119 vdd.n6665 vdd.n6664 35.2919
R38120 vdd.n6664 vdd.n6663 35.2919
R38121 vdd.n6591 vdd.n6586 35.2919
R38122 vdd.n6604 vdd.n6586 35.2919
R38123 vdd.n6605 vdd.n6604 35.2919
R38124 vdd.n6617 vdd.n6605 35.2919
R38125 vdd.n6617 vdd.n6616 35.2919
R38126 vdd.n6616 vdd.n6615 35.2919
R38127 vdd.n6688 vdd.n6683 35.2919
R38128 vdd.n6701 vdd.n6683 35.2919
R38129 vdd.n6702 vdd.n6701 35.2919
R38130 vdd.n6714 vdd.n6702 35.2919
R38131 vdd.n6714 vdd.n6713 35.2919
R38132 vdd.n6713 vdd.n6712 35.2919
R38133 vdd.n6738 vdd.n6733 35.2919
R38134 vdd.n6751 vdd.n6733 35.2919
R38135 vdd.n6752 vdd.n6751 35.2919
R38136 vdd.n6764 vdd.n6752 35.2919
R38137 vdd.n6764 vdd.n6763 35.2919
R38138 vdd.n6763 vdd.n6762 35.2919
R38139 vdd.n6786 vdd.n6781 35.2919
R38140 vdd.n6799 vdd.n6781 35.2919
R38141 vdd.n6800 vdd.n6799 35.2919
R38142 vdd.n6812 vdd.n6800 35.2919
R38143 vdd.n6812 vdd.n6811 35.2919
R38144 vdd.n6811 vdd.n6810 35.2919
R38145 vdd.n698 vdd.n693 35.2919
R38146 vdd.n711 vdd.n693 35.2919
R38147 vdd.n712 vdd.n711 35.2919
R38148 vdd.n724 vdd.n712 35.2919
R38149 vdd.n724 vdd.n723 35.2919
R38150 vdd.n723 vdd.n722 35.2919
R38151 vdd.n746 vdd.n741 35.2919
R38152 vdd.n759 vdd.n741 35.2919
R38153 vdd.n760 vdd.n759 35.2919
R38154 vdd.n772 vdd.n760 35.2919
R38155 vdd.n772 vdd.n771 35.2919
R38156 vdd.n771 vdd.n770 35.2919
R38157 vdd.n848 vdd.n843 35.2919
R38158 vdd.n861 vdd.n843 35.2919
R38159 vdd.n862 vdd.n861 35.2919
R38160 vdd.n874 vdd.n862 35.2919
R38161 vdd.n874 vdd.n873 35.2919
R38162 vdd.n873 vdd.n872 35.2919
R38163 vdd.n896 vdd.n891 35.2919
R38164 vdd.n909 vdd.n891 35.2919
R38165 vdd.n910 vdd.n909 35.2919
R38166 vdd.n922 vdd.n910 35.2919
R38167 vdd.n922 vdd.n921 35.2919
R38168 vdd.n921 vdd.n920 35.2919
R38169 vdd.n944 vdd.n939 35.2919
R38170 vdd.n957 vdd.n939 35.2919
R38171 vdd.n958 vdd.n957 35.2919
R38172 vdd.n970 vdd.n958 35.2919
R38173 vdd.n970 vdd.n969 35.2919
R38174 vdd.n969 vdd.n968 35.2919
R38175 vdd.n992 vdd.n987 35.2919
R38176 vdd.n1005 vdd.n987 35.2919
R38177 vdd.n1006 vdd.n1005 35.2919
R38178 vdd.n1018 vdd.n1006 35.2919
R38179 vdd.n1018 vdd.n1017 35.2919
R38180 vdd.n1017 vdd.n1016 35.2919
R38181 vdd.n1094 vdd.n1089 35.2919
R38182 vdd.n1107 vdd.n1089 35.2919
R38183 vdd.n1108 vdd.n1107 35.2919
R38184 vdd.n1120 vdd.n1108 35.2919
R38185 vdd.n1120 vdd.n1119 35.2919
R38186 vdd.n1119 vdd.n1118 35.2919
R38187 vdd.n2614 vdd.n2609 35.2919
R38188 vdd.n2627 vdd.n2609 35.2919
R38189 vdd.n2628 vdd.n2627 35.2919
R38190 vdd.n2640 vdd.n2628 35.2919
R38191 vdd.n2640 vdd.n2639 35.2919
R38192 vdd.n2639 vdd.n2638 35.2919
R38193 vdd.n1146 vdd.n1137 35.2919
R38194 vdd.n1155 vdd.n1137 35.2919
R38195 vdd.n1156 vdd.n1155 35.2919
R38196 vdd.n1168 vdd.n1156 35.2919
R38197 vdd.n1168 vdd.n1167 35.2919
R38198 vdd.n1167 vdd.n1166 35.2919
R38199 vdd.n1194 vdd.n1185 35.2919
R38200 vdd.n1203 vdd.n1185 35.2919
R38201 vdd.n1204 vdd.n1203 35.2919
R38202 vdd.n1216 vdd.n1204 35.2919
R38203 vdd.n1216 vdd.n1215 35.2919
R38204 vdd.n1215 vdd.n1214 35.2919
R38205 vdd.n1295 vdd.n1286 35.2919
R38206 vdd.n1304 vdd.n1286 35.2919
R38207 vdd.n1305 vdd.n1304 35.2919
R38208 vdd.n1317 vdd.n1305 35.2919
R38209 vdd.n1317 vdd.n1316 35.2919
R38210 vdd.n1316 vdd.n1315 35.2919
R38211 vdd.n1343 vdd.n1334 35.2919
R38212 vdd.n1352 vdd.n1334 35.2919
R38213 vdd.n1353 vdd.n1352 35.2919
R38214 vdd.n1365 vdd.n1353 35.2919
R38215 vdd.n1365 vdd.n1364 35.2919
R38216 vdd.n1364 vdd.n1363 35.2919
R38217 vdd.n1391 vdd.n1382 35.2919
R38218 vdd.n1400 vdd.n1382 35.2919
R38219 vdd.n1401 vdd.n1400 35.2919
R38220 vdd.n1413 vdd.n1401 35.2919
R38221 vdd.n1413 vdd.n1412 35.2919
R38222 vdd.n1412 vdd.n1411 35.2919
R38223 vdd.n1439 vdd.n1430 35.2919
R38224 vdd.n1448 vdd.n1430 35.2919
R38225 vdd.n1449 vdd.n1448 35.2919
R38226 vdd.n1461 vdd.n1449 35.2919
R38227 vdd.n1461 vdd.n1460 35.2919
R38228 vdd.n1460 vdd.n1459 35.2919
R38229 vdd.n1540 vdd.n1531 35.2919
R38230 vdd.n1549 vdd.n1531 35.2919
R38231 vdd.n1550 vdd.n1549 35.2919
R38232 vdd.n1562 vdd.n1550 35.2919
R38233 vdd.n1562 vdd.n1561 35.2919
R38234 vdd.n1561 vdd.n1560 35.2919
R38235 vdd.n653 vdd.n644 35.2919
R38236 vdd.n662 vdd.n644 35.2919
R38237 vdd.n663 vdd.n662 35.2919
R38238 vdd.n675 vdd.n663 35.2919
R38239 vdd.n675 vdd.n674 35.2919
R38240 vdd.n674 vdd.n673 35.2919
R38241 vdd.n1588 vdd.n1579 35.2919
R38242 vdd.n1597 vdd.n1579 35.2919
R38243 vdd.n1598 vdd.n1597 35.2919
R38244 vdd.n1610 vdd.n1598 35.2919
R38245 vdd.n1610 vdd.n1609 35.2919
R38246 vdd.n1609 vdd.n1608 35.2919
R38247 vdd.n1635 vdd.n1626 35.2919
R38248 vdd.n1644 vdd.n1626 35.2919
R38249 vdd.n1645 vdd.n1644 35.2919
R38250 vdd.n1657 vdd.n1645 35.2919
R38251 vdd.n1657 vdd.n1656 35.2919
R38252 vdd.n1656 vdd.n1655 35.2919
R38253 vdd.n1685 vdd.n1676 35.2919
R38254 vdd.n1694 vdd.n1676 35.2919
R38255 vdd.n1695 vdd.n1694 35.2919
R38256 vdd.n1707 vdd.n1695 35.2919
R38257 vdd.n1707 vdd.n1706 35.2919
R38258 vdd.n1706 vdd.n1705 35.2919
R38259 vdd.n1735 vdd.n1726 35.2919
R38260 vdd.n1744 vdd.n1726 35.2919
R38261 vdd.n1745 vdd.n1744 35.2919
R38262 vdd.n1757 vdd.n1745 35.2919
R38263 vdd.n1757 vdd.n1756 35.2919
R38264 vdd.n1756 vdd.n1755 35.2919
R38265 vdd.n1783 vdd.n1774 35.2919
R38266 vdd.n1792 vdd.n1774 35.2919
R38267 vdd.n1793 vdd.n1792 35.2919
R38268 vdd.n1805 vdd.n1793 35.2919
R38269 vdd.n1805 vdd.n1804 35.2919
R38270 vdd.n1804 vdd.n1803 35.2919
R38271 vdd.n1511 vdd.n1510 35.2919
R38272 vdd.n1510 vdd.n1509 35.2919
R38273 vdd.n1509 vdd.n1478 35.2919
R38274 vdd.n1497 vdd.n1478 35.2919
R38275 vdd.n1497 vdd.n1496 35.2919
R38276 vdd.n1496 vdd.n1495 35.2919
R38277 vdd.n1834 vdd.n1825 35.2919
R38278 vdd.n1843 vdd.n1825 35.2919
R38279 vdd.n1844 vdd.n1843 35.2919
R38280 vdd.n1856 vdd.n1844 35.2919
R38281 vdd.n1856 vdd.n1855 35.2919
R38282 vdd.n1855 vdd.n1854 35.2919
R38283 vdd.n1881 vdd.n1872 35.2919
R38284 vdd.n1890 vdd.n1872 35.2919
R38285 vdd.n1891 vdd.n1890 35.2919
R38286 vdd.n1903 vdd.n1891 35.2919
R38287 vdd.n1903 vdd.n1902 35.2919
R38288 vdd.n1902 vdd.n1901 35.2919
R38289 vdd.n1929 vdd.n1920 35.2919
R38290 vdd.n1938 vdd.n1920 35.2919
R38291 vdd.n1939 vdd.n1938 35.2919
R38292 vdd.n1951 vdd.n1939 35.2919
R38293 vdd.n1951 vdd.n1950 35.2919
R38294 vdd.n1950 vdd.n1949 35.2919
R38295 vdd.n1980 vdd.n1971 35.2919
R38296 vdd.n1989 vdd.n1971 35.2919
R38297 vdd.n1990 vdd.n1989 35.2919
R38298 vdd.n2002 vdd.n1990 35.2919
R38299 vdd.n2002 vdd.n2001 35.2919
R38300 vdd.n2001 vdd.n2000 35.2919
R38301 vdd.n2030 vdd.n2021 35.2919
R38302 vdd.n2039 vdd.n2021 35.2919
R38303 vdd.n2040 vdd.n2039 35.2919
R38304 vdd.n2052 vdd.n2040 35.2919
R38305 vdd.n2052 vdd.n2051 35.2919
R38306 vdd.n2051 vdd.n2050 35.2919
R38307 vdd.n2078 vdd.n2069 35.2919
R38308 vdd.n2087 vdd.n2069 35.2919
R38309 vdd.n2088 vdd.n2087 35.2919
R38310 vdd.n2100 vdd.n2088 35.2919
R38311 vdd.n2100 vdd.n2099 35.2919
R38312 vdd.n2099 vdd.n2098 35.2919
R38313 vdd.n2128 vdd.n2119 35.2919
R38314 vdd.n2137 vdd.n2119 35.2919
R38315 vdd.n2138 vdd.n2137 35.2919
R38316 vdd.n2150 vdd.n2138 35.2919
R38317 vdd.n2150 vdd.n2149 35.2919
R38318 vdd.n2149 vdd.n2148 35.2919
R38319 vdd.n2175 vdd.n2166 35.2919
R38320 vdd.n2184 vdd.n2166 35.2919
R38321 vdd.n2185 vdd.n2184 35.2919
R38322 vdd.n2197 vdd.n2185 35.2919
R38323 vdd.n2197 vdd.n2196 35.2919
R38324 vdd.n2196 vdd.n2195 35.2919
R38325 vdd.n2225 vdd.n2216 35.2919
R38326 vdd.n2234 vdd.n2216 35.2919
R38327 vdd.n2235 vdd.n2234 35.2919
R38328 vdd.n2247 vdd.n2235 35.2919
R38329 vdd.n2247 vdd.n2246 35.2919
R38330 vdd.n2246 vdd.n2245 35.2919
R38331 vdd.n2275 vdd.n2266 35.2919
R38332 vdd.n2284 vdd.n2266 35.2919
R38333 vdd.n2285 vdd.n2284 35.2919
R38334 vdd.n2297 vdd.n2285 35.2919
R38335 vdd.n2297 vdd.n2296 35.2919
R38336 vdd.n2296 vdd.n2295 35.2919
R38337 vdd.n2323 vdd.n2314 35.2919
R38338 vdd.n2332 vdd.n2314 35.2919
R38339 vdd.n2333 vdd.n2332 35.2919
R38340 vdd.n2345 vdd.n2333 35.2919
R38341 vdd.n2345 vdd.n2344 35.2919
R38342 vdd.n2344 vdd.n2343 35.2919
R38343 vdd.n1266 vdd.n1265 35.2919
R38344 vdd.n1265 vdd.n1264 35.2919
R38345 vdd.n1264 vdd.n1233 35.2919
R38346 vdd.n1252 vdd.n1233 35.2919
R38347 vdd.n1252 vdd.n1251 35.2919
R38348 vdd.n1251 vdd.n1250 35.2919
R38349 vdd.n2374 vdd.n2365 35.2919
R38350 vdd.n2383 vdd.n2365 35.2919
R38351 vdd.n2384 vdd.n2383 35.2919
R38352 vdd.n2396 vdd.n2384 35.2919
R38353 vdd.n2396 vdd.n2395 35.2919
R38354 vdd.n2395 vdd.n2394 35.2919
R38355 vdd.n2421 vdd.n2412 35.2919
R38356 vdd.n2430 vdd.n2412 35.2919
R38357 vdd.n2431 vdd.n2430 35.2919
R38358 vdd.n2443 vdd.n2431 35.2919
R38359 vdd.n2443 vdd.n2442 35.2919
R38360 vdd.n2442 vdd.n2441 35.2919
R38361 vdd.n2471 vdd.n2462 35.2919
R38362 vdd.n2480 vdd.n2462 35.2919
R38363 vdd.n2481 vdd.n2480 35.2919
R38364 vdd.n2493 vdd.n2481 35.2919
R38365 vdd.n2493 vdd.n2492 35.2919
R38366 vdd.n2492 vdd.n2491 35.2919
R38367 vdd.n2521 vdd.n2512 35.2919
R38368 vdd.n2530 vdd.n2512 35.2919
R38369 vdd.n2531 vdd.n2530 35.2919
R38370 vdd.n2543 vdd.n2531 35.2919
R38371 vdd.n2543 vdd.n2542 35.2919
R38372 vdd.n2542 vdd.n2541 35.2919
R38373 vdd.n2569 vdd.n2560 35.2919
R38374 vdd.n2578 vdd.n2560 35.2919
R38375 vdd.n2579 vdd.n2578 35.2919
R38376 vdd.n2591 vdd.n2579 35.2919
R38377 vdd.n2591 vdd.n2590 35.2919
R38378 vdd.n2590 vdd.n2589 35.2919
R38379 vdd.n2711 vdd.n2706 35.2919
R38380 vdd.n2724 vdd.n2706 35.2919
R38381 vdd.n2725 vdd.n2724 35.2919
R38382 vdd.n2737 vdd.n2725 35.2919
R38383 vdd.n2737 vdd.n2736 35.2919
R38384 vdd.n2736 vdd.n2735 35.2919
R38385 vdd.n2663 vdd.n2658 35.2919
R38386 vdd.n2676 vdd.n2658 35.2919
R38387 vdd.n2677 vdd.n2676 35.2919
R38388 vdd.n2689 vdd.n2677 35.2919
R38389 vdd.n2689 vdd.n2688 35.2919
R38390 vdd.n2688 vdd.n2687 35.2919
R38391 vdd.n2760 vdd.n2755 35.2919
R38392 vdd.n2773 vdd.n2755 35.2919
R38393 vdd.n2774 vdd.n2773 35.2919
R38394 vdd.n2786 vdd.n2774 35.2919
R38395 vdd.n2786 vdd.n2785 35.2919
R38396 vdd.n2785 vdd.n2784 35.2919
R38397 vdd.n2810 vdd.n2805 35.2919
R38398 vdd.n2823 vdd.n2805 35.2919
R38399 vdd.n2824 vdd.n2823 35.2919
R38400 vdd.n2836 vdd.n2824 35.2919
R38401 vdd.n2836 vdd.n2835 35.2919
R38402 vdd.n2835 vdd.n2834 35.2919
R38403 vdd.n2858 vdd.n2853 35.2919
R38404 vdd.n2871 vdd.n2853 35.2919
R38405 vdd.n2872 vdd.n2871 35.2919
R38406 vdd.n2884 vdd.n2872 35.2919
R38407 vdd.n2884 vdd.n2883 35.2919
R38408 vdd.n2883 vdd.n2882 35.2919
R38409 vdd.n1046 vdd.n1045 35.2919
R38410 vdd.n1045 vdd.n1044 35.2919
R38411 vdd.n1044 vdd.n1033 35.2919
R38412 vdd.n1056 vdd.n1033 35.2919
R38413 vdd.n1056 vdd.n1029 35.2919
R38414 vdd.n1072 vdd.n1029 35.2919
R38415 vdd.n3006 vdd.n3001 35.2919
R38416 vdd.n3019 vdd.n3001 35.2919
R38417 vdd.n3020 vdd.n3019 35.2919
R38418 vdd.n3032 vdd.n3020 35.2919
R38419 vdd.n3032 vdd.n3031 35.2919
R38420 vdd.n3031 vdd.n3030 35.2919
R38421 vdd.n2957 vdd.n2952 35.2919
R38422 vdd.n2970 vdd.n2952 35.2919
R38423 vdd.n2971 vdd.n2970 35.2919
R38424 vdd.n2983 vdd.n2971 35.2919
R38425 vdd.n2983 vdd.n2982 35.2919
R38426 vdd.n2982 vdd.n2981 35.2919
R38427 vdd.n2909 vdd.n2904 35.2919
R38428 vdd.n2922 vdd.n2904 35.2919
R38429 vdd.n2923 vdd.n2922 35.2919
R38430 vdd.n2935 vdd.n2923 35.2919
R38431 vdd.n2935 vdd.n2934 35.2919
R38432 vdd.n2934 vdd.n2933 35.2919
R38433 vdd.n3055 vdd.n3050 35.2919
R38434 vdd.n3068 vdd.n3050 35.2919
R38435 vdd.n3069 vdd.n3068 35.2919
R38436 vdd.n3081 vdd.n3069 35.2919
R38437 vdd.n3081 vdd.n3080 35.2919
R38438 vdd.n3080 vdd.n3079 35.2919
R38439 vdd.n3105 vdd.n3100 35.2919
R38440 vdd.n3118 vdd.n3100 35.2919
R38441 vdd.n3119 vdd.n3118 35.2919
R38442 vdd.n3131 vdd.n3119 35.2919
R38443 vdd.n3131 vdd.n3130 35.2919
R38444 vdd.n3130 vdd.n3129 35.2919
R38445 vdd.n3153 vdd.n3148 35.2919
R38446 vdd.n3166 vdd.n3148 35.2919
R38447 vdd.n3167 vdd.n3166 35.2919
R38448 vdd.n3179 vdd.n3167 35.2919
R38449 vdd.n3179 vdd.n3178 35.2919
R38450 vdd.n3178 vdd.n3177 35.2919
R38451 vdd.n3251 vdd.n3246 35.2919
R38452 vdd.n3264 vdd.n3246 35.2919
R38453 vdd.n3265 vdd.n3264 35.2919
R38454 vdd.n3277 vdd.n3265 35.2919
R38455 vdd.n3277 vdd.n3276 35.2919
R38456 vdd.n3276 vdd.n3275 35.2919
R38457 vdd.n3203 vdd.n3198 35.2919
R38458 vdd.n3216 vdd.n3198 35.2919
R38459 vdd.n3217 vdd.n3216 35.2919
R38460 vdd.n3229 vdd.n3217 35.2919
R38461 vdd.n3229 vdd.n3228 35.2919
R38462 vdd.n3228 vdd.n3227 35.2919
R38463 vdd.n3300 vdd.n3295 35.2919
R38464 vdd.n3313 vdd.n3295 35.2919
R38465 vdd.n3314 vdd.n3313 35.2919
R38466 vdd.n3326 vdd.n3314 35.2919
R38467 vdd.n3326 vdd.n3325 35.2919
R38468 vdd.n3325 vdd.n3324 35.2919
R38469 vdd.n3350 vdd.n3345 35.2919
R38470 vdd.n3363 vdd.n3345 35.2919
R38471 vdd.n3364 vdd.n3363 35.2919
R38472 vdd.n3376 vdd.n3364 35.2919
R38473 vdd.n3376 vdd.n3375 35.2919
R38474 vdd.n3375 vdd.n3374 35.2919
R38475 vdd.n3398 vdd.n3393 35.2919
R38476 vdd.n3411 vdd.n3393 35.2919
R38477 vdd.n3412 vdd.n3411 35.2919
R38478 vdd.n3424 vdd.n3412 35.2919
R38479 vdd.n3424 vdd.n3423 35.2919
R38480 vdd.n3423 vdd.n3422 35.2919
R38481 vdd.n800 vdd.n799 35.2919
R38482 vdd.n799 vdd.n798 35.2919
R38483 vdd.n798 vdd.n787 35.2919
R38484 vdd.n810 vdd.n787 35.2919
R38485 vdd.n810 vdd.n783 35.2919
R38486 vdd.n826 vdd.n783 35.2919
R38487 vdd.n3497 vdd.n3492 35.2919
R38488 vdd.n3510 vdd.n3492 35.2919
R38489 vdd.n3511 vdd.n3510 35.2919
R38490 vdd.n3523 vdd.n3511 35.2919
R38491 vdd.n3523 vdd.n3522 35.2919
R38492 vdd.n3522 vdd.n3521 35.2919
R38493 vdd.n3449 vdd.n3444 35.2919
R38494 vdd.n3462 vdd.n3444 35.2919
R38495 vdd.n3463 vdd.n3462 35.2919
R38496 vdd.n3475 vdd.n3463 35.2919
R38497 vdd.n3475 vdd.n3474 35.2919
R38498 vdd.n3474 vdd.n3473 35.2919
R38499 vdd.n3546 vdd.n3541 35.2919
R38500 vdd.n3559 vdd.n3541 35.2919
R38501 vdd.n3560 vdd.n3559 35.2919
R38502 vdd.n3572 vdd.n3560 35.2919
R38503 vdd.n3572 vdd.n3571 35.2919
R38504 vdd.n3571 vdd.n3570 35.2919
R38505 vdd.n3596 vdd.n3591 35.2919
R38506 vdd.n3609 vdd.n3591 35.2919
R38507 vdd.n3610 vdd.n3609 35.2919
R38508 vdd.n3622 vdd.n3610 35.2919
R38509 vdd.n3622 vdd.n3621 35.2919
R38510 vdd.n3621 vdd.n3620 35.2919
R38511 vdd.n3644 vdd.n3639 35.2919
R38512 vdd.n3657 vdd.n3639 35.2919
R38513 vdd.n3658 vdd.n3657 35.2919
R38514 vdd.n3670 vdd.n3658 35.2919
R38515 vdd.n3670 vdd.n3669 35.2919
R38516 vdd.n3669 vdd.n3668 35.2919
R38517 vdd.n602 vdd.n597 35.2919
R38518 vdd.n615 vdd.n597 35.2919
R38519 vdd.n616 vdd.n615 35.2919
R38520 vdd.n628 vdd.n616 35.2919
R38521 vdd.n628 vdd.n627 35.2919
R38522 vdd.n627 vdd.n626 35.2919
R38523 vdd.n3743 vdd.n3738 35.2919
R38524 vdd.n3756 vdd.n3738 35.2919
R38525 vdd.n3757 vdd.n3756 35.2919
R38526 vdd.n3769 vdd.n3757 35.2919
R38527 vdd.n3769 vdd.n3768 35.2919
R38528 vdd.n3768 vdd.n3767 35.2919
R38529 vdd.n3695 vdd.n3690 35.2919
R38530 vdd.n3708 vdd.n3690 35.2919
R38531 vdd.n3709 vdd.n3708 35.2919
R38532 vdd.n3721 vdd.n3709 35.2919
R38533 vdd.n3721 vdd.n3720 35.2919
R38534 vdd.n3720 vdd.n3719 35.2919
R38535 vdd.n6885 vdd.n6880 35.2919
R38536 vdd.n6898 vdd.n6880 35.2919
R38537 vdd.n6899 vdd.n6898 35.2919
R38538 vdd.n6911 vdd.n6899 35.2919
R38539 vdd.n6911 vdd.n6910 35.2919
R38540 vdd.n6910 vdd.n6909 35.2919
R38541 vdd.n6837 vdd.n6832 35.2919
R38542 vdd.n6850 vdd.n6832 35.2919
R38543 vdd.n6851 vdd.n6850 35.2919
R38544 vdd.n6863 vdd.n6851 35.2919
R38545 vdd.n6863 vdd.n6862 35.2919
R38546 vdd.n6862 vdd.n6861 35.2919
R38547 vdd.n10027 vdd.n10022 35.2919
R38548 vdd.n10040 vdd.n10022 35.2919
R38549 vdd.n10041 vdd.n10040 35.2919
R38550 vdd.n10053 vdd.n10041 35.2919
R38551 vdd.n10053 vdd.n10052 35.2919
R38552 vdd.n10052 vdd.n10051 35.2919
R38553 vdd.n9979 vdd.n9974 35.2919
R38554 vdd.n9992 vdd.n9974 35.2919
R38555 vdd.n9993 vdd.n9992 35.2919
R38556 vdd.n10005 vdd.n9993 35.2919
R38557 vdd.n10005 vdd.n10004 35.2919
R38558 vdd.n10004 vdd.n10003 35.2919
R38559 vdd.n10075 vdd.n10070 35.2919
R38560 vdd.n10088 vdd.n10070 35.2919
R38561 vdd.n10089 vdd.n10088 35.2919
R38562 vdd.n10101 vdd.n10089 35.2919
R38563 vdd.n10101 vdd.n10100 35.2919
R38564 vdd.n10100 vdd.n10099 35.2919
R38565 vdd.n10123 vdd.n10118 35.2919
R38566 vdd.n10136 vdd.n10118 35.2919
R38567 vdd.n10137 vdd.n10136 35.2919
R38568 vdd.n10149 vdd.n10137 35.2919
R38569 vdd.n10149 vdd.n10148 35.2919
R38570 vdd.n10148 vdd.n10147 35.2919
R38571 vdd.n10225 vdd.n10220 35.2919
R38572 vdd.n10238 vdd.n10220 35.2919
R38573 vdd.n10239 vdd.n10238 35.2919
R38574 vdd.n10251 vdd.n10239 35.2919
R38575 vdd.n10251 vdd.n10250 35.2919
R38576 vdd.n10250 vdd.n10249 35.2919
R38577 vdd.n10273 vdd.n10268 35.2919
R38578 vdd.n10286 vdd.n10268 35.2919
R38579 vdd.n10287 vdd.n10286 35.2919
R38580 vdd.n10299 vdd.n10287 35.2919
R38581 vdd.n10299 vdd.n10298 35.2919
R38582 vdd.n10298 vdd.n10297 35.2919
R38583 vdd.n10321 vdd.n10316 35.2919
R38584 vdd.n10334 vdd.n10316 35.2919
R38585 vdd.n10335 vdd.n10334 35.2919
R38586 vdd.n10347 vdd.n10335 35.2919
R38587 vdd.n10347 vdd.n10346 35.2919
R38588 vdd.n10346 vdd.n10345 35.2919
R38589 vdd.n10369 vdd.n10364 35.2919
R38590 vdd.n10382 vdd.n10364 35.2919
R38591 vdd.n10383 vdd.n10382 35.2919
R38592 vdd.n10395 vdd.n10383 35.2919
R38593 vdd.n10395 vdd.n10394 35.2919
R38594 vdd.n10394 vdd.n10393 35.2919
R38595 vdd.n10471 vdd.n10466 35.2919
R38596 vdd.n10484 vdd.n10466 35.2919
R38597 vdd.n10485 vdd.n10484 35.2919
R38598 vdd.n10497 vdd.n10485 35.2919
R38599 vdd.n10497 vdd.n10496 35.2919
R38600 vdd.n10496 vdd.n10495 35.2919
R38601 vdd.n63 vdd.n58 35.2919
R38602 vdd.n76 vdd.n58 35.2919
R38603 vdd.n77 vdd.n76 35.2919
R38604 vdd.n89 vdd.n77 35.2919
R38605 vdd.n89 vdd.n88 35.2919
R38606 vdd.n88 vdd.n87 35.2919
R38607 vdd.n15 vdd.n10 35.2919
R38608 vdd.n28 vdd.n10 35.2919
R38609 vdd.n29 vdd.n28 35.2919
R38610 vdd.n41 vdd.n29 35.2919
R38611 vdd.n41 vdd.n40 35.2919
R38612 vdd.n40 vdd.n39 35.2919
R38613 vdd.n10519 vdd.n10514 35.2919
R38614 vdd.n10532 vdd.n10514 35.2919
R38615 vdd.n10533 vdd.n10532 35.2919
R38616 vdd.n10545 vdd.n10533 35.2919
R38617 vdd.n10545 vdd.n10544 35.2919
R38618 vdd.n10544 vdd.n10543 35.2919
R38619 vdd.n10569 vdd.n10564 35.2919
R38620 vdd.n10582 vdd.n10564 35.2919
R38621 vdd.n10583 vdd.n10582 35.2919
R38622 vdd.n10595 vdd.n10583 35.2919
R38623 vdd.n10595 vdd.n10594 35.2919
R38624 vdd.n10594 vdd.n10593 35.2919
R38625 vdd.n10617 vdd.n10612 35.2919
R38626 vdd.n10630 vdd.n10612 35.2919
R38627 vdd.n10631 vdd.n10630 35.2919
R38628 vdd.n10643 vdd.n10631 35.2919
R38629 vdd.n10643 vdd.n10642 35.2919
R38630 vdd.n10642 vdd.n10641 35.2919
R38631 vdd.n10423 vdd.n10422 35.2919
R38632 vdd.n10422 vdd.n10421 35.2919
R38633 vdd.n10421 vdd.n10410 35.2919
R38634 vdd.n10433 vdd.n10410 35.2919
R38635 vdd.n10433 vdd.n10406 35.2919
R38636 vdd.n10449 vdd.n10406 35.2919
R38637 vdd.n10765 vdd.n10760 35.2919
R38638 vdd.n10778 vdd.n10760 35.2919
R38639 vdd.n10779 vdd.n10778 35.2919
R38640 vdd.n10791 vdd.n10779 35.2919
R38641 vdd.n10791 vdd.n10790 35.2919
R38642 vdd.n10790 vdd.n10789 35.2919
R38643 vdd.n10716 vdd.n10711 35.2919
R38644 vdd.n10729 vdd.n10711 35.2919
R38645 vdd.n10730 vdd.n10729 35.2919
R38646 vdd.n10742 vdd.n10730 35.2919
R38647 vdd.n10742 vdd.n10741 35.2919
R38648 vdd.n10741 vdd.n10740 35.2919
R38649 vdd.n10668 vdd.n10663 35.2919
R38650 vdd.n10681 vdd.n10663 35.2919
R38651 vdd.n10682 vdd.n10681 35.2919
R38652 vdd.n10694 vdd.n10682 35.2919
R38653 vdd.n10694 vdd.n10693 35.2919
R38654 vdd.n10693 vdd.n10692 35.2919
R38655 vdd.n10814 vdd.n10809 35.2919
R38656 vdd.n10827 vdd.n10809 35.2919
R38657 vdd.n10828 vdd.n10827 35.2919
R38658 vdd.n10840 vdd.n10828 35.2919
R38659 vdd.n10840 vdd.n10839 35.2919
R38660 vdd.n10839 vdd.n10838 35.2919
R38661 vdd.n10864 vdd.n10859 35.2919
R38662 vdd.n10877 vdd.n10859 35.2919
R38663 vdd.n10878 vdd.n10877 35.2919
R38664 vdd.n10890 vdd.n10878 35.2919
R38665 vdd.n10890 vdd.n10889 35.2919
R38666 vdd.n10889 vdd.n10888 35.2919
R38667 vdd.n10912 vdd.n10907 35.2919
R38668 vdd.n10925 vdd.n10907 35.2919
R38669 vdd.n10926 vdd.n10925 35.2919
R38670 vdd.n10938 vdd.n10926 35.2919
R38671 vdd.n10938 vdd.n10937 35.2919
R38672 vdd.n10937 vdd.n10936 35.2919
R38673 vdd.n11010 vdd.n11005 35.2919
R38674 vdd.n11023 vdd.n11005 35.2919
R38675 vdd.n11024 vdd.n11023 35.2919
R38676 vdd.n11036 vdd.n11024 35.2919
R38677 vdd.n11036 vdd.n11035 35.2919
R38678 vdd.n11035 vdd.n11034 35.2919
R38679 vdd.n10962 vdd.n10957 35.2919
R38680 vdd.n10975 vdd.n10957 35.2919
R38681 vdd.n10976 vdd.n10975 35.2919
R38682 vdd.n10988 vdd.n10976 35.2919
R38683 vdd.n10988 vdd.n10987 35.2919
R38684 vdd.n10987 vdd.n10986 35.2919
R38685 vdd.n11059 vdd.n11054 35.2919
R38686 vdd.n11072 vdd.n11054 35.2919
R38687 vdd.n11073 vdd.n11072 35.2919
R38688 vdd.n11085 vdd.n11073 35.2919
R38689 vdd.n11085 vdd.n11084 35.2919
R38690 vdd.n11084 vdd.n11083 35.2919
R38691 vdd.n11109 vdd.n11104 35.2919
R38692 vdd.n11122 vdd.n11104 35.2919
R38693 vdd.n11123 vdd.n11122 35.2919
R38694 vdd.n11135 vdd.n11123 35.2919
R38695 vdd.n11135 vdd.n11134 35.2919
R38696 vdd.n11134 vdd.n11133 35.2919
R38697 vdd.n11157 vdd.n11152 35.2919
R38698 vdd.n11170 vdd.n11152 35.2919
R38699 vdd.n11171 vdd.n11170 35.2919
R38700 vdd.n11183 vdd.n11171 35.2919
R38701 vdd.n11183 vdd.n11182 35.2919
R38702 vdd.n11182 vdd.n11181 35.2919
R38703 vdd.n10177 vdd.n10176 35.2919
R38704 vdd.n10176 vdd.n10175 35.2919
R38705 vdd.n10175 vdd.n10164 35.2919
R38706 vdd.n10187 vdd.n10164 35.2919
R38707 vdd.n10187 vdd.n10160 35.2919
R38708 vdd.n10203 vdd.n10160 35.2919
R38709 vdd.n11256 vdd.n11251 35.2919
R38710 vdd.n11269 vdd.n11251 35.2919
R38711 vdd.n11270 vdd.n11269 35.2919
R38712 vdd.n11282 vdd.n11270 35.2919
R38713 vdd.n11282 vdd.n11281 35.2919
R38714 vdd.n11281 vdd.n11280 35.2919
R38715 vdd.n11208 vdd.n11203 35.2919
R38716 vdd.n11221 vdd.n11203 35.2919
R38717 vdd.n11222 vdd.n11221 35.2919
R38718 vdd.n11234 vdd.n11222 35.2919
R38719 vdd.n11234 vdd.n11233 35.2919
R38720 vdd.n11233 vdd.n11232 35.2919
R38721 vdd.n11305 vdd.n11300 35.2919
R38722 vdd.n11318 vdd.n11300 35.2919
R38723 vdd.n11319 vdd.n11318 35.2919
R38724 vdd.n11331 vdd.n11319 35.2919
R38725 vdd.n11331 vdd.n11330 35.2919
R38726 vdd.n11330 vdd.n11329 35.2919
R38727 vdd.n11355 vdd.n11350 35.2919
R38728 vdd.n11368 vdd.n11350 35.2919
R38729 vdd.n11369 vdd.n11368 35.2919
R38730 vdd.n11381 vdd.n11369 35.2919
R38731 vdd.n11381 vdd.n11380 35.2919
R38732 vdd.n11380 vdd.n11379 35.2919
R38733 vdd.n11403 vdd.n11398 35.2919
R38734 vdd.n11416 vdd.n11398 35.2919
R38735 vdd.n11417 vdd.n11416 35.2919
R38736 vdd.n11429 vdd.n11417 35.2919
R38737 vdd.n11429 vdd.n11428 35.2919
R38738 vdd.n11428 vdd.n11427 35.2919
R38739 vdd.n11458 vdd.n11449 35.2919
R38740 vdd.n11467 vdd.n11449 35.2919
R38741 vdd.n11468 vdd.n11467 35.2919
R38742 vdd.n11480 vdd.n11468 35.2919
R38743 vdd.n11480 vdd.n11479 35.2919
R38744 vdd.n11479 vdd.n11478 35.2919
R38745 vdd.n11505 vdd.n11496 35.2919
R38746 vdd.n11514 vdd.n11496 35.2919
R38747 vdd.n11515 vdd.n11514 35.2919
R38748 vdd.n11527 vdd.n11515 35.2919
R38749 vdd.n11527 vdd.n11526 35.2919
R38750 vdd.n11526 vdd.n11525 35.2919
R38751 vdd.n11555 vdd.n11546 35.2919
R38752 vdd.n11564 vdd.n11546 35.2919
R38753 vdd.n11565 vdd.n11564 35.2919
R38754 vdd.n11577 vdd.n11565 35.2919
R38755 vdd.n11577 vdd.n11576 35.2919
R38756 vdd.n11576 vdd.n11575 35.2919
R38757 vdd.n11605 vdd.n11596 35.2919
R38758 vdd.n11614 vdd.n11596 35.2919
R38759 vdd.n11615 vdd.n11614 35.2919
R38760 vdd.n11627 vdd.n11615 35.2919
R38761 vdd.n11627 vdd.n11626 35.2919
R38762 vdd.n11626 vdd.n11625 35.2919
R38763 vdd.n11653 vdd.n11644 35.2919
R38764 vdd.n11662 vdd.n11644 35.2919
R38765 vdd.n11663 vdd.n11662 35.2919
R38766 vdd.n11675 vdd.n11663 35.2919
R38767 vdd.n11675 vdd.n11674 35.2919
R38768 vdd.n11674 vdd.n11673 35.2919
R38769 vdd.n481 vdd.n480 35.2919
R38770 vdd.n480 vdd.n479 35.2919
R38771 vdd.n479 vdd.n448 35.2919
R38772 vdd.n467 vdd.n448 35.2919
R38773 vdd.n467 vdd.n466 35.2919
R38774 vdd.n466 vdd.n465 35.2919
R38775 vdd.n11704 vdd.n11695 35.2919
R38776 vdd.n11713 vdd.n11695 35.2919
R38777 vdd.n11714 vdd.n11713 35.2919
R38778 vdd.n11726 vdd.n11714 35.2919
R38779 vdd.n11726 vdd.n11725 35.2919
R38780 vdd.n11725 vdd.n11724 35.2919
R38781 vdd.n11751 vdd.n11742 35.2919
R38782 vdd.n11760 vdd.n11742 35.2919
R38783 vdd.n11761 vdd.n11760 35.2919
R38784 vdd.n11773 vdd.n11761 35.2919
R38785 vdd.n11773 vdd.n11772 35.2919
R38786 vdd.n11772 vdd.n11771 35.2919
R38787 vdd.n11799 vdd.n11790 35.2919
R38788 vdd.n11808 vdd.n11790 35.2919
R38789 vdd.n11809 vdd.n11808 35.2919
R38790 vdd.n11821 vdd.n11809 35.2919
R38791 vdd.n11821 vdd.n11820 35.2919
R38792 vdd.n11820 vdd.n11819 35.2919
R38793 vdd.n11850 vdd.n11841 35.2919
R38794 vdd.n11859 vdd.n11841 35.2919
R38795 vdd.n11860 vdd.n11859 35.2919
R38796 vdd.n11872 vdd.n11860 35.2919
R38797 vdd.n11872 vdd.n11871 35.2919
R38798 vdd.n11871 vdd.n11870 35.2919
R38799 vdd.n11900 vdd.n11891 35.2919
R38800 vdd.n11909 vdd.n11891 35.2919
R38801 vdd.n11910 vdd.n11909 35.2919
R38802 vdd.n11922 vdd.n11910 35.2919
R38803 vdd.n11922 vdd.n11921 35.2919
R38804 vdd.n11921 vdd.n11920 35.2919
R38805 vdd.n11948 vdd.n11939 35.2919
R38806 vdd.n11957 vdd.n11939 35.2919
R38807 vdd.n11958 vdd.n11957 35.2919
R38808 vdd.n11970 vdd.n11958 35.2919
R38809 vdd.n11970 vdd.n11969 35.2919
R38810 vdd.n11969 vdd.n11968 35.2919
R38811 vdd.n11998 vdd.n11989 35.2919
R38812 vdd.n12007 vdd.n11989 35.2919
R38813 vdd.n12008 vdd.n12007 35.2919
R38814 vdd.n12020 vdd.n12008 35.2919
R38815 vdd.n12020 vdd.n12019 35.2919
R38816 vdd.n12019 vdd.n12018 35.2919
R38817 vdd.n12045 vdd.n12036 35.2919
R38818 vdd.n12054 vdd.n12036 35.2919
R38819 vdd.n12055 vdd.n12054 35.2919
R38820 vdd.n12067 vdd.n12055 35.2919
R38821 vdd.n12067 vdd.n12066 35.2919
R38822 vdd.n12066 vdd.n12065 35.2919
R38823 vdd.n12095 vdd.n12086 35.2919
R38824 vdd.n12104 vdd.n12086 35.2919
R38825 vdd.n12105 vdd.n12104 35.2919
R38826 vdd.n12117 vdd.n12105 35.2919
R38827 vdd.n12117 vdd.n12116 35.2919
R38828 vdd.n12116 vdd.n12115 35.2919
R38829 vdd.n12145 vdd.n12136 35.2919
R38830 vdd.n12154 vdd.n12136 35.2919
R38831 vdd.n12155 vdd.n12154 35.2919
R38832 vdd.n12167 vdd.n12155 35.2919
R38833 vdd.n12167 vdd.n12166 35.2919
R38834 vdd.n12166 vdd.n12165 35.2919
R38835 vdd.n12193 vdd.n12184 35.2919
R38836 vdd.n12202 vdd.n12184 35.2919
R38837 vdd.n12203 vdd.n12202 35.2919
R38838 vdd.n12215 vdd.n12203 35.2919
R38839 vdd.n12215 vdd.n12214 35.2919
R38840 vdd.n12214 vdd.n12213 35.2919
R38841 vdd.n236 vdd.n235 35.2919
R38842 vdd.n235 vdd.n234 35.2919
R38843 vdd.n234 vdd.n203 35.2919
R38844 vdd.n222 vdd.n203 35.2919
R38845 vdd.n222 vdd.n221 35.2919
R38846 vdd.n221 vdd.n220 35.2919
R38847 vdd.n12244 vdd.n12235 35.2919
R38848 vdd.n12253 vdd.n12235 35.2919
R38849 vdd.n12254 vdd.n12253 35.2919
R38850 vdd.n12266 vdd.n12254 35.2919
R38851 vdd.n12266 vdd.n12265 35.2919
R38852 vdd.n12265 vdd.n12264 35.2919
R38853 vdd.n12291 vdd.n12282 35.2919
R38854 vdd.n12300 vdd.n12282 35.2919
R38855 vdd.n12301 vdd.n12300 35.2919
R38856 vdd.n12313 vdd.n12301 35.2919
R38857 vdd.n12313 vdd.n12312 35.2919
R38858 vdd.n12312 vdd.n12311 35.2919
R38859 vdd.n12341 vdd.n12332 35.2919
R38860 vdd.n12350 vdd.n12332 35.2919
R38861 vdd.n12351 vdd.n12350 35.2919
R38862 vdd.n12363 vdd.n12351 35.2919
R38863 vdd.n12363 vdd.n12362 35.2919
R38864 vdd.n12362 vdd.n12361 35.2919
R38865 vdd.n12391 vdd.n12382 35.2919
R38866 vdd.n12400 vdd.n12382 35.2919
R38867 vdd.n12401 vdd.n12400 35.2919
R38868 vdd.n12413 vdd.n12401 35.2919
R38869 vdd.n12413 vdd.n12412 35.2919
R38870 vdd.n12412 vdd.n12411 35.2919
R38871 vdd.n12439 vdd.n12430 35.2919
R38872 vdd.n12448 vdd.n12430 35.2919
R38873 vdd.n12449 vdd.n12448 35.2919
R38874 vdd.n12461 vdd.n12449 35.2919
R38875 vdd.n12461 vdd.n12460 35.2919
R38876 vdd.n12460 vdd.n12459 35.2919
R38877 vdd.n12484 vdd.n12483 16.2531
R38878 vdd.n12495 vdd.n12484 16.2531
R38879 vdd.n12516 vdd.n12495 16.2531
R38880 vdd.n12516 vdd.n12515 16.2531
R38881 vdd.n12515 vdd.n12507 16.2531
R38882 vdd.n12507 vdd.n12506 16.2531
R38883 vdd.n114 vdd.n113 16.2531
R38884 vdd.n113 vdd.n98 16.2531
R38885 vdd.n143 vdd.n98 16.2531
R38886 vdd.n143 vdd.n142 16.2531
R38887 vdd.n142 vdd.n99 16.2531
R38888 vdd.n131 vdd.n99 16.2531
R38889 vdd.n162 vdd.n161 16.2531
R38890 vdd.n161 vdd.n146 16.2531
R38891 vdd.n191 vdd.n146 16.2531
R38892 vdd.n191 vdd.n190 16.2531
R38893 vdd.n190 vdd.n147 16.2531
R38894 vdd.n179 vdd.n147 16.2531
R38895 vdd.n263 vdd.n262 16.2531
R38896 vdd.n262 vdd.n247 16.2531
R38897 vdd.n292 vdd.n247 16.2531
R38898 vdd.n292 vdd.n291 16.2531
R38899 vdd.n291 vdd.n248 16.2531
R38900 vdd.n280 vdd.n248 16.2531
R38901 vdd.n311 vdd.n310 16.2531
R38902 vdd.n310 vdd.n295 16.2531
R38903 vdd.n340 vdd.n295 16.2531
R38904 vdd.n340 vdd.n339 16.2531
R38905 vdd.n339 vdd.n296 16.2531
R38906 vdd.n328 vdd.n296 16.2531
R38907 vdd.n359 vdd.n358 16.2531
R38908 vdd.n358 vdd.n343 16.2531
R38909 vdd.n388 vdd.n343 16.2531
R38910 vdd.n388 vdd.n387 16.2531
R38911 vdd.n387 vdd.n344 16.2531
R38912 vdd.n376 vdd.n344 16.2531
R38913 vdd.n407 vdd.n406 16.2531
R38914 vdd.n406 vdd.n391 16.2531
R38915 vdd.n436 vdd.n391 16.2531
R38916 vdd.n436 vdd.n435 16.2531
R38917 vdd.n435 vdd.n392 16.2531
R38918 vdd.n424 vdd.n392 16.2531
R38919 vdd.n508 vdd.n507 16.2531
R38920 vdd.n507 vdd.n492 16.2531
R38921 vdd.n537 vdd.n492 16.2531
R38922 vdd.n537 vdd.n536 16.2531
R38923 vdd.n536 vdd.n493 16.2531
R38924 vdd.n525 vdd.n493 16.2531
R38925 vdd.n556 vdd.n555 16.2531
R38926 vdd.n555 vdd.n540 16.2531
R38927 vdd.n585 vdd.n540 16.2531
R38928 vdd.n585 vdd.n584 16.2531
R38929 vdd.n584 vdd.n541 16.2531
R38930 vdd.n573 vdd.n541 16.2531
R38931 vdd.n6989 vdd.n6988 16.2531
R38932 vdd.n6988 vdd.n6968 16.2531
R38933 vdd.n7013 vdd.n6968 16.2531
R38934 vdd.n7013 vdd.n7012 16.2531
R38935 vdd.n7012 vdd.n6969 16.2531
R38936 vdd.n7001 vdd.n6969 16.2531
R38937 vdd.n7037 vdd.n7036 16.2531
R38938 vdd.n7036 vdd.n7016 16.2531
R38939 vdd.n7061 vdd.n7016 16.2531
R38940 vdd.n7061 vdd.n7060 16.2531
R38941 vdd.n7060 vdd.n7017 16.2531
R38942 vdd.n7049 vdd.n7017 16.2531
R38943 vdd.n7139 vdd.n7138 16.2531
R38944 vdd.n7138 vdd.n7118 16.2531
R38945 vdd.n7163 vdd.n7118 16.2531
R38946 vdd.n7163 vdd.n7162 16.2531
R38947 vdd.n7162 vdd.n7119 16.2531
R38948 vdd.n7151 vdd.n7119 16.2531
R38949 vdd.n7187 vdd.n7186 16.2531
R38950 vdd.n7186 vdd.n7166 16.2531
R38951 vdd.n7211 vdd.n7166 16.2531
R38952 vdd.n7211 vdd.n7210 16.2531
R38953 vdd.n7210 vdd.n7167 16.2531
R38954 vdd.n7199 vdd.n7167 16.2531
R38955 vdd.n7235 vdd.n7234 16.2531
R38956 vdd.n7234 vdd.n7214 16.2531
R38957 vdd.n7259 vdd.n7214 16.2531
R38958 vdd.n7259 vdd.n7258 16.2531
R38959 vdd.n7258 vdd.n7215 16.2531
R38960 vdd.n7247 vdd.n7215 16.2531
R38961 vdd.n7283 vdd.n7282 16.2531
R38962 vdd.n7282 vdd.n7262 16.2531
R38963 vdd.n7307 vdd.n7262 16.2531
R38964 vdd.n7307 vdd.n7306 16.2531
R38965 vdd.n7306 vdd.n7263 16.2531
R38966 vdd.n7295 vdd.n7263 16.2531
R38967 vdd.n7385 vdd.n7384 16.2531
R38968 vdd.n7384 vdd.n7364 16.2531
R38969 vdd.n7409 vdd.n7364 16.2531
R38970 vdd.n7409 vdd.n7408 16.2531
R38971 vdd.n7408 vdd.n7365 16.2531
R38972 vdd.n7397 vdd.n7365 16.2531
R38973 vdd.n8905 vdd.n8904 16.2531
R38974 vdd.n8904 vdd.n8884 16.2531
R38975 vdd.n8929 vdd.n8884 16.2531
R38976 vdd.n8929 vdd.n8928 16.2531
R38977 vdd.n8928 vdd.n8885 16.2531
R38978 vdd.n8917 vdd.n8885 16.2531
R38979 vdd.n7428 vdd.n7427 16.2531
R38980 vdd.n7427 vdd.n7412 16.2531
R38981 vdd.n7457 vdd.n7412 16.2531
R38982 vdd.n7457 vdd.n7456 16.2531
R38983 vdd.n7456 vdd.n7413 16.2531
R38984 vdd.n7445 vdd.n7413 16.2531
R38985 vdd.n7476 vdd.n7475 16.2531
R38986 vdd.n7475 vdd.n7460 16.2531
R38987 vdd.n7505 vdd.n7460 16.2531
R38988 vdd.n7505 vdd.n7504 16.2531
R38989 vdd.n7504 vdd.n7461 16.2531
R38990 vdd.n7493 vdd.n7461 16.2531
R38991 vdd.n7577 vdd.n7576 16.2531
R38992 vdd.n7576 vdd.n7561 16.2531
R38993 vdd.n7606 vdd.n7561 16.2531
R38994 vdd.n7606 vdd.n7605 16.2531
R38995 vdd.n7605 vdd.n7562 16.2531
R38996 vdd.n7594 vdd.n7562 16.2531
R38997 vdd.n7625 vdd.n7624 16.2531
R38998 vdd.n7624 vdd.n7609 16.2531
R38999 vdd.n7654 vdd.n7609 16.2531
R39000 vdd.n7654 vdd.n7653 16.2531
R39001 vdd.n7653 vdd.n7610 16.2531
R39002 vdd.n7642 vdd.n7610 16.2531
R39003 vdd.n7673 vdd.n7672 16.2531
R39004 vdd.n7672 vdd.n7657 16.2531
R39005 vdd.n7702 vdd.n7657 16.2531
R39006 vdd.n7702 vdd.n7701 16.2531
R39007 vdd.n7701 vdd.n7658 16.2531
R39008 vdd.n7690 vdd.n7658 16.2531
R39009 vdd.n7721 vdd.n7720 16.2531
R39010 vdd.n7720 vdd.n7705 16.2531
R39011 vdd.n7750 vdd.n7705 16.2531
R39012 vdd.n7750 vdd.n7749 16.2531
R39013 vdd.n7749 vdd.n7706 16.2531
R39014 vdd.n7738 vdd.n7706 16.2531
R39015 vdd.n7822 vdd.n7821 16.2531
R39016 vdd.n7821 vdd.n7806 16.2531
R39017 vdd.n7851 vdd.n7806 16.2531
R39018 vdd.n7851 vdd.n7850 16.2531
R39019 vdd.n7850 vdd.n7807 16.2531
R39020 vdd.n7839 vdd.n7807 16.2531
R39021 vdd.n6935 vdd.n6934 16.2531
R39022 vdd.n6934 vdd.n6919 16.2531
R39023 vdd.n6964 vdd.n6919 16.2531
R39024 vdd.n6964 vdd.n6963 16.2531
R39025 vdd.n6963 vdd.n6920 16.2531
R39026 vdd.n6952 vdd.n6920 16.2531
R39027 vdd.n7870 vdd.n7869 16.2531
R39028 vdd.n7869 vdd.n7854 16.2531
R39029 vdd.n7899 vdd.n7854 16.2531
R39030 vdd.n7899 vdd.n7898 16.2531
R39031 vdd.n7898 vdd.n7855 16.2531
R39032 vdd.n7887 vdd.n7855 16.2531
R39033 vdd.n7917 vdd.n7916 16.2531
R39034 vdd.n7916 vdd.n7901 16.2531
R39035 vdd.n7946 vdd.n7901 16.2531
R39036 vdd.n7946 vdd.n7945 16.2531
R39037 vdd.n7945 vdd.n7902 16.2531
R39038 vdd.n7934 vdd.n7902 16.2531
R39039 vdd.n7967 vdd.n7966 16.2531
R39040 vdd.n7966 vdd.n7951 16.2531
R39041 vdd.n7996 vdd.n7951 16.2531
R39042 vdd.n7996 vdd.n7995 16.2531
R39043 vdd.n7995 vdd.n7952 16.2531
R39044 vdd.n7984 vdd.n7952 16.2531
R39045 vdd.n8017 vdd.n8016 16.2531
R39046 vdd.n8016 vdd.n8001 16.2531
R39047 vdd.n8046 vdd.n8001 16.2531
R39048 vdd.n8046 vdd.n8045 16.2531
R39049 vdd.n8045 vdd.n8002 16.2531
R39050 vdd.n8034 vdd.n8002 16.2531
R39051 vdd.n8065 vdd.n8064 16.2531
R39052 vdd.n8064 vdd.n8049 16.2531
R39053 vdd.n8094 vdd.n8049 16.2531
R39054 vdd.n8094 vdd.n8093 16.2531
R39055 vdd.n8093 vdd.n8050 16.2531
R39056 vdd.n8082 vdd.n8050 16.2531
R39057 vdd.n7800 vdd.n7755 16.2531
R39058 vdd.n7789 vdd.n7755 16.2531
R39059 vdd.n7789 vdd.n7788 16.2531
R39060 vdd.n7773 vdd.n7766 16.2531
R39061 vdd.n7774 vdd.n7773 16.2531
R39062 vdd.n8116 vdd.n8115 16.2531
R39063 vdd.n8115 vdd.n8100 16.2531
R39064 vdd.n8145 vdd.n8100 16.2531
R39065 vdd.n8145 vdd.n8144 16.2531
R39066 vdd.n8144 vdd.n8101 16.2531
R39067 vdd.n8133 vdd.n8101 16.2531
R39068 vdd.n8163 vdd.n8162 16.2531
R39069 vdd.n8162 vdd.n8147 16.2531
R39070 vdd.n8192 vdd.n8147 16.2531
R39071 vdd.n8192 vdd.n8191 16.2531
R39072 vdd.n8191 vdd.n8148 16.2531
R39073 vdd.n8180 vdd.n8148 16.2531
R39074 vdd.n8211 vdd.n8210 16.2531
R39075 vdd.n8210 vdd.n8195 16.2531
R39076 vdd.n8240 vdd.n8195 16.2531
R39077 vdd.n8240 vdd.n8239 16.2531
R39078 vdd.n8239 vdd.n8196 16.2531
R39079 vdd.n8228 vdd.n8196 16.2531
R39080 vdd.n8262 vdd.n8261 16.2531
R39081 vdd.n8261 vdd.n8246 16.2531
R39082 vdd.n8291 vdd.n8246 16.2531
R39083 vdd.n8291 vdd.n8290 16.2531
R39084 vdd.n8290 vdd.n8247 16.2531
R39085 vdd.n8279 vdd.n8247 16.2531
R39086 vdd.n8312 vdd.n8311 16.2531
R39087 vdd.n8311 vdd.n8296 16.2531
R39088 vdd.n8341 vdd.n8296 16.2531
R39089 vdd.n8341 vdd.n8340 16.2531
R39090 vdd.n8340 vdd.n8297 16.2531
R39091 vdd.n8329 vdd.n8297 16.2531
R39092 vdd.n8360 vdd.n8359 16.2531
R39093 vdd.n8359 vdd.n8344 16.2531
R39094 vdd.n8389 vdd.n8344 16.2531
R39095 vdd.n8389 vdd.n8388 16.2531
R39096 vdd.n8388 vdd.n8345 16.2531
R39097 vdd.n8377 vdd.n8345 16.2531
R39098 vdd.n8410 vdd.n8409 16.2531
R39099 vdd.n8409 vdd.n8394 16.2531
R39100 vdd.n8439 vdd.n8394 16.2531
R39101 vdd.n8439 vdd.n8438 16.2531
R39102 vdd.n8438 vdd.n8395 16.2531
R39103 vdd.n8427 vdd.n8395 16.2531
R39104 vdd.n8457 vdd.n8456 16.2531
R39105 vdd.n8456 vdd.n8441 16.2531
R39106 vdd.n8486 vdd.n8441 16.2531
R39107 vdd.n8486 vdd.n8485 16.2531
R39108 vdd.n8485 vdd.n8442 16.2531
R39109 vdd.n8474 vdd.n8442 16.2531
R39110 vdd.n8507 vdd.n8506 16.2531
R39111 vdd.n8506 vdd.n8491 16.2531
R39112 vdd.n8536 vdd.n8491 16.2531
R39113 vdd.n8536 vdd.n8535 16.2531
R39114 vdd.n8535 vdd.n8492 16.2531
R39115 vdd.n8524 vdd.n8492 16.2531
R39116 vdd.n8557 vdd.n8556 16.2531
R39117 vdd.n8556 vdd.n8541 16.2531
R39118 vdd.n8586 vdd.n8541 16.2531
R39119 vdd.n8586 vdd.n8585 16.2531
R39120 vdd.n8585 vdd.n8542 16.2531
R39121 vdd.n8574 vdd.n8542 16.2531
R39122 vdd.n8605 vdd.n8604 16.2531
R39123 vdd.n8604 vdd.n8589 16.2531
R39124 vdd.n8634 vdd.n8589 16.2531
R39125 vdd.n8634 vdd.n8633 16.2531
R39126 vdd.n8633 vdd.n8590 16.2531
R39127 vdd.n8622 vdd.n8590 16.2531
R39128 vdd.n7555 vdd.n7510 16.2531
R39129 vdd.n7544 vdd.n7510 16.2531
R39130 vdd.n7544 vdd.n7543 16.2531
R39131 vdd.n7528 vdd.n7521 16.2531
R39132 vdd.n7529 vdd.n7528 16.2531
R39133 vdd.n8656 vdd.n8655 16.2531
R39134 vdd.n8655 vdd.n8640 16.2531
R39135 vdd.n8685 vdd.n8640 16.2531
R39136 vdd.n8685 vdd.n8684 16.2531
R39137 vdd.n8684 vdd.n8641 16.2531
R39138 vdd.n8673 vdd.n8641 16.2531
R39139 vdd.n8703 vdd.n8702 16.2531
R39140 vdd.n8702 vdd.n8687 16.2531
R39141 vdd.n8732 vdd.n8687 16.2531
R39142 vdd.n8732 vdd.n8731 16.2531
R39143 vdd.n8731 vdd.n8688 16.2531
R39144 vdd.n8720 vdd.n8688 16.2531
R39145 vdd.n8753 vdd.n8752 16.2531
R39146 vdd.n8752 vdd.n8737 16.2531
R39147 vdd.n8782 vdd.n8737 16.2531
R39148 vdd.n8782 vdd.n8781 16.2531
R39149 vdd.n8781 vdd.n8738 16.2531
R39150 vdd.n8770 vdd.n8738 16.2531
R39151 vdd.n8803 vdd.n8802 16.2531
R39152 vdd.n8802 vdd.n8787 16.2531
R39153 vdd.n8832 vdd.n8787 16.2531
R39154 vdd.n8832 vdd.n8831 16.2531
R39155 vdd.n8831 vdd.n8788 16.2531
R39156 vdd.n8820 vdd.n8788 16.2531
R39157 vdd.n8851 vdd.n8850 16.2531
R39158 vdd.n8850 vdd.n8835 16.2531
R39159 vdd.n8880 vdd.n8835 16.2531
R39160 vdd.n8880 vdd.n8879 16.2531
R39161 vdd.n8879 vdd.n8836 16.2531
R39162 vdd.n8868 vdd.n8836 16.2531
R39163 vdd.n9002 vdd.n9001 16.2531
R39164 vdd.n9001 vdd.n8981 16.2531
R39165 vdd.n9026 vdd.n8981 16.2531
R39166 vdd.n9026 vdd.n9025 16.2531
R39167 vdd.n9025 vdd.n8982 16.2531
R39168 vdd.n9014 vdd.n8982 16.2531
R39169 vdd.n8954 vdd.n8953 16.2531
R39170 vdd.n8953 vdd.n8933 16.2531
R39171 vdd.n8978 vdd.n8933 16.2531
R39172 vdd.n8978 vdd.n8977 16.2531
R39173 vdd.n8977 vdd.n8934 16.2531
R39174 vdd.n8966 vdd.n8934 16.2531
R39175 vdd.n9051 vdd.n9050 16.2531
R39176 vdd.n9050 vdd.n9030 16.2531
R39177 vdd.n9075 vdd.n9030 16.2531
R39178 vdd.n9075 vdd.n9074 16.2531
R39179 vdd.n9074 vdd.n9031 16.2531
R39180 vdd.n9063 vdd.n9031 16.2531
R39181 vdd.n9101 vdd.n9100 16.2531
R39182 vdd.n9100 vdd.n9080 16.2531
R39183 vdd.n9125 vdd.n9080 16.2531
R39184 vdd.n9125 vdd.n9124 16.2531
R39185 vdd.n9124 vdd.n9081 16.2531
R39186 vdd.n9113 vdd.n9081 16.2531
R39187 vdd.n9149 vdd.n9148 16.2531
R39188 vdd.n9148 vdd.n9128 16.2531
R39189 vdd.n9173 vdd.n9128 16.2531
R39190 vdd.n9173 vdd.n9172 16.2531
R39191 vdd.n9172 vdd.n9129 16.2531
R39192 vdd.n9161 vdd.n9129 16.2531
R39193 vdd.n7336 vdd.n7335 16.2531
R39194 vdd.n7337 vdd.n7336 16.2531
R39195 vdd.n7347 vdd.n7346 16.2531
R39196 vdd.n7348 vdd.n7347 16.2531
R39197 vdd.n7348 vdd.n7311 16.2531
R39198 vdd.n9297 vdd.n9296 16.2531
R39199 vdd.n9296 vdd.n9276 16.2531
R39200 vdd.n9321 vdd.n9276 16.2531
R39201 vdd.n9321 vdd.n9320 16.2531
R39202 vdd.n9320 vdd.n9277 16.2531
R39203 vdd.n9309 vdd.n9277 16.2531
R39204 vdd.n9248 vdd.n9247 16.2531
R39205 vdd.n9247 vdd.n9227 16.2531
R39206 vdd.n9272 vdd.n9227 16.2531
R39207 vdd.n9272 vdd.n9271 16.2531
R39208 vdd.n9271 vdd.n9228 16.2531
R39209 vdd.n9260 vdd.n9228 16.2531
R39210 vdd.n9200 vdd.n9199 16.2531
R39211 vdd.n9199 vdd.n9179 16.2531
R39212 vdd.n9224 vdd.n9179 16.2531
R39213 vdd.n9224 vdd.n9223 16.2531
R39214 vdd.n9223 vdd.n9180 16.2531
R39215 vdd.n9212 vdd.n9180 16.2531
R39216 vdd.n9346 vdd.n9345 16.2531
R39217 vdd.n9345 vdd.n9325 16.2531
R39218 vdd.n9370 vdd.n9325 16.2531
R39219 vdd.n9370 vdd.n9369 16.2531
R39220 vdd.n9369 vdd.n9326 16.2531
R39221 vdd.n9358 vdd.n9326 16.2531
R39222 vdd.n9396 vdd.n9395 16.2531
R39223 vdd.n9395 vdd.n9375 16.2531
R39224 vdd.n9420 vdd.n9375 16.2531
R39225 vdd.n9420 vdd.n9419 16.2531
R39226 vdd.n9419 vdd.n9376 16.2531
R39227 vdd.n9408 vdd.n9376 16.2531
R39228 vdd.n9444 vdd.n9443 16.2531
R39229 vdd.n9443 vdd.n9423 16.2531
R39230 vdd.n9468 vdd.n9423 16.2531
R39231 vdd.n9468 vdd.n9467 16.2531
R39232 vdd.n9467 vdd.n9424 16.2531
R39233 vdd.n9456 vdd.n9424 16.2531
R39234 vdd.n9542 vdd.n9541 16.2531
R39235 vdd.n9541 vdd.n9521 16.2531
R39236 vdd.n9566 vdd.n9521 16.2531
R39237 vdd.n9566 vdd.n9565 16.2531
R39238 vdd.n9565 vdd.n9522 16.2531
R39239 vdd.n9554 vdd.n9522 16.2531
R39240 vdd.n9494 vdd.n9493 16.2531
R39241 vdd.n9493 vdd.n9473 16.2531
R39242 vdd.n9518 vdd.n9473 16.2531
R39243 vdd.n9518 vdd.n9517 16.2531
R39244 vdd.n9517 vdd.n9474 16.2531
R39245 vdd.n9506 vdd.n9474 16.2531
R39246 vdd.n9591 vdd.n9590 16.2531
R39247 vdd.n9590 vdd.n9570 16.2531
R39248 vdd.n9615 vdd.n9570 16.2531
R39249 vdd.n9615 vdd.n9614 16.2531
R39250 vdd.n9614 vdd.n9571 16.2531
R39251 vdd.n9603 vdd.n9571 16.2531
R39252 vdd.n9641 vdd.n9640 16.2531
R39253 vdd.n9640 vdd.n9620 16.2531
R39254 vdd.n9665 vdd.n9620 16.2531
R39255 vdd.n9665 vdd.n9664 16.2531
R39256 vdd.n9664 vdd.n9621 16.2531
R39257 vdd.n9653 vdd.n9621 16.2531
R39258 vdd.n9689 vdd.n9688 16.2531
R39259 vdd.n9688 vdd.n9668 16.2531
R39260 vdd.n9713 vdd.n9668 16.2531
R39261 vdd.n9713 vdd.n9712 16.2531
R39262 vdd.n9712 vdd.n9669 16.2531
R39263 vdd.n9701 vdd.n9669 16.2531
R39264 vdd.n7090 vdd.n7089 16.2531
R39265 vdd.n7091 vdd.n7090 16.2531
R39266 vdd.n7101 vdd.n7100 16.2531
R39267 vdd.n7102 vdd.n7101 16.2531
R39268 vdd.n7102 vdd.n7065 16.2531
R39269 vdd.n9788 vdd.n9787 16.2531
R39270 vdd.n9787 vdd.n9767 16.2531
R39271 vdd.n9812 vdd.n9767 16.2531
R39272 vdd.n9812 vdd.n9811 16.2531
R39273 vdd.n9811 vdd.n9768 16.2531
R39274 vdd.n9800 vdd.n9768 16.2531
R39275 vdd.n9740 vdd.n9739 16.2531
R39276 vdd.n9739 vdd.n9719 16.2531
R39277 vdd.n9764 vdd.n9719 16.2531
R39278 vdd.n9764 vdd.n9763 16.2531
R39279 vdd.n9763 vdd.n9720 16.2531
R39280 vdd.n9752 vdd.n9720 16.2531
R39281 vdd.n9837 vdd.n9836 16.2531
R39282 vdd.n9836 vdd.n9816 16.2531
R39283 vdd.n9861 vdd.n9816 16.2531
R39284 vdd.n9861 vdd.n9860 16.2531
R39285 vdd.n9860 vdd.n9817 16.2531
R39286 vdd.n9849 vdd.n9817 16.2531
R39287 vdd.n9887 vdd.n9886 16.2531
R39288 vdd.n9886 vdd.n9866 16.2531
R39289 vdd.n9911 vdd.n9866 16.2531
R39290 vdd.n9911 vdd.n9910 16.2531
R39291 vdd.n9910 vdd.n9867 16.2531
R39292 vdd.n9899 vdd.n9867 16.2531
R39293 vdd.n9935 vdd.n9934 16.2531
R39294 vdd.n9934 vdd.n9914 16.2531
R39295 vdd.n9959 vdd.n9914 16.2531
R39296 vdd.n9959 vdd.n9958 16.2531
R39297 vdd.n9958 vdd.n9915 16.2531
R39298 vdd.n9947 vdd.n9915 16.2531
R39299 vdd.n3847 vdd.n3846 16.2531
R39300 vdd.n3846 vdd.n3826 16.2531
R39301 vdd.n3871 vdd.n3826 16.2531
R39302 vdd.n3871 vdd.n3870 16.2531
R39303 vdd.n3870 vdd.n3827 16.2531
R39304 vdd.n3859 vdd.n3827 16.2531
R39305 vdd.n3895 vdd.n3894 16.2531
R39306 vdd.n3894 vdd.n3874 16.2531
R39307 vdd.n3919 vdd.n3874 16.2531
R39308 vdd.n3919 vdd.n3918 16.2531
R39309 vdd.n3918 vdd.n3875 16.2531
R39310 vdd.n3907 vdd.n3875 16.2531
R39311 vdd.n3997 vdd.n3996 16.2531
R39312 vdd.n3996 vdd.n3976 16.2531
R39313 vdd.n4021 vdd.n3976 16.2531
R39314 vdd.n4021 vdd.n4020 16.2531
R39315 vdd.n4020 vdd.n3977 16.2531
R39316 vdd.n4009 vdd.n3977 16.2531
R39317 vdd.n4045 vdd.n4044 16.2531
R39318 vdd.n4044 vdd.n4024 16.2531
R39319 vdd.n4069 vdd.n4024 16.2531
R39320 vdd.n4069 vdd.n4068 16.2531
R39321 vdd.n4068 vdd.n4025 16.2531
R39322 vdd.n4057 vdd.n4025 16.2531
R39323 vdd.n4093 vdd.n4092 16.2531
R39324 vdd.n4092 vdd.n4072 16.2531
R39325 vdd.n4117 vdd.n4072 16.2531
R39326 vdd.n4117 vdd.n4116 16.2531
R39327 vdd.n4116 vdd.n4073 16.2531
R39328 vdd.n4105 vdd.n4073 16.2531
R39329 vdd.n4141 vdd.n4140 16.2531
R39330 vdd.n4140 vdd.n4120 16.2531
R39331 vdd.n4165 vdd.n4120 16.2531
R39332 vdd.n4165 vdd.n4164 16.2531
R39333 vdd.n4164 vdd.n4121 16.2531
R39334 vdd.n4153 vdd.n4121 16.2531
R39335 vdd.n4243 vdd.n4242 16.2531
R39336 vdd.n4242 vdd.n4222 16.2531
R39337 vdd.n4267 vdd.n4222 16.2531
R39338 vdd.n4267 vdd.n4266 16.2531
R39339 vdd.n4266 vdd.n4223 16.2531
R39340 vdd.n4255 vdd.n4223 16.2531
R39341 vdd.n5763 vdd.n5762 16.2531
R39342 vdd.n5762 vdd.n5742 16.2531
R39343 vdd.n5787 vdd.n5742 16.2531
R39344 vdd.n5787 vdd.n5786 16.2531
R39345 vdd.n5786 vdd.n5743 16.2531
R39346 vdd.n5775 vdd.n5743 16.2531
R39347 vdd.n4286 vdd.n4285 16.2531
R39348 vdd.n4285 vdd.n4270 16.2531
R39349 vdd.n4315 vdd.n4270 16.2531
R39350 vdd.n4315 vdd.n4314 16.2531
R39351 vdd.n4314 vdd.n4271 16.2531
R39352 vdd.n4303 vdd.n4271 16.2531
R39353 vdd.n4334 vdd.n4333 16.2531
R39354 vdd.n4333 vdd.n4318 16.2531
R39355 vdd.n4363 vdd.n4318 16.2531
R39356 vdd.n4363 vdd.n4362 16.2531
R39357 vdd.n4362 vdd.n4319 16.2531
R39358 vdd.n4351 vdd.n4319 16.2531
R39359 vdd.n4435 vdd.n4434 16.2531
R39360 vdd.n4434 vdd.n4419 16.2531
R39361 vdd.n4464 vdd.n4419 16.2531
R39362 vdd.n4464 vdd.n4463 16.2531
R39363 vdd.n4463 vdd.n4420 16.2531
R39364 vdd.n4452 vdd.n4420 16.2531
R39365 vdd.n4483 vdd.n4482 16.2531
R39366 vdd.n4482 vdd.n4467 16.2531
R39367 vdd.n4512 vdd.n4467 16.2531
R39368 vdd.n4512 vdd.n4511 16.2531
R39369 vdd.n4511 vdd.n4468 16.2531
R39370 vdd.n4500 vdd.n4468 16.2531
R39371 vdd.n4531 vdd.n4530 16.2531
R39372 vdd.n4530 vdd.n4515 16.2531
R39373 vdd.n4560 vdd.n4515 16.2531
R39374 vdd.n4560 vdd.n4559 16.2531
R39375 vdd.n4559 vdd.n4516 16.2531
R39376 vdd.n4548 vdd.n4516 16.2531
R39377 vdd.n4579 vdd.n4578 16.2531
R39378 vdd.n4578 vdd.n4563 16.2531
R39379 vdd.n4608 vdd.n4563 16.2531
R39380 vdd.n4608 vdd.n4607 16.2531
R39381 vdd.n4607 vdd.n4564 16.2531
R39382 vdd.n4596 vdd.n4564 16.2531
R39383 vdd.n4680 vdd.n4679 16.2531
R39384 vdd.n4679 vdd.n4664 16.2531
R39385 vdd.n4709 vdd.n4664 16.2531
R39386 vdd.n4709 vdd.n4708 16.2531
R39387 vdd.n4708 vdd.n4665 16.2531
R39388 vdd.n4697 vdd.n4665 16.2531
R39389 vdd.n3793 vdd.n3792 16.2531
R39390 vdd.n3792 vdd.n3777 16.2531
R39391 vdd.n3822 vdd.n3777 16.2531
R39392 vdd.n3822 vdd.n3821 16.2531
R39393 vdd.n3821 vdd.n3778 16.2531
R39394 vdd.n3810 vdd.n3778 16.2531
R39395 vdd.n4728 vdd.n4727 16.2531
R39396 vdd.n4727 vdd.n4712 16.2531
R39397 vdd.n4757 vdd.n4712 16.2531
R39398 vdd.n4757 vdd.n4756 16.2531
R39399 vdd.n4756 vdd.n4713 16.2531
R39400 vdd.n4745 vdd.n4713 16.2531
R39401 vdd.n4775 vdd.n4774 16.2531
R39402 vdd.n4774 vdd.n4759 16.2531
R39403 vdd.n4804 vdd.n4759 16.2531
R39404 vdd.n4804 vdd.n4803 16.2531
R39405 vdd.n4803 vdd.n4760 16.2531
R39406 vdd.n4792 vdd.n4760 16.2531
R39407 vdd.n4825 vdd.n4824 16.2531
R39408 vdd.n4824 vdd.n4809 16.2531
R39409 vdd.n4854 vdd.n4809 16.2531
R39410 vdd.n4854 vdd.n4853 16.2531
R39411 vdd.n4853 vdd.n4810 16.2531
R39412 vdd.n4842 vdd.n4810 16.2531
R39413 vdd.n4875 vdd.n4874 16.2531
R39414 vdd.n4874 vdd.n4859 16.2531
R39415 vdd.n4904 vdd.n4859 16.2531
R39416 vdd.n4904 vdd.n4903 16.2531
R39417 vdd.n4903 vdd.n4860 16.2531
R39418 vdd.n4892 vdd.n4860 16.2531
R39419 vdd.n4923 vdd.n4922 16.2531
R39420 vdd.n4922 vdd.n4907 16.2531
R39421 vdd.n4952 vdd.n4907 16.2531
R39422 vdd.n4952 vdd.n4951 16.2531
R39423 vdd.n4951 vdd.n4908 16.2531
R39424 vdd.n4940 vdd.n4908 16.2531
R39425 vdd.n4658 vdd.n4613 16.2531
R39426 vdd.n4647 vdd.n4613 16.2531
R39427 vdd.n4647 vdd.n4646 16.2531
R39428 vdd.n4631 vdd.n4624 16.2531
R39429 vdd.n4632 vdd.n4631 16.2531
R39430 vdd.n4974 vdd.n4973 16.2531
R39431 vdd.n4973 vdd.n4958 16.2531
R39432 vdd.n5003 vdd.n4958 16.2531
R39433 vdd.n5003 vdd.n5002 16.2531
R39434 vdd.n5002 vdd.n4959 16.2531
R39435 vdd.n4991 vdd.n4959 16.2531
R39436 vdd.n5021 vdd.n5020 16.2531
R39437 vdd.n5020 vdd.n5005 16.2531
R39438 vdd.n5050 vdd.n5005 16.2531
R39439 vdd.n5050 vdd.n5049 16.2531
R39440 vdd.n5049 vdd.n5006 16.2531
R39441 vdd.n5038 vdd.n5006 16.2531
R39442 vdd.n5069 vdd.n5068 16.2531
R39443 vdd.n5068 vdd.n5053 16.2531
R39444 vdd.n5098 vdd.n5053 16.2531
R39445 vdd.n5098 vdd.n5097 16.2531
R39446 vdd.n5097 vdd.n5054 16.2531
R39447 vdd.n5086 vdd.n5054 16.2531
R39448 vdd.n5120 vdd.n5119 16.2531
R39449 vdd.n5119 vdd.n5104 16.2531
R39450 vdd.n5149 vdd.n5104 16.2531
R39451 vdd.n5149 vdd.n5148 16.2531
R39452 vdd.n5148 vdd.n5105 16.2531
R39453 vdd.n5137 vdd.n5105 16.2531
R39454 vdd.n5170 vdd.n5169 16.2531
R39455 vdd.n5169 vdd.n5154 16.2531
R39456 vdd.n5199 vdd.n5154 16.2531
R39457 vdd.n5199 vdd.n5198 16.2531
R39458 vdd.n5198 vdd.n5155 16.2531
R39459 vdd.n5187 vdd.n5155 16.2531
R39460 vdd.n5218 vdd.n5217 16.2531
R39461 vdd.n5217 vdd.n5202 16.2531
R39462 vdd.n5247 vdd.n5202 16.2531
R39463 vdd.n5247 vdd.n5246 16.2531
R39464 vdd.n5246 vdd.n5203 16.2531
R39465 vdd.n5235 vdd.n5203 16.2531
R39466 vdd.n5268 vdd.n5267 16.2531
R39467 vdd.n5267 vdd.n5252 16.2531
R39468 vdd.n5297 vdd.n5252 16.2531
R39469 vdd.n5297 vdd.n5296 16.2531
R39470 vdd.n5296 vdd.n5253 16.2531
R39471 vdd.n5285 vdd.n5253 16.2531
R39472 vdd.n5315 vdd.n5314 16.2531
R39473 vdd.n5314 vdd.n5299 16.2531
R39474 vdd.n5344 vdd.n5299 16.2531
R39475 vdd.n5344 vdd.n5343 16.2531
R39476 vdd.n5343 vdd.n5300 16.2531
R39477 vdd.n5332 vdd.n5300 16.2531
R39478 vdd.n5365 vdd.n5364 16.2531
R39479 vdd.n5364 vdd.n5349 16.2531
R39480 vdd.n5394 vdd.n5349 16.2531
R39481 vdd.n5394 vdd.n5393 16.2531
R39482 vdd.n5393 vdd.n5350 16.2531
R39483 vdd.n5382 vdd.n5350 16.2531
R39484 vdd.n5415 vdd.n5414 16.2531
R39485 vdd.n5414 vdd.n5399 16.2531
R39486 vdd.n5444 vdd.n5399 16.2531
R39487 vdd.n5444 vdd.n5443 16.2531
R39488 vdd.n5443 vdd.n5400 16.2531
R39489 vdd.n5432 vdd.n5400 16.2531
R39490 vdd.n5463 vdd.n5462 16.2531
R39491 vdd.n5462 vdd.n5447 16.2531
R39492 vdd.n5492 vdd.n5447 16.2531
R39493 vdd.n5492 vdd.n5491 16.2531
R39494 vdd.n5491 vdd.n5448 16.2531
R39495 vdd.n5480 vdd.n5448 16.2531
R39496 vdd.n4413 vdd.n4368 16.2531
R39497 vdd.n4402 vdd.n4368 16.2531
R39498 vdd.n4402 vdd.n4401 16.2531
R39499 vdd.n4386 vdd.n4379 16.2531
R39500 vdd.n4387 vdd.n4386 16.2531
R39501 vdd.n5514 vdd.n5513 16.2531
R39502 vdd.n5513 vdd.n5498 16.2531
R39503 vdd.n5543 vdd.n5498 16.2531
R39504 vdd.n5543 vdd.n5542 16.2531
R39505 vdd.n5542 vdd.n5499 16.2531
R39506 vdd.n5531 vdd.n5499 16.2531
R39507 vdd.n5561 vdd.n5560 16.2531
R39508 vdd.n5560 vdd.n5545 16.2531
R39509 vdd.n5590 vdd.n5545 16.2531
R39510 vdd.n5590 vdd.n5589 16.2531
R39511 vdd.n5589 vdd.n5546 16.2531
R39512 vdd.n5578 vdd.n5546 16.2531
R39513 vdd.n5611 vdd.n5610 16.2531
R39514 vdd.n5610 vdd.n5595 16.2531
R39515 vdd.n5640 vdd.n5595 16.2531
R39516 vdd.n5640 vdd.n5639 16.2531
R39517 vdd.n5639 vdd.n5596 16.2531
R39518 vdd.n5628 vdd.n5596 16.2531
R39519 vdd.n5661 vdd.n5660 16.2531
R39520 vdd.n5660 vdd.n5645 16.2531
R39521 vdd.n5690 vdd.n5645 16.2531
R39522 vdd.n5690 vdd.n5689 16.2531
R39523 vdd.n5689 vdd.n5646 16.2531
R39524 vdd.n5678 vdd.n5646 16.2531
R39525 vdd.n5709 vdd.n5708 16.2531
R39526 vdd.n5708 vdd.n5693 16.2531
R39527 vdd.n5738 vdd.n5693 16.2531
R39528 vdd.n5738 vdd.n5737 16.2531
R39529 vdd.n5737 vdd.n5694 16.2531
R39530 vdd.n5726 vdd.n5694 16.2531
R39531 vdd.n5860 vdd.n5859 16.2531
R39532 vdd.n5859 vdd.n5839 16.2531
R39533 vdd.n5884 vdd.n5839 16.2531
R39534 vdd.n5884 vdd.n5883 16.2531
R39535 vdd.n5883 vdd.n5840 16.2531
R39536 vdd.n5872 vdd.n5840 16.2531
R39537 vdd.n5812 vdd.n5811 16.2531
R39538 vdd.n5811 vdd.n5791 16.2531
R39539 vdd.n5836 vdd.n5791 16.2531
R39540 vdd.n5836 vdd.n5835 16.2531
R39541 vdd.n5835 vdd.n5792 16.2531
R39542 vdd.n5824 vdd.n5792 16.2531
R39543 vdd.n5909 vdd.n5908 16.2531
R39544 vdd.n5908 vdd.n5888 16.2531
R39545 vdd.n5933 vdd.n5888 16.2531
R39546 vdd.n5933 vdd.n5932 16.2531
R39547 vdd.n5932 vdd.n5889 16.2531
R39548 vdd.n5921 vdd.n5889 16.2531
R39549 vdd.n5959 vdd.n5958 16.2531
R39550 vdd.n5958 vdd.n5938 16.2531
R39551 vdd.n5983 vdd.n5938 16.2531
R39552 vdd.n5983 vdd.n5982 16.2531
R39553 vdd.n5982 vdd.n5939 16.2531
R39554 vdd.n5971 vdd.n5939 16.2531
R39555 vdd.n6007 vdd.n6006 16.2531
R39556 vdd.n6006 vdd.n5986 16.2531
R39557 vdd.n6031 vdd.n5986 16.2531
R39558 vdd.n6031 vdd.n6030 16.2531
R39559 vdd.n6030 vdd.n5987 16.2531
R39560 vdd.n6019 vdd.n5987 16.2531
R39561 vdd.n4194 vdd.n4193 16.2531
R39562 vdd.n4195 vdd.n4194 16.2531
R39563 vdd.n4205 vdd.n4204 16.2531
R39564 vdd.n4206 vdd.n4205 16.2531
R39565 vdd.n4206 vdd.n4169 16.2531
R39566 vdd.n6155 vdd.n6154 16.2531
R39567 vdd.n6154 vdd.n6134 16.2531
R39568 vdd.n6179 vdd.n6134 16.2531
R39569 vdd.n6179 vdd.n6178 16.2531
R39570 vdd.n6178 vdd.n6135 16.2531
R39571 vdd.n6167 vdd.n6135 16.2531
R39572 vdd.n6106 vdd.n6105 16.2531
R39573 vdd.n6105 vdd.n6085 16.2531
R39574 vdd.n6130 vdd.n6085 16.2531
R39575 vdd.n6130 vdd.n6129 16.2531
R39576 vdd.n6129 vdd.n6086 16.2531
R39577 vdd.n6118 vdd.n6086 16.2531
R39578 vdd.n6058 vdd.n6057 16.2531
R39579 vdd.n6057 vdd.n6037 16.2531
R39580 vdd.n6082 vdd.n6037 16.2531
R39581 vdd.n6082 vdd.n6081 16.2531
R39582 vdd.n6081 vdd.n6038 16.2531
R39583 vdd.n6070 vdd.n6038 16.2531
R39584 vdd.n6204 vdd.n6203 16.2531
R39585 vdd.n6203 vdd.n6183 16.2531
R39586 vdd.n6228 vdd.n6183 16.2531
R39587 vdd.n6228 vdd.n6227 16.2531
R39588 vdd.n6227 vdd.n6184 16.2531
R39589 vdd.n6216 vdd.n6184 16.2531
R39590 vdd.n6254 vdd.n6253 16.2531
R39591 vdd.n6253 vdd.n6233 16.2531
R39592 vdd.n6278 vdd.n6233 16.2531
R39593 vdd.n6278 vdd.n6277 16.2531
R39594 vdd.n6277 vdd.n6234 16.2531
R39595 vdd.n6266 vdd.n6234 16.2531
R39596 vdd.n6302 vdd.n6301 16.2531
R39597 vdd.n6301 vdd.n6281 16.2531
R39598 vdd.n6326 vdd.n6281 16.2531
R39599 vdd.n6326 vdd.n6325 16.2531
R39600 vdd.n6325 vdd.n6282 16.2531
R39601 vdd.n6314 vdd.n6282 16.2531
R39602 vdd.n6400 vdd.n6399 16.2531
R39603 vdd.n6399 vdd.n6379 16.2531
R39604 vdd.n6424 vdd.n6379 16.2531
R39605 vdd.n6424 vdd.n6423 16.2531
R39606 vdd.n6423 vdd.n6380 16.2531
R39607 vdd.n6412 vdd.n6380 16.2531
R39608 vdd.n6352 vdd.n6351 16.2531
R39609 vdd.n6351 vdd.n6331 16.2531
R39610 vdd.n6376 vdd.n6331 16.2531
R39611 vdd.n6376 vdd.n6375 16.2531
R39612 vdd.n6375 vdd.n6332 16.2531
R39613 vdd.n6364 vdd.n6332 16.2531
R39614 vdd.n6449 vdd.n6448 16.2531
R39615 vdd.n6448 vdd.n6428 16.2531
R39616 vdd.n6473 vdd.n6428 16.2531
R39617 vdd.n6473 vdd.n6472 16.2531
R39618 vdd.n6472 vdd.n6429 16.2531
R39619 vdd.n6461 vdd.n6429 16.2531
R39620 vdd.n6499 vdd.n6498 16.2531
R39621 vdd.n6498 vdd.n6478 16.2531
R39622 vdd.n6523 vdd.n6478 16.2531
R39623 vdd.n6523 vdd.n6522 16.2531
R39624 vdd.n6522 vdd.n6479 16.2531
R39625 vdd.n6511 vdd.n6479 16.2531
R39626 vdd.n6547 vdd.n6546 16.2531
R39627 vdd.n6546 vdd.n6526 16.2531
R39628 vdd.n6571 vdd.n6526 16.2531
R39629 vdd.n6571 vdd.n6570 16.2531
R39630 vdd.n6570 vdd.n6527 16.2531
R39631 vdd.n6559 vdd.n6527 16.2531
R39632 vdd.n3948 vdd.n3947 16.2531
R39633 vdd.n3949 vdd.n3948 16.2531
R39634 vdd.n3959 vdd.n3958 16.2531
R39635 vdd.n3960 vdd.n3959 16.2531
R39636 vdd.n3960 vdd.n3923 16.2531
R39637 vdd.n6646 vdd.n6645 16.2531
R39638 vdd.n6645 vdd.n6625 16.2531
R39639 vdd.n6670 vdd.n6625 16.2531
R39640 vdd.n6670 vdd.n6669 16.2531
R39641 vdd.n6669 vdd.n6626 16.2531
R39642 vdd.n6658 vdd.n6626 16.2531
R39643 vdd.n6598 vdd.n6597 16.2531
R39644 vdd.n6597 vdd.n6577 16.2531
R39645 vdd.n6622 vdd.n6577 16.2531
R39646 vdd.n6622 vdd.n6621 16.2531
R39647 vdd.n6621 vdd.n6578 16.2531
R39648 vdd.n6610 vdd.n6578 16.2531
R39649 vdd.n6695 vdd.n6694 16.2531
R39650 vdd.n6694 vdd.n6674 16.2531
R39651 vdd.n6719 vdd.n6674 16.2531
R39652 vdd.n6719 vdd.n6718 16.2531
R39653 vdd.n6718 vdd.n6675 16.2531
R39654 vdd.n6707 vdd.n6675 16.2531
R39655 vdd.n6745 vdd.n6744 16.2531
R39656 vdd.n6744 vdd.n6724 16.2531
R39657 vdd.n6769 vdd.n6724 16.2531
R39658 vdd.n6769 vdd.n6768 16.2531
R39659 vdd.n6768 vdd.n6725 16.2531
R39660 vdd.n6757 vdd.n6725 16.2531
R39661 vdd.n6793 vdd.n6792 16.2531
R39662 vdd.n6792 vdd.n6772 16.2531
R39663 vdd.n6817 vdd.n6772 16.2531
R39664 vdd.n6817 vdd.n6816 16.2531
R39665 vdd.n6816 vdd.n6773 16.2531
R39666 vdd.n6805 vdd.n6773 16.2531
R39667 vdd.n705 vdd.n704 16.2531
R39668 vdd.n704 vdd.n684 16.2531
R39669 vdd.n729 vdd.n684 16.2531
R39670 vdd.n729 vdd.n728 16.2531
R39671 vdd.n728 vdd.n685 16.2531
R39672 vdd.n717 vdd.n685 16.2531
R39673 vdd.n753 vdd.n752 16.2531
R39674 vdd.n752 vdd.n732 16.2531
R39675 vdd.n777 vdd.n732 16.2531
R39676 vdd.n777 vdd.n776 16.2531
R39677 vdd.n776 vdd.n733 16.2531
R39678 vdd.n765 vdd.n733 16.2531
R39679 vdd.n855 vdd.n854 16.2531
R39680 vdd.n854 vdd.n834 16.2531
R39681 vdd.n879 vdd.n834 16.2531
R39682 vdd.n879 vdd.n878 16.2531
R39683 vdd.n878 vdd.n835 16.2531
R39684 vdd.n867 vdd.n835 16.2531
R39685 vdd.n903 vdd.n902 16.2531
R39686 vdd.n902 vdd.n882 16.2531
R39687 vdd.n927 vdd.n882 16.2531
R39688 vdd.n927 vdd.n926 16.2531
R39689 vdd.n926 vdd.n883 16.2531
R39690 vdd.n915 vdd.n883 16.2531
R39691 vdd.n951 vdd.n950 16.2531
R39692 vdd.n950 vdd.n930 16.2531
R39693 vdd.n975 vdd.n930 16.2531
R39694 vdd.n975 vdd.n974 16.2531
R39695 vdd.n974 vdd.n931 16.2531
R39696 vdd.n963 vdd.n931 16.2531
R39697 vdd.n999 vdd.n998 16.2531
R39698 vdd.n998 vdd.n978 16.2531
R39699 vdd.n1023 vdd.n978 16.2531
R39700 vdd.n1023 vdd.n1022 16.2531
R39701 vdd.n1022 vdd.n979 16.2531
R39702 vdd.n1011 vdd.n979 16.2531
R39703 vdd.n1101 vdd.n1100 16.2531
R39704 vdd.n1100 vdd.n1080 16.2531
R39705 vdd.n1125 vdd.n1080 16.2531
R39706 vdd.n1125 vdd.n1124 16.2531
R39707 vdd.n1124 vdd.n1081 16.2531
R39708 vdd.n1113 vdd.n1081 16.2531
R39709 vdd.n2621 vdd.n2620 16.2531
R39710 vdd.n2620 vdd.n2600 16.2531
R39711 vdd.n2645 vdd.n2600 16.2531
R39712 vdd.n2645 vdd.n2644 16.2531
R39713 vdd.n2644 vdd.n2601 16.2531
R39714 vdd.n2633 vdd.n2601 16.2531
R39715 vdd.n1144 vdd.n1143 16.2531
R39716 vdd.n1143 vdd.n1128 16.2531
R39717 vdd.n1173 vdd.n1128 16.2531
R39718 vdd.n1173 vdd.n1172 16.2531
R39719 vdd.n1172 vdd.n1129 16.2531
R39720 vdd.n1161 vdd.n1129 16.2531
R39721 vdd.n1192 vdd.n1191 16.2531
R39722 vdd.n1191 vdd.n1176 16.2531
R39723 vdd.n1221 vdd.n1176 16.2531
R39724 vdd.n1221 vdd.n1220 16.2531
R39725 vdd.n1220 vdd.n1177 16.2531
R39726 vdd.n1209 vdd.n1177 16.2531
R39727 vdd.n1293 vdd.n1292 16.2531
R39728 vdd.n1292 vdd.n1277 16.2531
R39729 vdd.n1322 vdd.n1277 16.2531
R39730 vdd.n1322 vdd.n1321 16.2531
R39731 vdd.n1321 vdd.n1278 16.2531
R39732 vdd.n1310 vdd.n1278 16.2531
R39733 vdd.n1341 vdd.n1340 16.2531
R39734 vdd.n1340 vdd.n1325 16.2531
R39735 vdd.n1370 vdd.n1325 16.2531
R39736 vdd.n1370 vdd.n1369 16.2531
R39737 vdd.n1369 vdd.n1326 16.2531
R39738 vdd.n1358 vdd.n1326 16.2531
R39739 vdd.n1389 vdd.n1388 16.2531
R39740 vdd.n1388 vdd.n1373 16.2531
R39741 vdd.n1418 vdd.n1373 16.2531
R39742 vdd.n1418 vdd.n1417 16.2531
R39743 vdd.n1417 vdd.n1374 16.2531
R39744 vdd.n1406 vdd.n1374 16.2531
R39745 vdd.n1437 vdd.n1436 16.2531
R39746 vdd.n1436 vdd.n1421 16.2531
R39747 vdd.n1466 vdd.n1421 16.2531
R39748 vdd.n1466 vdd.n1465 16.2531
R39749 vdd.n1465 vdd.n1422 16.2531
R39750 vdd.n1454 vdd.n1422 16.2531
R39751 vdd.n1538 vdd.n1537 16.2531
R39752 vdd.n1537 vdd.n1522 16.2531
R39753 vdd.n1567 vdd.n1522 16.2531
R39754 vdd.n1567 vdd.n1566 16.2531
R39755 vdd.n1566 vdd.n1523 16.2531
R39756 vdd.n1555 vdd.n1523 16.2531
R39757 vdd.n651 vdd.n650 16.2531
R39758 vdd.n650 vdd.n635 16.2531
R39759 vdd.n680 vdd.n635 16.2531
R39760 vdd.n680 vdd.n679 16.2531
R39761 vdd.n679 vdd.n636 16.2531
R39762 vdd.n668 vdd.n636 16.2531
R39763 vdd.n1586 vdd.n1585 16.2531
R39764 vdd.n1585 vdd.n1570 16.2531
R39765 vdd.n1615 vdd.n1570 16.2531
R39766 vdd.n1615 vdd.n1614 16.2531
R39767 vdd.n1614 vdd.n1571 16.2531
R39768 vdd.n1603 vdd.n1571 16.2531
R39769 vdd.n1633 vdd.n1632 16.2531
R39770 vdd.n1632 vdd.n1617 16.2531
R39771 vdd.n1662 vdd.n1617 16.2531
R39772 vdd.n1662 vdd.n1661 16.2531
R39773 vdd.n1661 vdd.n1618 16.2531
R39774 vdd.n1650 vdd.n1618 16.2531
R39775 vdd.n1683 vdd.n1682 16.2531
R39776 vdd.n1682 vdd.n1667 16.2531
R39777 vdd.n1712 vdd.n1667 16.2531
R39778 vdd.n1712 vdd.n1711 16.2531
R39779 vdd.n1711 vdd.n1668 16.2531
R39780 vdd.n1700 vdd.n1668 16.2531
R39781 vdd.n1733 vdd.n1732 16.2531
R39782 vdd.n1732 vdd.n1717 16.2531
R39783 vdd.n1762 vdd.n1717 16.2531
R39784 vdd.n1762 vdd.n1761 16.2531
R39785 vdd.n1761 vdd.n1718 16.2531
R39786 vdd.n1750 vdd.n1718 16.2531
R39787 vdd.n1781 vdd.n1780 16.2531
R39788 vdd.n1780 vdd.n1765 16.2531
R39789 vdd.n1810 vdd.n1765 16.2531
R39790 vdd.n1810 vdd.n1809 16.2531
R39791 vdd.n1809 vdd.n1766 16.2531
R39792 vdd.n1798 vdd.n1766 16.2531
R39793 vdd.n1516 vdd.n1471 16.2531
R39794 vdd.n1505 vdd.n1471 16.2531
R39795 vdd.n1505 vdd.n1504 16.2531
R39796 vdd.n1489 vdd.n1482 16.2531
R39797 vdd.n1490 vdd.n1489 16.2531
R39798 vdd.n1832 vdd.n1831 16.2531
R39799 vdd.n1831 vdd.n1816 16.2531
R39800 vdd.n1861 vdd.n1816 16.2531
R39801 vdd.n1861 vdd.n1860 16.2531
R39802 vdd.n1860 vdd.n1817 16.2531
R39803 vdd.n1849 vdd.n1817 16.2531
R39804 vdd.n1879 vdd.n1878 16.2531
R39805 vdd.n1878 vdd.n1863 16.2531
R39806 vdd.n1908 vdd.n1863 16.2531
R39807 vdd.n1908 vdd.n1907 16.2531
R39808 vdd.n1907 vdd.n1864 16.2531
R39809 vdd.n1896 vdd.n1864 16.2531
R39810 vdd.n1927 vdd.n1926 16.2531
R39811 vdd.n1926 vdd.n1911 16.2531
R39812 vdd.n1956 vdd.n1911 16.2531
R39813 vdd.n1956 vdd.n1955 16.2531
R39814 vdd.n1955 vdd.n1912 16.2531
R39815 vdd.n1944 vdd.n1912 16.2531
R39816 vdd.n1978 vdd.n1977 16.2531
R39817 vdd.n1977 vdd.n1962 16.2531
R39818 vdd.n2007 vdd.n1962 16.2531
R39819 vdd.n2007 vdd.n2006 16.2531
R39820 vdd.n2006 vdd.n1963 16.2531
R39821 vdd.n1995 vdd.n1963 16.2531
R39822 vdd.n2028 vdd.n2027 16.2531
R39823 vdd.n2027 vdd.n2012 16.2531
R39824 vdd.n2057 vdd.n2012 16.2531
R39825 vdd.n2057 vdd.n2056 16.2531
R39826 vdd.n2056 vdd.n2013 16.2531
R39827 vdd.n2045 vdd.n2013 16.2531
R39828 vdd.n2076 vdd.n2075 16.2531
R39829 vdd.n2075 vdd.n2060 16.2531
R39830 vdd.n2105 vdd.n2060 16.2531
R39831 vdd.n2105 vdd.n2104 16.2531
R39832 vdd.n2104 vdd.n2061 16.2531
R39833 vdd.n2093 vdd.n2061 16.2531
R39834 vdd.n2126 vdd.n2125 16.2531
R39835 vdd.n2125 vdd.n2110 16.2531
R39836 vdd.n2155 vdd.n2110 16.2531
R39837 vdd.n2155 vdd.n2154 16.2531
R39838 vdd.n2154 vdd.n2111 16.2531
R39839 vdd.n2143 vdd.n2111 16.2531
R39840 vdd.n2173 vdd.n2172 16.2531
R39841 vdd.n2172 vdd.n2157 16.2531
R39842 vdd.n2202 vdd.n2157 16.2531
R39843 vdd.n2202 vdd.n2201 16.2531
R39844 vdd.n2201 vdd.n2158 16.2531
R39845 vdd.n2190 vdd.n2158 16.2531
R39846 vdd.n2223 vdd.n2222 16.2531
R39847 vdd.n2222 vdd.n2207 16.2531
R39848 vdd.n2252 vdd.n2207 16.2531
R39849 vdd.n2252 vdd.n2251 16.2531
R39850 vdd.n2251 vdd.n2208 16.2531
R39851 vdd.n2240 vdd.n2208 16.2531
R39852 vdd.n2273 vdd.n2272 16.2531
R39853 vdd.n2272 vdd.n2257 16.2531
R39854 vdd.n2302 vdd.n2257 16.2531
R39855 vdd.n2302 vdd.n2301 16.2531
R39856 vdd.n2301 vdd.n2258 16.2531
R39857 vdd.n2290 vdd.n2258 16.2531
R39858 vdd.n2321 vdd.n2320 16.2531
R39859 vdd.n2320 vdd.n2305 16.2531
R39860 vdd.n2350 vdd.n2305 16.2531
R39861 vdd.n2350 vdd.n2349 16.2531
R39862 vdd.n2349 vdd.n2306 16.2531
R39863 vdd.n2338 vdd.n2306 16.2531
R39864 vdd.n1271 vdd.n1226 16.2531
R39865 vdd.n1260 vdd.n1226 16.2531
R39866 vdd.n1260 vdd.n1259 16.2531
R39867 vdd.n1244 vdd.n1237 16.2531
R39868 vdd.n1245 vdd.n1244 16.2531
R39869 vdd.n2372 vdd.n2371 16.2531
R39870 vdd.n2371 vdd.n2356 16.2531
R39871 vdd.n2401 vdd.n2356 16.2531
R39872 vdd.n2401 vdd.n2400 16.2531
R39873 vdd.n2400 vdd.n2357 16.2531
R39874 vdd.n2389 vdd.n2357 16.2531
R39875 vdd.n2419 vdd.n2418 16.2531
R39876 vdd.n2418 vdd.n2403 16.2531
R39877 vdd.n2448 vdd.n2403 16.2531
R39878 vdd.n2448 vdd.n2447 16.2531
R39879 vdd.n2447 vdd.n2404 16.2531
R39880 vdd.n2436 vdd.n2404 16.2531
R39881 vdd.n2469 vdd.n2468 16.2531
R39882 vdd.n2468 vdd.n2453 16.2531
R39883 vdd.n2498 vdd.n2453 16.2531
R39884 vdd.n2498 vdd.n2497 16.2531
R39885 vdd.n2497 vdd.n2454 16.2531
R39886 vdd.n2486 vdd.n2454 16.2531
R39887 vdd.n2519 vdd.n2518 16.2531
R39888 vdd.n2518 vdd.n2503 16.2531
R39889 vdd.n2548 vdd.n2503 16.2531
R39890 vdd.n2548 vdd.n2547 16.2531
R39891 vdd.n2547 vdd.n2504 16.2531
R39892 vdd.n2536 vdd.n2504 16.2531
R39893 vdd.n2567 vdd.n2566 16.2531
R39894 vdd.n2566 vdd.n2551 16.2531
R39895 vdd.n2596 vdd.n2551 16.2531
R39896 vdd.n2596 vdd.n2595 16.2531
R39897 vdd.n2595 vdd.n2552 16.2531
R39898 vdd.n2584 vdd.n2552 16.2531
R39899 vdd.n2718 vdd.n2717 16.2531
R39900 vdd.n2717 vdd.n2697 16.2531
R39901 vdd.n2742 vdd.n2697 16.2531
R39902 vdd.n2742 vdd.n2741 16.2531
R39903 vdd.n2741 vdd.n2698 16.2531
R39904 vdd.n2730 vdd.n2698 16.2531
R39905 vdd.n2670 vdd.n2669 16.2531
R39906 vdd.n2669 vdd.n2649 16.2531
R39907 vdd.n2694 vdd.n2649 16.2531
R39908 vdd.n2694 vdd.n2693 16.2531
R39909 vdd.n2693 vdd.n2650 16.2531
R39910 vdd.n2682 vdd.n2650 16.2531
R39911 vdd.n2767 vdd.n2766 16.2531
R39912 vdd.n2766 vdd.n2746 16.2531
R39913 vdd.n2791 vdd.n2746 16.2531
R39914 vdd.n2791 vdd.n2790 16.2531
R39915 vdd.n2790 vdd.n2747 16.2531
R39916 vdd.n2779 vdd.n2747 16.2531
R39917 vdd.n2817 vdd.n2816 16.2531
R39918 vdd.n2816 vdd.n2796 16.2531
R39919 vdd.n2841 vdd.n2796 16.2531
R39920 vdd.n2841 vdd.n2840 16.2531
R39921 vdd.n2840 vdd.n2797 16.2531
R39922 vdd.n2829 vdd.n2797 16.2531
R39923 vdd.n2865 vdd.n2864 16.2531
R39924 vdd.n2864 vdd.n2844 16.2531
R39925 vdd.n2889 vdd.n2844 16.2531
R39926 vdd.n2889 vdd.n2888 16.2531
R39927 vdd.n2888 vdd.n2845 16.2531
R39928 vdd.n2877 vdd.n2845 16.2531
R39929 vdd.n1052 vdd.n1051 16.2531
R39930 vdd.n1053 vdd.n1052 16.2531
R39931 vdd.n1063 vdd.n1062 16.2531
R39932 vdd.n1064 vdd.n1063 16.2531
R39933 vdd.n1064 vdd.n1027 16.2531
R39934 vdd.n3013 vdd.n3012 16.2531
R39935 vdd.n3012 vdd.n2992 16.2531
R39936 vdd.n3037 vdd.n2992 16.2531
R39937 vdd.n3037 vdd.n3036 16.2531
R39938 vdd.n3036 vdd.n2993 16.2531
R39939 vdd.n3025 vdd.n2993 16.2531
R39940 vdd.n2964 vdd.n2963 16.2531
R39941 vdd.n2963 vdd.n2943 16.2531
R39942 vdd.n2988 vdd.n2943 16.2531
R39943 vdd.n2988 vdd.n2987 16.2531
R39944 vdd.n2987 vdd.n2944 16.2531
R39945 vdd.n2976 vdd.n2944 16.2531
R39946 vdd.n2916 vdd.n2915 16.2531
R39947 vdd.n2915 vdd.n2895 16.2531
R39948 vdd.n2940 vdd.n2895 16.2531
R39949 vdd.n2940 vdd.n2939 16.2531
R39950 vdd.n2939 vdd.n2896 16.2531
R39951 vdd.n2928 vdd.n2896 16.2531
R39952 vdd.n3062 vdd.n3061 16.2531
R39953 vdd.n3061 vdd.n3041 16.2531
R39954 vdd.n3086 vdd.n3041 16.2531
R39955 vdd.n3086 vdd.n3085 16.2531
R39956 vdd.n3085 vdd.n3042 16.2531
R39957 vdd.n3074 vdd.n3042 16.2531
R39958 vdd.n3112 vdd.n3111 16.2531
R39959 vdd.n3111 vdd.n3091 16.2531
R39960 vdd.n3136 vdd.n3091 16.2531
R39961 vdd.n3136 vdd.n3135 16.2531
R39962 vdd.n3135 vdd.n3092 16.2531
R39963 vdd.n3124 vdd.n3092 16.2531
R39964 vdd.n3160 vdd.n3159 16.2531
R39965 vdd.n3159 vdd.n3139 16.2531
R39966 vdd.n3184 vdd.n3139 16.2531
R39967 vdd.n3184 vdd.n3183 16.2531
R39968 vdd.n3183 vdd.n3140 16.2531
R39969 vdd.n3172 vdd.n3140 16.2531
R39970 vdd.n3258 vdd.n3257 16.2531
R39971 vdd.n3257 vdd.n3237 16.2531
R39972 vdd.n3282 vdd.n3237 16.2531
R39973 vdd.n3282 vdd.n3281 16.2531
R39974 vdd.n3281 vdd.n3238 16.2531
R39975 vdd.n3270 vdd.n3238 16.2531
R39976 vdd.n3210 vdd.n3209 16.2531
R39977 vdd.n3209 vdd.n3189 16.2531
R39978 vdd.n3234 vdd.n3189 16.2531
R39979 vdd.n3234 vdd.n3233 16.2531
R39980 vdd.n3233 vdd.n3190 16.2531
R39981 vdd.n3222 vdd.n3190 16.2531
R39982 vdd.n3307 vdd.n3306 16.2531
R39983 vdd.n3306 vdd.n3286 16.2531
R39984 vdd.n3331 vdd.n3286 16.2531
R39985 vdd.n3331 vdd.n3330 16.2531
R39986 vdd.n3330 vdd.n3287 16.2531
R39987 vdd.n3319 vdd.n3287 16.2531
R39988 vdd.n3357 vdd.n3356 16.2531
R39989 vdd.n3356 vdd.n3336 16.2531
R39990 vdd.n3381 vdd.n3336 16.2531
R39991 vdd.n3381 vdd.n3380 16.2531
R39992 vdd.n3380 vdd.n3337 16.2531
R39993 vdd.n3369 vdd.n3337 16.2531
R39994 vdd.n3405 vdd.n3404 16.2531
R39995 vdd.n3404 vdd.n3384 16.2531
R39996 vdd.n3429 vdd.n3384 16.2531
R39997 vdd.n3429 vdd.n3428 16.2531
R39998 vdd.n3428 vdd.n3385 16.2531
R39999 vdd.n3417 vdd.n3385 16.2531
R40000 vdd.n806 vdd.n805 16.2531
R40001 vdd.n807 vdd.n806 16.2531
R40002 vdd.n817 vdd.n816 16.2531
R40003 vdd.n818 vdd.n817 16.2531
R40004 vdd.n818 vdd.n781 16.2531
R40005 vdd.n3504 vdd.n3503 16.2531
R40006 vdd.n3503 vdd.n3483 16.2531
R40007 vdd.n3528 vdd.n3483 16.2531
R40008 vdd.n3528 vdd.n3527 16.2531
R40009 vdd.n3527 vdd.n3484 16.2531
R40010 vdd.n3516 vdd.n3484 16.2531
R40011 vdd.n3456 vdd.n3455 16.2531
R40012 vdd.n3455 vdd.n3435 16.2531
R40013 vdd.n3480 vdd.n3435 16.2531
R40014 vdd.n3480 vdd.n3479 16.2531
R40015 vdd.n3479 vdd.n3436 16.2531
R40016 vdd.n3468 vdd.n3436 16.2531
R40017 vdd.n3553 vdd.n3552 16.2531
R40018 vdd.n3552 vdd.n3532 16.2531
R40019 vdd.n3577 vdd.n3532 16.2531
R40020 vdd.n3577 vdd.n3576 16.2531
R40021 vdd.n3576 vdd.n3533 16.2531
R40022 vdd.n3565 vdd.n3533 16.2531
R40023 vdd.n3603 vdd.n3602 16.2531
R40024 vdd.n3602 vdd.n3582 16.2531
R40025 vdd.n3627 vdd.n3582 16.2531
R40026 vdd.n3627 vdd.n3626 16.2531
R40027 vdd.n3626 vdd.n3583 16.2531
R40028 vdd.n3615 vdd.n3583 16.2531
R40029 vdd.n3651 vdd.n3650 16.2531
R40030 vdd.n3650 vdd.n3630 16.2531
R40031 vdd.n3675 vdd.n3630 16.2531
R40032 vdd.n3675 vdd.n3674 16.2531
R40033 vdd.n3674 vdd.n3631 16.2531
R40034 vdd.n3663 vdd.n3631 16.2531
R40035 vdd.n609 vdd.n608 16.2531
R40036 vdd.n608 vdd.n588 16.2531
R40037 vdd.n633 vdd.n588 16.2531
R40038 vdd.n633 vdd.n632 16.2531
R40039 vdd.n632 vdd.n589 16.2531
R40040 vdd.n621 vdd.n589 16.2531
R40041 vdd.n3750 vdd.n3749 16.2531
R40042 vdd.n3749 vdd.n3729 16.2531
R40043 vdd.n3774 vdd.n3729 16.2531
R40044 vdd.n3774 vdd.n3773 16.2531
R40045 vdd.n3773 vdd.n3730 16.2531
R40046 vdd.n3762 vdd.n3730 16.2531
R40047 vdd.n3702 vdd.n3701 16.2531
R40048 vdd.n3701 vdd.n3681 16.2531
R40049 vdd.n3726 vdd.n3681 16.2531
R40050 vdd.n3726 vdd.n3725 16.2531
R40051 vdd.n3725 vdd.n3682 16.2531
R40052 vdd.n3714 vdd.n3682 16.2531
R40053 vdd.n6892 vdd.n6891 16.2531
R40054 vdd.n6891 vdd.n6871 16.2531
R40055 vdd.n6916 vdd.n6871 16.2531
R40056 vdd.n6916 vdd.n6915 16.2531
R40057 vdd.n6915 vdd.n6872 16.2531
R40058 vdd.n6904 vdd.n6872 16.2531
R40059 vdd.n6844 vdd.n6843 16.2531
R40060 vdd.n6843 vdd.n6823 16.2531
R40061 vdd.n6868 vdd.n6823 16.2531
R40062 vdd.n6868 vdd.n6867 16.2531
R40063 vdd.n6867 vdd.n6824 16.2531
R40064 vdd.n6856 vdd.n6824 16.2531
R40065 vdd.n10034 vdd.n10033 16.2531
R40066 vdd.n10033 vdd.n10013 16.2531
R40067 vdd.n10058 vdd.n10013 16.2531
R40068 vdd.n10058 vdd.n10057 16.2531
R40069 vdd.n10057 vdd.n10014 16.2531
R40070 vdd.n10046 vdd.n10014 16.2531
R40071 vdd.n9986 vdd.n9985 16.2531
R40072 vdd.n9985 vdd.n9965 16.2531
R40073 vdd.n10010 vdd.n9965 16.2531
R40074 vdd.n10010 vdd.n10009 16.2531
R40075 vdd.n10009 vdd.n9966 16.2531
R40076 vdd.n9998 vdd.n9966 16.2531
R40077 vdd.n10082 vdd.n10081 16.2531
R40078 vdd.n10081 vdd.n10061 16.2531
R40079 vdd.n10106 vdd.n10061 16.2531
R40080 vdd.n10106 vdd.n10105 16.2531
R40081 vdd.n10105 vdd.n10062 16.2531
R40082 vdd.n10094 vdd.n10062 16.2531
R40083 vdd.n10130 vdd.n10129 16.2531
R40084 vdd.n10129 vdd.n10109 16.2531
R40085 vdd.n10154 vdd.n10109 16.2531
R40086 vdd.n10154 vdd.n10153 16.2531
R40087 vdd.n10153 vdd.n10110 16.2531
R40088 vdd.n10142 vdd.n10110 16.2531
R40089 vdd.n10232 vdd.n10231 16.2531
R40090 vdd.n10231 vdd.n10211 16.2531
R40091 vdd.n10256 vdd.n10211 16.2531
R40092 vdd.n10256 vdd.n10255 16.2531
R40093 vdd.n10255 vdd.n10212 16.2531
R40094 vdd.n10244 vdd.n10212 16.2531
R40095 vdd.n10280 vdd.n10279 16.2531
R40096 vdd.n10279 vdd.n10259 16.2531
R40097 vdd.n10304 vdd.n10259 16.2531
R40098 vdd.n10304 vdd.n10303 16.2531
R40099 vdd.n10303 vdd.n10260 16.2531
R40100 vdd.n10292 vdd.n10260 16.2531
R40101 vdd.n10328 vdd.n10327 16.2531
R40102 vdd.n10327 vdd.n10307 16.2531
R40103 vdd.n10352 vdd.n10307 16.2531
R40104 vdd.n10352 vdd.n10351 16.2531
R40105 vdd.n10351 vdd.n10308 16.2531
R40106 vdd.n10340 vdd.n10308 16.2531
R40107 vdd.n10376 vdd.n10375 16.2531
R40108 vdd.n10375 vdd.n10355 16.2531
R40109 vdd.n10400 vdd.n10355 16.2531
R40110 vdd.n10400 vdd.n10399 16.2531
R40111 vdd.n10399 vdd.n10356 16.2531
R40112 vdd.n10388 vdd.n10356 16.2531
R40113 vdd.n10478 vdd.n10477 16.2531
R40114 vdd.n10477 vdd.n10457 16.2531
R40115 vdd.n10502 vdd.n10457 16.2531
R40116 vdd.n10502 vdd.n10501 16.2531
R40117 vdd.n10501 vdd.n10458 16.2531
R40118 vdd.n10490 vdd.n10458 16.2531
R40119 vdd.n70 vdd.n69 16.2531
R40120 vdd.n69 vdd.n49 16.2531
R40121 vdd.n94 vdd.n49 16.2531
R40122 vdd.n94 vdd.n93 16.2531
R40123 vdd.n93 vdd.n50 16.2531
R40124 vdd.n82 vdd.n50 16.2531
R40125 vdd.n22 vdd.n21 16.2531
R40126 vdd.n21 vdd.n1 16.2531
R40127 vdd.n46 vdd.n1 16.2531
R40128 vdd.n46 vdd.n45 16.2531
R40129 vdd.n45 vdd.n2 16.2531
R40130 vdd.n34 vdd.n2 16.2531
R40131 vdd.n10526 vdd.n10525 16.2531
R40132 vdd.n10525 vdd.n10505 16.2531
R40133 vdd.n10550 vdd.n10505 16.2531
R40134 vdd.n10550 vdd.n10549 16.2531
R40135 vdd.n10549 vdd.n10506 16.2531
R40136 vdd.n10538 vdd.n10506 16.2531
R40137 vdd.n10576 vdd.n10575 16.2531
R40138 vdd.n10575 vdd.n10555 16.2531
R40139 vdd.n10600 vdd.n10555 16.2531
R40140 vdd.n10600 vdd.n10599 16.2531
R40141 vdd.n10599 vdd.n10556 16.2531
R40142 vdd.n10588 vdd.n10556 16.2531
R40143 vdd.n10624 vdd.n10623 16.2531
R40144 vdd.n10623 vdd.n10603 16.2531
R40145 vdd.n10648 vdd.n10603 16.2531
R40146 vdd.n10648 vdd.n10647 16.2531
R40147 vdd.n10647 vdd.n10604 16.2531
R40148 vdd.n10636 vdd.n10604 16.2531
R40149 vdd.n10429 vdd.n10428 16.2531
R40150 vdd.n10430 vdd.n10429 16.2531
R40151 vdd.n10440 vdd.n10439 16.2531
R40152 vdd.n10441 vdd.n10440 16.2531
R40153 vdd.n10441 vdd.n10404 16.2531
R40154 vdd.n10772 vdd.n10771 16.2531
R40155 vdd.n10771 vdd.n10751 16.2531
R40156 vdd.n10796 vdd.n10751 16.2531
R40157 vdd.n10796 vdd.n10795 16.2531
R40158 vdd.n10795 vdd.n10752 16.2531
R40159 vdd.n10784 vdd.n10752 16.2531
R40160 vdd.n10723 vdd.n10722 16.2531
R40161 vdd.n10722 vdd.n10702 16.2531
R40162 vdd.n10747 vdd.n10702 16.2531
R40163 vdd.n10747 vdd.n10746 16.2531
R40164 vdd.n10746 vdd.n10703 16.2531
R40165 vdd.n10735 vdd.n10703 16.2531
R40166 vdd.n10675 vdd.n10674 16.2531
R40167 vdd.n10674 vdd.n10654 16.2531
R40168 vdd.n10699 vdd.n10654 16.2531
R40169 vdd.n10699 vdd.n10698 16.2531
R40170 vdd.n10698 vdd.n10655 16.2531
R40171 vdd.n10687 vdd.n10655 16.2531
R40172 vdd.n10821 vdd.n10820 16.2531
R40173 vdd.n10820 vdd.n10800 16.2531
R40174 vdd.n10845 vdd.n10800 16.2531
R40175 vdd.n10845 vdd.n10844 16.2531
R40176 vdd.n10844 vdd.n10801 16.2531
R40177 vdd.n10833 vdd.n10801 16.2531
R40178 vdd.n10871 vdd.n10870 16.2531
R40179 vdd.n10870 vdd.n10850 16.2531
R40180 vdd.n10895 vdd.n10850 16.2531
R40181 vdd.n10895 vdd.n10894 16.2531
R40182 vdd.n10894 vdd.n10851 16.2531
R40183 vdd.n10883 vdd.n10851 16.2531
R40184 vdd.n10919 vdd.n10918 16.2531
R40185 vdd.n10918 vdd.n10898 16.2531
R40186 vdd.n10943 vdd.n10898 16.2531
R40187 vdd.n10943 vdd.n10942 16.2531
R40188 vdd.n10942 vdd.n10899 16.2531
R40189 vdd.n10931 vdd.n10899 16.2531
R40190 vdd.n11017 vdd.n11016 16.2531
R40191 vdd.n11016 vdd.n10996 16.2531
R40192 vdd.n11041 vdd.n10996 16.2531
R40193 vdd.n11041 vdd.n11040 16.2531
R40194 vdd.n11040 vdd.n10997 16.2531
R40195 vdd.n11029 vdd.n10997 16.2531
R40196 vdd.n10969 vdd.n10968 16.2531
R40197 vdd.n10968 vdd.n10948 16.2531
R40198 vdd.n10993 vdd.n10948 16.2531
R40199 vdd.n10993 vdd.n10992 16.2531
R40200 vdd.n10992 vdd.n10949 16.2531
R40201 vdd.n10981 vdd.n10949 16.2531
R40202 vdd.n11066 vdd.n11065 16.2531
R40203 vdd.n11065 vdd.n11045 16.2531
R40204 vdd.n11090 vdd.n11045 16.2531
R40205 vdd.n11090 vdd.n11089 16.2531
R40206 vdd.n11089 vdd.n11046 16.2531
R40207 vdd.n11078 vdd.n11046 16.2531
R40208 vdd.n11116 vdd.n11115 16.2531
R40209 vdd.n11115 vdd.n11095 16.2531
R40210 vdd.n11140 vdd.n11095 16.2531
R40211 vdd.n11140 vdd.n11139 16.2531
R40212 vdd.n11139 vdd.n11096 16.2531
R40213 vdd.n11128 vdd.n11096 16.2531
R40214 vdd.n11164 vdd.n11163 16.2531
R40215 vdd.n11163 vdd.n11143 16.2531
R40216 vdd.n11188 vdd.n11143 16.2531
R40217 vdd.n11188 vdd.n11187 16.2531
R40218 vdd.n11187 vdd.n11144 16.2531
R40219 vdd.n11176 vdd.n11144 16.2531
R40220 vdd.n10183 vdd.n10182 16.2531
R40221 vdd.n10184 vdd.n10183 16.2531
R40222 vdd.n10194 vdd.n10193 16.2531
R40223 vdd.n10195 vdd.n10194 16.2531
R40224 vdd.n10195 vdd.n10158 16.2531
R40225 vdd.n11263 vdd.n11262 16.2531
R40226 vdd.n11262 vdd.n11242 16.2531
R40227 vdd.n11287 vdd.n11242 16.2531
R40228 vdd.n11287 vdd.n11286 16.2531
R40229 vdd.n11286 vdd.n11243 16.2531
R40230 vdd.n11275 vdd.n11243 16.2531
R40231 vdd.n11215 vdd.n11214 16.2531
R40232 vdd.n11214 vdd.n11194 16.2531
R40233 vdd.n11239 vdd.n11194 16.2531
R40234 vdd.n11239 vdd.n11238 16.2531
R40235 vdd.n11238 vdd.n11195 16.2531
R40236 vdd.n11227 vdd.n11195 16.2531
R40237 vdd.n11312 vdd.n11311 16.2531
R40238 vdd.n11311 vdd.n11291 16.2531
R40239 vdd.n11336 vdd.n11291 16.2531
R40240 vdd.n11336 vdd.n11335 16.2531
R40241 vdd.n11335 vdd.n11292 16.2531
R40242 vdd.n11324 vdd.n11292 16.2531
R40243 vdd.n11362 vdd.n11361 16.2531
R40244 vdd.n11361 vdd.n11341 16.2531
R40245 vdd.n11386 vdd.n11341 16.2531
R40246 vdd.n11386 vdd.n11385 16.2531
R40247 vdd.n11385 vdd.n11342 16.2531
R40248 vdd.n11374 vdd.n11342 16.2531
R40249 vdd.n11410 vdd.n11409 16.2531
R40250 vdd.n11409 vdd.n11389 16.2531
R40251 vdd.n11434 vdd.n11389 16.2531
R40252 vdd.n11434 vdd.n11433 16.2531
R40253 vdd.n11433 vdd.n11390 16.2531
R40254 vdd.n11422 vdd.n11390 16.2531
R40255 vdd.n11456 vdd.n11455 16.2531
R40256 vdd.n11455 vdd.n11440 16.2531
R40257 vdd.n11485 vdd.n11440 16.2531
R40258 vdd.n11485 vdd.n11484 16.2531
R40259 vdd.n11484 vdd.n11441 16.2531
R40260 vdd.n11473 vdd.n11441 16.2531
R40261 vdd.n11503 vdd.n11502 16.2531
R40262 vdd.n11502 vdd.n11487 16.2531
R40263 vdd.n11532 vdd.n11487 16.2531
R40264 vdd.n11532 vdd.n11531 16.2531
R40265 vdd.n11531 vdd.n11488 16.2531
R40266 vdd.n11520 vdd.n11488 16.2531
R40267 vdd.n11553 vdd.n11552 16.2531
R40268 vdd.n11552 vdd.n11537 16.2531
R40269 vdd.n11582 vdd.n11537 16.2531
R40270 vdd.n11582 vdd.n11581 16.2531
R40271 vdd.n11581 vdd.n11538 16.2531
R40272 vdd.n11570 vdd.n11538 16.2531
R40273 vdd.n11603 vdd.n11602 16.2531
R40274 vdd.n11602 vdd.n11587 16.2531
R40275 vdd.n11632 vdd.n11587 16.2531
R40276 vdd.n11632 vdd.n11631 16.2531
R40277 vdd.n11631 vdd.n11588 16.2531
R40278 vdd.n11620 vdd.n11588 16.2531
R40279 vdd.n11651 vdd.n11650 16.2531
R40280 vdd.n11650 vdd.n11635 16.2531
R40281 vdd.n11680 vdd.n11635 16.2531
R40282 vdd.n11680 vdd.n11679 16.2531
R40283 vdd.n11679 vdd.n11636 16.2531
R40284 vdd.n11668 vdd.n11636 16.2531
R40285 vdd.n486 vdd.n441 16.2531
R40286 vdd.n475 vdd.n441 16.2531
R40287 vdd.n475 vdd.n474 16.2531
R40288 vdd.n459 vdd.n452 16.2531
R40289 vdd.n460 vdd.n459 16.2531
R40290 vdd.n11702 vdd.n11701 16.2531
R40291 vdd.n11701 vdd.n11686 16.2531
R40292 vdd.n11731 vdd.n11686 16.2531
R40293 vdd.n11731 vdd.n11730 16.2531
R40294 vdd.n11730 vdd.n11687 16.2531
R40295 vdd.n11719 vdd.n11687 16.2531
R40296 vdd.n11749 vdd.n11748 16.2531
R40297 vdd.n11748 vdd.n11733 16.2531
R40298 vdd.n11778 vdd.n11733 16.2531
R40299 vdd.n11778 vdd.n11777 16.2531
R40300 vdd.n11777 vdd.n11734 16.2531
R40301 vdd.n11766 vdd.n11734 16.2531
R40302 vdd.n11797 vdd.n11796 16.2531
R40303 vdd.n11796 vdd.n11781 16.2531
R40304 vdd.n11826 vdd.n11781 16.2531
R40305 vdd.n11826 vdd.n11825 16.2531
R40306 vdd.n11825 vdd.n11782 16.2531
R40307 vdd.n11814 vdd.n11782 16.2531
R40308 vdd.n11848 vdd.n11847 16.2531
R40309 vdd.n11847 vdd.n11832 16.2531
R40310 vdd.n11877 vdd.n11832 16.2531
R40311 vdd.n11877 vdd.n11876 16.2531
R40312 vdd.n11876 vdd.n11833 16.2531
R40313 vdd.n11865 vdd.n11833 16.2531
R40314 vdd.n11898 vdd.n11897 16.2531
R40315 vdd.n11897 vdd.n11882 16.2531
R40316 vdd.n11927 vdd.n11882 16.2531
R40317 vdd.n11927 vdd.n11926 16.2531
R40318 vdd.n11926 vdd.n11883 16.2531
R40319 vdd.n11915 vdd.n11883 16.2531
R40320 vdd.n11946 vdd.n11945 16.2531
R40321 vdd.n11945 vdd.n11930 16.2531
R40322 vdd.n11975 vdd.n11930 16.2531
R40323 vdd.n11975 vdd.n11974 16.2531
R40324 vdd.n11974 vdd.n11931 16.2531
R40325 vdd.n11963 vdd.n11931 16.2531
R40326 vdd.n11996 vdd.n11995 16.2531
R40327 vdd.n11995 vdd.n11980 16.2531
R40328 vdd.n12025 vdd.n11980 16.2531
R40329 vdd.n12025 vdd.n12024 16.2531
R40330 vdd.n12024 vdd.n11981 16.2531
R40331 vdd.n12013 vdd.n11981 16.2531
R40332 vdd.n12043 vdd.n12042 16.2531
R40333 vdd.n12042 vdd.n12027 16.2531
R40334 vdd.n12072 vdd.n12027 16.2531
R40335 vdd.n12072 vdd.n12071 16.2531
R40336 vdd.n12071 vdd.n12028 16.2531
R40337 vdd.n12060 vdd.n12028 16.2531
R40338 vdd.n12093 vdd.n12092 16.2531
R40339 vdd.n12092 vdd.n12077 16.2531
R40340 vdd.n12122 vdd.n12077 16.2531
R40341 vdd.n12122 vdd.n12121 16.2531
R40342 vdd.n12121 vdd.n12078 16.2531
R40343 vdd.n12110 vdd.n12078 16.2531
R40344 vdd.n12143 vdd.n12142 16.2531
R40345 vdd.n12142 vdd.n12127 16.2531
R40346 vdd.n12172 vdd.n12127 16.2531
R40347 vdd.n12172 vdd.n12171 16.2531
R40348 vdd.n12171 vdd.n12128 16.2531
R40349 vdd.n12160 vdd.n12128 16.2531
R40350 vdd.n12191 vdd.n12190 16.2531
R40351 vdd.n12190 vdd.n12175 16.2531
R40352 vdd.n12220 vdd.n12175 16.2531
R40353 vdd.n12220 vdd.n12219 16.2531
R40354 vdd.n12219 vdd.n12176 16.2531
R40355 vdd.n12208 vdd.n12176 16.2531
R40356 vdd.n241 vdd.n196 16.2531
R40357 vdd.n230 vdd.n196 16.2531
R40358 vdd.n230 vdd.n229 16.2531
R40359 vdd.n214 vdd.n207 16.2531
R40360 vdd.n215 vdd.n214 16.2531
R40361 vdd.n12242 vdd.n12241 16.2531
R40362 vdd.n12241 vdd.n12226 16.2531
R40363 vdd.n12271 vdd.n12226 16.2531
R40364 vdd.n12271 vdd.n12270 16.2531
R40365 vdd.n12270 vdd.n12227 16.2531
R40366 vdd.n12259 vdd.n12227 16.2531
R40367 vdd.n12289 vdd.n12288 16.2531
R40368 vdd.n12288 vdd.n12273 16.2531
R40369 vdd.n12318 vdd.n12273 16.2531
R40370 vdd.n12318 vdd.n12317 16.2531
R40371 vdd.n12317 vdd.n12274 16.2531
R40372 vdd.n12306 vdd.n12274 16.2531
R40373 vdd.n12339 vdd.n12338 16.2531
R40374 vdd.n12338 vdd.n12323 16.2531
R40375 vdd.n12368 vdd.n12323 16.2531
R40376 vdd.n12368 vdd.n12367 16.2531
R40377 vdd.n12367 vdd.n12324 16.2531
R40378 vdd.n12356 vdd.n12324 16.2531
R40379 vdd.n12389 vdd.n12388 16.2531
R40380 vdd.n12388 vdd.n12373 16.2531
R40381 vdd.n12418 vdd.n12373 16.2531
R40382 vdd.n12418 vdd.n12417 16.2531
R40383 vdd.n12417 vdd.n12374 16.2531
R40384 vdd.n12406 vdd.n12374 16.2531
R40385 vdd.n12437 vdd.n12436 16.2531
R40386 vdd.n12436 vdd.n12421 16.2531
R40387 vdd.n12466 vdd.n12421 16.2531
R40388 vdd.n12466 vdd.n12465 16.2531
R40389 vdd.n12465 vdd.n12422 16.2531
R40390 vdd.n12454 vdd.n12422 16.2531
R40391 vdd.n7766 vdd.n7753 13.9199
R40392 vdd.n7521 vdd.n7508 13.9199
R40393 vdd.n4624 vdd.n4611 13.9199
R40394 vdd.n4379 vdd.n4366 13.9199
R40395 vdd.n1482 vdd.n1469 13.9199
R40396 vdd.n1237 vdd.n1224 13.9199
R40397 vdd.n452 vdd.n439 13.9199
R40398 vdd.n207 vdd.n194 13.9199
R40399 vdd.n7337 vdd.n7310 13.9189
R40400 vdd.n7091 vdd.n7064 13.9189
R40401 vdd.n4195 vdd.n4168 13.9189
R40402 vdd.n3949 vdd.n3922 13.9189
R40403 vdd.n1053 vdd.n1026 13.9189
R40404 vdd.n807 vdd.n780 13.9189
R40405 vdd.n10430 vdd.n10403 13.9189
R40406 vdd.n10184 vdd.n10157 13.9189
R40407 vdd.n7801 vdd.n7800 12.4637
R40408 vdd.n7556 vdd.n7555 12.4637
R40409 vdd.n7358 vdd.n7311 12.4637
R40410 vdd.n7112 vdd.n7065 12.4637
R40411 vdd.n4659 vdd.n4658 12.4637
R40412 vdd.n4414 vdd.n4413 12.4637
R40413 vdd.n4216 vdd.n4169 12.4637
R40414 vdd.n3970 vdd.n3923 12.4637
R40415 vdd.n1517 vdd.n1516 12.4637
R40416 vdd.n1272 vdd.n1271 12.4637
R40417 vdd.n1074 vdd.n1027 12.4637
R40418 vdd.n828 vdd.n781 12.4637
R40419 vdd.n10451 vdd.n10404 12.4637
R40420 vdd.n10205 vdd.n10158 12.4637
R40421 vdd.n487 vdd.n486 12.4637
R40422 vdd.n242 vdd.n241 12.4637
R40423 vdd vdd.n7752 9.01037
R40424 vdd vdd.n7507 9.01037
R40425 vdd vdd.n4610 9.01037
R40426 vdd vdd.n4365 9.01037
R40427 vdd vdd.n1468 9.01037
R40428 vdd vdd.n1223 9.01037
R40429 vdd vdd.n438 9.01037
R40430 vdd vdd.n193 9.01037
R40431 vdd.n7360 vdd.n7309 9.0005
R40432 vdd.n7114 vdd.n7063 9.0005
R40433 vdd.n4218 vdd.n4167 9.0005
R40434 vdd.n3972 vdd.n3921 9.0005
R40435 vdd.n1076 vdd.n1025 9.0005
R40436 vdd.n830 vdd.n779 9.0005
R40437 vdd.n10453 vdd.n10402 9.0005
R40438 vdd.n10207 vdd.n10156 9.0005
R40439 vdd.n8931 vdd.n8882 6.24557
R40440 vdd.n5789 vdd.n5740 6.24557
R40441 vdd.n2647 vdd.n2598 6.24557
R40442 vdd.n12469 vdd.n12468 6.24557
R40443 vdd.n3775 vdd 5.95856
R40444 vdd.n10059 vdd 5.95856
R40445 vdd.n6917 vdd 5.76119
R40446 vdd.n9962 vdd.n6966 4.70938
R40447 vdd.n6820 vdd.n3824 4.70938
R40448 vdd.n3678 vdd.n682 4.70938
R40449 vdd.n11438 vdd.n11437 4.70938
R40450 vdd.n6869 vdd.n6821 4.23159
R40451 vdd.n8242 vdd.n8241 4.08685
R40452 vdd.n9274 vdd.n9225 4.08685
R40453 vdd.n5100 vdd.n5099 4.08685
R40454 vdd.n6132 vdd.n6083 4.08685
R40455 vdd.n1958 vdd.n1957 4.08685
R40456 vdd.n2990 vdd.n2941 4.08685
R40457 vdd.n10749 vdd.n10700 4.08685
R40458 vdd.n11828 vdd.n11827 4.08685
R40459 vdd.n3727 vdd.n3679 4.03422
R40460 vdd.n10011 vdd.n9963 4.03422
R40461 vdd.n7948 vdd.n7947 2.95445
R40462 vdd.n8488 vdd.n8487 2.95445
R40463 vdd.n8734 vdd.n8733 2.95445
R40464 vdd.n9027 vdd.n8979 2.95445
R40465 vdd.n9567 vdd.n9519 2.95445
R40466 vdd.n9813 vdd.n9765 2.95445
R40467 vdd.n4806 vdd.n4805 2.95445
R40468 vdd.n5346 vdd.n5345 2.95445
R40469 vdd.n5592 vdd.n5591 2.95445
R40470 vdd.n5885 vdd.n5837 2.95445
R40471 vdd.n6425 vdd.n6377 2.95445
R40472 vdd.n6671 vdd.n6623 2.95445
R40473 vdd.n1664 vdd.n1663 2.95445
R40474 vdd.n2204 vdd.n2203 2.95445
R40475 vdd.n2450 vdd.n2449 2.95445
R40476 vdd.n2743 vdd.n2695 2.95445
R40477 vdd.n3283 vdd.n3235 2.95445
R40478 vdd.n3529 vdd.n3481 2.95445
R40479 vdd.n95 vdd.n47 2.95445
R40480 vdd.n11042 vdd.n10994 2.95445
R40481 vdd.n11288 vdd.n11240 2.95445
R40482 vdd.n11534 vdd.n11533 2.95445
R40483 vdd.n12074 vdd.n12073 2.95445
R40484 vdd.n12320 vdd.n12319 2.95445
R40485 vdd.n8243 vdd.n8242 2.33849
R40486 vdd.n9322 vdd.n9274 2.33849
R40487 vdd.n5101 vdd.n5100 2.33849
R40488 vdd.n6180 vdd.n6132 2.33849
R40489 vdd.n1959 vdd.n1958 2.33849
R40490 vdd.n3038 vdd.n2990 2.33849
R40491 vdd.n10797 vdd.n10749 2.33849
R40492 vdd.n11829 vdd.n11828 2.33849
R40493 vdd.n11437 vdd 2.27025
R40494 vdd.n9963 vdd.n9962 1.54656
R40495 vdd.n6821 vdd.n6820 1.54656
R40496 vdd.n3679 vdd.n3678 1.54656
R40497 vdd.n9962 vdd.n9961 1.53669
R40498 vdd.n6820 vdd.n6819 1.53669
R40499 vdd.n3678 vdd.n3677 1.53669
R40500 vdd.n11437 vdd.n11436 1.53669
R40501 vdd.n7999 vdd.n7998 1.50544
R40502 vdd.n8294 vdd.n8293 1.50544
R40503 vdd.n8392 vdd.n8391 1.50544
R40504 vdd.n8539 vdd.n8538 1.50544
R40505 vdd.n8785 vdd.n8784 1.50544
R40506 vdd.n9078 vdd.n9077 1.50544
R40507 vdd.n9373 vdd.n9372 1.50544
R40508 vdd.n9471 vdd.n9470 1.50544
R40509 vdd.n9618 vdd.n9617 1.50544
R40510 vdd.n9864 vdd.n9863 1.50544
R40511 vdd.n4857 vdd.n4856 1.50544
R40512 vdd.n5152 vdd.n5151 1.50544
R40513 vdd.n5250 vdd.n5249 1.50544
R40514 vdd.n5397 vdd.n5396 1.50544
R40515 vdd.n5643 vdd.n5642 1.50544
R40516 vdd.n5936 vdd.n5935 1.50544
R40517 vdd.n6231 vdd.n6230 1.50544
R40518 vdd.n6329 vdd.n6328 1.50544
R40519 vdd.n6476 vdd.n6475 1.50544
R40520 vdd.n6722 vdd.n6721 1.50544
R40521 vdd.n1715 vdd.n1714 1.50544
R40522 vdd.n2010 vdd.n2009 1.50544
R40523 vdd.n2108 vdd.n2107 1.50544
R40524 vdd.n2255 vdd.n2254 1.50544
R40525 vdd.n2501 vdd.n2500 1.50544
R40526 vdd.n2794 vdd.n2793 1.50544
R40527 vdd.n3089 vdd.n3088 1.50544
R40528 vdd.n3187 vdd.n3186 1.50544
R40529 vdd.n3334 vdd.n3333 1.50544
R40530 vdd.n3580 vdd.n3579 1.50544
R40531 vdd.n10553 vdd.n10552 1.50544
R40532 vdd.n10848 vdd.n10847 1.50544
R40533 vdd.n10946 vdd.n10945 1.50544
R40534 vdd.n11093 vdd.n11092 1.50544
R40535 vdd.n11339 vdd.n11338 1.50544
R40536 vdd.n11585 vdd.n11584 1.50544
R40537 vdd.n11880 vdd.n11879 1.50544
R40538 vdd.n11978 vdd.n11977 1.50544
R40539 vdd.n12125 vdd.n12124 1.50544
R40540 vdd.n12371 vdd.n12370 1.50544
R40541 vdd.n7998 vdd.n7997 0.904283
R40542 vdd.n7999 vdd.n7852 0.904283
R40543 vdd.n8096 vdd.n8095 0.904283
R40544 vdd.n8293 vdd.n8292 0.904283
R40545 vdd.n8294 vdd.n7703 0.904283
R40546 vdd.n8391 vdd.n8390 0.904283
R40547 vdd.n8538 vdd.n8537 0.904283
R40548 vdd.n8539 vdd.n7607 0.904283
R40549 vdd.n8636 vdd.n8635 0.904283
R40550 vdd.n8784 vdd.n8783 0.904283
R40551 vdd.n8785 vdd.n7458 0.904283
R40552 vdd.n8882 vdd.n8881 0.904283
R40553 vdd.n9077 vdd.n9076 0.904283
R40554 vdd.n9078 vdd.n7410 0.904283
R40555 vdd.n9175 vdd.n9174 0.904283
R40556 vdd.n9372 vdd.n9371 0.904283
R40557 vdd.n9373 vdd.n7260 0.904283
R40558 vdd.n9470 vdd.n9469 0.904283
R40559 vdd.n9617 vdd.n9616 0.904283
R40560 vdd.n9618 vdd.n7164 0.904283
R40561 vdd.n9715 vdd.n9714 0.904283
R40562 vdd.n9863 vdd.n9862 0.904283
R40563 vdd.n9864 vdd.n7014 0.904283
R40564 vdd.n9961 vdd.n9960 0.904283
R40565 vdd.n4856 vdd.n4855 0.904283
R40566 vdd.n4857 vdd.n4710 0.904283
R40567 vdd.n4954 vdd.n4953 0.904283
R40568 vdd.n5151 vdd.n5150 0.904283
R40569 vdd.n5152 vdd.n4561 0.904283
R40570 vdd.n5249 vdd.n5248 0.904283
R40571 vdd.n5396 vdd.n5395 0.904283
R40572 vdd.n5397 vdd.n4465 0.904283
R40573 vdd.n5494 vdd.n5493 0.904283
R40574 vdd.n5642 vdd.n5641 0.904283
R40575 vdd.n5643 vdd.n4316 0.904283
R40576 vdd.n5740 vdd.n5739 0.904283
R40577 vdd.n5935 vdd.n5934 0.904283
R40578 vdd.n5936 vdd.n4268 0.904283
R40579 vdd.n6033 vdd.n6032 0.904283
R40580 vdd.n6230 vdd.n6229 0.904283
R40581 vdd.n6231 vdd.n4118 0.904283
R40582 vdd.n6328 vdd.n6327 0.904283
R40583 vdd.n6475 vdd.n6474 0.904283
R40584 vdd.n6476 vdd.n4022 0.904283
R40585 vdd.n6573 vdd.n6572 0.904283
R40586 vdd.n6721 vdd.n6720 0.904283
R40587 vdd.n6722 vdd.n3872 0.904283
R40588 vdd.n6819 vdd.n6818 0.904283
R40589 vdd.n1714 vdd.n1713 0.904283
R40590 vdd.n1715 vdd.n1568 0.904283
R40591 vdd.n1812 vdd.n1811 0.904283
R40592 vdd.n2009 vdd.n2008 0.904283
R40593 vdd.n2010 vdd.n1419 0.904283
R40594 vdd.n2107 vdd.n2106 0.904283
R40595 vdd.n2254 vdd.n2253 0.904283
R40596 vdd.n2255 vdd.n1323 0.904283
R40597 vdd.n2352 vdd.n2351 0.904283
R40598 vdd.n2500 vdd.n2499 0.904283
R40599 vdd.n2501 vdd.n1174 0.904283
R40600 vdd.n2598 vdd.n2597 0.904283
R40601 vdd.n2793 vdd.n2792 0.904283
R40602 vdd.n2794 vdd.n1126 0.904283
R40603 vdd.n2891 vdd.n2890 0.904283
R40604 vdd.n3088 vdd.n3087 0.904283
R40605 vdd.n3089 vdd.n976 0.904283
R40606 vdd.n3186 vdd.n3185 0.904283
R40607 vdd.n3333 vdd.n3332 0.904283
R40608 vdd.n3334 vdd.n880 0.904283
R40609 vdd.n3431 vdd.n3430 0.904283
R40610 vdd.n3579 vdd.n3578 0.904283
R40611 vdd.n3580 vdd.n730 0.904283
R40612 vdd.n3677 vdd.n3676 0.904283
R40613 vdd.n10552 vdd.n10551 0.904283
R40614 vdd.n10553 vdd.n10503 0.904283
R40615 vdd.n10650 vdd.n10649 0.904283
R40616 vdd.n10847 vdd.n10846 0.904283
R40617 vdd.n10848 vdd.n10353 0.904283
R40618 vdd.n10945 vdd.n10944 0.904283
R40619 vdd.n11092 vdd.n11091 0.904283
R40620 vdd.n11093 vdd.n10257 0.904283
R40621 vdd.n11190 vdd.n11189 0.904283
R40622 vdd.n11338 vdd.n11337 0.904283
R40623 vdd.n11339 vdd.n10107 0.904283
R40624 vdd.n11436 vdd.n11435 0.904283
R40625 vdd.n11584 vdd.n11583 0.904283
R40626 vdd.n11585 vdd.n538 0.904283
R40627 vdd.n11682 vdd.n11681 0.904283
R40628 vdd.n11879 vdd.n11878 0.904283
R40629 vdd.n11880 vdd.n389 0.904283
R40630 vdd.n11977 vdd.n11976 0.904283
R40631 vdd.n12124 vdd.n12123 0.904283
R40632 vdd.n12125 vdd.n293 0.904283
R40633 vdd.n12222 vdd.n12221 0.904283
R40634 vdd.n12370 vdd.n12369 0.904283
R40635 vdd.n12371 vdd.n144 0.904283
R40636 vdd.n12468 vdd.n12467 0.904283
R40637 vdd.n8097 vdd.n8096 0.854122
R40638 vdd.n8637 vdd.n8636 0.854122
R40639 vdd.n9176 vdd.n9175 0.854122
R40640 vdd.n9716 vdd.n9715 0.854122
R40641 vdd.n4955 vdd.n4954 0.854122
R40642 vdd.n5495 vdd.n5494 0.854122
R40643 vdd.n6034 vdd.n6033 0.854122
R40644 vdd.n6574 vdd.n6573 0.854122
R40645 vdd.n1813 vdd.n1812 0.854122
R40646 vdd.n2353 vdd.n2352 0.854122
R40647 vdd.n2892 vdd.n2891 0.854122
R40648 vdd.n3432 vdd.n3431 0.854122
R40649 vdd.n10651 vdd.n10650 0.854122
R40650 vdd.n11191 vdd.n11190 0.854122
R40651 vdd.n11683 vdd.n11682 0.854122
R40652 vdd.n12223 vdd.n12222 0.854122
R40653 vdd vdd.n7751 0.76448
R40654 vdd vdd.n7506 0.76448
R40655 vdd vdd.n4609 0.76448
R40656 vdd vdd.n4364 0.76448
R40657 vdd vdd.n1467 0.76448
R40658 vdd vdd.n1222 0.76448
R40659 vdd vdd.n437 0.76448
R40660 vdd vdd.n192 0.76448
R40661 vdd vdd.n6965 0.752967
R40662 vdd vdd.n7655 0.752967
R40663 vdd vdd.n3823 0.752967
R40664 vdd vdd.n4513 0.752967
R40665 vdd vdd.n681 0.752967
R40666 vdd vdd.n1371 0.752967
R40667 vdd vdd.n586 0.752967
R40668 vdd vdd.n341 0.752967
R40669 vdd.n3679 vdd 0.724184
R40670 vdd.n6821 vdd 0.724184
R40671 vdd.n9963 vdd 0.724184
R40672 vdd vdd.n12517 0.711849
R40673 vdd vdd.n8930 0.698691
R40674 vdd vdd.n7308 0.698691
R40675 vdd vdd.n7212 0.698691
R40676 vdd vdd.n7062 0.698691
R40677 vdd vdd.n5788 0.698691
R40678 vdd vdd.n4166 0.698691
R40679 vdd vdd.n4070 0.698691
R40680 vdd vdd.n3920 0.698691
R40681 vdd vdd.n2646 0.698691
R40682 vdd vdd.n1024 0.698691
R40683 vdd vdd.n928 0.698691
R40684 vdd vdd.n778 0.698691
R40685 vdd vdd.n10401 0.698691
R40686 vdd vdd.n10305 0.698691
R40687 vdd vdd.n10155 0.698691
R40688 vdd.n7998 vdd.n7949 0.697868
R40689 vdd.n8096 vdd.n8047 0.697868
R40690 vdd.n8293 vdd.n8244 0.697868
R40691 vdd.n8391 vdd.n8342 0.697868
R40692 vdd.n8538 vdd.n8489 0.697868
R40693 vdd.n8636 vdd.n8587 0.697868
R40694 vdd.n8784 vdd.n8735 0.697868
R40695 vdd.n8882 vdd.n8833 0.697868
R40696 vdd.n9077 vdd.n9028 0.697868
R40697 vdd.n9175 vdd.n9126 0.697868
R40698 vdd.n9372 vdd.n9323 0.697868
R40699 vdd.n9470 vdd.n9421 0.697868
R40700 vdd.n9617 vdd.n9568 0.697868
R40701 vdd.n9715 vdd.n9666 0.697868
R40702 vdd.n9863 vdd.n9814 0.697868
R40703 vdd.n9961 vdd.n9912 0.697868
R40704 vdd.n4856 vdd.n4807 0.697868
R40705 vdd.n4954 vdd.n4905 0.697868
R40706 vdd.n5151 vdd.n5102 0.697868
R40707 vdd.n5249 vdd.n5200 0.697868
R40708 vdd.n5396 vdd.n5347 0.697868
R40709 vdd.n5494 vdd.n5445 0.697868
R40710 vdd.n5642 vdd.n5593 0.697868
R40711 vdd.n5740 vdd.n5691 0.697868
R40712 vdd.n5935 vdd.n5886 0.697868
R40713 vdd.n6033 vdd.n5984 0.697868
R40714 vdd.n6230 vdd.n6181 0.697868
R40715 vdd.n6328 vdd.n6279 0.697868
R40716 vdd.n6475 vdd.n6426 0.697868
R40717 vdd.n6573 vdd.n6524 0.697868
R40718 vdd.n6721 vdd.n6672 0.697868
R40719 vdd.n6819 vdd.n6770 0.697868
R40720 vdd.n1714 vdd.n1665 0.697868
R40721 vdd.n1812 vdd.n1763 0.697868
R40722 vdd.n2009 vdd.n1960 0.697868
R40723 vdd.n2107 vdd.n2058 0.697868
R40724 vdd.n2254 vdd.n2205 0.697868
R40725 vdd.n2352 vdd.n2303 0.697868
R40726 vdd.n2500 vdd.n2451 0.697868
R40727 vdd.n2598 vdd.n2549 0.697868
R40728 vdd.n2793 vdd.n2744 0.697868
R40729 vdd.n2891 vdd.n2842 0.697868
R40730 vdd.n3088 vdd.n3039 0.697868
R40731 vdd.n3186 vdd.n3137 0.697868
R40732 vdd.n3333 vdd.n3284 0.697868
R40733 vdd.n3431 vdd.n3382 0.697868
R40734 vdd.n3579 vdd.n3530 0.697868
R40735 vdd.n3677 vdd.n3628 0.697868
R40736 vdd.n10552 vdd.n96 0.697868
R40737 vdd.n10650 vdd.n10601 0.697868
R40738 vdd.n10847 vdd.n10798 0.697868
R40739 vdd.n10945 vdd.n10896 0.697868
R40740 vdd.n11092 vdd.n11043 0.697868
R40741 vdd.n11190 vdd.n11141 0.697868
R40742 vdd.n11338 vdd.n11289 0.697868
R40743 vdd.n11436 vdd.n11387 0.697868
R40744 vdd.n11584 vdd.n11535 0.697868
R40745 vdd.n11682 vdd.n11633 0.697868
R40746 vdd.n11879 vdd.n11830 0.697868
R40747 vdd.n11977 vdd.n11928 0.697868
R40748 vdd.n12124 vdd.n12075 0.697868
R40749 vdd.n12222 vdd.n12173 0.697868
R40750 vdd.n12370 vdd.n12321 0.697868
R40751 vdd.n12468 vdd.n12419 0.697868
R40752 vdd vdd.n9125 0.662508
R40753 vdd vdd.n9420 0.662508
R40754 vdd vdd.n9665 0.662508
R40755 vdd vdd.n9911 0.662508
R40756 vdd vdd.n5983 0.662508
R40757 vdd vdd.n6278 0.662508
R40758 vdd vdd.n6523 0.662508
R40759 vdd vdd.n6769 0.662508
R40760 vdd vdd.n2841 0.662508
R40761 vdd vdd.n3136 0.662508
R40762 vdd vdd.n3381 0.662508
R40763 vdd vdd.n3627 0.662508
R40764 vdd vdd.n633 0.662508
R40765 vdd vdd.n10600 0.662508
R40766 vdd vdd.n10895 0.662508
R40767 vdd vdd.n11140 0.662508
R40768 vdd vdd.n11386 0.662508
R40769 vdd.n8930 vdd 0.662507
R40770 vdd.n8979 vdd 0.662507
R40771 vdd vdd.n9027 0.662507
R40772 vdd.n9076 vdd 0.662507
R40773 vdd.n7410 vdd 0.662507
R40774 vdd.n9174 vdd 0.662507
R40775 vdd.n7308 vdd 0.662507
R40776 vdd.n9225 vdd 0.662507
R40777 vdd.n9273 vdd 0.662507
R40778 vdd vdd.n9322 0.662507
R40779 vdd.n9371 vdd 0.662507
R40780 vdd.n7260 vdd 0.662507
R40781 vdd.n9469 vdd 0.662507
R40782 vdd.n7212 vdd 0.662507
R40783 vdd.n9519 vdd 0.662507
R40784 vdd vdd.n9567 0.662507
R40785 vdd.n9616 vdd 0.662507
R40786 vdd.n7164 vdd 0.662507
R40787 vdd.n9714 vdd 0.662507
R40788 vdd.n7062 vdd 0.662507
R40789 vdd.n9765 vdd 0.662507
R40790 vdd vdd.n9813 0.662507
R40791 vdd.n9862 vdd 0.662507
R40792 vdd.n7014 vdd 0.662507
R40793 vdd.n9960 vdd 0.662507
R40794 vdd.n5788 vdd 0.662507
R40795 vdd.n5837 vdd 0.662507
R40796 vdd vdd.n5885 0.662507
R40797 vdd.n5934 vdd 0.662507
R40798 vdd.n4268 vdd 0.662507
R40799 vdd.n6032 vdd 0.662507
R40800 vdd.n4166 vdd 0.662507
R40801 vdd.n6083 vdd 0.662507
R40802 vdd.n6131 vdd 0.662507
R40803 vdd vdd.n6180 0.662507
R40804 vdd.n6229 vdd 0.662507
R40805 vdd.n4118 vdd 0.662507
R40806 vdd.n6327 vdd 0.662507
R40807 vdd.n4070 vdd 0.662507
R40808 vdd.n6377 vdd 0.662507
R40809 vdd vdd.n6425 0.662507
R40810 vdd.n6474 vdd 0.662507
R40811 vdd.n4022 vdd 0.662507
R40812 vdd.n6572 vdd 0.662507
R40813 vdd.n3920 vdd 0.662507
R40814 vdd.n6623 vdd 0.662507
R40815 vdd vdd.n6671 0.662507
R40816 vdd.n6720 vdd 0.662507
R40817 vdd.n3872 vdd 0.662507
R40818 vdd.n6818 vdd 0.662507
R40819 vdd.n2646 vdd 0.662507
R40820 vdd.n2695 vdd 0.662507
R40821 vdd vdd.n2743 0.662507
R40822 vdd.n2792 vdd 0.662507
R40823 vdd.n1126 vdd 0.662507
R40824 vdd.n2890 vdd 0.662507
R40825 vdd.n1024 vdd 0.662507
R40826 vdd.n2941 vdd 0.662507
R40827 vdd.n2989 vdd 0.662507
R40828 vdd vdd.n3038 0.662507
R40829 vdd.n3087 vdd 0.662507
R40830 vdd.n976 vdd 0.662507
R40831 vdd.n3185 vdd 0.662507
R40832 vdd.n928 vdd 0.662507
R40833 vdd.n3235 vdd 0.662507
R40834 vdd vdd.n3283 0.662507
R40835 vdd.n3332 vdd 0.662507
R40836 vdd.n880 vdd 0.662507
R40837 vdd.n3430 vdd 0.662507
R40838 vdd.n778 vdd 0.662507
R40839 vdd.n3481 vdd 0.662507
R40840 vdd vdd.n3529 0.662507
R40841 vdd.n3578 vdd 0.662507
R40842 vdd.n730 vdd 0.662507
R40843 vdd.n3676 vdd 0.662507
R40844 vdd vdd.n3727 0.662507
R40845 vdd vdd.n3775 0.662507
R40846 vdd vdd.n6869 0.662507
R40847 vdd vdd.n6917 0.662507
R40848 vdd vdd.n10011 0.662507
R40849 vdd vdd.n10059 0.662507
R40850 vdd.n47 vdd 0.662507
R40851 vdd vdd.n95 0.662507
R40852 vdd.n10551 vdd 0.662507
R40853 vdd.n10503 vdd 0.662507
R40854 vdd.n10649 vdd 0.662507
R40855 vdd.n10401 vdd 0.662507
R40856 vdd.n10700 vdd 0.662507
R40857 vdd.n10748 vdd 0.662507
R40858 vdd vdd.n10797 0.662507
R40859 vdd.n10846 vdd 0.662507
R40860 vdd.n10353 vdd 0.662507
R40861 vdd.n10944 vdd 0.662507
R40862 vdd.n10305 vdd 0.662507
R40863 vdd.n10994 vdd 0.662507
R40864 vdd vdd.n11042 0.662507
R40865 vdd.n11091 vdd 0.662507
R40866 vdd.n10257 vdd 0.662507
R40867 vdd.n11189 vdd 0.662507
R40868 vdd.n10155 vdd 0.662507
R40869 vdd.n11240 vdd 0.662507
R40870 vdd vdd.n11288 0.662507
R40871 vdd.n11337 vdd 0.662507
R40872 vdd.n10107 vdd 0.662507
R40873 vdd.n11435 vdd 0.662507
R40874 vdd.n12517 vdd 0.662507
R40875 vdd vdd.n8046 0.629613
R40876 vdd vdd.n8341 0.629613
R40877 vdd vdd.n8586 0.629613
R40878 vdd vdd.n8832 0.629613
R40879 vdd vdd.n4904 0.629613
R40880 vdd vdd.n5199 0.629613
R40881 vdd vdd.n5444 0.629613
R40882 vdd vdd.n5690 0.629613
R40883 vdd vdd.n1762 0.629613
R40884 vdd vdd.n2057 0.629613
R40885 vdd vdd.n2302 0.629613
R40886 vdd vdd.n2548 0.629613
R40887 vdd vdd.n11632 0.629613
R40888 vdd vdd.n11927 0.629613
R40889 vdd vdd.n12172 0.629613
R40890 vdd vdd.n12418 0.629613
R40891 vdd.n7947 vdd 0.629612
R40892 vdd vdd.n7948 0.629612
R40893 vdd.n7997 vdd 0.629612
R40894 vdd.n7852 vdd 0.629612
R40895 vdd.n8095 vdd 0.629612
R40896 vdd.n7751 vdd 0.629612
R40897 vdd.n8241 vdd 0.629612
R40898 vdd.n8193 vdd 0.629612
R40899 vdd vdd.n8243 0.629612
R40900 vdd.n8292 vdd 0.629612
R40901 vdd.n7703 vdd 0.629612
R40902 vdd.n8390 vdd 0.629612
R40903 vdd.n7655 vdd 0.629612
R40904 vdd.n8487 vdd 0.629612
R40905 vdd vdd.n8488 0.629612
R40906 vdd.n8537 vdd 0.629612
R40907 vdd.n7607 vdd 0.629612
R40908 vdd.n8635 vdd 0.629612
R40909 vdd.n7506 vdd 0.629612
R40910 vdd.n8733 vdd 0.629612
R40911 vdd vdd.n8734 0.629612
R40912 vdd.n8783 vdd 0.629612
R40913 vdd.n7458 vdd 0.629612
R40914 vdd.n8881 vdd 0.629612
R40915 vdd.n4805 vdd 0.629612
R40916 vdd vdd.n4806 0.629612
R40917 vdd.n4855 vdd 0.629612
R40918 vdd.n4710 vdd 0.629612
R40919 vdd.n4953 vdd 0.629612
R40920 vdd.n4609 vdd 0.629612
R40921 vdd.n5099 vdd 0.629612
R40922 vdd.n5051 vdd 0.629612
R40923 vdd vdd.n5101 0.629612
R40924 vdd.n5150 vdd 0.629612
R40925 vdd.n4561 vdd 0.629612
R40926 vdd.n5248 vdd 0.629612
R40927 vdd.n4513 vdd 0.629612
R40928 vdd.n5345 vdd 0.629612
R40929 vdd vdd.n5346 0.629612
R40930 vdd.n5395 vdd 0.629612
R40931 vdd.n4465 vdd 0.629612
R40932 vdd.n5493 vdd 0.629612
R40933 vdd.n4364 vdd 0.629612
R40934 vdd.n5591 vdd 0.629612
R40935 vdd vdd.n5592 0.629612
R40936 vdd.n5641 vdd 0.629612
R40937 vdd.n4316 vdd 0.629612
R40938 vdd.n5739 vdd 0.629612
R40939 vdd.n1663 vdd 0.629612
R40940 vdd vdd.n1664 0.629612
R40941 vdd.n1713 vdd 0.629612
R40942 vdd.n1568 vdd 0.629612
R40943 vdd.n1811 vdd 0.629612
R40944 vdd.n1467 vdd 0.629612
R40945 vdd.n1957 vdd 0.629612
R40946 vdd.n1909 vdd 0.629612
R40947 vdd vdd.n1959 0.629612
R40948 vdd.n2008 vdd 0.629612
R40949 vdd.n1419 vdd 0.629612
R40950 vdd.n2106 vdd 0.629612
R40951 vdd.n1371 vdd 0.629612
R40952 vdd.n2203 vdd 0.629612
R40953 vdd vdd.n2204 0.629612
R40954 vdd.n2253 vdd 0.629612
R40955 vdd.n1323 vdd 0.629612
R40956 vdd.n2351 vdd 0.629612
R40957 vdd.n1222 vdd 0.629612
R40958 vdd.n2449 vdd 0.629612
R40959 vdd vdd.n2450 0.629612
R40960 vdd.n2499 vdd 0.629612
R40961 vdd.n1174 vdd 0.629612
R40962 vdd.n2597 vdd 0.629612
R40963 vdd.n11533 vdd 0.629612
R40964 vdd vdd.n11534 0.629612
R40965 vdd.n11583 vdd 0.629612
R40966 vdd.n538 vdd 0.629612
R40967 vdd.n11681 vdd 0.629612
R40968 vdd.n437 vdd 0.629612
R40969 vdd.n11827 vdd 0.629612
R40970 vdd.n11779 vdd 0.629612
R40971 vdd vdd.n11829 0.629612
R40972 vdd.n11878 vdd 0.629612
R40973 vdd.n389 vdd 0.629612
R40974 vdd.n11976 vdd 0.629612
R40975 vdd.n341 vdd 0.629612
R40976 vdd.n12073 vdd 0.629612
R40977 vdd vdd.n12074 0.629612
R40978 vdd.n12123 vdd 0.629612
R40979 vdd.n293 vdd 0.629612
R40980 vdd.n12221 vdd 0.629612
R40981 vdd.n192 vdd 0.629612
R40982 vdd.n12319 vdd 0.629612
R40983 vdd vdd.n12320 0.629612
R40984 vdd.n12369 vdd 0.629612
R40985 vdd.n144 vdd 0.629612
R40986 vdd.n12467 vdd 0.629612
R40987 vdd.n8097 vdd.n7804 0.628061
R40988 vdd.n8637 vdd.n7559 0.628061
R40989 vdd.n9176 vdd.n7362 0.628061
R40990 vdd.n9716 vdd.n7116 0.628061
R40991 vdd.n4955 vdd.n4662 0.628061
R40992 vdd.n5495 vdd.n4417 0.628061
R40993 vdd.n6034 vdd.n4220 0.628061
R40994 vdd.n6574 vdd.n3974 0.628061
R40995 vdd.n1813 vdd.n1520 0.628061
R40996 vdd.n2353 vdd.n1275 0.628061
R40997 vdd.n2892 vdd.n1078 0.628061
R40998 vdd.n3432 vdd.n832 0.628061
R40999 vdd.n10651 vdd.n10455 0.628061
R41000 vdd.n11191 vdd.n10209 0.628061
R41001 vdd.n11683 vdd.n490 0.628061
R41002 vdd.n12223 vdd.n245 0.628061
R41003 vdd.n7949 vdd.n6966 0.620566
R41004 vdd.n8047 vdd.n7999 0.620566
R41005 vdd.n8244 vdd.n8098 0.620566
R41006 vdd.n8342 vdd.n8294 0.620566
R41007 vdd.n8489 vdd.n8392 0.620566
R41008 vdd.n8587 vdd.n8539 0.620566
R41009 vdd.n8735 vdd.n8638 0.620566
R41010 vdd.n8833 vdd.n8785 0.620566
R41011 vdd.n9028 vdd.n8931 0.620566
R41012 vdd.n9126 vdd.n9078 0.620566
R41013 vdd.n9323 vdd.n9177 0.620566
R41014 vdd.n9421 vdd.n9373 0.620566
R41015 vdd.n9568 vdd.n9471 0.620566
R41016 vdd.n9666 vdd.n9618 0.620566
R41017 vdd.n9814 vdd.n9717 0.620566
R41018 vdd.n9912 vdd.n9864 0.620566
R41019 vdd.n4807 vdd.n3824 0.620566
R41020 vdd.n4905 vdd.n4857 0.620566
R41021 vdd.n5102 vdd.n4956 0.620566
R41022 vdd.n5200 vdd.n5152 0.620566
R41023 vdd.n5347 vdd.n5250 0.620566
R41024 vdd.n5445 vdd.n5397 0.620566
R41025 vdd.n5593 vdd.n5496 0.620566
R41026 vdd.n5691 vdd.n5643 0.620566
R41027 vdd.n5886 vdd.n5789 0.620566
R41028 vdd.n5984 vdd.n5936 0.620566
R41029 vdd.n6181 vdd.n6035 0.620566
R41030 vdd.n6279 vdd.n6231 0.620566
R41031 vdd.n6426 vdd.n6329 0.620566
R41032 vdd.n6524 vdd.n6476 0.620566
R41033 vdd.n6672 vdd.n6575 0.620566
R41034 vdd.n6770 vdd.n6722 0.620566
R41035 vdd.n1665 vdd.n682 0.620566
R41036 vdd.n1763 vdd.n1715 0.620566
R41037 vdd.n1960 vdd.n1814 0.620566
R41038 vdd.n2058 vdd.n2010 0.620566
R41039 vdd.n2205 vdd.n2108 0.620566
R41040 vdd.n2303 vdd.n2255 0.620566
R41041 vdd.n2451 vdd.n2354 0.620566
R41042 vdd.n2549 vdd.n2501 0.620566
R41043 vdd.n2744 vdd.n2647 0.620566
R41044 vdd.n2842 vdd.n2794 0.620566
R41045 vdd.n3039 vdd.n2893 0.620566
R41046 vdd.n3137 vdd.n3089 0.620566
R41047 vdd.n3284 vdd.n3187 0.620566
R41048 vdd.n3382 vdd.n3334 0.620566
R41049 vdd.n3530 vdd.n3433 0.620566
R41050 vdd.n3628 vdd.n3580 0.620566
R41051 vdd.n12469 vdd.n96 0.620566
R41052 vdd.n10601 vdd.n10553 0.620566
R41053 vdd.n10798 vdd.n10652 0.620566
R41054 vdd.n10896 vdd.n10848 0.620566
R41055 vdd.n11043 vdd.n10946 0.620566
R41056 vdd.n11141 vdd.n11093 0.620566
R41057 vdd.n11289 vdd.n11192 0.620566
R41058 vdd.n11387 vdd.n11339 0.620566
R41059 vdd.n11535 vdd.n11438 0.620566
R41060 vdd.n11633 vdd.n11585 0.620566
R41061 vdd.n11830 vdd.n11684 0.620566
R41062 vdd.n11928 vdd.n11880 0.620566
R41063 vdd.n12075 vdd.n11978 0.620566
R41064 vdd.n12173 vdd.n12125 0.620566
R41065 vdd.n12321 vdd.n12224 0.620566
R41066 vdd.n12419 vdd.n12371 0.620566
R41067 vdd.n8242 vdd.n8193 0.616454
R41068 vdd.n9274 vdd.n9273 0.616454
R41069 vdd.n5100 vdd.n5051 0.616454
R41070 vdd.n6132 vdd.n6131 0.616454
R41071 vdd.n1958 vdd.n1909 0.616454
R41072 vdd.n2990 vdd.n2989 0.616454
R41073 vdd.n10749 vdd.n10748 0.616454
R41074 vdd.n11828 vdd.n11779 0.616454
R41075 vdd.n6965 vdd 0.613164
R41076 vdd.n3823 vdd 0.613164
R41077 vdd.n681 vdd 0.613164
R41078 vdd.n586 vdd 0.613164
R41079 vdd.n7802 vdd.n7753 0.598862
R41080 vdd.n7557 vdd.n7508 0.598862
R41081 vdd.n7359 vdd.n7310 0.598862
R41082 vdd.n7113 vdd.n7064 0.598862
R41083 vdd.n4660 vdd.n4611 0.598862
R41084 vdd.n4415 vdd.n4366 0.598862
R41085 vdd.n4217 vdd.n4168 0.598862
R41086 vdd.n3971 vdd.n3922 0.598862
R41087 vdd.n1518 vdd.n1469 0.598862
R41088 vdd.n1273 vdd.n1224 0.598862
R41089 vdd.n1075 vdd.n1026 0.598862
R41090 vdd.n829 vdd.n780 0.598862
R41091 vdd.n10452 vdd.n10403 0.598862
R41092 vdd.n10206 vdd.n10157 0.598862
R41093 vdd.n488 vdd.n439 0.598862
R41094 vdd.n243 vdd.n194 0.598862
R41095 vdd.n8098 vdd.n8097 0.594253
R41096 vdd.n8638 vdd.n8637 0.594253
R41097 vdd.n9177 vdd.n9176 0.594253
R41098 vdd.n9717 vdd.n9716 0.594253
R41099 vdd.n4956 vdd.n4955 0.594253
R41100 vdd.n5496 vdd.n5495 0.594253
R41101 vdd.n6035 vdd.n6034 0.594253
R41102 vdd.n6575 vdd.n6574 0.594253
R41103 vdd.n1814 vdd.n1813 0.594253
R41104 vdd.n2354 vdd.n2353 0.594253
R41105 vdd.n2893 vdd.n2892 0.594253
R41106 vdd.n3433 vdd.n3432 0.594253
R41107 vdd.n10652 vdd.n10651 0.594253
R41108 vdd.n11192 vdd.n11191 0.594253
R41109 vdd.n11684 vdd.n11683 0.594253
R41110 vdd.n12224 vdd.n12223 0.594253
R41111 vdd.n7949 vdd 0.276816
R41112 vdd.n8047 vdd 0.276816
R41113 vdd.n8244 vdd 0.276816
R41114 vdd.n8342 vdd 0.276816
R41115 vdd.n8489 vdd 0.276816
R41116 vdd.n8587 vdd 0.276816
R41117 vdd.n8735 vdd 0.276816
R41118 vdd.n8833 vdd 0.276816
R41119 vdd.n4807 vdd 0.276816
R41120 vdd.n4905 vdd 0.276816
R41121 vdd.n5102 vdd 0.276816
R41122 vdd.n5200 vdd 0.276816
R41123 vdd.n5347 vdd 0.276816
R41124 vdd.n5445 vdd 0.276816
R41125 vdd.n5593 vdd 0.276816
R41126 vdd.n5691 vdd 0.276816
R41127 vdd.n1665 vdd 0.276816
R41128 vdd.n1763 vdd 0.276816
R41129 vdd.n1960 vdd 0.276816
R41130 vdd.n2058 vdd 0.276816
R41131 vdd.n2205 vdd 0.276816
R41132 vdd.n2303 vdd 0.276816
R41133 vdd.n2451 vdd 0.276816
R41134 vdd.n2549 vdd 0.276816
R41135 vdd.n11535 vdd 0.276816
R41136 vdd.n11633 vdd 0.276816
R41137 vdd.n11830 vdd 0.276816
R41138 vdd.n11928 vdd 0.276816
R41139 vdd.n12075 vdd 0.276816
R41140 vdd.n12173 vdd 0.276816
R41141 vdd.n12321 vdd 0.276816
R41142 vdd.n12419 vdd 0.276816
R41143 vdd.n9028 vdd 0.243921
R41144 vdd.n9126 vdd 0.243921
R41145 vdd.n9323 vdd 0.243921
R41146 vdd.n9421 vdd 0.243921
R41147 vdd.n9568 vdd 0.243921
R41148 vdd.n9666 vdd 0.243921
R41149 vdd.n9814 vdd 0.243921
R41150 vdd.n9912 vdd 0.243921
R41151 vdd.n5886 vdd 0.243921
R41152 vdd.n5984 vdd 0.243921
R41153 vdd.n6181 vdd 0.243921
R41154 vdd.n6279 vdd 0.243921
R41155 vdd.n6426 vdd 0.243921
R41156 vdd.n6524 vdd 0.243921
R41157 vdd.n6672 vdd 0.243921
R41158 vdd.n6770 vdd 0.243921
R41159 vdd.n2744 vdd 0.243921
R41160 vdd.n2842 vdd 0.243921
R41161 vdd.n3039 vdd 0.243921
R41162 vdd.n3137 vdd 0.243921
R41163 vdd.n3284 vdd 0.243921
R41164 vdd.n3382 vdd 0.243921
R41165 vdd.n3530 vdd 0.243921
R41166 vdd.n3628 vdd 0.243921
R41167 vdd.n96 vdd 0.243921
R41168 vdd.n10601 vdd 0.243921
R41169 vdd.n10798 vdd 0.243921
R41170 vdd.n10896 vdd 0.243921
R41171 vdd.n11043 vdd 0.243921
R41172 vdd.n11141 vdd 0.243921
R41173 vdd.n11289 vdd 0.243921
R41174 vdd.n11387 vdd 0.243921
R41175 vdd.n9177 vdd 0.206092
R41176 vdd.n9717 vdd 0.206092
R41177 vdd.n6035 vdd 0.206092
R41178 vdd.n6575 vdd 0.206092
R41179 vdd.n2893 vdd 0.206092
R41180 vdd.n3433 vdd 0.206092
R41181 vdd.n10652 vdd 0.206092
R41182 vdd.n11192 vdd 0.206092
R41183 vdd.n8931 vdd 0.184711
R41184 vdd.n9471 vdd 0.184711
R41185 vdd.n5789 vdd 0.184711
R41186 vdd.n6329 vdd 0.184711
R41187 vdd.n2647 vdd 0.184711
R41188 vdd.n3187 vdd 0.184711
R41189 vdd.n10946 vdd 0.184711
R41190 vdd vdd.n12469 0.183066
R41191 vdd.n6966 vdd 0.140303
R41192 vdd.n8098 vdd 0.140303
R41193 vdd.n8392 vdd 0.140303
R41194 vdd.n8638 vdd 0.140303
R41195 vdd.n3824 vdd 0.140303
R41196 vdd.n4956 vdd 0.140303
R41197 vdd.n5250 vdd 0.140303
R41198 vdd.n5496 vdd 0.140303
R41199 vdd.n682 vdd 0.140303
R41200 vdd.n1814 vdd 0.140303
R41201 vdd.n2108 vdd 0.140303
R41202 vdd.n2354 vdd 0.140303
R41203 vdd.n11438 vdd 0.140303
R41204 vdd.n11684 vdd 0.140303
R41205 vdd.n11978 vdd 0.140303
R41206 vdd.n12224 vdd 0.140303
R41207 vdd.n7804 vdd.n7752 0.02926
R41208 vdd.n7559 vdd.n7507 0.02926
R41209 vdd.n7362 vdd.n7309 0.02926
R41210 vdd.n7116 vdd.n7063 0.02926
R41211 vdd.n4662 vdd.n4610 0.02926
R41212 vdd.n4417 vdd.n4365 0.02926
R41213 vdd.n4220 vdd.n4167 0.02926
R41214 vdd.n3974 vdd.n3921 0.02926
R41215 vdd.n1520 vdd.n1468 0.02926
R41216 vdd.n1275 vdd.n1223 0.02926
R41217 vdd.n1078 vdd.n1025 0.02926
R41218 vdd.n832 vdd.n779 0.02926
R41219 vdd.n10455 vdd.n10402 0.02926
R41220 vdd.n10209 vdd.n10156 0.02926
R41221 vdd.n490 vdd.n438 0.02926
R41222 vdd.n245 vdd.n193 0.02926
R41223 vdd.n7361 vdd.n7360 0.0235263
R41224 vdd.n7360 vdd 0.0235263
R41225 vdd.n7115 vdd.n7114 0.0235263
R41226 vdd.n7114 vdd 0.0235263
R41227 vdd.n4219 vdd.n4218 0.0235263
R41228 vdd.n4218 vdd 0.0235263
R41229 vdd.n3973 vdd.n3972 0.0235263
R41230 vdd.n3972 vdd 0.0235263
R41231 vdd.n1077 vdd.n1076 0.0235263
R41232 vdd.n1076 vdd 0.0235263
R41233 vdd.n831 vdd.n830 0.0235263
R41234 vdd.n830 vdd 0.0235263
R41235 vdd.n10454 vdd.n10453 0.0235263
R41236 vdd.n10453 vdd 0.0235263
R41237 vdd.n10208 vdd.n10207 0.0235263
R41238 vdd.n10207 vdd 0.0235263
R41239 vdd.n12479 vdd.n12478 0.0225448
R41240 vdd.n12480 vdd.n12479 0.0225448
R41241 vdd.n12492 vdd.n12491 0.0225448
R41242 vdd.n12493 vdd.n12492 0.0225448
R41243 vdd.n12512 vdd.n12511 0.0225448
R41244 vdd.n12513 vdd.n12512 0.0225448
R41245 vdd.n12502 vdd.n12501 0.0225448
R41246 vdd.n12483 vdd.n12482 0.0225448
R41247 vdd.n12495 vdd.n12494 0.0225448
R41248 vdd.n12494 vdd.n12493 0.0225448
R41249 vdd.n12515 vdd.n12514 0.0225448
R41250 vdd.n12514 vdd.n12513 0.0225448
R41251 vdd.n12506 vdd.n12505 0.0225448
R41252 vdd.n12505 vdd.n12504 0.0225448
R41253 vdd.n117 vdd.n116 0.0225448
R41254 vdd.n125 vdd.n124 0.0225448
R41255 vdd.n124 vdd.n123 0.0225448
R41256 vdd.n139 vdd.n138 0.0225448
R41257 vdd.n140 vdd.n139 0.0225448
R41258 vdd.n136 vdd.n135 0.0225448
R41259 vdd.n135 vdd.n134 0.0225448
R41260 vdd.n132 vdd.n131 0.0225448
R41261 vdd.n142 vdd.n141 0.0225448
R41262 vdd.n141 vdd.n140 0.0225448
R41263 vdd.n122 vdd.n98 0.0225448
R41264 vdd.n123 vdd.n122 0.0225448
R41265 vdd.n120 vdd.n114 0.0225448
R41266 vdd.n120 vdd.n119 0.0225448
R41267 vdd.n165 vdd.n164 0.0225448
R41268 vdd.n173 vdd.n172 0.0225448
R41269 vdd.n172 vdd.n171 0.0225448
R41270 vdd.n187 vdd.n186 0.0225448
R41271 vdd.n188 vdd.n187 0.0225448
R41272 vdd.n184 vdd.n183 0.0225448
R41273 vdd.n183 vdd.n182 0.0225448
R41274 vdd.n180 vdd.n179 0.0225448
R41275 vdd.n190 vdd.n189 0.0225448
R41276 vdd.n189 vdd.n188 0.0225448
R41277 vdd.n170 vdd.n146 0.0225448
R41278 vdd.n171 vdd.n170 0.0225448
R41279 vdd.n168 vdd.n162 0.0225448
R41280 vdd.n168 vdd.n167 0.0225448
R41281 vdd.n266 vdd.n265 0.0225448
R41282 vdd.n274 vdd.n273 0.0225448
R41283 vdd.n273 vdd.n272 0.0225448
R41284 vdd.n288 vdd.n287 0.0225448
R41285 vdd.n289 vdd.n288 0.0225448
R41286 vdd.n285 vdd.n284 0.0225448
R41287 vdd.n284 vdd.n283 0.0225448
R41288 vdd.n281 vdd.n280 0.0225448
R41289 vdd.n291 vdd.n290 0.0225448
R41290 vdd.n290 vdd.n289 0.0225448
R41291 vdd.n271 vdd.n247 0.0225448
R41292 vdd.n272 vdd.n271 0.0225448
R41293 vdd.n269 vdd.n263 0.0225448
R41294 vdd.n269 vdd.n268 0.0225448
R41295 vdd.n314 vdd.n313 0.0225448
R41296 vdd.n322 vdd.n321 0.0225448
R41297 vdd.n321 vdd.n320 0.0225448
R41298 vdd.n336 vdd.n335 0.0225448
R41299 vdd.n337 vdd.n336 0.0225448
R41300 vdd.n333 vdd.n332 0.0225448
R41301 vdd.n332 vdd.n331 0.0225448
R41302 vdd.n329 vdd.n328 0.0225448
R41303 vdd.n339 vdd.n338 0.0225448
R41304 vdd.n338 vdd.n337 0.0225448
R41305 vdd.n319 vdd.n295 0.0225448
R41306 vdd.n320 vdd.n319 0.0225448
R41307 vdd.n317 vdd.n311 0.0225448
R41308 vdd.n317 vdd.n316 0.0225448
R41309 vdd.n362 vdd.n361 0.0225448
R41310 vdd.n370 vdd.n369 0.0225448
R41311 vdd.n369 vdd.n368 0.0225448
R41312 vdd.n384 vdd.n383 0.0225448
R41313 vdd.n385 vdd.n384 0.0225448
R41314 vdd.n381 vdd.n380 0.0225448
R41315 vdd.n380 vdd.n379 0.0225448
R41316 vdd.n377 vdd.n376 0.0225448
R41317 vdd.n387 vdd.n386 0.0225448
R41318 vdd.n386 vdd.n385 0.0225448
R41319 vdd.n367 vdd.n343 0.0225448
R41320 vdd.n368 vdd.n367 0.0225448
R41321 vdd.n365 vdd.n359 0.0225448
R41322 vdd.n365 vdd.n364 0.0225448
R41323 vdd.n410 vdd.n409 0.0225448
R41324 vdd.n418 vdd.n417 0.0225448
R41325 vdd.n417 vdd.n416 0.0225448
R41326 vdd.n432 vdd.n431 0.0225448
R41327 vdd.n433 vdd.n432 0.0225448
R41328 vdd.n429 vdd.n428 0.0225448
R41329 vdd.n428 vdd.n427 0.0225448
R41330 vdd.n425 vdd.n424 0.0225448
R41331 vdd.n435 vdd.n434 0.0225448
R41332 vdd.n434 vdd.n433 0.0225448
R41333 vdd.n415 vdd.n391 0.0225448
R41334 vdd.n416 vdd.n415 0.0225448
R41335 vdd.n413 vdd.n407 0.0225448
R41336 vdd.n413 vdd.n412 0.0225448
R41337 vdd.n511 vdd.n510 0.0225448
R41338 vdd.n519 vdd.n518 0.0225448
R41339 vdd.n518 vdd.n517 0.0225448
R41340 vdd.n533 vdd.n532 0.0225448
R41341 vdd.n534 vdd.n533 0.0225448
R41342 vdd.n530 vdd.n529 0.0225448
R41343 vdd.n529 vdd.n528 0.0225448
R41344 vdd.n526 vdd.n525 0.0225448
R41345 vdd.n536 vdd.n535 0.0225448
R41346 vdd.n535 vdd.n534 0.0225448
R41347 vdd.n516 vdd.n492 0.0225448
R41348 vdd.n517 vdd.n516 0.0225448
R41349 vdd.n514 vdd.n508 0.0225448
R41350 vdd.n514 vdd.n513 0.0225448
R41351 vdd.n559 vdd.n558 0.0225448
R41352 vdd.n567 vdd.n566 0.0225448
R41353 vdd.n566 vdd.n565 0.0225448
R41354 vdd.n581 vdd.n580 0.0225448
R41355 vdd.n582 vdd.n581 0.0225448
R41356 vdd.n578 vdd.n577 0.0225448
R41357 vdd.n577 vdd.n576 0.0225448
R41358 vdd.n574 vdd.n573 0.0225448
R41359 vdd.n584 vdd.n583 0.0225448
R41360 vdd.n583 vdd.n582 0.0225448
R41361 vdd.n564 vdd.n540 0.0225448
R41362 vdd.n565 vdd.n564 0.0225448
R41363 vdd.n562 vdd.n556 0.0225448
R41364 vdd.n562 vdd.n561 0.0225448
R41365 vdd.n6984 vdd.n6982 0.0225448
R41366 vdd.n6984 vdd.n6983 0.0225448
R41367 vdd.n6995 vdd.n6994 0.0225448
R41368 vdd.n6994 vdd.n6993 0.0225448
R41369 vdd.n7009 vdd.n7008 0.0225448
R41370 vdd.n7010 vdd.n7009 0.0225448
R41371 vdd.n7006 vdd.n7005 0.0225448
R41372 vdd.n7002 vdd.n7001 0.0225448
R41373 vdd.n7003 vdd.n7002 0.0225448
R41374 vdd.n7012 vdd.n7011 0.0225448
R41375 vdd.n7011 vdd.n7010 0.0225448
R41376 vdd.n6992 vdd.n6968 0.0225448
R41377 vdd.n6993 vdd.n6992 0.0225448
R41378 vdd.n6990 vdd.n6989 0.0225448
R41379 vdd.n7032 vdd.n7030 0.0225448
R41380 vdd.n7032 vdd.n7031 0.0225448
R41381 vdd.n7043 vdd.n7042 0.0225448
R41382 vdd.n7042 vdd.n7041 0.0225448
R41383 vdd.n7057 vdd.n7056 0.0225448
R41384 vdd.n7058 vdd.n7057 0.0225448
R41385 vdd.n7054 vdd.n7053 0.0225448
R41386 vdd.n7050 vdd.n7049 0.0225448
R41387 vdd.n7051 vdd.n7050 0.0225448
R41388 vdd.n7060 vdd.n7059 0.0225448
R41389 vdd.n7059 vdd.n7058 0.0225448
R41390 vdd.n7040 vdd.n7016 0.0225448
R41391 vdd.n7041 vdd.n7040 0.0225448
R41392 vdd.n7038 vdd.n7037 0.0225448
R41393 vdd.n7134 vdd.n7132 0.0225448
R41394 vdd.n7134 vdd.n7133 0.0225448
R41395 vdd.n7145 vdd.n7144 0.0225448
R41396 vdd.n7144 vdd.n7143 0.0225448
R41397 vdd.n7159 vdd.n7158 0.0225448
R41398 vdd.n7160 vdd.n7159 0.0225448
R41399 vdd.n7156 vdd.n7155 0.0225448
R41400 vdd.n7152 vdd.n7151 0.0225448
R41401 vdd.n7153 vdd.n7152 0.0225448
R41402 vdd.n7162 vdd.n7161 0.0225448
R41403 vdd.n7161 vdd.n7160 0.0225448
R41404 vdd.n7142 vdd.n7118 0.0225448
R41405 vdd.n7143 vdd.n7142 0.0225448
R41406 vdd.n7140 vdd.n7139 0.0225448
R41407 vdd.n7182 vdd.n7180 0.0225448
R41408 vdd.n7182 vdd.n7181 0.0225448
R41409 vdd.n7193 vdd.n7192 0.0225448
R41410 vdd.n7192 vdd.n7191 0.0225448
R41411 vdd.n7207 vdd.n7206 0.0225448
R41412 vdd.n7208 vdd.n7207 0.0225448
R41413 vdd.n7204 vdd.n7203 0.0225448
R41414 vdd.n7200 vdd.n7199 0.0225448
R41415 vdd.n7201 vdd.n7200 0.0225448
R41416 vdd.n7210 vdd.n7209 0.0225448
R41417 vdd.n7209 vdd.n7208 0.0225448
R41418 vdd.n7190 vdd.n7166 0.0225448
R41419 vdd.n7191 vdd.n7190 0.0225448
R41420 vdd.n7188 vdd.n7187 0.0225448
R41421 vdd.n7230 vdd.n7228 0.0225448
R41422 vdd.n7230 vdd.n7229 0.0225448
R41423 vdd.n7241 vdd.n7240 0.0225448
R41424 vdd.n7240 vdd.n7239 0.0225448
R41425 vdd.n7255 vdd.n7254 0.0225448
R41426 vdd.n7256 vdd.n7255 0.0225448
R41427 vdd.n7252 vdd.n7251 0.0225448
R41428 vdd.n7248 vdd.n7247 0.0225448
R41429 vdd.n7249 vdd.n7248 0.0225448
R41430 vdd.n7258 vdd.n7257 0.0225448
R41431 vdd.n7257 vdd.n7256 0.0225448
R41432 vdd.n7238 vdd.n7214 0.0225448
R41433 vdd.n7239 vdd.n7238 0.0225448
R41434 vdd.n7236 vdd.n7235 0.0225448
R41435 vdd.n7278 vdd.n7276 0.0225448
R41436 vdd.n7278 vdd.n7277 0.0225448
R41437 vdd.n7289 vdd.n7288 0.0225448
R41438 vdd.n7288 vdd.n7287 0.0225448
R41439 vdd.n7303 vdd.n7302 0.0225448
R41440 vdd.n7304 vdd.n7303 0.0225448
R41441 vdd.n7300 vdd.n7299 0.0225448
R41442 vdd.n7296 vdd.n7295 0.0225448
R41443 vdd.n7297 vdd.n7296 0.0225448
R41444 vdd.n7306 vdd.n7305 0.0225448
R41445 vdd.n7305 vdd.n7304 0.0225448
R41446 vdd.n7286 vdd.n7262 0.0225448
R41447 vdd.n7287 vdd.n7286 0.0225448
R41448 vdd.n7284 vdd.n7283 0.0225448
R41449 vdd.n7380 vdd.n7378 0.0225448
R41450 vdd.n7380 vdd.n7379 0.0225448
R41451 vdd.n7391 vdd.n7390 0.0225448
R41452 vdd.n7390 vdd.n7389 0.0225448
R41453 vdd.n7405 vdd.n7404 0.0225448
R41454 vdd.n7406 vdd.n7405 0.0225448
R41455 vdd.n7402 vdd.n7401 0.0225448
R41456 vdd.n7398 vdd.n7397 0.0225448
R41457 vdd.n7399 vdd.n7398 0.0225448
R41458 vdd.n7408 vdd.n7407 0.0225448
R41459 vdd.n7407 vdd.n7406 0.0225448
R41460 vdd.n7388 vdd.n7364 0.0225448
R41461 vdd.n7389 vdd.n7388 0.0225448
R41462 vdd.n7386 vdd.n7385 0.0225448
R41463 vdd.n8900 vdd.n8898 0.0225448
R41464 vdd.n8900 vdd.n8899 0.0225448
R41465 vdd.n8911 vdd.n8910 0.0225448
R41466 vdd.n8910 vdd.n8909 0.0225448
R41467 vdd.n8925 vdd.n8924 0.0225448
R41468 vdd.n8926 vdd.n8925 0.0225448
R41469 vdd.n8922 vdd.n8921 0.0225448
R41470 vdd.n8918 vdd.n8917 0.0225448
R41471 vdd.n8919 vdd.n8918 0.0225448
R41472 vdd.n8928 vdd.n8927 0.0225448
R41473 vdd.n8927 vdd.n8926 0.0225448
R41474 vdd.n8908 vdd.n8884 0.0225448
R41475 vdd.n8909 vdd.n8908 0.0225448
R41476 vdd.n8906 vdd.n8905 0.0225448
R41477 vdd.n7431 vdd.n7430 0.0225448
R41478 vdd.n7439 vdd.n7438 0.0225448
R41479 vdd.n7438 vdd.n7437 0.0225448
R41480 vdd.n7453 vdd.n7452 0.0225448
R41481 vdd.n7454 vdd.n7453 0.0225448
R41482 vdd.n7450 vdd.n7449 0.0225448
R41483 vdd.n7449 vdd.n7448 0.0225448
R41484 vdd.n7446 vdd.n7445 0.0225448
R41485 vdd.n7456 vdd.n7455 0.0225448
R41486 vdd.n7455 vdd.n7454 0.0225448
R41487 vdd.n7436 vdd.n7412 0.0225448
R41488 vdd.n7437 vdd.n7436 0.0225448
R41489 vdd.n7434 vdd.n7428 0.0225448
R41490 vdd.n7434 vdd.n7433 0.0225448
R41491 vdd.n7479 vdd.n7478 0.0225448
R41492 vdd.n7487 vdd.n7486 0.0225448
R41493 vdd.n7486 vdd.n7485 0.0225448
R41494 vdd.n7501 vdd.n7500 0.0225448
R41495 vdd.n7502 vdd.n7501 0.0225448
R41496 vdd.n7498 vdd.n7497 0.0225448
R41497 vdd.n7497 vdd.n7496 0.0225448
R41498 vdd.n7494 vdd.n7493 0.0225448
R41499 vdd.n7504 vdd.n7503 0.0225448
R41500 vdd.n7503 vdd.n7502 0.0225448
R41501 vdd.n7484 vdd.n7460 0.0225448
R41502 vdd.n7485 vdd.n7484 0.0225448
R41503 vdd.n7482 vdd.n7476 0.0225448
R41504 vdd.n7482 vdd.n7481 0.0225448
R41505 vdd.n7580 vdd.n7579 0.0225448
R41506 vdd.n7588 vdd.n7587 0.0225448
R41507 vdd.n7587 vdd.n7586 0.0225448
R41508 vdd.n7602 vdd.n7601 0.0225448
R41509 vdd.n7603 vdd.n7602 0.0225448
R41510 vdd.n7599 vdd.n7598 0.0225448
R41511 vdd.n7598 vdd.n7597 0.0225448
R41512 vdd.n7595 vdd.n7594 0.0225448
R41513 vdd.n7605 vdd.n7604 0.0225448
R41514 vdd.n7604 vdd.n7603 0.0225448
R41515 vdd.n7585 vdd.n7561 0.0225448
R41516 vdd.n7586 vdd.n7585 0.0225448
R41517 vdd.n7583 vdd.n7577 0.0225448
R41518 vdd.n7583 vdd.n7582 0.0225448
R41519 vdd.n7628 vdd.n7627 0.0225448
R41520 vdd.n7636 vdd.n7635 0.0225448
R41521 vdd.n7635 vdd.n7634 0.0225448
R41522 vdd.n7650 vdd.n7649 0.0225448
R41523 vdd.n7651 vdd.n7650 0.0225448
R41524 vdd.n7647 vdd.n7646 0.0225448
R41525 vdd.n7646 vdd.n7645 0.0225448
R41526 vdd.n7643 vdd.n7642 0.0225448
R41527 vdd.n7653 vdd.n7652 0.0225448
R41528 vdd.n7652 vdd.n7651 0.0225448
R41529 vdd.n7633 vdd.n7609 0.0225448
R41530 vdd.n7634 vdd.n7633 0.0225448
R41531 vdd.n7631 vdd.n7625 0.0225448
R41532 vdd.n7631 vdd.n7630 0.0225448
R41533 vdd.n7676 vdd.n7675 0.0225448
R41534 vdd.n7684 vdd.n7683 0.0225448
R41535 vdd.n7683 vdd.n7682 0.0225448
R41536 vdd.n7698 vdd.n7697 0.0225448
R41537 vdd.n7699 vdd.n7698 0.0225448
R41538 vdd.n7695 vdd.n7694 0.0225448
R41539 vdd.n7694 vdd.n7693 0.0225448
R41540 vdd.n7691 vdd.n7690 0.0225448
R41541 vdd.n7701 vdd.n7700 0.0225448
R41542 vdd.n7700 vdd.n7699 0.0225448
R41543 vdd.n7681 vdd.n7657 0.0225448
R41544 vdd.n7682 vdd.n7681 0.0225448
R41545 vdd.n7679 vdd.n7673 0.0225448
R41546 vdd.n7679 vdd.n7678 0.0225448
R41547 vdd.n7724 vdd.n7723 0.0225448
R41548 vdd.n7732 vdd.n7731 0.0225448
R41549 vdd.n7731 vdd.n7730 0.0225448
R41550 vdd.n7746 vdd.n7745 0.0225448
R41551 vdd.n7747 vdd.n7746 0.0225448
R41552 vdd.n7743 vdd.n7742 0.0225448
R41553 vdd.n7742 vdd.n7741 0.0225448
R41554 vdd.n7739 vdd.n7738 0.0225448
R41555 vdd.n7749 vdd.n7748 0.0225448
R41556 vdd.n7748 vdd.n7747 0.0225448
R41557 vdd.n7729 vdd.n7705 0.0225448
R41558 vdd.n7730 vdd.n7729 0.0225448
R41559 vdd.n7727 vdd.n7721 0.0225448
R41560 vdd.n7727 vdd.n7726 0.0225448
R41561 vdd.n7825 vdd.n7824 0.0225448
R41562 vdd.n7833 vdd.n7832 0.0225448
R41563 vdd.n7832 vdd.n7831 0.0225448
R41564 vdd.n7847 vdd.n7846 0.0225448
R41565 vdd.n7848 vdd.n7847 0.0225448
R41566 vdd.n7844 vdd.n7843 0.0225448
R41567 vdd.n7843 vdd.n7842 0.0225448
R41568 vdd.n7840 vdd.n7839 0.0225448
R41569 vdd.n7850 vdd.n7849 0.0225448
R41570 vdd.n7849 vdd.n7848 0.0225448
R41571 vdd.n7830 vdd.n7806 0.0225448
R41572 vdd.n7831 vdd.n7830 0.0225448
R41573 vdd.n7828 vdd.n7822 0.0225448
R41574 vdd.n7828 vdd.n7827 0.0225448
R41575 vdd.n6938 vdd.n6937 0.0225448
R41576 vdd.n6946 vdd.n6945 0.0225448
R41577 vdd.n6945 vdd.n6944 0.0225448
R41578 vdd.n6960 vdd.n6959 0.0225448
R41579 vdd.n6961 vdd.n6960 0.0225448
R41580 vdd.n6957 vdd.n6956 0.0225448
R41581 vdd.n6956 vdd.n6955 0.0225448
R41582 vdd.n6953 vdd.n6952 0.0225448
R41583 vdd.n6963 vdd.n6962 0.0225448
R41584 vdd.n6962 vdd.n6961 0.0225448
R41585 vdd.n6943 vdd.n6919 0.0225448
R41586 vdd.n6944 vdd.n6943 0.0225448
R41587 vdd.n6941 vdd.n6935 0.0225448
R41588 vdd.n6941 vdd.n6940 0.0225448
R41589 vdd.n7873 vdd.n7872 0.0225448
R41590 vdd.n7881 vdd.n7880 0.0225448
R41591 vdd.n7880 vdd.n7879 0.0225448
R41592 vdd.n7895 vdd.n7894 0.0225448
R41593 vdd.n7896 vdd.n7895 0.0225448
R41594 vdd.n7892 vdd.n7891 0.0225448
R41595 vdd.n7891 vdd.n7890 0.0225448
R41596 vdd.n7888 vdd.n7887 0.0225448
R41597 vdd.n7898 vdd.n7897 0.0225448
R41598 vdd.n7897 vdd.n7896 0.0225448
R41599 vdd.n7878 vdd.n7854 0.0225448
R41600 vdd.n7879 vdd.n7878 0.0225448
R41601 vdd.n7876 vdd.n7870 0.0225448
R41602 vdd.n7876 vdd.n7875 0.0225448
R41603 vdd.n7920 vdd.n7919 0.0225448
R41604 vdd.n7928 vdd.n7927 0.0225448
R41605 vdd.n7927 vdd.n7926 0.0225448
R41606 vdd.n7942 vdd.n7941 0.0225448
R41607 vdd.n7943 vdd.n7942 0.0225448
R41608 vdd.n7939 vdd.n7938 0.0225448
R41609 vdd.n7938 vdd.n7937 0.0225448
R41610 vdd.n7935 vdd.n7934 0.0225448
R41611 vdd.n7945 vdd.n7944 0.0225448
R41612 vdd.n7944 vdd.n7943 0.0225448
R41613 vdd.n7925 vdd.n7901 0.0225448
R41614 vdd.n7926 vdd.n7925 0.0225448
R41615 vdd.n7923 vdd.n7917 0.0225448
R41616 vdd.n7923 vdd.n7922 0.0225448
R41617 vdd.n7970 vdd.n7969 0.0225448
R41618 vdd.n7978 vdd.n7977 0.0225448
R41619 vdd.n7977 vdd.n7976 0.0225448
R41620 vdd.n7992 vdd.n7991 0.0225448
R41621 vdd.n7993 vdd.n7992 0.0225448
R41622 vdd.n7989 vdd.n7988 0.0225448
R41623 vdd.n7988 vdd.n7987 0.0225448
R41624 vdd.n7985 vdd.n7984 0.0225448
R41625 vdd.n7995 vdd.n7994 0.0225448
R41626 vdd.n7994 vdd.n7993 0.0225448
R41627 vdd.n7975 vdd.n7951 0.0225448
R41628 vdd.n7976 vdd.n7975 0.0225448
R41629 vdd.n7973 vdd.n7967 0.0225448
R41630 vdd.n7973 vdd.n7972 0.0225448
R41631 vdd.n8020 vdd.n8019 0.0225448
R41632 vdd.n8028 vdd.n8027 0.0225448
R41633 vdd.n8027 vdd.n8026 0.0225448
R41634 vdd.n8042 vdd.n8041 0.0225448
R41635 vdd.n8043 vdd.n8042 0.0225448
R41636 vdd.n8039 vdd.n8038 0.0225448
R41637 vdd.n8038 vdd.n8037 0.0225448
R41638 vdd.n8035 vdd.n8034 0.0225448
R41639 vdd.n8045 vdd.n8044 0.0225448
R41640 vdd.n8044 vdd.n8043 0.0225448
R41641 vdd.n8025 vdd.n8001 0.0225448
R41642 vdd.n8026 vdd.n8025 0.0225448
R41643 vdd.n8023 vdd.n8017 0.0225448
R41644 vdd.n8023 vdd.n8022 0.0225448
R41645 vdd.n8068 vdd.n8067 0.0225448
R41646 vdd.n8076 vdd.n8075 0.0225448
R41647 vdd.n8075 vdd.n8074 0.0225448
R41648 vdd.n8090 vdd.n8089 0.0225448
R41649 vdd.n8091 vdd.n8090 0.0225448
R41650 vdd.n8087 vdd.n8086 0.0225448
R41651 vdd.n8086 vdd.n8085 0.0225448
R41652 vdd.n8083 vdd.n8082 0.0225448
R41653 vdd.n8093 vdd.n8092 0.0225448
R41654 vdd.n8092 vdd.n8091 0.0225448
R41655 vdd.n8073 vdd.n8049 0.0225448
R41656 vdd.n8074 vdd.n8073 0.0225448
R41657 vdd.n8071 vdd.n8065 0.0225448
R41658 vdd.n8071 vdd.n8070 0.0225448
R41659 vdd.n7796 vdd.n7795 0.0225448
R41660 vdd.n7793 vdd.n7792 0.0225448
R41661 vdd.n7792 vdd.n7791 0.0225448
R41662 vdd.n7782 vdd.n7781 0.0225448
R41663 vdd.n7783 vdd.n7782 0.0225448
R41664 vdd.n7779 vdd.n7778 0.0225448
R41665 vdd.n7778 vdd.n7777 0.0225448
R41666 vdd.n7775 vdd.n7774 0.0225448
R41667 vdd.n7784 vdd.n7766 0.0225448
R41668 vdd.n7784 vdd.n7783 0.0225448
R41669 vdd.n7790 vdd.n7789 0.0225448
R41670 vdd.n7791 vdd.n7790 0.0225448
R41671 vdd.n7800 vdd.n7799 0.0225448
R41672 vdd.n7799 vdd.n7798 0.0225448
R41673 vdd.n8119 vdd.n8118 0.0225448
R41674 vdd.n8127 vdd.n8126 0.0225448
R41675 vdd.n8126 vdd.n8125 0.0225448
R41676 vdd.n8141 vdd.n8140 0.0225448
R41677 vdd.n8142 vdd.n8141 0.0225448
R41678 vdd.n8138 vdd.n8137 0.0225448
R41679 vdd.n8137 vdd.n8136 0.0225448
R41680 vdd.n8134 vdd.n8133 0.0225448
R41681 vdd.n8144 vdd.n8143 0.0225448
R41682 vdd.n8143 vdd.n8142 0.0225448
R41683 vdd.n8124 vdd.n8100 0.0225448
R41684 vdd.n8125 vdd.n8124 0.0225448
R41685 vdd.n8122 vdd.n8116 0.0225448
R41686 vdd.n8122 vdd.n8121 0.0225448
R41687 vdd.n8166 vdd.n8165 0.0225448
R41688 vdd.n8174 vdd.n8173 0.0225448
R41689 vdd.n8173 vdd.n8172 0.0225448
R41690 vdd.n8188 vdd.n8187 0.0225448
R41691 vdd.n8189 vdd.n8188 0.0225448
R41692 vdd.n8185 vdd.n8184 0.0225448
R41693 vdd.n8184 vdd.n8183 0.0225448
R41694 vdd.n8181 vdd.n8180 0.0225448
R41695 vdd.n8191 vdd.n8190 0.0225448
R41696 vdd.n8190 vdd.n8189 0.0225448
R41697 vdd.n8171 vdd.n8147 0.0225448
R41698 vdd.n8172 vdd.n8171 0.0225448
R41699 vdd.n8169 vdd.n8163 0.0225448
R41700 vdd.n8169 vdd.n8168 0.0225448
R41701 vdd.n8214 vdd.n8213 0.0225448
R41702 vdd.n8222 vdd.n8221 0.0225448
R41703 vdd.n8221 vdd.n8220 0.0225448
R41704 vdd.n8236 vdd.n8235 0.0225448
R41705 vdd.n8237 vdd.n8236 0.0225448
R41706 vdd.n8233 vdd.n8232 0.0225448
R41707 vdd.n8232 vdd.n8231 0.0225448
R41708 vdd.n8229 vdd.n8228 0.0225448
R41709 vdd.n8239 vdd.n8238 0.0225448
R41710 vdd.n8238 vdd.n8237 0.0225448
R41711 vdd.n8219 vdd.n8195 0.0225448
R41712 vdd.n8220 vdd.n8219 0.0225448
R41713 vdd.n8217 vdd.n8211 0.0225448
R41714 vdd.n8217 vdd.n8216 0.0225448
R41715 vdd.n8265 vdd.n8264 0.0225448
R41716 vdd.n8273 vdd.n8272 0.0225448
R41717 vdd.n8272 vdd.n8271 0.0225448
R41718 vdd.n8287 vdd.n8286 0.0225448
R41719 vdd.n8288 vdd.n8287 0.0225448
R41720 vdd.n8284 vdd.n8283 0.0225448
R41721 vdd.n8283 vdd.n8282 0.0225448
R41722 vdd.n8280 vdd.n8279 0.0225448
R41723 vdd.n8290 vdd.n8289 0.0225448
R41724 vdd.n8289 vdd.n8288 0.0225448
R41725 vdd.n8270 vdd.n8246 0.0225448
R41726 vdd.n8271 vdd.n8270 0.0225448
R41727 vdd.n8268 vdd.n8262 0.0225448
R41728 vdd.n8268 vdd.n8267 0.0225448
R41729 vdd.n8315 vdd.n8314 0.0225448
R41730 vdd.n8323 vdd.n8322 0.0225448
R41731 vdd.n8322 vdd.n8321 0.0225448
R41732 vdd.n8337 vdd.n8336 0.0225448
R41733 vdd.n8338 vdd.n8337 0.0225448
R41734 vdd.n8334 vdd.n8333 0.0225448
R41735 vdd.n8333 vdd.n8332 0.0225448
R41736 vdd.n8330 vdd.n8329 0.0225448
R41737 vdd.n8340 vdd.n8339 0.0225448
R41738 vdd.n8339 vdd.n8338 0.0225448
R41739 vdd.n8320 vdd.n8296 0.0225448
R41740 vdd.n8321 vdd.n8320 0.0225448
R41741 vdd.n8318 vdd.n8312 0.0225448
R41742 vdd.n8318 vdd.n8317 0.0225448
R41743 vdd.n8363 vdd.n8362 0.0225448
R41744 vdd.n8371 vdd.n8370 0.0225448
R41745 vdd.n8370 vdd.n8369 0.0225448
R41746 vdd.n8385 vdd.n8384 0.0225448
R41747 vdd.n8386 vdd.n8385 0.0225448
R41748 vdd.n8382 vdd.n8381 0.0225448
R41749 vdd.n8381 vdd.n8380 0.0225448
R41750 vdd.n8378 vdd.n8377 0.0225448
R41751 vdd.n8388 vdd.n8387 0.0225448
R41752 vdd.n8387 vdd.n8386 0.0225448
R41753 vdd.n8368 vdd.n8344 0.0225448
R41754 vdd.n8369 vdd.n8368 0.0225448
R41755 vdd.n8366 vdd.n8360 0.0225448
R41756 vdd.n8366 vdd.n8365 0.0225448
R41757 vdd.n8413 vdd.n8412 0.0225448
R41758 vdd.n8421 vdd.n8420 0.0225448
R41759 vdd.n8420 vdd.n8419 0.0225448
R41760 vdd.n8435 vdd.n8434 0.0225448
R41761 vdd.n8436 vdd.n8435 0.0225448
R41762 vdd.n8432 vdd.n8431 0.0225448
R41763 vdd.n8431 vdd.n8430 0.0225448
R41764 vdd.n8428 vdd.n8427 0.0225448
R41765 vdd.n8438 vdd.n8437 0.0225448
R41766 vdd.n8437 vdd.n8436 0.0225448
R41767 vdd.n8418 vdd.n8394 0.0225448
R41768 vdd.n8419 vdd.n8418 0.0225448
R41769 vdd.n8416 vdd.n8410 0.0225448
R41770 vdd.n8416 vdd.n8415 0.0225448
R41771 vdd.n8460 vdd.n8459 0.0225448
R41772 vdd.n8468 vdd.n8467 0.0225448
R41773 vdd.n8467 vdd.n8466 0.0225448
R41774 vdd.n8482 vdd.n8481 0.0225448
R41775 vdd.n8483 vdd.n8482 0.0225448
R41776 vdd.n8479 vdd.n8478 0.0225448
R41777 vdd.n8478 vdd.n8477 0.0225448
R41778 vdd.n8475 vdd.n8474 0.0225448
R41779 vdd.n8485 vdd.n8484 0.0225448
R41780 vdd.n8484 vdd.n8483 0.0225448
R41781 vdd.n8465 vdd.n8441 0.0225448
R41782 vdd.n8466 vdd.n8465 0.0225448
R41783 vdd.n8463 vdd.n8457 0.0225448
R41784 vdd.n8463 vdd.n8462 0.0225448
R41785 vdd.n8510 vdd.n8509 0.0225448
R41786 vdd.n8518 vdd.n8517 0.0225448
R41787 vdd.n8517 vdd.n8516 0.0225448
R41788 vdd.n8532 vdd.n8531 0.0225448
R41789 vdd.n8533 vdd.n8532 0.0225448
R41790 vdd.n8529 vdd.n8528 0.0225448
R41791 vdd.n8528 vdd.n8527 0.0225448
R41792 vdd.n8525 vdd.n8524 0.0225448
R41793 vdd.n8535 vdd.n8534 0.0225448
R41794 vdd.n8534 vdd.n8533 0.0225448
R41795 vdd.n8515 vdd.n8491 0.0225448
R41796 vdd.n8516 vdd.n8515 0.0225448
R41797 vdd.n8513 vdd.n8507 0.0225448
R41798 vdd.n8513 vdd.n8512 0.0225448
R41799 vdd.n8560 vdd.n8559 0.0225448
R41800 vdd.n8568 vdd.n8567 0.0225448
R41801 vdd.n8567 vdd.n8566 0.0225448
R41802 vdd.n8582 vdd.n8581 0.0225448
R41803 vdd.n8583 vdd.n8582 0.0225448
R41804 vdd.n8579 vdd.n8578 0.0225448
R41805 vdd.n8578 vdd.n8577 0.0225448
R41806 vdd.n8575 vdd.n8574 0.0225448
R41807 vdd.n8585 vdd.n8584 0.0225448
R41808 vdd.n8584 vdd.n8583 0.0225448
R41809 vdd.n8565 vdd.n8541 0.0225448
R41810 vdd.n8566 vdd.n8565 0.0225448
R41811 vdd.n8563 vdd.n8557 0.0225448
R41812 vdd.n8563 vdd.n8562 0.0225448
R41813 vdd.n8608 vdd.n8607 0.0225448
R41814 vdd.n8616 vdd.n8615 0.0225448
R41815 vdd.n8615 vdd.n8614 0.0225448
R41816 vdd.n8630 vdd.n8629 0.0225448
R41817 vdd.n8631 vdd.n8630 0.0225448
R41818 vdd.n8627 vdd.n8626 0.0225448
R41819 vdd.n8626 vdd.n8625 0.0225448
R41820 vdd.n8623 vdd.n8622 0.0225448
R41821 vdd.n8633 vdd.n8632 0.0225448
R41822 vdd.n8632 vdd.n8631 0.0225448
R41823 vdd.n8613 vdd.n8589 0.0225448
R41824 vdd.n8614 vdd.n8613 0.0225448
R41825 vdd.n8611 vdd.n8605 0.0225448
R41826 vdd.n8611 vdd.n8610 0.0225448
R41827 vdd.n7551 vdd.n7550 0.0225448
R41828 vdd.n7548 vdd.n7547 0.0225448
R41829 vdd.n7547 vdd.n7546 0.0225448
R41830 vdd.n7537 vdd.n7536 0.0225448
R41831 vdd.n7538 vdd.n7537 0.0225448
R41832 vdd.n7534 vdd.n7533 0.0225448
R41833 vdd.n7533 vdd.n7532 0.0225448
R41834 vdd.n7530 vdd.n7529 0.0225448
R41835 vdd.n7539 vdd.n7521 0.0225448
R41836 vdd.n7539 vdd.n7538 0.0225448
R41837 vdd.n7545 vdd.n7544 0.0225448
R41838 vdd.n7546 vdd.n7545 0.0225448
R41839 vdd.n7555 vdd.n7554 0.0225448
R41840 vdd.n7554 vdd.n7553 0.0225448
R41841 vdd.n8659 vdd.n8658 0.0225448
R41842 vdd.n8667 vdd.n8666 0.0225448
R41843 vdd.n8666 vdd.n8665 0.0225448
R41844 vdd.n8681 vdd.n8680 0.0225448
R41845 vdd.n8682 vdd.n8681 0.0225448
R41846 vdd.n8678 vdd.n8677 0.0225448
R41847 vdd.n8677 vdd.n8676 0.0225448
R41848 vdd.n8674 vdd.n8673 0.0225448
R41849 vdd.n8684 vdd.n8683 0.0225448
R41850 vdd.n8683 vdd.n8682 0.0225448
R41851 vdd.n8664 vdd.n8640 0.0225448
R41852 vdd.n8665 vdd.n8664 0.0225448
R41853 vdd.n8662 vdd.n8656 0.0225448
R41854 vdd.n8662 vdd.n8661 0.0225448
R41855 vdd.n8706 vdd.n8705 0.0225448
R41856 vdd.n8714 vdd.n8713 0.0225448
R41857 vdd.n8713 vdd.n8712 0.0225448
R41858 vdd.n8728 vdd.n8727 0.0225448
R41859 vdd.n8729 vdd.n8728 0.0225448
R41860 vdd.n8725 vdd.n8724 0.0225448
R41861 vdd.n8724 vdd.n8723 0.0225448
R41862 vdd.n8721 vdd.n8720 0.0225448
R41863 vdd.n8731 vdd.n8730 0.0225448
R41864 vdd.n8730 vdd.n8729 0.0225448
R41865 vdd.n8711 vdd.n8687 0.0225448
R41866 vdd.n8712 vdd.n8711 0.0225448
R41867 vdd.n8709 vdd.n8703 0.0225448
R41868 vdd.n8709 vdd.n8708 0.0225448
R41869 vdd.n8756 vdd.n8755 0.0225448
R41870 vdd.n8764 vdd.n8763 0.0225448
R41871 vdd.n8763 vdd.n8762 0.0225448
R41872 vdd.n8778 vdd.n8777 0.0225448
R41873 vdd.n8779 vdd.n8778 0.0225448
R41874 vdd.n8775 vdd.n8774 0.0225448
R41875 vdd.n8774 vdd.n8773 0.0225448
R41876 vdd.n8771 vdd.n8770 0.0225448
R41877 vdd.n8781 vdd.n8780 0.0225448
R41878 vdd.n8780 vdd.n8779 0.0225448
R41879 vdd.n8761 vdd.n8737 0.0225448
R41880 vdd.n8762 vdd.n8761 0.0225448
R41881 vdd.n8759 vdd.n8753 0.0225448
R41882 vdd.n8759 vdd.n8758 0.0225448
R41883 vdd.n8806 vdd.n8805 0.0225448
R41884 vdd.n8814 vdd.n8813 0.0225448
R41885 vdd.n8813 vdd.n8812 0.0225448
R41886 vdd.n8828 vdd.n8827 0.0225448
R41887 vdd.n8829 vdd.n8828 0.0225448
R41888 vdd.n8825 vdd.n8824 0.0225448
R41889 vdd.n8824 vdd.n8823 0.0225448
R41890 vdd.n8821 vdd.n8820 0.0225448
R41891 vdd.n8831 vdd.n8830 0.0225448
R41892 vdd.n8830 vdd.n8829 0.0225448
R41893 vdd.n8811 vdd.n8787 0.0225448
R41894 vdd.n8812 vdd.n8811 0.0225448
R41895 vdd.n8809 vdd.n8803 0.0225448
R41896 vdd.n8809 vdd.n8808 0.0225448
R41897 vdd.n8854 vdd.n8853 0.0225448
R41898 vdd.n8862 vdd.n8861 0.0225448
R41899 vdd.n8861 vdd.n8860 0.0225448
R41900 vdd.n8876 vdd.n8875 0.0225448
R41901 vdd.n8877 vdd.n8876 0.0225448
R41902 vdd.n8873 vdd.n8872 0.0225448
R41903 vdd.n8872 vdd.n8871 0.0225448
R41904 vdd.n8869 vdd.n8868 0.0225448
R41905 vdd.n8879 vdd.n8878 0.0225448
R41906 vdd.n8878 vdd.n8877 0.0225448
R41907 vdd.n8859 vdd.n8835 0.0225448
R41908 vdd.n8860 vdd.n8859 0.0225448
R41909 vdd.n8857 vdd.n8851 0.0225448
R41910 vdd.n8857 vdd.n8856 0.0225448
R41911 vdd.n8997 vdd.n8995 0.0225448
R41912 vdd.n8997 vdd.n8996 0.0225448
R41913 vdd.n9008 vdd.n9007 0.0225448
R41914 vdd.n9007 vdd.n9006 0.0225448
R41915 vdd.n9022 vdd.n9021 0.0225448
R41916 vdd.n9023 vdd.n9022 0.0225448
R41917 vdd.n9019 vdd.n9018 0.0225448
R41918 vdd.n9015 vdd.n9014 0.0225448
R41919 vdd.n9016 vdd.n9015 0.0225448
R41920 vdd.n9025 vdd.n9024 0.0225448
R41921 vdd.n9024 vdd.n9023 0.0225448
R41922 vdd.n9005 vdd.n8981 0.0225448
R41923 vdd.n9006 vdd.n9005 0.0225448
R41924 vdd.n9003 vdd.n9002 0.0225448
R41925 vdd.n8949 vdd.n8947 0.0225448
R41926 vdd.n8949 vdd.n8948 0.0225448
R41927 vdd.n8960 vdd.n8959 0.0225448
R41928 vdd.n8959 vdd.n8958 0.0225448
R41929 vdd.n8974 vdd.n8973 0.0225448
R41930 vdd.n8975 vdd.n8974 0.0225448
R41931 vdd.n8971 vdd.n8970 0.0225448
R41932 vdd.n8967 vdd.n8966 0.0225448
R41933 vdd.n8968 vdd.n8967 0.0225448
R41934 vdd.n8977 vdd.n8976 0.0225448
R41935 vdd.n8976 vdd.n8975 0.0225448
R41936 vdd.n8957 vdd.n8933 0.0225448
R41937 vdd.n8958 vdd.n8957 0.0225448
R41938 vdd.n8955 vdd.n8954 0.0225448
R41939 vdd.n9046 vdd.n9044 0.0225448
R41940 vdd.n9046 vdd.n9045 0.0225448
R41941 vdd.n9057 vdd.n9056 0.0225448
R41942 vdd.n9056 vdd.n9055 0.0225448
R41943 vdd.n9071 vdd.n9070 0.0225448
R41944 vdd.n9072 vdd.n9071 0.0225448
R41945 vdd.n9068 vdd.n9067 0.0225448
R41946 vdd.n9064 vdd.n9063 0.0225448
R41947 vdd.n9065 vdd.n9064 0.0225448
R41948 vdd.n9074 vdd.n9073 0.0225448
R41949 vdd.n9073 vdd.n9072 0.0225448
R41950 vdd.n9054 vdd.n9030 0.0225448
R41951 vdd.n9055 vdd.n9054 0.0225448
R41952 vdd.n9052 vdd.n9051 0.0225448
R41953 vdd.n9096 vdd.n9094 0.0225448
R41954 vdd.n9096 vdd.n9095 0.0225448
R41955 vdd.n9107 vdd.n9106 0.0225448
R41956 vdd.n9106 vdd.n9105 0.0225448
R41957 vdd.n9121 vdd.n9120 0.0225448
R41958 vdd.n9122 vdd.n9121 0.0225448
R41959 vdd.n9118 vdd.n9117 0.0225448
R41960 vdd.n9114 vdd.n9113 0.0225448
R41961 vdd.n9115 vdd.n9114 0.0225448
R41962 vdd.n9124 vdd.n9123 0.0225448
R41963 vdd.n9123 vdd.n9122 0.0225448
R41964 vdd.n9104 vdd.n9080 0.0225448
R41965 vdd.n9105 vdd.n9104 0.0225448
R41966 vdd.n9102 vdd.n9101 0.0225448
R41967 vdd.n9144 vdd.n9142 0.0225448
R41968 vdd.n9144 vdd.n9143 0.0225448
R41969 vdd.n9155 vdd.n9154 0.0225448
R41970 vdd.n9154 vdd.n9153 0.0225448
R41971 vdd.n9169 vdd.n9168 0.0225448
R41972 vdd.n9170 vdd.n9169 0.0225448
R41973 vdd.n9166 vdd.n9165 0.0225448
R41974 vdd.n9162 vdd.n9161 0.0225448
R41975 vdd.n9163 vdd.n9162 0.0225448
R41976 vdd.n9172 vdd.n9171 0.0225448
R41977 vdd.n9171 vdd.n9170 0.0225448
R41978 vdd.n9152 vdd.n9128 0.0225448
R41979 vdd.n9153 vdd.n9152 0.0225448
R41980 vdd.n9150 vdd.n9149 0.0225448
R41981 vdd.n7331 vdd.n7330 0.0225448
R41982 vdd.n7332 vdd.n7331 0.0225448
R41983 vdd.n7328 vdd.n7321 0.0225448
R41984 vdd.n7339 vdd.n7321 0.0225448
R41985 vdd.n7341 vdd.n7340 0.0225448
R41986 vdd.n7342 vdd.n7341 0.0225448
R41987 vdd.n7356 vdd.n7355 0.0225448
R41988 vdd.n7352 vdd.n7311 0.0225448
R41989 vdd.n7353 vdd.n7352 0.0225448
R41990 vdd.n7347 vdd.n7316 0.0225448
R41991 vdd.n7342 vdd.n7316 0.0225448
R41992 vdd.n7338 vdd.n7337 0.0225448
R41993 vdd.n7339 vdd.n7338 0.0225448
R41994 vdd.n7335 vdd.n7334 0.0225448
R41995 vdd.n9292 vdd.n9290 0.0225448
R41996 vdd.n9292 vdd.n9291 0.0225448
R41997 vdd.n9303 vdd.n9302 0.0225448
R41998 vdd.n9302 vdd.n9301 0.0225448
R41999 vdd.n9317 vdd.n9316 0.0225448
R42000 vdd.n9318 vdd.n9317 0.0225448
R42001 vdd.n9314 vdd.n9313 0.0225448
R42002 vdd.n9310 vdd.n9309 0.0225448
R42003 vdd.n9311 vdd.n9310 0.0225448
R42004 vdd.n9320 vdd.n9319 0.0225448
R42005 vdd.n9319 vdd.n9318 0.0225448
R42006 vdd.n9300 vdd.n9276 0.0225448
R42007 vdd.n9301 vdd.n9300 0.0225448
R42008 vdd.n9298 vdd.n9297 0.0225448
R42009 vdd.n9243 vdd.n9241 0.0225448
R42010 vdd.n9243 vdd.n9242 0.0225448
R42011 vdd.n9254 vdd.n9253 0.0225448
R42012 vdd.n9253 vdd.n9252 0.0225448
R42013 vdd.n9268 vdd.n9267 0.0225448
R42014 vdd.n9269 vdd.n9268 0.0225448
R42015 vdd.n9265 vdd.n9264 0.0225448
R42016 vdd.n9261 vdd.n9260 0.0225448
R42017 vdd.n9262 vdd.n9261 0.0225448
R42018 vdd.n9271 vdd.n9270 0.0225448
R42019 vdd.n9270 vdd.n9269 0.0225448
R42020 vdd.n9251 vdd.n9227 0.0225448
R42021 vdd.n9252 vdd.n9251 0.0225448
R42022 vdd.n9249 vdd.n9248 0.0225448
R42023 vdd.n9195 vdd.n9193 0.0225448
R42024 vdd.n9195 vdd.n9194 0.0225448
R42025 vdd.n9206 vdd.n9205 0.0225448
R42026 vdd.n9205 vdd.n9204 0.0225448
R42027 vdd.n9220 vdd.n9219 0.0225448
R42028 vdd.n9221 vdd.n9220 0.0225448
R42029 vdd.n9217 vdd.n9216 0.0225448
R42030 vdd.n9213 vdd.n9212 0.0225448
R42031 vdd.n9214 vdd.n9213 0.0225448
R42032 vdd.n9223 vdd.n9222 0.0225448
R42033 vdd.n9222 vdd.n9221 0.0225448
R42034 vdd.n9203 vdd.n9179 0.0225448
R42035 vdd.n9204 vdd.n9203 0.0225448
R42036 vdd.n9201 vdd.n9200 0.0225448
R42037 vdd.n9341 vdd.n9339 0.0225448
R42038 vdd.n9341 vdd.n9340 0.0225448
R42039 vdd.n9352 vdd.n9351 0.0225448
R42040 vdd.n9351 vdd.n9350 0.0225448
R42041 vdd.n9366 vdd.n9365 0.0225448
R42042 vdd.n9367 vdd.n9366 0.0225448
R42043 vdd.n9363 vdd.n9362 0.0225448
R42044 vdd.n9359 vdd.n9358 0.0225448
R42045 vdd.n9360 vdd.n9359 0.0225448
R42046 vdd.n9369 vdd.n9368 0.0225448
R42047 vdd.n9368 vdd.n9367 0.0225448
R42048 vdd.n9349 vdd.n9325 0.0225448
R42049 vdd.n9350 vdd.n9349 0.0225448
R42050 vdd.n9347 vdd.n9346 0.0225448
R42051 vdd.n9391 vdd.n9389 0.0225448
R42052 vdd.n9391 vdd.n9390 0.0225448
R42053 vdd.n9402 vdd.n9401 0.0225448
R42054 vdd.n9401 vdd.n9400 0.0225448
R42055 vdd.n9416 vdd.n9415 0.0225448
R42056 vdd.n9417 vdd.n9416 0.0225448
R42057 vdd.n9413 vdd.n9412 0.0225448
R42058 vdd.n9409 vdd.n9408 0.0225448
R42059 vdd.n9410 vdd.n9409 0.0225448
R42060 vdd.n9419 vdd.n9418 0.0225448
R42061 vdd.n9418 vdd.n9417 0.0225448
R42062 vdd.n9399 vdd.n9375 0.0225448
R42063 vdd.n9400 vdd.n9399 0.0225448
R42064 vdd.n9397 vdd.n9396 0.0225448
R42065 vdd.n9439 vdd.n9437 0.0225448
R42066 vdd.n9439 vdd.n9438 0.0225448
R42067 vdd.n9450 vdd.n9449 0.0225448
R42068 vdd.n9449 vdd.n9448 0.0225448
R42069 vdd.n9464 vdd.n9463 0.0225448
R42070 vdd.n9465 vdd.n9464 0.0225448
R42071 vdd.n9461 vdd.n9460 0.0225448
R42072 vdd.n9457 vdd.n9456 0.0225448
R42073 vdd.n9458 vdd.n9457 0.0225448
R42074 vdd.n9467 vdd.n9466 0.0225448
R42075 vdd.n9466 vdd.n9465 0.0225448
R42076 vdd.n9447 vdd.n9423 0.0225448
R42077 vdd.n9448 vdd.n9447 0.0225448
R42078 vdd.n9445 vdd.n9444 0.0225448
R42079 vdd.n9537 vdd.n9535 0.0225448
R42080 vdd.n9537 vdd.n9536 0.0225448
R42081 vdd.n9548 vdd.n9547 0.0225448
R42082 vdd.n9547 vdd.n9546 0.0225448
R42083 vdd.n9562 vdd.n9561 0.0225448
R42084 vdd.n9563 vdd.n9562 0.0225448
R42085 vdd.n9559 vdd.n9558 0.0225448
R42086 vdd.n9555 vdd.n9554 0.0225448
R42087 vdd.n9556 vdd.n9555 0.0225448
R42088 vdd.n9565 vdd.n9564 0.0225448
R42089 vdd.n9564 vdd.n9563 0.0225448
R42090 vdd.n9545 vdd.n9521 0.0225448
R42091 vdd.n9546 vdd.n9545 0.0225448
R42092 vdd.n9543 vdd.n9542 0.0225448
R42093 vdd.n9489 vdd.n9487 0.0225448
R42094 vdd.n9489 vdd.n9488 0.0225448
R42095 vdd.n9500 vdd.n9499 0.0225448
R42096 vdd.n9499 vdd.n9498 0.0225448
R42097 vdd.n9514 vdd.n9513 0.0225448
R42098 vdd.n9515 vdd.n9514 0.0225448
R42099 vdd.n9511 vdd.n9510 0.0225448
R42100 vdd.n9507 vdd.n9506 0.0225448
R42101 vdd.n9508 vdd.n9507 0.0225448
R42102 vdd.n9517 vdd.n9516 0.0225448
R42103 vdd.n9516 vdd.n9515 0.0225448
R42104 vdd.n9497 vdd.n9473 0.0225448
R42105 vdd.n9498 vdd.n9497 0.0225448
R42106 vdd.n9495 vdd.n9494 0.0225448
R42107 vdd.n9586 vdd.n9584 0.0225448
R42108 vdd.n9586 vdd.n9585 0.0225448
R42109 vdd.n9597 vdd.n9596 0.0225448
R42110 vdd.n9596 vdd.n9595 0.0225448
R42111 vdd.n9611 vdd.n9610 0.0225448
R42112 vdd.n9612 vdd.n9611 0.0225448
R42113 vdd.n9608 vdd.n9607 0.0225448
R42114 vdd.n9604 vdd.n9603 0.0225448
R42115 vdd.n9605 vdd.n9604 0.0225448
R42116 vdd.n9614 vdd.n9613 0.0225448
R42117 vdd.n9613 vdd.n9612 0.0225448
R42118 vdd.n9594 vdd.n9570 0.0225448
R42119 vdd.n9595 vdd.n9594 0.0225448
R42120 vdd.n9592 vdd.n9591 0.0225448
R42121 vdd.n9636 vdd.n9634 0.0225448
R42122 vdd.n9636 vdd.n9635 0.0225448
R42123 vdd.n9647 vdd.n9646 0.0225448
R42124 vdd.n9646 vdd.n9645 0.0225448
R42125 vdd.n9661 vdd.n9660 0.0225448
R42126 vdd.n9662 vdd.n9661 0.0225448
R42127 vdd.n9658 vdd.n9657 0.0225448
R42128 vdd.n9654 vdd.n9653 0.0225448
R42129 vdd.n9655 vdd.n9654 0.0225448
R42130 vdd.n9664 vdd.n9663 0.0225448
R42131 vdd.n9663 vdd.n9662 0.0225448
R42132 vdd.n9644 vdd.n9620 0.0225448
R42133 vdd.n9645 vdd.n9644 0.0225448
R42134 vdd.n9642 vdd.n9641 0.0225448
R42135 vdd.n9684 vdd.n9682 0.0225448
R42136 vdd.n9684 vdd.n9683 0.0225448
R42137 vdd.n9695 vdd.n9694 0.0225448
R42138 vdd.n9694 vdd.n9693 0.0225448
R42139 vdd.n9709 vdd.n9708 0.0225448
R42140 vdd.n9710 vdd.n9709 0.0225448
R42141 vdd.n9706 vdd.n9705 0.0225448
R42142 vdd.n9702 vdd.n9701 0.0225448
R42143 vdd.n9703 vdd.n9702 0.0225448
R42144 vdd.n9712 vdd.n9711 0.0225448
R42145 vdd.n9711 vdd.n9710 0.0225448
R42146 vdd.n9692 vdd.n9668 0.0225448
R42147 vdd.n9693 vdd.n9692 0.0225448
R42148 vdd.n9690 vdd.n9689 0.0225448
R42149 vdd.n7085 vdd.n7084 0.0225448
R42150 vdd.n7086 vdd.n7085 0.0225448
R42151 vdd.n7082 vdd.n7075 0.0225448
R42152 vdd.n7093 vdd.n7075 0.0225448
R42153 vdd.n7095 vdd.n7094 0.0225448
R42154 vdd.n7096 vdd.n7095 0.0225448
R42155 vdd.n7110 vdd.n7109 0.0225448
R42156 vdd.n7106 vdd.n7065 0.0225448
R42157 vdd.n7107 vdd.n7106 0.0225448
R42158 vdd.n7101 vdd.n7070 0.0225448
R42159 vdd.n7096 vdd.n7070 0.0225448
R42160 vdd.n7092 vdd.n7091 0.0225448
R42161 vdd.n7093 vdd.n7092 0.0225448
R42162 vdd.n7089 vdd.n7088 0.0225448
R42163 vdd.n9783 vdd.n9781 0.0225448
R42164 vdd.n9783 vdd.n9782 0.0225448
R42165 vdd.n9794 vdd.n9793 0.0225448
R42166 vdd.n9793 vdd.n9792 0.0225448
R42167 vdd.n9808 vdd.n9807 0.0225448
R42168 vdd.n9809 vdd.n9808 0.0225448
R42169 vdd.n9805 vdd.n9804 0.0225448
R42170 vdd.n9801 vdd.n9800 0.0225448
R42171 vdd.n9802 vdd.n9801 0.0225448
R42172 vdd.n9811 vdd.n9810 0.0225448
R42173 vdd.n9810 vdd.n9809 0.0225448
R42174 vdd.n9791 vdd.n9767 0.0225448
R42175 vdd.n9792 vdd.n9791 0.0225448
R42176 vdd.n9789 vdd.n9788 0.0225448
R42177 vdd.n9735 vdd.n9733 0.0225448
R42178 vdd.n9735 vdd.n9734 0.0225448
R42179 vdd.n9746 vdd.n9745 0.0225448
R42180 vdd.n9745 vdd.n9744 0.0225448
R42181 vdd.n9760 vdd.n9759 0.0225448
R42182 vdd.n9761 vdd.n9760 0.0225448
R42183 vdd.n9757 vdd.n9756 0.0225448
R42184 vdd.n9753 vdd.n9752 0.0225448
R42185 vdd.n9754 vdd.n9753 0.0225448
R42186 vdd.n9763 vdd.n9762 0.0225448
R42187 vdd.n9762 vdd.n9761 0.0225448
R42188 vdd.n9743 vdd.n9719 0.0225448
R42189 vdd.n9744 vdd.n9743 0.0225448
R42190 vdd.n9741 vdd.n9740 0.0225448
R42191 vdd.n9832 vdd.n9830 0.0225448
R42192 vdd.n9832 vdd.n9831 0.0225448
R42193 vdd.n9843 vdd.n9842 0.0225448
R42194 vdd.n9842 vdd.n9841 0.0225448
R42195 vdd.n9857 vdd.n9856 0.0225448
R42196 vdd.n9858 vdd.n9857 0.0225448
R42197 vdd.n9854 vdd.n9853 0.0225448
R42198 vdd.n9850 vdd.n9849 0.0225448
R42199 vdd.n9851 vdd.n9850 0.0225448
R42200 vdd.n9860 vdd.n9859 0.0225448
R42201 vdd.n9859 vdd.n9858 0.0225448
R42202 vdd.n9840 vdd.n9816 0.0225448
R42203 vdd.n9841 vdd.n9840 0.0225448
R42204 vdd.n9838 vdd.n9837 0.0225448
R42205 vdd.n9882 vdd.n9880 0.0225448
R42206 vdd.n9882 vdd.n9881 0.0225448
R42207 vdd.n9893 vdd.n9892 0.0225448
R42208 vdd.n9892 vdd.n9891 0.0225448
R42209 vdd.n9907 vdd.n9906 0.0225448
R42210 vdd.n9908 vdd.n9907 0.0225448
R42211 vdd.n9904 vdd.n9903 0.0225448
R42212 vdd.n9900 vdd.n9899 0.0225448
R42213 vdd.n9901 vdd.n9900 0.0225448
R42214 vdd.n9910 vdd.n9909 0.0225448
R42215 vdd.n9909 vdd.n9908 0.0225448
R42216 vdd.n9890 vdd.n9866 0.0225448
R42217 vdd.n9891 vdd.n9890 0.0225448
R42218 vdd.n9888 vdd.n9887 0.0225448
R42219 vdd.n9930 vdd.n9928 0.0225448
R42220 vdd.n9930 vdd.n9929 0.0225448
R42221 vdd.n9941 vdd.n9940 0.0225448
R42222 vdd.n9940 vdd.n9939 0.0225448
R42223 vdd.n9955 vdd.n9954 0.0225448
R42224 vdd.n9956 vdd.n9955 0.0225448
R42225 vdd.n9952 vdd.n9951 0.0225448
R42226 vdd.n9948 vdd.n9947 0.0225448
R42227 vdd.n9949 vdd.n9948 0.0225448
R42228 vdd.n9958 vdd.n9957 0.0225448
R42229 vdd.n9957 vdd.n9956 0.0225448
R42230 vdd.n9938 vdd.n9914 0.0225448
R42231 vdd.n9939 vdd.n9938 0.0225448
R42232 vdd.n9936 vdd.n9935 0.0225448
R42233 vdd.n3842 vdd.n3840 0.0225448
R42234 vdd.n3842 vdd.n3841 0.0225448
R42235 vdd.n3853 vdd.n3852 0.0225448
R42236 vdd.n3852 vdd.n3851 0.0225448
R42237 vdd.n3867 vdd.n3866 0.0225448
R42238 vdd.n3868 vdd.n3867 0.0225448
R42239 vdd.n3864 vdd.n3863 0.0225448
R42240 vdd.n3860 vdd.n3859 0.0225448
R42241 vdd.n3861 vdd.n3860 0.0225448
R42242 vdd.n3870 vdd.n3869 0.0225448
R42243 vdd.n3869 vdd.n3868 0.0225448
R42244 vdd.n3850 vdd.n3826 0.0225448
R42245 vdd.n3851 vdd.n3850 0.0225448
R42246 vdd.n3848 vdd.n3847 0.0225448
R42247 vdd.n3890 vdd.n3888 0.0225448
R42248 vdd.n3890 vdd.n3889 0.0225448
R42249 vdd.n3901 vdd.n3900 0.0225448
R42250 vdd.n3900 vdd.n3899 0.0225448
R42251 vdd.n3915 vdd.n3914 0.0225448
R42252 vdd.n3916 vdd.n3915 0.0225448
R42253 vdd.n3912 vdd.n3911 0.0225448
R42254 vdd.n3908 vdd.n3907 0.0225448
R42255 vdd.n3909 vdd.n3908 0.0225448
R42256 vdd.n3918 vdd.n3917 0.0225448
R42257 vdd.n3917 vdd.n3916 0.0225448
R42258 vdd.n3898 vdd.n3874 0.0225448
R42259 vdd.n3899 vdd.n3898 0.0225448
R42260 vdd.n3896 vdd.n3895 0.0225448
R42261 vdd.n3992 vdd.n3990 0.0225448
R42262 vdd.n3992 vdd.n3991 0.0225448
R42263 vdd.n4003 vdd.n4002 0.0225448
R42264 vdd.n4002 vdd.n4001 0.0225448
R42265 vdd.n4017 vdd.n4016 0.0225448
R42266 vdd.n4018 vdd.n4017 0.0225448
R42267 vdd.n4014 vdd.n4013 0.0225448
R42268 vdd.n4010 vdd.n4009 0.0225448
R42269 vdd.n4011 vdd.n4010 0.0225448
R42270 vdd.n4020 vdd.n4019 0.0225448
R42271 vdd.n4019 vdd.n4018 0.0225448
R42272 vdd.n4000 vdd.n3976 0.0225448
R42273 vdd.n4001 vdd.n4000 0.0225448
R42274 vdd.n3998 vdd.n3997 0.0225448
R42275 vdd.n4040 vdd.n4038 0.0225448
R42276 vdd.n4040 vdd.n4039 0.0225448
R42277 vdd.n4051 vdd.n4050 0.0225448
R42278 vdd.n4050 vdd.n4049 0.0225448
R42279 vdd.n4065 vdd.n4064 0.0225448
R42280 vdd.n4066 vdd.n4065 0.0225448
R42281 vdd.n4062 vdd.n4061 0.0225448
R42282 vdd.n4058 vdd.n4057 0.0225448
R42283 vdd.n4059 vdd.n4058 0.0225448
R42284 vdd.n4068 vdd.n4067 0.0225448
R42285 vdd.n4067 vdd.n4066 0.0225448
R42286 vdd.n4048 vdd.n4024 0.0225448
R42287 vdd.n4049 vdd.n4048 0.0225448
R42288 vdd.n4046 vdd.n4045 0.0225448
R42289 vdd.n4088 vdd.n4086 0.0225448
R42290 vdd.n4088 vdd.n4087 0.0225448
R42291 vdd.n4099 vdd.n4098 0.0225448
R42292 vdd.n4098 vdd.n4097 0.0225448
R42293 vdd.n4113 vdd.n4112 0.0225448
R42294 vdd.n4114 vdd.n4113 0.0225448
R42295 vdd.n4110 vdd.n4109 0.0225448
R42296 vdd.n4106 vdd.n4105 0.0225448
R42297 vdd.n4107 vdd.n4106 0.0225448
R42298 vdd.n4116 vdd.n4115 0.0225448
R42299 vdd.n4115 vdd.n4114 0.0225448
R42300 vdd.n4096 vdd.n4072 0.0225448
R42301 vdd.n4097 vdd.n4096 0.0225448
R42302 vdd.n4094 vdd.n4093 0.0225448
R42303 vdd.n4136 vdd.n4134 0.0225448
R42304 vdd.n4136 vdd.n4135 0.0225448
R42305 vdd.n4147 vdd.n4146 0.0225448
R42306 vdd.n4146 vdd.n4145 0.0225448
R42307 vdd.n4161 vdd.n4160 0.0225448
R42308 vdd.n4162 vdd.n4161 0.0225448
R42309 vdd.n4158 vdd.n4157 0.0225448
R42310 vdd.n4154 vdd.n4153 0.0225448
R42311 vdd.n4155 vdd.n4154 0.0225448
R42312 vdd.n4164 vdd.n4163 0.0225448
R42313 vdd.n4163 vdd.n4162 0.0225448
R42314 vdd.n4144 vdd.n4120 0.0225448
R42315 vdd.n4145 vdd.n4144 0.0225448
R42316 vdd.n4142 vdd.n4141 0.0225448
R42317 vdd.n4238 vdd.n4236 0.0225448
R42318 vdd.n4238 vdd.n4237 0.0225448
R42319 vdd.n4249 vdd.n4248 0.0225448
R42320 vdd.n4248 vdd.n4247 0.0225448
R42321 vdd.n4263 vdd.n4262 0.0225448
R42322 vdd.n4264 vdd.n4263 0.0225448
R42323 vdd.n4260 vdd.n4259 0.0225448
R42324 vdd.n4256 vdd.n4255 0.0225448
R42325 vdd.n4257 vdd.n4256 0.0225448
R42326 vdd.n4266 vdd.n4265 0.0225448
R42327 vdd.n4265 vdd.n4264 0.0225448
R42328 vdd.n4246 vdd.n4222 0.0225448
R42329 vdd.n4247 vdd.n4246 0.0225448
R42330 vdd.n4244 vdd.n4243 0.0225448
R42331 vdd.n5758 vdd.n5756 0.0225448
R42332 vdd.n5758 vdd.n5757 0.0225448
R42333 vdd.n5769 vdd.n5768 0.0225448
R42334 vdd.n5768 vdd.n5767 0.0225448
R42335 vdd.n5783 vdd.n5782 0.0225448
R42336 vdd.n5784 vdd.n5783 0.0225448
R42337 vdd.n5780 vdd.n5779 0.0225448
R42338 vdd.n5776 vdd.n5775 0.0225448
R42339 vdd.n5777 vdd.n5776 0.0225448
R42340 vdd.n5786 vdd.n5785 0.0225448
R42341 vdd.n5785 vdd.n5784 0.0225448
R42342 vdd.n5766 vdd.n5742 0.0225448
R42343 vdd.n5767 vdd.n5766 0.0225448
R42344 vdd.n5764 vdd.n5763 0.0225448
R42345 vdd.n4289 vdd.n4288 0.0225448
R42346 vdd.n4297 vdd.n4296 0.0225448
R42347 vdd.n4296 vdd.n4295 0.0225448
R42348 vdd.n4311 vdd.n4310 0.0225448
R42349 vdd.n4312 vdd.n4311 0.0225448
R42350 vdd.n4308 vdd.n4307 0.0225448
R42351 vdd.n4307 vdd.n4306 0.0225448
R42352 vdd.n4304 vdd.n4303 0.0225448
R42353 vdd.n4314 vdd.n4313 0.0225448
R42354 vdd.n4313 vdd.n4312 0.0225448
R42355 vdd.n4294 vdd.n4270 0.0225448
R42356 vdd.n4295 vdd.n4294 0.0225448
R42357 vdd.n4292 vdd.n4286 0.0225448
R42358 vdd.n4292 vdd.n4291 0.0225448
R42359 vdd.n4337 vdd.n4336 0.0225448
R42360 vdd.n4345 vdd.n4344 0.0225448
R42361 vdd.n4344 vdd.n4343 0.0225448
R42362 vdd.n4359 vdd.n4358 0.0225448
R42363 vdd.n4360 vdd.n4359 0.0225448
R42364 vdd.n4356 vdd.n4355 0.0225448
R42365 vdd.n4355 vdd.n4354 0.0225448
R42366 vdd.n4352 vdd.n4351 0.0225448
R42367 vdd.n4362 vdd.n4361 0.0225448
R42368 vdd.n4361 vdd.n4360 0.0225448
R42369 vdd.n4342 vdd.n4318 0.0225448
R42370 vdd.n4343 vdd.n4342 0.0225448
R42371 vdd.n4340 vdd.n4334 0.0225448
R42372 vdd.n4340 vdd.n4339 0.0225448
R42373 vdd.n4438 vdd.n4437 0.0225448
R42374 vdd.n4446 vdd.n4445 0.0225448
R42375 vdd.n4445 vdd.n4444 0.0225448
R42376 vdd.n4460 vdd.n4459 0.0225448
R42377 vdd.n4461 vdd.n4460 0.0225448
R42378 vdd.n4457 vdd.n4456 0.0225448
R42379 vdd.n4456 vdd.n4455 0.0225448
R42380 vdd.n4453 vdd.n4452 0.0225448
R42381 vdd.n4463 vdd.n4462 0.0225448
R42382 vdd.n4462 vdd.n4461 0.0225448
R42383 vdd.n4443 vdd.n4419 0.0225448
R42384 vdd.n4444 vdd.n4443 0.0225448
R42385 vdd.n4441 vdd.n4435 0.0225448
R42386 vdd.n4441 vdd.n4440 0.0225448
R42387 vdd.n4486 vdd.n4485 0.0225448
R42388 vdd.n4494 vdd.n4493 0.0225448
R42389 vdd.n4493 vdd.n4492 0.0225448
R42390 vdd.n4508 vdd.n4507 0.0225448
R42391 vdd.n4509 vdd.n4508 0.0225448
R42392 vdd.n4505 vdd.n4504 0.0225448
R42393 vdd.n4504 vdd.n4503 0.0225448
R42394 vdd.n4501 vdd.n4500 0.0225448
R42395 vdd.n4511 vdd.n4510 0.0225448
R42396 vdd.n4510 vdd.n4509 0.0225448
R42397 vdd.n4491 vdd.n4467 0.0225448
R42398 vdd.n4492 vdd.n4491 0.0225448
R42399 vdd.n4489 vdd.n4483 0.0225448
R42400 vdd.n4489 vdd.n4488 0.0225448
R42401 vdd.n4534 vdd.n4533 0.0225448
R42402 vdd.n4542 vdd.n4541 0.0225448
R42403 vdd.n4541 vdd.n4540 0.0225448
R42404 vdd.n4556 vdd.n4555 0.0225448
R42405 vdd.n4557 vdd.n4556 0.0225448
R42406 vdd.n4553 vdd.n4552 0.0225448
R42407 vdd.n4552 vdd.n4551 0.0225448
R42408 vdd.n4549 vdd.n4548 0.0225448
R42409 vdd.n4559 vdd.n4558 0.0225448
R42410 vdd.n4558 vdd.n4557 0.0225448
R42411 vdd.n4539 vdd.n4515 0.0225448
R42412 vdd.n4540 vdd.n4539 0.0225448
R42413 vdd.n4537 vdd.n4531 0.0225448
R42414 vdd.n4537 vdd.n4536 0.0225448
R42415 vdd.n4582 vdd.n4581 0.0225448
R42416 vdd.n4590 vdd.n4589 0.0225448
R42417 vdd.n4589 vdd.n4588 0.0225448
R42418 vdd.n4604 vdd.n4603 0.0225448
R42419 vdd.n4605 vdd.n4604 0.0225448
R42420 vdd.n4601 vdd.n4600 0.0225448
R42421 vdd.n4600 vdd.n4599 0.0225448
R42422 vdd.n4597 vdd.n4596 0.0225448
R42423 vdd.n4607 vdd.n4606 0.0225448
R42424 vdd.n4606 vdd.n4605 0.0225448
R42425 vdd.n4587 vdd.n4563 0.0225448
R42426 vdd.n4588 vdd.n4587 0.0225448
R42427 vdd.n4585 vdd.n4579 0.0225448
R42428 vdd.n4585 vdd.n4584 0.0225448
R42429 vdd.n4683 vdd.n4682 0.0225448
R42430 vdd.n4691 vdd.n4690 0.0225448
R42431 vdd.n4690 vdd.n4689 0.0225448
R42432 vdd.n4705 vdd.n4704 0.0225448
R42433 vdd.n4706 vdd.n4705 0.0225448
R42434 vdd.n4702 vdd.n4701 0.0225448
R42435 vdd.n4701 vdd.n4700 0.0225448
R42436 vdd.n4698 vdd.n4697 0.0225448
R42437 vdd.n4708 vdd.n4707 0.0225448
R42438 vdd.n4707 vdd.n4706 0.0225448
R42439 vdd.n4688 vdd.n4664 0.0225448
R42440 vdd.n4689 vdd.n4688 0.0225448
R42441 vdd.n4686 vdd.n4680 0.0225448
R42442 vdd.n4686 vdd.n4685 0.0225448
R42443 vdd.n3796 vdd.n3795 0.0225448
R42444 vdd.n3804 vdd.n3803 0.0225448
R42445 vdd.n3803 vdd.n3802 0.0225448
R42446 vdd.n3818 vdd.n3817 0.0225448
R42447 vdd.n3819 vdd.n3818 0.0225448
R42448 vdd.n3815 vdd.n3814 0.0225448
R42449 vdd.n3814 vdd.n3813 0.0225448
R42450 vdd.n3811 vdd.n3810 0.0225448
R42451 vdd.n3821 vdd.n3820 0.0225448
R42452 vdd.n3820 vdd.n3819 0.0225448
R42453 vdd.n3801 vdd.n3777 0.0225448
R42454 vdd.n3802 vdd.n3801 0.0225448
R42455 vdd.n3799 vdd.n3793 0.0225448
R42456 vdd.n3799 vdd.n3798 0.0225448
R42457 vdd.n4731 vdd.n4730 0.0225448
R42458 vdd.n4739 vdd.n4738 0.0225448
R42459 vdd.n4738 vdd.n4737 0.0225448
R42460 vdd.n4753 vdd.n4752 0.0225448
R42461 vdd.n4754 vdd.n4753 0.0225448
R42462 vdd.n4750 vdd.n4749 0.0225448
R42463 vdd.n4749 vdd.n4748 0.0225448
R42464 vdd.n4746 vdd.n4745 0.0225448
R42465 vdd.n4756 vdd.n4755 0.0225448
R42466 vdd.n4755 vdd.n4754 0.0225448
R42467 vdd.n4736 vdd.n4712 0.0225448
R42468 vdd.n4737 vdd.n4736 0.0225448
R42469 vdd.n4734 vdd.n4728 0.0225448
R42470 vdd.n4734 vdd.n4733 0.0225448
R42471 vdd.n4778 vdd.n4777 0.0225448
R42472 vdd.n4786 vdd.n4785 0.0225448
R42473 vdd.n4785 vdd.n4784 0.0225448
R42474 vdd.n4800 vdd.n4799 0.0225448
R42475 vdd.n4801 vdd.n4800 0.0225448
R42476 vdd.n4797 vdd.n4796 0.0225448
R42477 vdd.n4796 vdd.n4795 0.0225448
R42478 vdd.n4793 vdd.n4792 0.0225448
R42479 vdd.n4803 vdd.n4802 0.0225448
R42480 vdd.n4802 vdd.n4801 0.0225448
R42481 vdd.n4783 vdd.n4759 0.0225448
R42482 vdd.n4784 vdd.n4783 0.0225448
R42483 vdd.n4781 vdd.n4775 0.0225448
R42484 vdd.n4781 vdd.n4780 0.0225448
R42485 vdd.n4828 vdd.n4827 0.0225448
R42486 vdd.n4836 vdd.n4835 0.0225448
R42487 vdd.n4835 vdd.n4834 0.0225448
R42488 vdd.n4850 vdd.n4849 0.0225448
R42489 vdd.n4851 vdd.n4850 0.0225448
R42490 vdd.n4847 vdd.n4846 0.0225448
R42491 vdd.n4846 vdd.n4845 0.0225448
R42492 vdd.n4843 vdd.n4842 0.0225448
R42493 vdd.n4853 vdd.n4852 0.0225448
R42494 vdd.n4852 vdd.n4851 0.0225448
R42495 vdd.n4833 vdd.n4809 0.0225448
R42496 vdd.n4834 vdd.n4833 0.0225448
R42497 vdd.n4831 vdd.n4825 0.0225448
R42498 vdd.n4831 vdd.n4830 0.0225448
R42499 vdd.n4878 vdd.n4877 0.0225448
R42500 vdd.n4886 vdd.n4885 0.0225448
R42501 vdd.n4885 vdd.n4884 0.0225448
R42502 vdd.n4900 vdd.n4899 0.0225448
R42503 vdd.n4901 vdd.n4900 0.0225448
R42504 vdd.n4897 vdd.n4896 0.0225448
R42505 vdd.n4896 vdd.n4895 0.0225448
R42506 vdd.n4893 vdd.n4892 0.0225448
R42507 vdd.n4903 vdd.n4902 0.0225448
R42508 vdd.n4902 vdd.n4901 0.0225448
R42509 vdd.n4883 vdd.n4859 0.0225448
R42510 vdd.n4884 vdd.n4883 0.0225448
R42511 vdd.n4881 vdd.n4875 0.0225448
R42512 vdd.n4881 vdd.n4880 0.0225448
R42513 vdd.n4926 vdd.n4925 0.0225448
R42514 vdd.n4934 vdd.n4933 0.0225448
R42515 vdd.n4933 vdd.n4932 0.0225448
R42516 vdd.n4948 vdd.n4947 0.0225448
R42517 vdd.n4949 vdd.n4948 0.0225448
R42518 vdd.n4945 vdd.n4944 0.0225448
R42519 vdd.n4944 vdd.n4943 0.0225448
R42520 vdd.n4941 vdd.n4940 0.0225448
R42521 vdd.n4951 vdd.n4950 0.0225448
R42522 vdd.n4950 vdd.n4949 0.0225448
R42523 vdd.n4931 vdd.n4907 0.0225448
R42524 vdd.n4932 vdd.n4931 0.0225448
R42525 vdd.n4929 vdd.n4923 0.0225448
R42526 vdd.n4929 vdd.n4928 0.0225448
R42527 vdd.n4654 vdd.n4653 0.0225448
R42528 vdd.n4651 vdd.n4650 0.0225448
R42529 vdd.n4650 vdd.n4649 0.0225448
R42530 vdd.n4640 vdd.n4639 0.0225448
R42531 vdd.n4641 vdd.n4640 0.0225448
R42532 vdd.n4637 vdd.n4636 0.0225448
R42533 vdd.n4636 vdd.n4635 0.0225448
R42534 vdd.n4633 vdd.n4632 0.0225448
R42535 vdd.n4642 vdd.n4624 0.0225448
R42536 vdd.n4642 vdd.n4641 0.0225448
R42537 vdd.n4648 vdd.n4647 0.0225448
R42538 vdd.n4649 vdd.n4648 0.0225448
R42539 vdd.n4658 vdd.n4657 0.0225448
R42540 vdd.n4657 vdd.n4656 0.0225448
R42541 vdd.n4977 vdd.n4976 0.0225448
R42542 vdd.n4985 vdd.n4984 0.0225448
R42543 vdd.n4984 vdd.n4983 0.0225448
R42544 vdd.n4999 vdd.n4998 0.0225448
R42545 vdd.n5000 vdd.n4999 0.0225448
R42546 vdd.n4996 vdd.n4995 0.0225448
R42547 vdd.n4995 vdd.n4994 0.0225448
R42548 vdd.n4992 vdd.n4991 0.0225448
R42549 vdd.n5002 vdd.n5001 0.0225448
R42550 vdd.n5001 vdd.n5000 0.0225448
R42551 vdd.n4982 vdd.n4958 0.0225448
R42552 vdd.n4983 vdd.n4982 0.0225448
R42553 vdd.n4980 vdd.n4974 0.0225448
R42554 vdd.n4980 vdd.n4979 0.0225448
R42555 vdd.n5024 vdd.n5023 0.0225448
R42556 vdd.n5032 vdd.n5031 0.0225448
R42557 vdd.n5031 vdd.n5030 0.0225448
R42558 vdd.n5046 vdd.n5045 0.0225448
R42559 vdd.n5047 vdd.n5046 0.0225448
R42560 vdd.n5043 vdd.n5042 0.0225448
R42561 vdd.n5042 vdd.n5041 0.0225448
R42562 vdd.n5039 vdd.n5038 0.0225448
R42563 vdd.n5049 vdd.n5048 0.0225448
R42564 vdd.n5048 vdd.n5047 0.0225448
R42565 vdd.n5029 vdd.n5005 0.0225448
R42566 vdd.n5030 vdd.n5029 0.0225448
R42567 vdd.n5027 vdd.n5021 0.0225448
R42568 vdd.n5027 vdd.n5026 0.0225448
R42569 vdd.n5072 vdd.n5071 0.0225448
R42570 vdd.n5080 vdd.n5079 0.0225448
R42571 vdd.n5079 vdd.n5078 0.0225448
R42572 vdd.n5094 vdd.n5093 0.0225448
R42573 vdd.n5095 vdd.n5094 0.0225448
R42574 vdd.n5091 vdd.n5090 0.0225448
R42575 vdd.n5090 vdd.n5089 0.0225448
R42576 vdd.n5087 vdd.n5086 0.0225448
R42577 vdd.n5097 vdd.n5096 0.0225448
R42578 vdd.n5096 vdd.n5095 0.0225448
R42579 vdd.n5077 vdd.n5053 0.0225448
R42580 vdd.n5078 vdd.n5077 0.0225448
R42581 vdd.n5075 vdd.n5069 0.0225448
R42582 vdd.n5075 vdd.n5074 0.0225448
R42583 vdd.n5123 vdd.n5122 0.0225448
R42584 vdd.n5131 vdd.n5130 0.0225448
R42585 vdd.n5130 vdd.n5129 0.0225448
R42586 vdd.n5145 vdd.n5144 0.0225448
R42587 vdd.n5146 vdd.n5145 0.0225448
R42588 vdd.n5142 vdd.n5141 0.0225448
R42589 vdd.n5141 vdd.n5140 0.0225448
R42590 vdd.n5138 vdd.n5137 0.0225448
R42591 vdd.n5148 vdd.n5147 0.0225448
R42592 vdd.n5147 vdd.n5146 0.0225448
R42593 vdd.n5128 vdd.n5104 0.0225448
R42594 vdd.n5129 vdd.n5128 0.0225448
R42595 vdd.n5126 vdd.n5120 0.0225448
R42596 vdd.n5126 vdd.n5125 0.0225448
R42597 vdd.n5173 vdd.n5172 0.0225448
R42598 vdd.n5181 vdd.n5180 0.0225448
R42599 vdd.n5180 vdd.n5179 0.0225448
R42600 vdd.n5195 vdd.n5194 0.0225448
R42601 vdd.n5196 vdd.n5195 0.0225448
R42602 vdd.n5192 vdd.n5191 0.0225448
R42603 vdd.n5191 vdd.n5190 0.0225448
R42604 vdd.n5188 vdd.n5187 0.0225448
R42605 vdd.n5198 vdd.n5197 0.0225448
R42606 vdd.n5197 vdd.n5196 0.0225448
R42607 vdd.n5178 vdd.n5154 0.0225448
R42608 vdd.n5179 vdd.n5178 0.0225448
R42609 vdd.n5176 vdd.n5170 0.0225448
R42610 vdd.n5176 vdd.n5175 0.0225448
R42611 vdd.n5221 vdd.n5220 0.0225448
R42612 vdd.n5229 vdd.n5228 0.0225448
R42613 vdd.n5228 vdd.n5227 0.0225448
R42614 vdd.n5243 vdd.n5242 0.0225448
R42615 vdd.n5244 vdd.n5243 0.0225448
R42616 vdd.n5240 vdd.n5239 0.0225448
R42617 vdd.n5239 vdd.n5238 0.0225448
R42618 vdd.n5236 vdd.n5235 0.0225448
R42619 vdd.n5246 vdd.n5245 0.0225448
R42620 vdd.n5245 vdd.n5244 0.0225448
R42621 vdd.n5226 vdd.n5202 0.0225448
R42622 vdd.n5227 vdd.n5226 0.0225448
R42623 vdd.n5224 vdd.n5218 0.0225448
R42624 vdd.n5224 vdd.n5223 0.0225448
R42625 vdd.n5271 vdd.n5270 0.0225448
R42626 vdd.n5279 vdd.n5278 0.0225448
R42627 vdd.n5278 vdd.n5277 0.0225448
R42628 vdd.n5293 vdd.n5292 0.0225448
R42629 vdd.n5294 vdd.n5293 0.0225448
R42630 vdd.n5290 vdd.n5289 0.0225448
R42631 vdd.n5289 vdd.n5288 0.0225448
R42632 vdd.n5286 vdd.n5285 0.0225448
R42633 vdd.n5296 vdd.n5295 0.0225448
R42634 vdd.n5295 vdd.n5294 0.0225448
R42635 vdd.n5276 vdd.n5252 0.0225448
R42636 vdd.n5277 vdd.n5276 0.0225448
R42637 vdd.n5274 vdd.n5268 0.0225448
R42638 vdd.n5274 vdd.n5273 0.0225448
R42639 vdd.n5318 vdd.n5317 0.0225448
R42640 vdd.n5326 vdd.n5325 0.0225448
R42641 vdd.n5325 vdd.n5324 0.0225448
R42642 vdd.n5340 vdd.n5339 0.0225448
R42643 vdd.n5341 vdd.n5340 0.0225448
R42644 vdd.n5337 vdd.n5336 0.0225448
R42645 vdd.n5336 vdd.n5335 0.0225448
R42646 vdd.n5333 vdd.n5332 0.0225448
R42647 vdd.n5343 vdd.n5342 0.0225448
R42648 vdd.n5342 vdd.n5341 0.0225448
R42649 vdd.n5323 vdd.n5299 0.0225448
R42650 vdd.n5324 vdd.n5323 0.0225448
R42651 vdd.n5321 vdd.n5315 0.0225448
R42652 vdd.n5321 vdd.n5320 0.0225448
R42653 vdd.n5368 vdd.n5367 0.0225448
R42654 vdd.n5376 vdd.n5375 0.0225448
R42655 vdd.n5375 vdd.n5374 0.0225448
R42656 vdd.n5390 vdd.n5389 0.0225448
R42657 vdd.n5391 vdd.n5390 0.0225448
R42658 vdd.n5387 vdd.n5386 0.0225448
R42659 vdd.n5386 vdd.n5385 0.0225448
R42660 vdd.n5383 vdd.n5382 0.0225448
R42661 vdd.n5393 vdd.n5392 0.0225448
R42662 vdd.n5392 vdd.n5391 0.0225448
R42663 vdd.n5373 vdd.n5349 0.0225448
R42664 vdd.n5374 vdd.n5373 0.0225448
R42665 vdd.n5371 vdd.n5365 0.0225448
R42666 vdd.n5371 vdd.n5370 0.0225448
R42667 vdd.n5418 vdd.n5417 0.0225448
R42668 vdd.n5426 vdd.n5425 0.0225448
R42669 vdd.n5425 vdd.n5424 0.0225448
R42670 vdd.n5440 vdd.n5439 0.0225448
R42671 vdd.n5441 vdd.n5440 0.0225448
R42672 vdd.n5437 vdd.n5436 0.0225448
R42673 vdd.n5436 vdd.n5435 0.0225448
R42674 vdd.n5433 vdd.n5432 0.0225448
R42675 vdd.n5443 vdd.n5442 0.0225448
R42676 vdd.n5442 vdd.n5441 0.0225448
R42677 vdd.n5423 vdd.n5399 0.0225448
R42678 vdd.n5424 vdd.n5423 0.0225448
R42679 vdd.n5421 vdd.n5415 0.0225448
R42680 vdd.n5421 vdd.n5420 0.0225448
R42681 vdd.n5466 vdd.n5465 0.0225448
R42682 vdd.n5474 vdd.n5473 0.0225448
R42683 vdd.n5473 vdd.n5472 0.0225448
R42684 vdd.n5488 vdd.n5487 0.0225448
R42685 vdd.n5489 vdd.n5488 0.0225448
R42686 vdd.n5485 vdd.n5484 0.0225448
R42687 vdd.n5484 vdd.n5483 0.0225448
R42688 vdd.n5481 vdd.n5480 0.0225448
R42689 vdd.n5491 vdd.n5490 0.0225448
R42690 vdd.n5490 vdd.n5489 0.0225448
R42691 vdd.n5471 vdd.n5447 0.0225448
R42692 vdd.n5472 vdd.n5471 0.0225448
R42693 vdd.n5469 vdd.n5463 0.0225448
R42694 vdd.n5469 vdd.n5468 0.0225448
R42695 vdd.n4409 vdd.n4408 0.0225448
R42696 vdd.n4406 vdd.n4405 0.0225448
R42697 vdd.n4405 vdd.n4404 0.0225448
R42698 vdd.n4395 vdd.n4394 0.0225448
R42699 vdd.n4396 vdd.n4395 0.0225448
R42700 vdd.n4392 vdd.n4391 0.0225448
R42701 vdd.n4391 vdd.n4390 0.0225448
R42702 vdd.n4388 vdd.n4387 0.0225448
R42703 vdd.n4397 vdd.n4379 0.0225448
R42704 vdd.n4397 vdd.n4396 0.0225448
R42705 vdd.n4403 vdd.n4402 0.0225448
R42706 vdd.n4404 vdd.n4403 0.0225448
R42707 vdd.n4413 vdd.n4412 0.0225448
R42708 vdd.n4412 vdd.n4411 0.0225448
R42709 vdd.n5517 vdd.n5516 0.0225448
R42710 vdd.n5525 vdd.n5524 0.0225448
R42711 vdd.n5524 vdd.n5523 0.0225448
R42712 vdd.n5539 vdd.n5538 0.0225448
R42713 vdd.n5540 vdd.n5539 0.0225448
R42714 vdd.n5536 vdd.n5535 0.0225448
R42715 vdd.n5535 vdd.n5534 0.0225448
R42716 vdd.n5532 vdd.n5531 0.0225448
R42717 vdd.n5542 vdd.n5541 0.0225448
R42718 vdd.n5541 vdd.n5540 0.0225448
R42719 vdd.n5522 vdd.n5498 0.0225448
R42720 vdd.n5523 vdd.n5522 0.0225448
R42721 vdd.n5520 vdd.n5514 0.0225448
R42722 vdd.n5520 vdd.n5519 0.0225448
R42723 vdd.n5564 vdd.n5563 0.0225448
R42724 vdd.n5572 vdd.n5571 0.0225448
R42725 vdd.n5571 vdd.n5570 0.0225448
R42726 vdd.n5586 vdd.n5585 0.0225448
R42727 vdd.n5587 vdd.n5586 0.0225448
R42728 vdd.n5583 vdd.n5582 0.0225448
R42729 vdd.n5582 vdd.n5581 0.0225448
R42730 vdd.n5579 vdd.n5578 0.0225448
R42731 vdd.n5589 vdd.n5588 0.0225448
R42732 vdd.n5588 vdd.n5587 0.0225448
R42733 vdd.n5569 vdd.n5545 0.0225448
R42734 vdd.n5570 vdd.n5569 0.0225448
R42735 vdd.n5567 vdd.n5561 0.0225448
R42736 vdd.n5567 vdd.n5566 0.0225448
R42737 vdd.n5614 vdd.n5613 0.0225448
R42738 vdd.n5622 vdd.n5621 0.0225448
R42739 vdd.n5621 vdd.n5620 0.0225448
R42740 vdd.n5636 vdd.n5635 0.0225448
R42741 vdd.n5637 vdd.n5636 0.0225448
R42742 vdd.n5633 vdd.n5632 0.0225448
R42743 vdd.n5632 vdd.n5631 0.0225448
R42744 vdd.n5629 vdd.n5628 0.0225448
R42745 vdd.n5639 vdd.n5638 0.0225448
R42746 vdd.n5638 vdd.n5637 0.0225448
R42747 vdd.n5619 vdd.n5595 0.0225448
R42748 vdd.n5620 vdd.n5619 0.0225448
R42749 vdd.n5617 vdd.n5611 0.0225448
R42750 vdd.n5617 vdd.n5616 0.0225448
R42751 vdd.n5664 vdd.n5663 0.0225448
R42752 vdd.n5672 vdd.n5671 0.0225448
R42753 vdd.n5671 vdd.n5670 0.0225448
R42754 vdd.n5686 vdd.n5685 0.0225448
R42755 vdd.n5687 vdd.n5686 0.0225448
R42756 vdd.n5683 vdd.n5682 0.0225448
R42757 vdd.n5682 vdd.n5681 0.0225448
R42758 vdd.n5679 vdd.n5678 0.0225448
R42759 vdd.n5689 vdd.n5688 0.0225448
R42760 vdd.n5688 vdd.n5687 0.0225448
R42761 vdd.n5669 vdd.n5645 0.0225448
R42762 vdd.n5670 vdd.n5669 0.0225448
R42763 vdd.n5667 vdd.n5661 0.0225448
R42764 vdd.n5667 vdd.n5666 0.0225448
R42765 vdd.n5712 vdd.n5711 0.0225448
R42766 vdd.n5720 vdd.n5719 0.0225448
R42767 vdd.n5719 vdd.n5718 0.0225448
R42768 vdd.n5734 vdd.n5733 0.0225448
R42769 vdd.n5735 vdd.n5734 0.0225448
R42770 vdd.n5731 vdd.n5730 0.0225448
R42771 vdd.n5730 vdd.n5729 0.0225448
R42772 vdd.n5727 vdd.n5726 0.0225448
R42773 vdd.n5737 vdd.n5736 0.0225448
R42774 vdd.n5736 vdd.n5735 0.0225448
R42775 vdd.n5717 vdd.n5693 0.0225448
R42776 vdd.n5718 vdd.n5717 0.0225448
R42777 vdd.n5715 vdd.n5709 0.0225448
R42778 vdd.n5715 vdd.n5714 0.0225448
R42779 vdd.n5855 vdd.n5853 0.0225448
R42780 vdd.n5855 vdd.n5854 0.0225448
R42781 vdd.n5866 vdd.n5865 0.0225448
R42782 vdd.n5865 vdd.n5864 0.0225448
R42783 vdd.n5880 vdd.n5879 0.0225448
R42784 vdd.n5881 vdd.n5880 0.0225448
R42785 vdd.n5877 vdd.n5876 0.0225448
R42786 vdd.n5873 vdd.n5872 0.0225448
R42787 vdd.n5874 vdd.n5873 0.0225448
R42788 vdd.n5883 vdd.n5882 0.0225448
R42789 vdd.n5882 vdd.n5881 0.0225448
R42790 vdd.n5863 vdd.n5839 0.0225448
R42791 vdd.n5864 vdd.n5863 0.0225448
R42792 vdd.n5861 vdd.n5860 0.0225448
R42793 vdd.n5807 vdd.n5805 0.0225448
R42794 vdd.n5807 vdd.n5806 0.0225448
R42795 vdd.n5818 vdd.n5817 0.0225448
R42796 vdd.n5817 vdd.n5816 0.0225448
R42797 vdd.n5832 vdd.n5831 0.0225448
R42798 vdd.n5833 vdd.n5832 0.0225448
R42799 vdd.n5829 vdd.n5828 0.0225448
R42800 vdd.n5825 vdd.n5824 0.0225448
R42801 vdd.n5826 vdd.n5825 0.0225448
R42802 vdd.n5835 vdd.n5834 0.0225448
R42803 vdd.n5834 vdd.n5833 0.0225448
R42804 vdd.n5815 vdd.n5791 0.0225448
R42805 vdd.n5816 vdd.n5815 0.0225448
R42806 vdd.n5813 vdd.n5812 0.0225448
R42807 vdd.n5904 vdd.n5902 0.0225448
R42808 vdd.n5904 vdd.n5903 0.0225448
R42809 vdd.n5915 vdd.n5914 0.0225448
R42810 vdd.n5914 vdd.n5913 0.0225448
R42811 vdd.n5929 vdd.n5928 0.0225448
R42812 vdd.n5930 vdd.n5929 0.0225448
R42813 vdd.n5926 vdd.n5925 0.0225448
R42814 vdd.n5922 vdd.n5921 0.0225448
R42815 vdd.n5923 vdd.n5922 0.0225448
R42816 vdd.n5932 vdd.n5931 0.0225448
R42817 vdd.n5931 vdd.n5930 0.0225448
R42818 vdd.n5912 vdd.n5888 0.0225448
R42819 vdd.n5913 vdd.n5912 0.0225448
R42820 vdd.n5910 vdd.n5909 0.0225448
R42821 vdd.n5954 vdd.n5952 0.0225448
R42822 vdd.n5954 vdd.n5953 0.0225448
R42823 vdd.n5965 vdd.n5964 0.0225448
R42824 vdd.n5964 vdd.n5963 0.0225448
R42825 vdd.n5979 vdd.n5978 0.0225448
R42826 vdd.n5980 vdd.n5979 0.0225448
R42827 vdd.n5976 vdd.n5975 0.0225448
R42828 vdd.n5972 vdd.n5971 0.0225448
R42829 vdd.n5973 vdd.n5972 0.0225448
R42830 vdd.n5982 vdd.n5981 0.0225448
R42831 vdd.n5981 vdd.n5980 0.0225448
R42832 vdd.n5962 vdd.n5938 0.0225448
R42833 vdd.n5963 vdd.n5962 0.0225448
R42834 vdd.n5960 vdd.n5959 0.0225448
R42835 vdd.n6002 vdd.n6000 0.0225448
R42836 vdd.n6002 vdd.n6001 0.0225448
R42837 vdd.n6013 vdd.n6012 0.0225448
R42838 vdd.n6012 vdd.n6011 0.0225448
R42839 vdd.n6027 vdd.n6026 0.0225448
R42840 vdd.n6028 vdd.n6027 0.0225448
R42841 vdd.n6024 vdd.n6023 0.0225448
R42842 vdd.n6020 vdd.n6019 0.0225448
R42843 vdd.n6021 vdd.n6020 0.0225448
R42844 vdd.n6030 vdd.n6029 0.0225448
R42845 vdd.n6029 vdd.n6028 0.0225448
R42846 vdd.n6010 vdd.n5986 0.0225448
R42847 vdd.n6011 vdd.n6010 0.0225448
R42848 vdd.n6008 vdd.n6007 0.0225448
R42849 vdd.n4189 vdd.n4188 0.0225448
R42850 vdd.n4190 vdd.n4189 0.0225448
R42851 vdd.n4186 vdd.n4179 0.0225448
R42852 vdd.n4197 vdd.n4179 0.0225448
R42853 vdd.n4199 vdd.n4198 0.0225448
R42854 vdd.n4200 vdd.n4199 0.0225448
R42855 vdd.n4214 vdd.n4213 0.0225448
R42856 vdd.n4210 vdd.n4169 0.0225448
R42857 vdd.n4211 vdd.n4210 0.0225448
R42858 vdd.n4205 vdd.n4174 0.0225448
R42859 vdd.n4200 vdd.n4174 0.0225448
R42860 vdd.n4196 vdd.n4195 0.0225448
R42861 vdd.n4197 vdd.n4196 0.0225448
R42862 vdd.n4193 vdd.n4192 0.0225448
R42863 vdd.n6150 vdd.n6148 0.0225448
R42864 vdd.n6150 vdd.n6149 0.0225448
R42865 vdd.n6161 vdd.n6160 0.0225448
R42866 vdd.n6160 vdd.n6159 0.0225448
R42867 vdd.n6175 vdd.n6174 0.0225448
R42868 vdd.n6176 vdd.n6175 0.0225448
R42869 vdd.n6172 vdd.n6171 0.0225448
R42870 vdd.n6168 vdd.n6167 0.0225448
R42871 vdd.n6169 vdd.n6168 0.0225448
R42872 vdd.n6178 vdd.n6177 0.0225448
R42873 vdd.n6177 vdd.n6176 0.0225448
R42874 vdd.n6158 vdd.n6134 0.0225448
R42875 vdd.n6159 vdd.n6158 0.0225448
R42876 vdd.n6156 vdd.n6155 0.0225448
R42877 vdd.n6101 vdd.n6099 0.0225448
R42878 vdd.n6101 vdd.n6100 0.0225448
R42879 vdd.n6112 vdd.n6111 0.0225448
R42880 vdd.n6111 vdd.n6110 0.0225448
R42881 vdd.n6126 vdd.n6125 0.0225448
R42882 vdd.n6127 vdd.n6126 0.0225448
R42883 vdd.n6123 vdd.n6122 0.0225448
R42884 vdd.n6119 vdd.n6118 0.0225448
R42885 vdd.n6120 vdd.n6119 0.0225448
R42886 vdd.n6129 vdd.n6128 0.0225448
R42887 vdd.n6128 vdd.n6127 0.0225448
R42888 vdd.n6109 vdd.n6085 0.0225448
R42889 vdd.n6110 vdd.n6109 0.0225448
R42890 vdd.n6107 vdd.n6106 0.0225448
R42891 vdd.n6053 vdd.n6051 0.0225448
R42892 vdd.n6053 vdd.n6052 0.0225448
R42893 vdd.n6064 vdd.n6063 0.0225448
R42894 vdd.n6063 vdd.n6062 0.0225448
R42895 vdd.n6078 vdd.n6077 0.0225448
R42896 vdd.n6079 vdd.n6078 0.0225448
R42897 vdd.n6075 vdd.n6074 0.0225448
R42898 vdd.n6071 vdd.n6070 0.0225448
R42899 vdd.n6072 vdd.n6071 0.0225448
R42900 vdd.n6081 vdd.n6080 0.0225448
R42901 vdd.n6080 vdd.n6079 0.0225448
R42902 vdd.n6061 vdd.n6037 0.0225448
R42903 vdd.n6062 vdd.n6061 0.0225448
R42904 vdd.n6059 vdd.n6058 0.0225448
R42905 vdd.n6199 vdd.n6197 0.0225448
R42906 vdd.n6199 vdd.n6198 0.0225448
R42907 vdd.n6210 vdd.n6209 0.0225448
R42908 vdd.n6209 vdd.n6208 0.0225448
R42909 vdd.n6224 vdd.n6223 0.0225448
R42910 vdd.n6225 vdd.n6224 0.0225448
R42911 vdd.n6221 vdd.n6220 0.0225448
R42912 vdd.n6217 vdd.n6216 0.0225448
R42913 vdd.n6218 vdd.n6217 0.0225448
R42914 vdd.n6227 vdd.n6226 0.0225448
R42915 vdd.n6226 vdd.n6225 0.0225448
R42916 vdd.n6207 vdd.n6183 0.0225448
R42917 vdd.n6208 vdd.n6207 0.0225448
R42918 vdd.n6205 vdd.n6204 0.0225448
R42919 vdd.n6249 vdd.n6247 0.0225448
R42920 vdd.n6249 vdd.n6248 0.0225448
R42921 vdd.n6260 vdd.n6259 0.0225448
R42922 vdd.n6259 vdd.n6258 0.0225448
R42923 vdd.n6274 vdd.n6273 0.0225448
R42924 vdd.n6275 vdd.n6274 0.0225448
R42925 vdd.n6271 vdd.n6270 0.0225448
R42926 vdd.n6267 vdd.n6266 0.0225448
R42927 vdd.n6268 vdd.n6267 0.0225448
R42928 vdd.n6277 vdd.n6276 0.0225448
R42929 vdd.n6276 vdd.n6275 0.0225448
R42930 vdd.n6257 vdd.n6233 0.0225448
R42931 vdd.n6258 vdd.n6257 0.0225448
R42932 vdd.n6255 vdd.n6254 0.0225448
R42933 vdd.n6297 vdd.n6295 0.0225448
R42934 vdd.n6297 vdd.n6296 0.0225448
R42935 vdd.n6308 vdd.n6307 0.0225448
R42936 vdd.n6307 vdd.n6306 0.0225448
R42937 vdd.n6322 vdd.n6321 0.0225448
R42938 vdd.n6323 vdd.n6322 0.0225448
R42939 vdd.n6319 vdd.n6318 0.0225448
R42940 vdd.n6315 vdd.n6314 0.0225448
R42941 vdd.n6316 vdd.n6315 0.0225448
R42942 vdd.n6325 vdd.n6324 0.0225448
R42943 vdd.n6324 vdd.n6323 0.0225448
R42944 vdd.n6305 vdd.n6281 0.0225448
R42945 vdd.n6306 vdd.n6305 0.0225448
R42946 vdd.n6303 vdd.n6302 0.0225448
R42947 vdd.n6395 vdd.n6393 0.0225448
R42948 vdd.n6395 vdd.n6394 0.0225448
R42949 vdd.n6406 vdd.n6405 0.0225448
R42950 vdd.n6405 vdd.n6404 0.0225448
R42951 vdd.n6420 vdd.n6419 0.0225448
R42952 vdd.n6421 vdd.n6420 0.0225448
R42953 vdd.n6417 vdd.n6416 0.0225448
R42954 vdd.n6413 vdd.n6412 0.0225448
R42955 vdd.n6414 vdd.n6413 0.0225448
R42956 vdd.n6423 vdd.n6422 0.0225448
R42957 vdd.n6422 vdd.n6421 0.0225448
R42958 vdd.n6403 vdd.n6379 0.0225448
R42959 vdd.n6404 vdd.n6403 0.0225448
R42960 vdd.n6401 vdd.n6400 0.0225448
R42961 vdd.n6347 vdd.n6345 0.0225448
R42962 vdd.n6347 vdd.n6346 0.0225448
R42963 vdd.n6358 vdd.n6357 0.0225448
R42964 vdd.n6357 vdd.n6356 0.0225448
R42965 vdd.n6372 vdd.n6371 0.0225448
R42966 vdd.n6373 vdd.n6372 0.0225448
R42967 vdd.n6369 vdd.n6368 0.0225448
R42968 vdd.n6365 vdd.n6364 0.0225448
R42969 vdd.n6366 vdd.n6365 0.0225448
R42970 vdd.n6375 vdd.n6374 0.0225448
R42971 vdd.n6374 vdd.n6373 0.0225448
R42972 vdd.n6355 vdd.n6331 0.0225448
R42973 vdd.n6356 vdd.n6355 0.0225448
R42974 vdd.n6353 vdd.n6352 0.0225448
R42975 vdd.n6444 vdd.n6442 0.0225448
R42976 vdd.n6444 vdd.n6443 0.0225448
R42977 vdd.n6455 vdd.n6454 0.0225448
R42978 vdd.n6454 vdd.n6453 0.0225448
R42979 vdd.n6469 vdd.n6468 0.0225448
R42980 vdd.n6470 vdd.n6469 0.0225448
R42981 vdd.n6466 vdd.n6465 0.0225448
R42982 vdd.n6462 vdd.n6461 0.0225448
R42983 vdd.n6463 vdd.n6462 0.0225448
R42984 vdd.n6472 vdd.n6471 0.0225448
R42985 vdd.n6471 vdd.n6470 0.0225448
R42986 vdd.n6452 vdd.n6428 0.0225448
R42987 vdd.n6453 vdd.n6452 0.0225448
R42988 vdd.n6450 vdd.n6449 0.0225448
R42989 vdd.n6494 vdd.n6492 0.0225448
R42990 vdd.n6494 vdd.n6493 0.0225448
R42991 vdd.n6505 vdd.n6504 0.0225448
R42992 vdd.n6504 vdd.n6503 0.0225448
R42993 vdd.n6519 vdd.n6518 0.0225448
R42994 vdd.n6520 vdd.n6519 0.0225448
R42995 vdd.n6516 vdd.n6515 0.0225448
R42996 vdd.n6512 vdd.n6511 0.0225448
R42997 vdd.n6513 vdd.n6512 0.0225448
R42998 vdd.n6522 vdd.n6521 0.0225448
R42999 vdd.n6521 vdd.n6520 0.0225448
R43000 vdd.n6502 vdd.n6478 0.0225448
R43001 vdd.n6503 vdd.n6502 0.0225448
R43002 vdd.n6500 vdd.n6499 0.0225448
R43003 vdd.n6542 vdd.n6540 0.0225448
R43004 vdd.n6542 vdd.n6541 0.0225448
R43005 vdd.n6553 vdd.n6552 0.0225448
R43006 vdd.n6552 vdd.n6551 0.0225448
R43007 vdd.n6567 vdd.n6566 0.0225448
R43008 vdd.n6568 vdd.n6567 0.0225448
R43009 vdd.n6564 vdd.n6563 0.0225448
R43010 vdd.n6560 vdd.n6559 0.0225448
R43011 vdd.n6561 vdd.n6560 0.0225448
R43012 vdd.n6570 vdd.n6569 0.0225448
R43013 vdd.n6569 vdd.n6568 0.0225448
R43014 vdd.n6550 vdd.n6526 0.0225448
R43015 vdd.n6551 vdd.n6550 0.0225448
R43016 vdd.n6548 vdd.n6547 0.0225448
R43017 vdd.n3943 vdd.n3942 0.0225448
R43018 vdd.n3944 vdd.n3943 0.0225448
R43019 vdd.n3940 vdd.n3933 0.0225448
R43020 vdd.n3951 vdd.n3933 0.0225448
R43021 vdd.n3953 vdd.n3952 0.0225448
R43022 vdd.n3954 vdd.n3953 0.0225448
R43023 vdd.n3968 vdd.n3967 0.0225448
R43024 vdd.n3964 vdd.n3923 0.0225448
R43025 vdd.n3965 vdd.n3964 0.0225448
R43026 vdd.n3959 vdd.n3928 0.0225448
R43027 vdd.n3954 vdd.n3928 0.0225448
R43028 vdd.n3950 vdd.n3949 0.0225448
R43029 vdd.n3951 vdd.n3950 0.0225448
R43030 vdd.n3947 vdd.n3946 0.0225448
R43031 vdd.n6641 vdd.n6639 0.0225448
R43032 vdd.n6641 vdd.n6640 0.0225448
R43033 vdd.n6652 vdd.n6651 0.0225448
R43034 vdd.n6651 vdd.n6650 0.0225448
R43035 vdd.n6666 vdd.n6665 0.0225448
R43036 vdd.n6667 vdd.n6666 0.0225448
R43037 vdd.n6663 vdd.n6662 0.0225448
R43038 vdd.n6659 vdd.n6658 0.0225448
R43039 vdd.n6660 vdd.n6659 0.0225448
R43040 vdd.n6669 vdd.n6668 0.0225448
R43041 vdd.n6668 vdd.n6667 0.0225448
R43042 vdd.n6649 vdd.n6625 0.0225448
R43043 vdd.n6650 vdd.n6649 0.0225448
R43044 vdd.n6647 vdd.n6646 0.0225448
R43045 vdd.n6593 vdd.n6591 0.0225448
R43046 vdd.n6593 vdd.n6592 0.0225448
R43047 vdd.n6604 vdd.n6603 0.0225448
R43048 vdd.n6603 vdd.n6602 0.0225448
R43049 vdd.n6618 vdd.n6617 0.0225448
R43050 vdd.n6619 vdd.n6618 0.0225448
R43051 vdd.n6615 vdd.n6614 0.0225448
R43052 vdd.n6611 vdd.n6610 0.0225448
R43053 vdd.n6612 vdd.n6611 0.0225448
R43054 vdd.n6621 vdd.n6620 0.0225448
R43055 vdd.n6620 vdd.n6619 0.0225448
R43056 vdd.n6601 vdd.n6577 0.0225448
R43057 vdd.n6602 vdd.n6601 0.0225448
R43058 vdd.n6599 vdd.n6598 0.0225448
R43059 vdd.n6690 vdd.n6688 0.0225448
R43060 vdd.n6690 vdd.n6689 0.0225448
R43061 vdd.n6701 vdd.n6700 0.0225448
R43062 vdd.n6700 vdd.n6699 0.0225448
R43063 vdd.n6715 vdd.n6714 0.0225448
R43064 vdd.n6716 vdd.n6715 0.0225448
R43065 vdd.n6712 vdd.n6711 0.0225448
R43066 vdd.n6708 vdd.n6707 0.0225448
R43067 vdd.n6709 vdd.n6708 0.0225448
R43068 vdd.n6718 vdd.n6717 0.0225448
R43069 vdd.n6717 vdd.n6716 0.0225448
R43070 vdd.n6698 vdd.n6674 0.0225448
R43071 vdd.n6699 vdd.n6698 0.0225448
R43072 vdd.n6696 vdd.n6695 0.0225448
R43073 vdd.n6740 vdd.n6738 0.0225448
R43074 vdd.n6740 vdd.n6739 0.0225448
R43075 vdd.n6751 vdd.n6750 0.0225448
R43076 vdd.n6750 vdd.n6749 0.0225448
R43077 vdd.n6765 vdd.n6764 0.0225448
R43078 vdd.n6766 vdd.n6765 0.0225448
R43079 vdd.n6762 vdd.n6761 0.0225448
R43080 vdd.n6758 vdd.n6757 0.0225448
R43081 vdd.n6759 vdd.n6758 0.0225448
R43082 vdd.n6768 vdd.n6767 0.0225448
R43083 vdd.n6767 vdd.n6766 0.0225448
R43084 vdd.n6748 vdd.n6724 0.0225448
R43085 vdd.n6749 vdd.n6748 0.0225448
R43086 vdd.n6746 vdd.n6745 0.0225448
R43087 vdd.n6788 vdd.n6786 0.0225448
R43088 vdd.n6788 vdd.n6787 0.0225448
R43089 vdd.n6799 vdd.n6798 0.0225448
R43090 vdd.n6798 vdd.n6797 0.0225448
R43091 vdd.n6813 vdd.n6812 0.0225448
R43092 vdd.n6814 vdd.n6813 0.0225448
R43093 vdd.n6810 vdd.n6809 0.0225448
R43094 vdd.n6806 vdd.n6805 0.0225448
R43095 vdd.n6807 vdd.n6806 0.0225448
R43096 vdd.n6816 vdd.n6815 0.0225448
R43097 vdd.n6815 vdd.n6814 0.0225448
R43098 vdd.n6796 vdd.n6772 0.0225448
R43099 vdd.n6797 vdd.n6796 0.0225448
R43100 vdd.n6794 vdd.n6793 0.0225448
R43101 vdd.n700 vdd.n698 0.0225448
R43102 vdd.n700 vdd.n699 0.0225448
R43103 vdd.n711 vdd.n710 0.0225448
R43104 vdd.n710 vdd.n709 0.0225448
R43105 vdd.n725 vdd.n724 0.0225448
R43106 vdd.n726 vdd.n725 0.0225448
R43107 vdd.n722 vdd.n721 0.0225448
R43108 vdd.n718 vdd.n717 0.0225448
R43109 vdd.n719 vdd.n718 0.0225448
R43110 vdd.n728 vdd.n727 0.0225448
R43111 vdd.n727 vdd.n726 0.0225448
R43112 vdd.n708 vdd.n684 0.0225448
R43113 vdd.n709 vdd.n708 0.0225448
R43114 vdd.n706 vdd.n705 0.0225448
R43115 vdd.n748 vdd.n746 0.0225448
R43116 vdd.n748 vdd.n747 0.0225448
R43117 vdd.n759 vdd.n758 0.0225448
R43118 vdd.n758 vdd.n757 0.0225448
R43119 vdd.n773 vdd.n772 0.0225448
R43120 vdd.n774 vdd.n773 0.0225448
R43121 vdd.n770 vdd.n769 0.0225448
R43122 vdd.n766 vdd.n765 0.0225448
R43123 vdd.n767 vdd.n766 0.0225448
R43124 vdd.n776 vdd.n775 0.0225448
R43125 vdd.n775 vdd.n774 0.0225448
R43126 vdd.n756 vdd.n732 0.0225448
R43127 vdd.n757 vdd.n756 0.0225448
R43128 vdd.n754 vdd.n753 0.0225448
R43129 vdd.n850 vdd.n848 0.0225448
R43130 vdd.n850 vdd.n849 0.0225448
R43131 vdd.n861 vdd.n860 0.0225448
R43132 vdd.n860 vdd.n859 0.0225448
R43133 vdd.n875 vdd.n874 0.0225448
R43134 vdd.n876 vdd.n875 0.0225448
R43135 vdd.n872 vdd.n871 0.0225448
R43136 vdd.n868 vdd.n867 0.0225448
R43137 vdd.n869 vdd.n868 0.0225448
R43138 vdd.n878 vdd.n877 0.0225448
R43139 vdd.n877 vdd.n876 0.0225448
R43140 vdd.n858 vdd.n834 0.0225448
R43141 vdd.n859 vdd.n858 0.0225448
R43142 vdd.n856 vdd.n855 0.0225448
R43143 vdd.n898 vdd.n896 0.0225448
R43144 vdd.n898 vdd.n897 0.0225448
R43145 vdd.n909 vdd.n908 0.0225448
R43146 vdd.n908 vdd.n907 0.0225448
R43147 vdd.n923 vdd.n922 0.0225448
R43148 vdd.n924 vdd.n923 0.0225448
R43149 vdd.n920 vdd.n919 0.0225448
R43150 vdd.n916 vdd.n915 0.0225448
R43151 vdd.n917 vdd.n916 0.0225448
R43152 vdd.n926 vdd.n925 0.0225448
R43153 vdd.n925 vdd.n924 0.0225448
R43154 vdd.n906 vdd.n882 0.0225448
R43155 vdd.n907 vdd.n906 0.0225448
R43156 vdd.n904 vdd.n903 0.0225448
R43157 vdd.n946 vdd.n944 0.0225448
R43158 vdd.n946 vdd.n945 0.0225448
R43159 vdd.n957 vdd.n956 0.0225448
R43160 vdd.n956 vdd.n955 0.0225448
R43161 vdd.n971 vdd.n970 0.0225448
R43162 vdd.n972 vdd.n971 0.0225448
R43163 vdd.n968 vdd.n967 0.0225448
R43164 vdd.n964 vdd.n963 0.0225448
R43165 vdd.n965 vdd.n964 0.0225448
R43166 vdd.n974 vdd.n973 0.0225448
R43167 vdd.n973 vdd.n972 0.0225448
R43168 vdd.n954 vdd.n930 0.0225448
R43169 vdd.n955 vdd.n954 0.0225448
R43170 vdd.n952 vdd.n951 0.0225448
R43171 vdd.n994 vdd.n992 0.0225448
R43172 vdd.n994 vdd.n993 0.0225448
R43173 vdd.n1005 vdd.n1004 0.0225448
R43174 vdd.n1004 vdd.n1003 0.0225448
R43175 vdd.n1019 vdd.n1018 0.0225448
R43176 vdd.n1020 vdd.n1019 0.0225448
R43177 vdd.n1016 vdd.n1015 0.0225448
R43178 vdd.n1012 vdd.n1011 0.0225448
R43179 vdd.n1013 vdd.n1012 0.0225448
R43180 vdd.n1022 vdd.n1021 0.0225448
R43181 vdd.n1021 vdd.n1020 0.0225448
R43182 vdd.n1002 vdd.n978 0.0225448
R43183 vdd.n1003 vdd.n1002 0.0225448
R43184 vdd.n1000 vdd.n999 0.0225448
R43185 vdd.n1096 vdd.n1094 0.0225448
R43186 vdd.n1096 vdd.n1095 0.0225448
R43187 vdd.n1107 vdd.n1106 0.0225448
R43188 vdd.n1106 vdd.n1105 0.0225448
R43189 vdd.n1121 vdd.n1120 0.0225448
R43190 vdd.n1122 vdd.n1121 0.0225448
R43191 vdd.n1118 vdd.n1117 0.0225448
R43192 vdd.n1114 vdd.n1113 0.0225448
R43193 vdd.n1115 vdd.n1114 0.0225448
R43194 vdd.n1124 vdd.n1123 0.0225448
R43195 vdd.n1123 vdd.n1122 0.0225448
R43196 vdd.n1104 vdd.n1080 0.0225448
R43197 vdd.n1105 vdd.n1104 0.0225448
R43198 vdd.n1102 vdd.n1101 0.0225448
R43199 vdd.n2616 vdd.n2614 0.0225448
R43200 vdd.n2616 vdd.n2615 0.0225448
R43201 vdd.n2627 vdd.n2626 0.0225448
R43202 vdd.n2626 vdd.n2625 0.0225448
R43203 vdd.n2641 vdd.n2640 0.0225448
R43204 vdd.n2642 vdd.n2641 0.0225448
R43205 vdd.n2638 vdd.n2637 0.0225448
R43206 vdd.n2634 vdd.n2633 0.0225448
R43207 vdd.n2635 vdd.n2634 0.0225448
R43208 vdd.n2644 vdd.n2643 0.0225448
R43209 vdd.n2643 vdd.n2642 0.0225448
R43210 vdd.n2624 vdd.n2600 0.0225448
R43211 vdd.n2625 vdd.n2624 0.0225448
R43212 vdd.n2622 vdd.n2621 0.0225448
R43213 vdd.n1147 vdd.n1146 0.0225448
R43214 vdd.n1155 vdd.n1154 0.0225448
R43215 vdd.n1154 vdd.n1153 0.0225448
R43216 vdd.n1169 vdd.n1168 0.0225448
R43217 vdd.n1170 vdd.n1169 0.0225448
R43218 vdd.n1166 vdd.n1165 0.0225448
R43219 vdd.n1165 vdd.n1164 0.0225448
R43220 vdd.n1162 vdd.n1161 0.0225448
R43221 vdd.n1172 vdd.n1171 0.0225448
R43222 vdd.n1171 vdd.n1170 0.0225448
R43223 vdd.n1152 vdd.n1128 0.0225448
R43224 vdd.n1153 vdd.n1152 0.0225448
R43225 vdd.n1150 vdd.n1144 0.0225448
R43226 vdd.n1150 vdd.n1149 0.0225448
R43227 vdd.n1195 vdd.n1194 0.0225448
R43228 vdd.n1203 vdd.n1202 0.0225448
R43229 vdd.n1202 vdd.n1201 0.0225448
R43230 vdd.n1217 vdd.n1216 0.0225448
R43231 vdd.n1218 vdd.n1217 0.0225448
R43232 vdd.n1214 vdd.n1213 0.0225448
R43233 vdd.n1213 vdd.n1212 0.0225448
R43234 vdd.n1210 vdd.n1209 0.0225448
R43235 vdd.n1220 vdd.n1219 0.0225448
R43236 vdd.n1219 vdd.n1218 0.0225448
R43237 vdd.n1200 vdd.n1176 0.0225448
R43238 vdd.n1201 vdd.n1200 0.0225448
R43239 vdd.n1198 vdd.n1192 0.0225448
R43240 vdd.n1198 vdd.n1197 0.0225448
R43241 vdd.n1296 vdd.n1295 0.0225448
R43242 vdd.n1304 vdd.n1303 0.0225448
R43243 vdd.n1303 vdd.n1302 0.0225448
R43244 vdd.n1318 vdd.n1317 0.0225448
R43245 vdd.n1319 vdd.n1318 0.0225448
R43246 vdd.n1315 vdd.n1314 0.0225448
R43247 vdd.n1314 vdd.n1313 0.0225448
R43248 vdd.n1311 vdd.n1310 0.0225448
R43249 vdd.n1321 vdd.n1320 0.0225448
R43250 vdd.n1320 vdd.n1319 0.0225448
R43251 vdd.n1301 vdd.n1277 0.0225448
R43252 vdd.n1302 vdd.n1301 0.0225448
R43253 vdd.n1299 vdd.n1293 0.0225448
R43254 vdd.n1299 vdd.n1298 0.0225448
R43255 vdd.n1344 vdd.n1343 0.0225448
R43256 vdd.n1352 vdd.n1351 0.0225448
R43257 vdd.n1351 vdd.n1350 0.0225448
R43258 vdd.n1366 vdd.n1365 0.0225448
R43259 vdd.n1367 vdd.n1366 0.0225448
R43260 vdd.n1363 vdd.n1362 0.0225448
R43261 vdd.n1362 vdd.n1361 0.0225448
R43262 vdd.n1359 vdd.n1358 0.0225448
R43263 vdd.n1369 vdd.n1368 0.0225448
R43264 vdd.n1368 vdd.n1367 0.0225448
R43265 vdd.n1349 vdd.n1325 0.0225448
R43266 vdd.n1350 vdd.n1349 0.0225448
R43267 vdd.n1347 vdd.n1341 0.0225448
R43268 vdd.n1347 vdd.n1346 0.0225448
R43269 vdd.n1392 vdd.n1391 0.0225448
R43270 vdd.n1400 vdd.n1399 0.0225448
R43271 vdd.n1399 vdd.n1398 0.0225448
R43272 vdd.n1414 vdd.n1413 0.0225448
R43273 vdd.n1415 vdd.n1414 0.0225448
R43274 vdd.n1411 vdd.n1410 0.0225448
R43275 vdd.n1410 vdd.n1409 0.0225448
R43276 vdd.n1407 vdd.n1406 0.0225448
R43277 vdd.n1417 vdd.n1416 0.0225448
R43278 vdd.n1416 vdd.n1415 0.0225448
R43279 vdd.n1397 vdd.n1373 0.0225448
R43280 vdd.n1398 vdd.n1397 0.0225448
R43281 vdd.n1395 vdd.n1389 0.0225448
R43282 vdd.n1395 vdd.n1394 0.0225448
R43283 vdd.n1440 vdd.n1439 0.0225448
R43284 vdd.n1448 vdd.n1447 0.0225448
R43285 vdd.n1447 vdd.n1446 0.0225448
R43286 vdd.n1462 vdd.n1461 0.0225448
R43287 vdd.n1463 vdd.n1462 0.0225448
R43288 vdd.n1459 vdd.n1458 0.0225448
R43289 vdd.n1458 vdd.n1457 0.0225448
R43290 vdd.n1455 vdd.n1454 0.0225448
R43291 vdd.n1465 vdd.n1464 0.0225448
R43292 vdd.n1464 vdd.n1463 0.0225448
R43293 vdd.n1445 vdd.n1421 0.0225448
R43294 vdd.n1446 vdd.n1445 0.0225448
R43295 vdd.n1443 vdd.n1437 0.0225448
R43296 vdd.n1443 vdd.n1442 0.0225448
R43297 vdd.n1541 vdd.n1540 0.0225448
R43298 vdd.n1549 vdd.n1548 0.0225448
R43299 vdd.n1548 vdd.n1547 0.0225448
R43300 vdd.n1563 vdd.n1562 0.0225448
R43301 vdd.n1564 vdd.n1563 0.0225448
R43302 vdd.n1560 vdd.n1559 0.0225448
R43303 vdd.n1559 vdd.n1558 0.0225448
R43304 vdd.n1556 vdd.n1555 0.0225448
R43305 vdd.n1566 vdd.n1565 0.0225448
R43306 vdd.n1565 vdd.n1564 0.0225448
R43307 vdd.n1546 vdd.n1522 0.0225448
R43308 vdd.n1547 vdd.n1546 0.0225448
R43309 vdd.n1544 vdd.n1538 0.0225448
R43310 vdd.n1544 vdd.n1543 0.0225448
R43311 vdd.n654 vdd.n653 0.0225448
R43312 vdd.n662 vdd.n661 0.0225448
R43313 vdd.n661 vdd.n660 0.0225448
R43314 vdd.n676 vdd.n675 0.0225448
R43315 vdd.n677 vdd.n676 0.0225448
R43316 vdd.n673 vdd.n672 0.0225448
R43317 vdd.n672 vdd.n671 0.0225448
R43318 vdd.n669 vdd.n668 0.0225448
R43319 vdd.n679 vdd.n678 0.0225448
R43320 vdd.n678 vdd.n677 0.0225448
R43321 vdd.n659 vdd.n635 0.0225448
R43322 vdd.n660 vdd.n659 0.0225448
R43323 vdd.n657 vdd.n651 0.0225448
R43324 vdd.n657 vdd.n656 0.0225448
R43325 vdd.n1589 vdd.n1588 0.0225448
R43326 vdd.n1597 vdd.n1596 0.0225448
R43327 vdd.n1596 vdd.n1595 0.0225448
R43328 vdd.n1611 vdd.n1610 0.0225448
R43329 vdd.n1612 vdd.n1611 0.0225448
R43330 vdd.n1608 vdd.n1607 0.0225448
R43331 vdd.n1607 vdd.n1606 0.0225448
R43332 vdd.n1604 vdd.n1603 0.0225448
R43333 vdd.n1614 vdd.n1613 0.0225448
R43334 vdd.n1613 vdd.n1612 0.0225448
R43335 vdd.n1594 vdd.n1570 0.0225448
R43336 vdd.n1595 vdd.n1594 0.0225448
R43337 vdd.n1592 vdd.n1586 0.0225448
R43338 vdd.n1592 vdd.n1591 0.0225448
R43339 vdd.n1636 vdd.n1635 0.0225448
R43340 vdd.n1644 vdd.n1643 0.0225448
R43341 vdd.n1643 vdd.n1642 0.0225448
R43342 vdd.n1658 vdd.n1657 0.0225448
R43343 vdd.n1659 vdd.n1658 0.0225448
R43344 vdd.n1655 vdd.n1654 0.0225448
R43345 vdd.n1654 vdd.n1653 0.0225448
R43346 vdd.n1651 vdd.n1650 0.0225448
R43347 vdd.n1661 vdd.n1660 0.0225448
R43348 vdd.n1660 vdd.n1659 0.0225448
R43349 vdd.n1641 vdd.n1617 0.0225448
R43350 vdd.n1642 vdd.n1641 0.0225448
R43351 vdd.n1639 vdd.n1633 0.0225448
R43352 vdd.n1639 vdd.n1638 0.0225448
R43353 vdd.n1686 vdd.n1685 0.0225448
R43354 vdd.n1694 vdd.n1693 0.0225448
R43355 vdd.n1693 vdd.n1692 0.0225448
R43356 vdd.n1708 vdd.n1707 0.0225448
R43357 vdd.n1709 vdd.n1708 0.0225448
R43358 vdd.n1705 vdd.n1704 0.0225448
R43359 vdd.n1704 vdd.n1703 0.0225448
R43360 vdd.n1701 vdd.n1700 0.0225448
R43361 vdd.n1711 vdd.n1710 0.0225448
R43362 vdd.n1710 vdd.n1709 0.0225448
R43363 vdd.n1691 vdd.n1667 0.0225448
R43364 vdd.n1692 vdd.n1691 0.0225448
R43365 vdd.n1689 vdd.n1683 0.0225448
R43366 vdd.n1689 vdd.n1688 0.0225448
R43367 vdd.n1736 vdd.n1735 0.0225448
R43368 vdd.n1744 vdd.n1743 0.0225448
R43369 vdd.n1743 vdd.n1742 0.0225448
R43370 vdd.n1758 vdd.n1757 0.0225448
R43371 vdd.n1759 vdd.n1758 0.0225448
R43372 vdd.n1755 vdd.n1754 0.0225448
R43373 vdd.n1754 vdd.n1753 0.0225448
R43374 vdd.n1751 vdd.n1750 0.0225448
R43375 vdd.n1761 vdd.n1760 0.0225448
R43376 vdd.n1760 vdd.n1759 0.0225448
R43377 vdd.n1741 vdd.n1717 0.0225448
R43378 vdd.n1742 vdd.n1741 0.0225448
R43379 vdd.n1739 vdd.n1733 0.0225448
R43380 vdd.n1739 vdd.n1738 0.0225448
R43381 vdd.n1784 vdd.n1783 0.0225448
R43382 vdd.n1792 vdd.n1791 0.0225448
R43383 vdd.n1791 vdd.n1790 0.0225448
R43384 vdd.n1806 vdd.n1805 0.0225448
R43385 vdd.n1807 vdd.n1806 0.0225448
R43386 vdd.n1803 vdd.n1802 0.0225448
R43387 vdd.n1802 vdd.n1801 0.0225448
R43388 vdd.n1799 vdd.n1798 0.0225448
R43389 vdd.n1809 vdd.n1808 0.0225448
R43390 vdd.n1808 vdd.n1807 0.0225448
R43391 vdd.n1789 vdd.n1765 0.0225448
R43392 vdd.n1790 vdd.n1789 0.0225448
R43393 vdd.n1787 vdd.n1781 0.0225448
R43394 vdd.n1787 vdd.n1786 0.0225448
R43395 vdd.n1512 vdd.n1511 0.0225448
R43396 vdd.n1509 vdd.n1508 0.0225448
R43397 vdd.n1508 vdd.n1507 0.0225448
R43398 vdd.n1498 vdd.n1497 0.0225448
R43399 vdd.n1499 vdd.n1498 0.0225448
R43400 vdd.n1495 vdd.n1494 0.0225448
R43401 vdd.n1494 vdd.n1493 0.0225448
R43402 vdd.n1491 vdd.n1490 0.0225448
R43403 vdd.n1500 vdd.n1482 0.0225448
R43404 vdd.n1500 vdd.n1499 0.0225448
R43405 vdd.n1506 vdd.n1505 0.0225448
R43406 vdd.n1507 vdd.n1506 0.0225448
R43407 vdd.n1516 vdd.n1515 0.0225448
R43408 vdd.n1515 vdd.n1514 0.0225448
R43409 vdd.n1835 vdd.n1834 0.0225448
R43410 vdd.n1843 vdd.n1842 0.0225448
R43411 vdd.n1842 vdd.n1841 0.0225448
R43412 vdd.n1857 vdd.n1856 0.0225448
R43413 vdd.n1858 vdd.n1857 0.0225448
R43414 vdd.n1854 vdd.n1853 0.0225448
R43415 vdd.n1853 vdd.n1852 0.0225448
R43416 vdd.n1850 vdd.n1849 0.0225448
R43417 vdd.n1860 vdd.n1859 0.0225448
R43418 vdd.n1859 vdd.n1858 0.0225448
R43419 vdd.n1840 vdd.n1816 0.0225448
R43420 vdd.n1841 vdd.n1840 0.0225448
R43421 vdd.n1838 vdd.n1832 0.0225448
R43422 vdd.n1838 vdd.n1837 0.0225448
R43423 vdd.n1882 vdd.n1881 0.0225448
R43424 vdd.n1890 vdd.n1889 0.0225448
R43425 vdd.n1889 vdd.n1888 0.0225448
R43426 vdd.n1904 vdd.n1903 0.0225448
R43427 vdd.n1905 vdd.n1904 0.0225448
R43428 vdd.n1901 vdd.n1900 0.0225448
R43429 vdd.n1900 vdd.n1899 0.0225448
R43430 vdd.n1897 vdd.n1896 0.0225448
R43431 vdd.n1907 vdd.n1906 0.0225448
R43432 vdd.n1906 vdd.n1905 0.0225448
R43433 vdd.n1887 vdd.n1863 0.0225448
R43434 vdd.n1888 vdd.n1887 0.0225448
R43435 vdd.n1885 vdd.n1879 0.0225448
R43436 vdd.n1885 vdd.n1884 0.0225448
R43437 vdd.n1930 vdd.n1929 0.0225448
R43438 vdd.n1938 vdd.n1937 0.0225448
R43439 vdd.n1937 vdd.n1936 0.0225448
R43440 vdd.n1952 vdd.n1951 0.0225448
R43441 vdd.n1953 vdd.n1952 0.0225448
R43442 vdd.n1949 vdd.n1948 0.0225448
R43443 vdd.n1948 vdd.n1947 0.0225448
R43444 vdd.n1945 vdd.n1944 0.0225448
R43445 vdd.n1955 vdd.n1954 0.0225448
R43446 vdd.n1954 vdd.n1953 0.0225448
R43447 vdd.n1935 vdd.n1911 0.0225448
R43448 vdd.n1936 vdd.n1935 0.0225448
R43449 vdd.n1933 vdd.n1927 0.0225448
R43450 vdd.n1933 vdd.n1932 0.0225448
R43451 vdd.n1981 vdd.n1980 0.0225448
R43452 vdd.n1989 vdd.n1988 0.0225448
R43453 vdd.n1988 vdd.n1987 0.0225448
R43454 vdd.n2003 vdd.n2002 0.0225448
R43455 vdd.n2004 vdd.n2003 0.0225448
R43456 vdd.n2000 vdd.n1999 0.0225448
R43457 vdd.n1999 vdd.n1998 0.0225448
R43458 vdd.n1996 vdd.n1995 0.0225448
R43459 vdd.n2006 vdd.n2005 0.0225448
R43460 vdd.n2005 vdd.n2004 0.0225448
R43461 vdd.n1986 vdd.n1962 0.0225448
R43462 vdd.n1987 vdd.n1986 0.0225448
R43463 vdd.n1984 vdd.n1978 0.0225448
R43464 vdd.n1984 vdd.n1983 0.0225448
R43465 vdd.n2031 vdd.n2030 0.0225448
R43466 vdd.n2039 vdd.n2038 0.0225448
R43467 vdd.n2038 vdd.n2037 0.0225448
R43468 vdd.n2053 vdd.n2052 0.0225448
R43469 vdd.n2054 vdd.n2053 0.0225448
R43470 vdd.n2050 vdd.n2049 0.0225448
R43471 vdd.n2049 vdd.n2048 0.0225448
R43472 vdd.n2046 vdd.n2045 0.0225448
R43473 vdd.n2056 vdd.n2055 0.0225448
R43474 vdd.n2055 vdd.n2054 0.0225448
R43475 vdd.n2036 vdd.n2012 0.0225448
R43476 vdd.n2037 vdd.n2036 0.0225448
R43477 vdd.n2034 vdd.n2028 0.0225448
R43478 vdd.n2034 vdd.n2033 0.0225448
R43479 vdd.n2079 vdd.n2078 0.0225448
R43480 vdd.n2087 vdd.n2086 0.0225448
R43481 vdd.n2086 vdd.n2085 0.0225448
R43482 vdd.n2101 vdd.n2100 0.0225448
R43483 vdd.n2102 vdd.n2101 0.0225448
R43484 vdd.n2098 vdd.n2097 0.0225448
R43485 vdd.n2097 vdd.n2096 0.0225448
R43486 vdd.n2094 vdd.n2093 0.0225448
R43487 vdd.n2104 vdd.n2103 0.0225448
R43488 vdd.n2103 vdd.n2102 0.0225448
R43489 vdd.n2084 vdd.n2060 0.0225448
R43490 vdd.n2085 vdd.n2084 0.0225448
R43491 vdd.n2082 vdd.n2076 0.0225448
R43492 vdd.n2082 vdd.n2081 0.0225448
R43493 vdd.n2129 vdd.n2128 0.0225448
R43494 vdd.n2137 vdd.n2136 0.0225448
R43495 vdd.n2136 vdd.n2135 0.0225448
R43496 vdd.n2151 vdd.n2150 0.0225448
R43497 vdd.n2152 vdd.n2151 0.0225448
R43498 vdd.n2148 vdd.n2147 0.0225448
R43499 vdd.n2147 vdd.n2146 0.0225448
R43500 vdd.n2144 vdd.n2143 0.0225448
R43501 vdd.n2154 vdd.n2153 0.0225448
R43502 vdd.n2153 vdd.n2152 0.0225448
R43503 vdd.n2134 vdd.n2110 0.0225448
R43504 vdd.n2135 vdd.n2134 0.0225448
R43505 vdd.n2132 vdd.n2126 0.0225448
R43506 vdd.n2132 vdd.n2131 0.0225448
R43507 vdd.n2176 vdd.n2175 0.0225448
R43508 vdd.n2184 vdd.n2183 0.0225448
R43509 vdd.n2183 vdd.n2182 0.0225448
R43510 vdd.n2198 vdd.n2197 0.0225448
R43511 vdd.n2199 vdd.n2198 0.0225448
R43512 vdd.n2195 vdd.n2194 0.0225448
R43513 vdd.n2194 vdd.n2193 0.0225448
R43514 vdd.n2191 vdd.n2190 0.0225448
R43515 vdd.n2201 vdd.n2200 0.0225448
R43516 vdd.n2200 vdd.n2199 0.0225448
R43517 vdd.n2181 vdd.n2157 0.0225448
R43518 vdd.n2182 vdd.n2181 0.0225448
R43519 vdd.n2179 vdd.n2173 0.0225448
R43520 vdd.n2179 vdd.n2178 0.0225448
R43521 vdd.n2226 vdd.n2225 0.0225448
R43522 vdd.n2234 vdd.n2233 0.0225448
R43523 vdd.n2233 vdd.n2232 0.0225448
R43524 vdd.n2248 vdd.n2247 0.0225448
R43525 vdd.n2249 vdd.n2248 0.0225448
R43526 vdd.n2245 vdd.n2244 0.0225448
R43527 vdd.n2244 vdd.n2243 0.0225448
R43528 vdd.n2241 vdd.n2240 0.0225448
R43529 vdd.n2251 vdd.n2250 0.0225448
R43530 vdd.n2250 vdd.n2249 0.0225448
R43531 vdd.n2231 vdd.n2207 0.0225448
R43532 vdd.n2232 vdd.n2231 0.0225448
R43533 vdd.n2229 vdd.n2223 0.0225448
R43534 vdd.n2229 vdd.n2228 0.0225448
R43535 vdd.n2276 vdd.n2275 0.0225448
R43536 vdd.n2284 vdd.n2283 0.0225448
R43537 vdd.n2283 vdd.n2282 0.0225448
R43538 vdd.n2298 vdd.n2297 0.0225448
R43539 vdd.n2299 vdd.n2298 0.0225448
R43540 vdd.n2295 vdd.n2294 0.0225448
R43541 vdd.n2294 vdd.n2293 0.0225448
R43542 vdd.n2291 vdd.n2290 0.0225448
R43543 vdd.n2301 vdd.n2300 0.0225448
R43544 vdd.n2300 vdd.n2299 0.0225448
R43545 vdd.n2281 vdd.n2257 0.0225448
R43546 vdd.n2282 vdd.n2281 0.0225448
R43547 vdd.n2279 vdd.n2273 0.0225448
R43548 vdd.n2279 vdd.n2278 0.0225448
R43549 vdd.n2324 vdd.n2323 0.0225448
R43550 vdd.n2332 vdd.n2331 0.0225448
R43551 vdd.n2331 vdd.n2330 0.0225448
R43552 vdd.n2346 vdd.n2345 0.0225448
R43553 vdd.n2347 vdd.n2346 0.0225448
R43554 vdd.n2343 vdd.n2342 0.0225448
R43555 vdd.n2342 vdd.n2341 0.0225448
R43556 vdd.n2339 vdd.n2338 0.0225448
R43557 vdd.n2349 vdd.n2348 0.0225448
R43558 vdd.n2348 vdd.n2347 0.0225448
R43559 vdd.n2329 vdd.n2305 0.0225448
R43560 vdd.n2330 vdd.n2329 0.0225448
R43561 vdd.n2327 vdd.n2321 0.0225448
R43562 vdd.n2327 vdd.n2326 0.0225448
R43563 vdd.n1267 vdd.n1266 0.0225448
R43564 vdd.n1264 vdd.n1263 0.0225448
R43565 vdd.n1263 vdd.n1262 0.0225448
R43566 vdd.n1253 vdd.n1252 0.0225448
R43567 vdd.n1254 vdd.n1253 0.0225448
R43568 vdd.n1250 vdd.n1249 0.0225448
R43569 vdd.n1249 vdd.n1248 0.0225448
R43570 vdd.n1246 vdd.n1245 0.0225448
R43571 vdd.n1255 vdd.n1237 0.0225448
R43572 vdd.n1255 vdd.n1254 0.0225448
R43573 vdd.n1261 vdd.n1260 0.0225448
R43574 vdd.n1262 vdd.n1261 0.0225448
R43575 vdd.n1271 vdd.n1270 0.0225448
R43576 vdd.n1270 vdd.n1269 0.0225448
R43577 vdd.n2375 vdd.n2374 0.0225448
R43578 vdd.n2383 vdd.n2382 0.0225448
R43579 vdd.n2382 vdd.n2381 0.0225448
R43580 vdd.n2397 vdd.n2396 0.0225448
R43581 vdd.n2398 vdd.n2397 0.0225448
R43582 vdd.n2394 vdd.n2393 0.0225448
R43583 vdd.n2393 vdd.n2392 0.0225448
R43584 vdd.n2390 vdd.n2389 0.0225448
R43585 vdd.n2400 vdd.n2399 0.0225448
R43586 vdd.n2399 vdd.n2398 0.0225448
R43587 vdd.n2380 vdd.n2356 0.0225448
R43588 vdd.n2381 vdd.n2380 0.0225448
R43589 vdd.n2378 vdd.n2372 0.0225448
R43590 vdd.n2378 vdd.n2377 0.0225448
R43591 vdd.n2422 vdd.n2421 0.0225448
R43592 vdd.n2430 vdd.n2429 0.0225448
R43593 vdd.n2429 vdd.n2428 0.0225448
R43594 vdd.n2444 vdd.n2443 0.0225448
R43595 vdd.n2445 vdd.n2444 0.0225448
R43596 vdd.n2441 vdd.n2440 0.0225448
R43597 vdd.n2440 vdd.n2439 0.0225448
R43598 vdd.n2437 vdd.n2436 0.0225448
R43599 vdd.n2447 vdd.n2446 0.0225448
R43600 vdd.n2446 vdd.n2445 0.0225448
R43601 vdd.n2427 vdd.n2403 0.0225448
R43602 vdd.n2428 vdd.n2427 0.0225448
R43603 vdd.n2425 vdd.n2419 0.0225448
R43604 vdd.n2425 vdd.n2424 0.0225448
R43605 vdd.n2472 vdd.n2471 0.0225448
R43606 vdd.n2480 vdd.n2479 0.0225448
R43607 vdd.n2479 vdd.n2478 0.0225448
R43608 vdd.n2494 vdd.n2493 0.0225448
R43609 vdd.n2495 vdd.n2494 0.0225448
R43610 vdd.n2491 vdd.n2490 0.0225448
R43611 vdd.n2490 vdd.n2489 0.0225448
R43612 vdd.n2487 vdd.n2486 0.0225448
R43613 vdd.n2497 vdd.n2496 0.0225448
R43614 vdd.n2496 vdd.n2495 0.0225448
R43615 vdd.n2477 vdd.n2453 0.0225448
R43616 vdd.n2478 vdd.n2477 0.0225448
R43617 vdd.n2475 vdd.n2469 0.0225448
R43618 vdd.n2475 vdd.n2474 0.0225448
R43619 vdd.n2522 vdd.n2521 0.0225448
R43620 vdd.n2530 vdd.n2529 0.0225448
R43621 vdd.n2529 vdd.n2528 0.0225448
R43622 vdd.n2544 vdd.n2543 0.0225448
R43623 vdd.n2545 vdd.n2544 0.0225448
R43624 vdd.n2541 vdd.n2540 0.0225448
R43625 vdd.n2540 vdd.n2539 0.0225448
R43626 vdd.n2537 vdd.n2536 0.0225448
R43627 vdd.n2547 vdd.n2546 0.0225448
R43628 vdd.n2546 vdd.n2545 0.0225448
R43629 vdd.n2527 vdd.n2503 0.0225448
R43630 vdd.n2528 vdd.n2527 0.0225448
R43631 vdd.n2525 vdd.n2519 0.0225448
R43632 vdd.n2525 vdd.n2524 0.0225448
R43633 vdd.n2570 vdd.n2569 0.0225448
R43634 vdd.n2578 vdd.n2577 0.0225448
R43635 vdd.n2577 vdd.n2576 0.0225448
R43636 vdd.n2592 vdd.n2591 0.0225448
R43637 vdd.n2593 vdd.n2592 0.0225448
R43638 vdd.n2589 vdd.n2588 0.0225448
R43639 vdd.n2588 vdd.n2587 0.0225448
R43640 vdd.n2585 vdd.n2584 0.0225448
R43641 vdd.n2595 vdd.n2594 0.0225448
R43642 vdd.n2594 vdd.n2593 0.0225448
R43643 vdd.n2575 vdd.n2551 0.0225448
R43644 vdd.n2576 vdd.n2575 0.0225448
R43645 vdd.n2573 vdd.n2567 0.0225448
R43646 vdd.n2573 vdd.n2572 0.0225448
R43647 vdd.n2713 vdd.n2711 0.0225448
R43648 vdd.n2713 vdd.n2712 0.0225448
R43649 vdd.n2724 vdd.n2723 0.0225448
R43650 vdd.n2723 vdd.n2722 0.0225448
R43651 vdd.n2738 vdd.n2737 0.0225448
R43652 vdd.n2739 vdd.n2738 0.0225448
R43653 vdd.n2735 vdd.n2734 0.0225448
R43654 vdd.n2731 vdd.n2730 0.0225448
R43655 vdd.n2732 vdd.n2731 0.0225448
R43656 vdd.n2741 vdd.n2740 0.0225448
R43657 vdd.n2740 vdd.n2739 0.0225448
R43658 vdd.n2721 vdd.n2697 0.0225448
R43659 vdd.n2722 vdd.n2721 0.0225448
R43660 vdd.n2719 vdd.n2718 0.0225448
R43661 vdd.n2665 vdd.n2663 0.0225448
R43662 vdd.n2665 vdd.n2664 0.0225448
R43663 vdd.n2676 vdd.n2675 0.0225448
R43664 vdd.n2675 vdd.n2674 0.0225448
R43665 vdd.n2690 vdd.n2689 0.0225448
R43666 vdd.n2691 vdd.n2690 0.0225448
R43667 vdd.n2687 vdd.n2686 0.0225448
R43668 vdd.n2683 vdd.n2682 0.0225448
R43669 vdd.n2684 vdd.n2683 0.0225448
R43670 vdd.n2693 vdd.n2692 0.0225448
R43671 vdd.n2692 vdd.n2691 0.0225448
R43672 vdd.n2673 vdd.n2649 0.0225448
R43673 vdd.n2674 vdd.n2673 0.0225448
R43674 vdd.n2671 vdd.n2670 0.0225448
R43675 vdd.n2762 vdd.n2760 0.0225448
R43676 vdd.n2762 vdd.n2761 0.0225448
R43677 vdd.n2773 vdd.n2772 0.0225448
R43678 vdd.n2772 vdd.n2771 0.0225448
R43679 vdd.n2787 vdd.n2786 0.0225448
R43680 vdd.n2788 vdd.n2787 0.0225448
R43681 vdd.n2784 vdd.n2783 0.0225448
R43682 vdd.n2780 vdd.n2779 0.0225448
R43683 vdd.n2781 vdd.n2780 0.0225448
R43684 vdd.n2790 vdd.n2789 0.0225448
R43685 vdd.n2789 vdd.n2788 0.0225448
R43686 vdd.n2770 vdd.n2746 0.0225448
R43687 vdd.n2771 vdd.n2770 0.0225448
R43688 vdd.n2768 vdd.n2767 0.0225448
R43689 vdd.n2812 vdd.n2810 0.0225448
R43690 vdd.n2812 vdd.n2811 0.0225448
R43691 vdd.n2823 vdd.n2822 0.0225448
R43692 vdd.n2822 vdd.n2821 0.0225448
R43693 vdd.n2837 vdd.n2836 0.0225448
R43694 vdd.n2838 vdd.n2837 0.0225448
R43695 vdd.n2834 vdd.n2833 0.0225448
R43696 vdd.n2830 vdd.n2829 0.0225448
R43697 vdd.n2831 vdd.n2830 0.0225448
R43698 vdd.n2840 vdd.n2839 0.0225448
R43699 vdd.n2839 vdd.n2838 0.0225448
R43700 vdd.n2820 vdd.n2796 0.0225448
R43701 vdd.n2821 vdd.n2820 0.0225448
R43702 vdd.n2818 vdd.n2817 0.0225448
R43703 vdd.n2860 vdd.n2858 0.0225448
R43704 vdd.n2860 vdd.n2859 0.0225448
R43705 vdd.n2871 vdd.n2870 0.0225448
R43706 vdd.n2870 vdd.n2869 0.0225448
R43707 vdd.n2885 vdd.n2884 0.0225448
R43708 vdd.n2886 vdd.n2885 0.0225448
R43709 vdd.n2882 vdd.n2881 0.0225448
R43710 vdd.n2878 vdd.n2877 0.0225448
R43711 vdd.n2879 vdd.n2878 0.0225448
R43712 vdd.n2888 vdd.n2887 0.0225448
R43713 vdd.n2887 vdd.n2886 0.0225448
R43714 vdd.n2868 vdd.n2844 0.0225448
R43715 vdd.n2869 vdd.n2868 0.0225448
R43716 vdd.n2866 vdd.n2865 0.0225448
R43717 vdd.n1047 vdd.n1046 0.0225448
R43718 vdd.n1048 vdd.n1047 0.0225448
R43719 vdd.n1044 vdd.n1037 0.0225448
R43720 vdd.n1055 vdd.n1037 0.0225448
R43721 vdd.n1057 vdd.n1056 0.0225448
R43722 vdd.n1058 vdd.n1057 0.0225448
R43723 vdd.n1072 vdd.n1071 0.0225448
R43724 vdd.n1068 vdd.n1027 0.0225448
R43725 vdd.n1069 vdd.n1068 0.0225448
R43726 vdd.n1063 vdd.n1032 0.0225448
R43727 vdd.n1058 vdd.n1032 0.0225448
R43728 vdd.n1054 vdd.n1053 0.0225448
R43729 vdd.n1055 vdd.n1054 0.0225448
R43730 vdd.n1051 vdd.n1050 0.0225448
R43731 vdd.n3008 vdd.n3006 0.0225448
R43732 vdd.n3008 vdd.n3007 0.0225448
R43733 vdd.n3019 vdd.n3018 0.0225448
R43734 vdd.n3018 vdd.n3017 0.0225448
R43735 vdd.n3033 vdd.n3032 0.0225448
R43736 vdd.n3034 vdd.n3033 0.0225448
R43737 vdd.n3030 vdd.n3029 0.0225448
R43738 vdd.n3026 vdd.n3025 0.0225448
R43739 vdd.n3027 vdd.n3026 0.0225448
R43740 vdd.n3036 vdd.n3035 0.0225448
R43741 vdd.n3035 vdd.n3034 0.0225448
R43742 vdd.n3016 vdd.n2992 0.0225448
R43743 vdd.n3017 vdd.n3016 0.0225448
R43744 vdd.n3014 vdd.n3013 0.0225448
R43745 vdd.n2959 vdd.n2957 0.0225448
R43746 vdd.n2959 vdd.n2958 0.0225448
R43747 vdd.n2970 vdd.n2969 0.0225448
R43748 vdd.n2969 vdd.n2968 0.0225448
R43749 vdd.n2984 vdd.n2983 0.0225448
R43750 vdd.n2985 vdd.n2984 0.0225448
R43751 vdd.n2981 vdd.n2980 0.0225448
R43752 vdd.n2977 vdd.n2976 0.0225448
R43753 vdd.n2978 vdd.n2977 0.0225448
R43754 vdd.n2987 vdd.n2986 0.0225448
R43755 vdd.n2986 vdd.n2985 0.0225448
R43756 vdd.n2967 vdd.n2943 0.0225448
R43757 vdd.n2968 vdd.n2967 0.0225448
R43758 vdd.n2965 vdd.n2964 0.0225448
R43759 vdd.n2911 vdd.n2909 0.0225448
R43760 vdd.n2911 vdd.n2910 0.0225448
R43761 vdd.n2922 vdd.n2921 0.0225448
R43762 vdd.n2921 vdd.n2920 0.0225448
R43763 vdd.n2936 vdd.n2935 0.0225448
R43764 vdd.n2937 vdd.n2936 0.0225448
R43765 vdd.n2933 vdd.n2932 0.0225448
R43766 vdd.n2929 vdd.n2928 0.0225448
R43767 vdd.n2930 vdd.n2929 0.0225448
R43768 vdd.n2939 vdd.n2938 0.0225448
R43769 vdd.n2938 vdd.n2937 0.0225448
R43770 vdd.n2919 vdd.n2895 0.0225448
R43771 vdd.n2920 vdd.n2919 0.0225448
R43772 vdd.n2917 vdd.n2916 0.0225448
R43773 vdd.n3057 vdd.n3055 0.0225448
R43774 vdd.n3057 vdd.n3056 0.0225448
R43775 vdd.n3068 vdd.n3067 0.0225448
R43776 vdd.n3067 vdd.n3066 0.0225448
R43777 vdd.n3082 vdd.n3081 0.0225448
R43778 vdd.n3083 vdd.n3082 0.0225448
R43779 vdd.n3079 vdd.n3078 0.0225448
R43780 vdd.n3075 vdd.n3074 0.0225448
R43781 vdd.n3076 vdd.n3075 0.0225448
R43782 vdd.n3085 vdd.n3084 0.0225448
R43783 vdd.n3084 vdd.n3083 0.0225448
R43784 vdd.n3065 vdd.n3041 0.0225448
R43785 vdd.n3066 vdd.n3065 0.0225448
R43786 vdd.n3063 vdd.n3062 0.0225448
R43787 vdd.n3107 vdd.n3105 0.0225448
R43788 vdd.n3107 vdd.n3106 0.0225448
R43789 vdd.n3118 vdd.n3117 0.0225448
R43790 vdd.n3117 vdd.n3116 0.0225448
R43791 vdd.n3132 vdd.n3131 0.0225448
R43792 vdd.n3133 vdd.n3132 0.0225448
R43793 vdd.n3129 vdd.n3128 0.0225448
R43794 vdd.n3125 vdd.n3124 0.0225448
R43795 vdd.n3126 vdd.n3125 0.0225448
R43796 vdd.n3135 vdd.n3134 0.0225448
R43797 vdd.n3134 vdd.n3133 0.0225448
R43798 vdd.n3115 vdd.n3091 0.0225448
R43799 vdd.n3116 vdd.n3115 0.0225448
R43800 vdd.n3113 vdd.n3112 0.0225448
R43801 vdd.n3155 vdd.n3153 0.0225448
R43802 vdd.n3155 vdd.n3154 0.0225448
R43803 vdd.n3166 vdd.n3165 0.0225448
R43804 vdd.n3165 vdd.n3164 0.0225448
R43805 vdd.n3180 vdd.n3179 0.0225448
R43806 vdd.n3181 vdd.n3180 0.0225448
R43807 vdd.n3177 vdd.n3176 0.0225448
R43808 vdd.n3173 vdd.n3172 0.0225448
R43809 vdd.n3174 vdd.n3173 0.0225448
R43810 vdd.n3183 vdd.n3182 0.0225448
R43811 vdd.n3182 vdd.n3181 0.0225448
R43812 vdd.n3163 vdd.n3139 0.0225448
R43813 vdd.n3164 vdd.n3163 0.0225448
R43814 vdd.n3161 vdd.n3160 0.0225448
R43815 vdd.n3253 vdd.n3251 0.0225448
R43816 vdd.n3253 vdd.n3252 0.0225448
R43817 vdd.n3264 vdd.n3263 0.0225448
R43818 vdd.n3263 vdd.n3262 0.0225448
R43819 vdd.n3278 vdd.n3277 0.0225448
R43820 vdd.n3279 vdd.n3278 0.0225448
R43821 vdd.n3275 vdd.n3274 0.0225448
R43822 vdd.n3271 vdd.n3270 0.0225448
R43823 vdd.n3272 vdd.n3271 0.0225448
R43824 vdd.n3281 vdd.n3280 0.0225448
R43825 vdd.n3280 vdd.n3279 0.0225448
R43826 vdd.n3261 vdd.n3237 0.0225448
R43827 vdd.n3262 vdd.n3261 0.0225448
R43828 vdd.n3259 vdd.n3258 0.0225448
R43829 vdd.n3205 vdd.n3203 0.0225448
R43830 vdd.n3205 vdd.n3204 0.0225448
R43831 vdd.n3216 vdd.n3215 0.0225448
R43832 vdd.n3215 vdd.n3214 0.0225448
R43833 vdd.n3230 vdd.n3229 0.0225448
R43834 vdd.n3231 vdd.n3230 0.0225448
R43835 vdd.n3227 vdd.n3226 0.0225448
R43836 vdd.n3223 vdd.n3222 0.0225448
R43837 vdd.n3224 vdd.n3223 0.0225448
R43838 vdd.n3233 vdd.n3232 0.0225448
R43839 vdd.n3232 vdd.n3231 0.0225448
R43840 vdd.n3213 vdd.n3189 0.0225448
R43841 vdd.n3214 vdd.n3213 0.0225448
R43842 vdd.n3211 vdd.n3210 0.0225448
R43843 vdd.n3302 vdd.n3300 0.0225448
R43844 vdd.n3302 vdd.n3301 0.0225448
R43845 vdd.n3313 vdd.n3312 0.0225448
R43846 vdd.n3312 vdd.n3311 0.0225448
R43847 vdd.n3327 vdd.n3326 0.0225448
R43848 vdd.n3328 vdd.n3327 0.0225448
R43849 vdd.n3324 vdd.n3323 0.0225448
R43850 vdd.n3320 vdd.n3319 0.0225448
R43851 vdd.n3321 vdd.n3320 0.0225448
R43852 vdd.n3330 vdd.n3329 0.0225448
R43853 vdd.n3329 vdd.n3328 0.0225448
R43854 vdd.n3310 vdd.n3286 0.0225448
R43855 vdd.n3311 vdd.n3310 0.0225448
R43856 vdd.n3308 vdd.n3307 0.0225448
R43857 vdd.n3352 vdd.n3350 0.0225448
R43858 vdd.n3352 vdd.n3351 0.0225448
R43859 vdd.n3363 vdd.n3362 0.0225448
R43860 vdd.n3362 vdd.n3361 0.0225448
R43861 vdd.n3377 vdd.n3376 0.0225448
R43862 vdd.n3378 vdd.n3377 0.0225448
R43863 vdd.n3374 vdd.n3373 0.0225448
R43864 vdd.n3370 vdd.n3369 0.0225448
R43865 vdd.n3371 vdd.n3370 0.0225448
R43866 vdd.n3380 vdd.n3379 0.0225448
R43867 vdd.n3379 vdd.n3378 0.0225448
R43868 vdd.n3360 vdd.n3336 0.0225448
R43869 vdd.n3361 vdd.n3360 0.0225448
R43870 vdd.n3358 vdd.n3357 0.0225448
R43871 vdd.n3400 vdd.n3398 0.0225448
R43872 vdd.n3400 vdd.n3399 0.0225448
R43873 vdd.n3411 vdd.n3410 0.0225448
R43874 vdd.n3410 vdd.n3409 0.0225448
R43875 vdd.n3425 vdd.n3424 0.0225448
R43876 vdd.n3426 vdd.n3425 0.0225448
R43877 vdd.n3422 vdd.n3421 0.0225448
R43878 vdd.n3418 vdd.n3417 0.0225448
R43879 vdd.n3419 vdd.n3418 0.0225448
R43880 vdd.n3428 vdd.n3427 0.0225448
R43881 vdd.n3427 vdd.n3426 0.0225448
R43882 vdd.n3408 vdd.n3384 0.0225448
R43883 vdd.n3409 vdd.n3408 0.0225448
R43884 vdd.n3406 vdd.n3405 0.0225448
R43885 vdd.n801 vdd.n800 0.0225448
R43886 vdd.n802 vdd.n801 0.0225448
R43887 vdd.n798 vdd.n791 0.0225448
R43888 vdd.n809 vdd.n791 0.0225448
R43889 vdd.n811 vdd.n810 0.0225448
R43890 vdd.n812 vdd.n811 0.0225448
R43891 vdd.n826 vdd.n825 0.0225448
R43892 vdd.n822 vdd.n781 0.0225448
R43893 vdd.n823 vdd.n822 0.0225448
R43894 vdd.n817 vdd.n786 0.0225448
R43895 vdd.n812 vdd.n786 0.0225448
R43896 vdd.n808 vdd.n807 0.0225448
R43897 vdd.n809 vdd.n808 0.0225448
R43898 vdd.n805 vdd.n804 0.0225448
R43899 vdd.n3499 vdd.n3497 0.0225448
R43900 vdd.n3499 vdd.n3498 0.0225448
R43901 vdd.n3510 vdd.n3509 0.0225448
R43902 vdd.n3509 vdd.n3508 0.0225448
R43903 vdd.n3524 vdd.n3523 0.0225448
R43904 vdd.n3525 vdd.n3524 0.0225448
R43905 vdd.n3521 vdd.n3520 0.0225448
R43906 vdd.n3517 vdd.n3516 0.0225448
R43907 vdd.n3518 vdd.n3517 0.0225448
R43908 vdd.n3527 vdd.n3526 0.0225448
R43909 vdd.n3526 vdd.n3525 0.0225448
R43910 vdd.n3507 vdd.n3483 0.0225448
R43911 vdd.n3508 vdd.n3507 0.0225448
R43912 vdd.n3505 vdd.n3504 0.0225448
R43913 vdd.n3451 vdd.n3449 0.0225448
R43914 vdd.n3451 vdd.n3450 0.0225448
R43915 vdd.n3462 vdd.n3461 0.0225448
R43916 vdd.n3461 vdd.n3460 0.0225448
R43917 vdd.n3476 vdd.n3475 0.0225448
R43918 vdd.n3477 vdd.n3476 0.0225448
R43919 vdd.n3473 vdd.n3472 0.0225448
R43920 vdd.n3469 vdd.n3468 0.0225448
R43921 vdd.n3470 vdd.n3469 0.0225448
R43922 vdd.n3479 vdd.n3478 0.0225448
R43923 vdd.n3478 vdd.n3477 0.0225448
R43924 vdd.n3459 vdd.n3435 0.0225448
R43925 vdd.n3460 vdd.n3459 0.0225448
R43926 vdd.n3457 vdd.n3456 0.0225448
R43927 vdd.n3548 vdd.n3546 0.0225448
R43928 vdd.n3548 vdd.n3547 0.0225448
R43929 vdd.n3559 vdd.n3558 0.0225448
R43930 vdd.n3558 vdd.n3557 0.0225448
R43931 vdd.n3573 vdd.n3572 0.0225448
R43932 vdd.n3574 vdd.n3573 0.0225448
R43933 vdd.n3570 vdd.n3569 0.0225448
R43934 vdd.n3566 vdd.n3565 0.0225448
R43935 vdd.n3567 vdd.n3566 0.0225448
R43936 vdd.n3576 vdd.n3575 0.0225448
R43937 vdd.n3575 vdd.n3574 0.0225448
R43938 vdd.n3556 vdd.n3532 0.0225448
R43939 vdd.n3557 vdd.n3556 0.0225448
R43940 vdd.n3554 vdd.n3553 0.0225448
R43941 vdd.n3598 vdd.n3596 0.0225448
R43942 vdd.n3598 vdd.n3597 0.0225448
R43943 vdd.n3609 vdd.n3608 0.0225448
R43944 vdd.n3608 vdd.n3607 0.0225448
R43945 vdd.n3623 vdd.n3622 0.0225448
R43946 vdd.n3624 vdd.n3623 0.0225448
R43947 vdd.n3620 vdd.n3619 0.0225448
R43948 vdd.n3616 vdd.n3615 0.0225448
R43949 vdd.n3617 vdd.n3616 0.0225448
R43950 vdd.n3626 vdd.n3625 0.0225448
R43951 vdd.n3625 vdd.n3624 0.0225448
R43952 vdd.n3606 vdd.n3582 0.0225448
R43953 vdd.n3607 vdd.n3606 0.0225448
R43954 vdd.n3604 vdd.n3603 0.0225448
R43955 vdd.n3646 vdd.n3644 0.0225448
R43956 vdd.n3646 vdd.n3645 0.0225448
R43957 vdd.n3657 vdd.n3656 0.0225448
R43958 vdd.n3656 vdd.n3655 0.0225448
R43959 vdd.n3671 vdd.n3670 0.0225448
R43960 vdd.n3672 vdd.n3671 0.0225448
R43961 vdd.n3668 vdd.n3667 0.0225448
R43962 vdd.n3664 vdd.n3663 0.0225448
R43963 vdd.n3665 vdd.n3664 0.0225448
R43964 vdd.n3674 vdd.n3673 0.0225448
R43965 vdd.n3673 vdd.n3672 0.0225448
R43966 vdd.n3654 vdd.n3630 0.0225448
R43967 vdd.n3655 vdd.n3654 0.0225448
R43968 vdd.n3652 vdd.n3651 0.0225448
R43969 vdd.n604 vdd.n602 0.0225448
R43970 vdd.n604 vdd.n603 0.0225448
R43971 vdd.n615 vdd.n614 0.0225448
R43972 vdd.n614 vdd.n613 0.0225448
R43973 vdd.n629 vdd.n628 0.0225448
R43974 vdd.n630 vdd.n629 0.0225448
R43975 vdd.n626 vdd.n625 0.0225448
R43976 vdd.n622 vdd.n621 0.0225448
R43977 vdd.n623 vdd.n622 0.0225448
R43978 vdd.n632 vdd.n631 0.0225448
R43979 vdd.n631 vdd.n630 0.0225448
R43980 vdd.n612 vdd.n588 0.0225448
R43981 vdd.n613 vdd.n612 0.0225448
R43982 vdd.n610 vdd.n609 0.0225448
R43983 vdd.n3745 vdd.n3743 0.0225448
R43984 vdd.n3745 vdd.n3744 0.0225448
R43985 vdd.n3756 vdd.n3755 0.0225448
R43986 vdd.n3755 vdd.n3754 0.0225448
R43987 vdd.n3770 vdd.n3769 0.0225448
R43988 vdd.n3771 vdd.n3770 0.0225448
R43989 vdd.n3767 vdd.n3766 0.0225448
R43990 vdd.n3763 vdd.n3762 0.0225448
R43991 vdd.n3764 vdd.n3763 0.0225448
R43992 vdd.n3773 vdd.n3772 0.0225448
R43993 vdd.n3772 vdd.n3771 0.0225448
R43994 vdd.n3753 vdd.n3729 0.0225448
R43995 vdd.n3754 vdd.n3753 0.0225448
R43996 vdd.n3751 vdd.n3750 0.0225448
R43997 vdd.n3697 vdd.n3695 0.0225448
R43998 vdd.n3697 vdd.n3696 0.0225448
R43999 vdd.n3708 vdd.n3707 0.0225448
R44000 vdd.n3707 vdd.n3706 0.0225448
R44001 vdd.n3722 vdd.n3721 0.0225448
R44002 vdd.n3723 vdd.n3722 0.0225448
R44003 vdd.n3719 vdd.n3718 0.0225448
R44004 vdd.n3715 vdd.n3714 0.0225448
R44005 vdd.n3716 vdd.n3715 0.0225448
R44006 vdd.n3725 vdd.n3724 0.0225448
R44007 vdd.n3724 vdd.n3723 0.0225448
R44008 vdd.n3705 vdd.n3681 0.0225448
R44009 vdd.n3706 vdd.n3705 0.0225448
R44010 vdd.n3703 vdd.n3702 0.0225448
R44011 vdd.n6887 vdd.n6885 0.0225448
R44012 vdd.n6887 vdd.n6886 0.0225448
R44013 vdd.n6898 vdd.n6897 0.0225448
R44014 vdd.n6897 vdd.n6896 0.0225448
R44015 vdd.n6912 vdd.n6911 0.0225448
R44016 vdd.n6913 vdd.n6912 0.0225448
R44017 vdd.n6909 vdd.n6908 0.0225448
R44018 vdd.n6905 vdd.n6904 0.0225448
R44019 vdd.n6906 vdd.n6905 0.0225448
R44020 vdd.n6915 vdd.n6914 0.0225448
R44021 vdd.n6914 vdd.n6913 0.0225448
R44022 vdd.n6895 vdd.n6871 0.0225448
R44023 vdd.n6896 vdd.n6895 0.0225448
R44024 vdd.n6893 vdd.n6892 0.0225448
R44025 vdd.n6839 vdd.n6837 0.0225448
R44026 vdd.n6839 vdd.n6838 0.0225448
R44027 vdd.n6850 vdd.n6849 0.0225448
R44028 vdd.n6849 vdd.n6848 0.0225448
R44029 vdd.n6864 vdd.n6863 0.0225448
R44030 vdd.n6865 vdd.n6864 0.0225448
R44031 vdd.n6861 vdd.n6860 0.0225448
R44032 vdd.n6857 vdd.n6856 0.0225448
R44033 vdd.n6858 vdd.n6857 0.0225448
R44034 vdd.n6867 vdd.n6866 0.0225448
R44035 vdd.n6866 vdd.n6865 0.0225448
R44036 vdd.n6847 vdd.n6823 0.0225448
R44037 vdd.n6848 vdd.n6847 0.0225448
R44038 vdd.n6845 vdd.n6844 0.0225448
R44039 vdd.n10029 vdd.n10027 0.0225448
R44040 vdd.n10029 vdd.n10028 0.0225448
R44041 vdd.n10040 vdd.n10039 0.0225448
R44042 vdd.n10039 vdd.n10038 0.0225448
R44043 vdd.n10054 vdd.n10053 0.0225448
R44044 vdd.n10055 vdd.n10054 0.0225448
R44045 vdd.n10051 vdd.n10050 0.0225448
R44046 vdd.n10047 vdd.n10046 0.0225448
R44047 vdd.n10048 vdd.n10047 0.0225448
R44048 vdd.n10057 vdd.n10056 0.0225448
R44049 vdd.n10056 vdd.n10055 0.0225448
R44050 vdd.n10037 vdd.n10013 0.0225448
R44051 vdd.n10038 vdd.n10037 0.0225448
R44052 vdd.n10035 vdd.n10034 0.0225448
R44053 vdd.n9981 vdd.n9979 0.0225448
R44054 vdd.n9981 vdd.n9980 0.0225448
R44055 vdd.n9992 vdd.n9991 0.0225448
R44056 vdd.n9991 vdd.n9990 0.0225448
R44057 vdd.n10006 vdd.n10005 0.0225448
R44058 vdd.n10007 vdd.n10006 0.0225448
R44059 vdd.n10003 vdd.n10002 0.0225448
R44060 vdd.n9999 vdd.n9998 0.0225448
R44061 vdd.n10000 vdd.n9999 0.0225448
R44062 vdd.n10009 vdd.n10008 0.0225448
R44063 vdd.n10008 vdd.n10007 0.0225448
R44064 vdd.n9989 vdd.n9965 0.0225448
R44065 vdd.n9990 vdd.n9989 0.0225448
R44066 vdd.n9987 vdd.n9986 0.0225448
R44067 vdd.n10077 vdd.n10075 0.0225448
R44068 vdd.n10077 vdd.n10076 0.0225448
R44069 vdd.n10088 vdd.n10087 0.0225448
R44070 vdd.n10087 vdd.n10086 0.0225448
R44071 vdd.n10102 vdd.n10101 0.0225448
R44072 vdd.n10103 vdd.n10102 0.0225448
R44073 vdd.n10099 vdd.n10098 0.0225448
R44074 vdd.n10095 vdd.n10094 0.0225448
R44075 vdd.n10096 vdd.n10095 0.0225448
R44076 vdd.n10105 vdd.n10104 0.0225448
R44077 vdd.n10104 vdd.n10103 0.0225448
R44078 vdd.n10085 vdd.n10061 0.0225448
R44079 vdd.n10086 vdd.n10085 0.0225448
R44080 vdd.n10083 vdd.n10082 0.0225448
R44081 vdd.n10125 vdd.n10123 0.0225448
R44082 vdd.n10125 vdd.n10124 0.0225448
R44083 vdd.n10136 vdd.n10135 0.0225448
R44084 vdd.n10135 vdd.n10134 0.0225448
R44085 vdd.n10150 vdd.n10149 0.0225448
R44086 vdd.n10151 vdd.n10150 0.0225448
R44087 vdd.n10147 vdd.n10146 0.0225448
R44088 vdd.n10143 vdd.n10142 0.0225448
R44089 vdd.n10144 vdd.n10143 0.0225448
R44090 vdd.n10153 vdd.n10152 0.0225448
R44091 vdd.n10152 vdd.n10151 0.0225448
R44092 vdd.n10133 vdd.n10109 0.0225448
R44093 vdd.n10134 vdd.n10133 0.0225448
R44094 vdd.n10131 vdd.n10130 0.0225448
R44095 vdd.n10227 vdd.n10225 0.0225448
R44096 vdd.n10227 vdd.n10226 0.0225448
R44097 vdd.n10238 vdd.n10237 0.0225448
R44098 vdd.n10237 vdd.n10236 0.0225448
R44099 vdd.n10252 vdd.n10251 0.0225448
R44100 vdd.n10253 vdd.n10252 0.0225448
R44101 vdd.n10249 vdd.n10248 0.0225448
R44102 vdd.n10245 vdd.n10244 0.0225448
R44103 vdd.n10246 vdd.n10245 0.0225448
R44104 vdd.n10255 vdd.n10254 0.0225448
R44105 vdd.n10254 vdd.n10253 0.0225448
R44106 vdd.n10235 vdd.n10211 0.0225448
R44107 vdd.n10236 vdd.n10235 0.0225448
R44108 vdd.n10233 vdd.n10232 0.0225448
R44109 vdd.n10275 vdd.n10273 0.0225448
R44110 vdd.n10275 vdd.n10274 0.0225448
R44111 vdd.n10286 vdd.n10285 0.0225448
R44112 vdd.n10285 vdd.n10284 0.0225448
R44113 vdd.n10300 vdd.n10299 0.0225448
R44114 vdd.n10301 vdd.n10300 0.0225448
R44115 vdd.n10297 vdd.n10296 0.0225448
R44116 vdd.n10293 vdd.n10292 0.0225448
R44117 vdd.n10294 vdd.n10293 0.0225448
R44118 vdd.n10303 vdd.n10302 0.0225448
R44119 vdd.n10302 vdd.n10301 0.0225448
R44120 vdd.n10283 vdd.n10259 0.0225448
R44121 vdd.n10284 vdd.n10283 0.0225448
R44122 vdd.n10281 vdd.n10280 0.0225448
R44123 vdd.n10323 vdd.n10321 0.0225448
R44124 vdd.n10323 vdd.n10322 0.0225448
R44125 vdd.n10334 vdd.n10333 0.0225448
R44126 vdd.n10333 vdd.n10332 0.0225448
R44127 vdd.n10348 vdd.n10347 0.0225448
R44128 vdd.n10349 vdd.n10348 0.0225448
R44129 vdd.n10345 vdd.n10344 0.0225448
R44130 vdd.n10341 vdd.n10340 0.0225448
R44131 vdd.n10342 vdd.n10341 0.0225448
R44132 vdd.n10351 vdd.n10350 0.0225448
R44133 vdd.n10350 vdd.n10349 0.0225448
R44134 vdd.n10331 vdd.n10307 0.0225448
R44135 vdd.n10332 vdd.n10331 0.0225448
R44136 vdd.n10329 vdd.n10328 0.0225448
R44137 vdd.n10371 vdd.n10369 0.0225448
R44138 vdd.n10371 vdd.n10370 0.0225448
R44139 vdd.n10382 vdd.n10381 0.0225448
R44140 vdd.n10381 vdd.n10380 0.0225448
R44141 vdd.n10396 vdd.n10395 0.0225448
R44142 vdd.n10397 vdd.n10396 0.0225448
R44143 vdd.n10393 vdd.n10392 0.0225448
R44144 vdd.n10389 vdd.n10388 0.0225448
R44145 vdd.n10390 vdd.n10389 0.0225448
R44146 vdd.n10399 vdd.n10398 0.0225448
R44147 vdd.n10398 vdd.n10397 0.0225448
R44148 vdd.n10379 vdd.n10355 0.0225448
R44149 vdd.n10380 vdd.n10379 0.0225448
R44150 vdd.n10377 vdd.n10376 0.0225448
R44151 vdd.n10473 vdd.n10471 0.0225448
R44152 vdd.n10473 vdd.n10472 0.0225448
R44153 vdd.n10484 vdd.n10483 0.0225448
R44154 vdd.n10483 vdd.n10482 0.0225448
R44155 vdd.n10498 vdd.n10497 0.0225448
R44156 vdd.n10499 vdd.n10498 0.0225448
R44157 vdd.n10495 vdd.n10494 0.0225448
R44158 vdd.n10491 vdd.n10490 0.0225448
R44159 vdd.n10492 vdd.n10491 0.0225448
R44160 vdd.n10501 vdd.n10500 0.0225448
R44161 vdd.n10500 vdd.n10499 0.0225448
R44162 vdd.n10481 vdd.n10457 0.0225448
R44163 vdd.n10482 vdd.n10481 0.0225448
R44164 vdd.n10479 vdd.n10478 0.0225448
R44165 vdd.n65 vdd.n63 0.0225448
R44166 vdd.n65 vdd.n64 0.0225448
R44167 vdd.n76 vdd.n75 0.0225448
R44168 vdd.n75 vdd.n74 0.0225448
R44169 vdd.n90 vdd.n89 0.0225448
R44170 vdd.n91 vdd.n90 0.0225448
R44171 vdd.n87 vdd.n86 0.0225448
R44172 vdd.n83 vdd.n82 0.0225448
R44173 vdd.n84 vdd.n83 0.0225448
R44174 vdd.n93 vdd.n92 0.0225448
R44175 vdd.n92 vdd.n91 0.0225448
R44176 vdd.n73 vdd.n49 0.0225448
R44177 vdd.n74 vdd.n73 0.0225448
R44178 vdd.n71 vdd.n70 0.0225448
R44179 vdd.n17 vdd.n15 0.0225448
R44180 vdd.n17 vdd.n16 0.0225448
R44181 vdd.n28 vdd.n27 0.0225448
R44182 vdd.n27 vdd.n26 0.0225448
R44183 vdd.n42 vdd.n41 0.0225448
R44184 vdd.n43 vdd.n42 0.0225448
R44185 vdd.n39 vdd.n38 0.0225448
R44186 vdd.n35 vdd.n34 0.0225448
R44187 vdd.n36 vdd.n35 0.0225448
R44188 vdd.n45 vdd.n44 0.0225448
R44189 vdd.n44 vdd.n43 0.0225448
R44190 vdd.n25 vdd.n1 0.0225448
R44191 vdd.n26 vdd.n25 0.0225448
R44192 vdd.n23 vdd.n22 0.0225448
R44193 vdd.n10521 vdd.n10519 0.0225448
R44194 vdd.n10521 vdd.n10520 0.0225448
R44195 vdd.n10532 vdd.n10531 0.0225448
R44196 vdd.n10531 vdd.n10530 0.0225448
R44197 vdd.n10546 vdd.n10545 0.0225448
R44198 vdd.n10547 vdd.n10546 0.0225448
R44199 vdd.n10543 vdd.n10542 0.0225448
R44200 vdd.n10539 vdd.n10538 0.0225448
R44201 vdd.n10540 vdd.n10539 0.0225448
R44202 vdd.n10549 vdd.n10548 0.0225448
R44203 vdd.n10548 vdd.n10547 0.0225448
R44204 vdd.n10529 vdd.n10505 0.0225448
R44205 vdd.n10530 vdd.n10529 0.0225448
R44206 vdd.n10527 vdd.n10526 0.0225448
R44207 vdd.n10571 vdd.n10569 0.0225448
R44208 vdd.n10571 vdd.n10570 0.0225448
R44209 vdd.n10582 vdd.n10581 0.0225448
R44210 vdd.n10581 vdd.n10580 0.0225448
R44211 vdd.n10596 vdd.n10595 0.0225448
R44212 vdd.n10597 vdd.n10596 0.0225448
R44213 vdd.n10593 vdd.n10592 0.0225448
R44214 vdd.n10589 vdd.n10588 0.0225448
R44215 vdd.n10590 vdd.n10589 0.0225448
R44216 vdd.n10599 vdd.n10598 0.0225448
R44217 vdd.n10598 vdd.n10597 0.0225448
R44218 vdd.n10579 vdd.n10555 0.0225448
R44219 vdd.n10580 vdd.n10579 0.0225448
R44220 vdd.n10577 vdd.n10576 0.0225448
R44221 vdd.n10619 vdd.n10617 0.0225448
R44222 vdd.n10619 vdd.n10618 0.0225448
R44223 vdd.n10630 vdd.n10629 0.0225448
R44224 vdd.n10629 vdd.n10628 0.0225448
R44225 vdd.n10644 vdd.n10643 0.0225448
R44226 vdd.n10645 vdd.n10644 0.0225448
R44227 vdd.n10641 vdd.n10640 0.0225448
R44228 vdd.n10637 vdd.n10636 0.0225448
R44229 vdd.n10638 vdd.n10637 0.0225448
R44230 vdd.n10647 vdd.n10646 0.0225448
R44231 vdd.n10646 vdd.n10645 0.0225448
R44232 vdd.n10627 vdd.n10603 0.0225448
R44233 vdd.n10628 vdd.n10627 0.0225448
R44234 vdd.n10625 vdd.n10624 0.0225448
R44235 vdd.n10424 vdd.n10423 0.0225448
R44236 vdd.n10425 vdd.n10424 0.0225448
R44237 vdd.n10421 vdd.n10414 0.0225448
R44238 vdd.n10432 vdd.n10414 0.0225448
R44239 vdd.n10434 vdd.n10433 0.0225448
R44240 vdd.n10435 vdd.n10434 0.0225448
R44241 vdd.n10449 vdd.n10448 0.0225448
R44242 vdd.n10445 vdd.n10404 0.0225448
R44243 vdd.n10446 vdd.n10445 0.0225448
R44244 vdd.n10440 vdd.n10409 0.0225448
R44245 vdd.n10435 vdd.n10409 0.0225448
R44246 vdd.n10431 vdd.n10430 0.0225448
R44247 vdd.n10432 vdd.n10431 0.0225448
R44248 vdd.n10428 vdd.n10427 0.0225448
R44249 vdd.n10767 vdd.n10765 0.0225448
R44250 vdd.n10767 vdd.n10766 0.0225448
R44251 vdd.n10778 vdd.n10777 0.0225448
R44252 vdd.n10777 vdd.n10776 0.0225448
R44253 vdd.n10792 vdd.n10791 0.0225448
R44254 vdd.n10793 vdd.n10792 0.0225448
R44255 vdd.n10789 vdd.n10788 0.0225448
R44256 vdd.n10785 vdd.n10784 0.0225448
R44257 vdd.n10786 vdd.n10785 0.0225448
R44258 vdd.n10795 vdd.n10794 0.0225448
R44259 vdd.n10794 vdd.n10793 0.0225448
R44260 vdd.n10775 vdd.n10751 0.0225448
R44261 vdd.n10776 vdd.n10775 0.0225448
R44262 vdd.n10773 vdd.n10772 0.0225448
R44263 vdd.n10718 vdd.n10716 0.0225448
R44264 vdd.n10718 vdd.n10717 0.0225448
R44265 vdd.n10729 vdd.n10728 0.0225448
R44266 vdd.n10728 vdd.n10727 0.0225448
R44267 vdd.n10743 vdd.n10742 0.0225448
R44268 vdd.n10744 vdd.n10743 0.0225448
R44269 vdd.n10740 vdd.n10739 0.0225448
R44270 vdd.n10736 vdd.n10735 0.0225448
R44271 vdd.n10737 vdd.n10736 0.0225448
R44272 vdd.n10746 vdd.n10745 0.0225448
R44273 vdd.n10745 vdd.n10744 0.0225448
R44274 vdd.n10726 vdd.n10702 0.0225448
R44275 vdd.n10727 vdd.n10726 0.0225448
R44276 vdd.n10724 vdd.n10723 0.0225448
R44277 vdd.n10670 vdd.n10668 0.0225448
R44278 vdd.n10670 vdd.n10669 0.0225448
R44279 vdd.n10681 vdd.n10680 0.0225448
R44280 vdd.n10680 vdd.n10679 0.0225448
R44281 vdd.n10695 vdd.n10694 0.0225448
R44282 vdd.n10696 vdd.n10695 0.0225448
R44283 vdd.n10692 vdd.n10691 0.0225448
R44284 vdd.n10688 vdd.n10687 0.0225448
R44285 vdd.n10689 vdd.n10688 0.0225448
R44286 vdd.n10698 vdd.n10697 0.0225448
R44287 vdd.n10697 vdd.n10696 0.0225448
R44288 vdd.n10678 vdd.n10654 0.0225448
R44289 vdd.n10679 vdd.n10678 0.0225448
R44290 vdd.n10676 vdd.n10675 0.0225448
R44291 vdd.n10816 vdd.n10814 0.0225448
R44292 vdd.n10816 vdd.n10815 0.0225448
R44293 vdd.n10827 vdd.n10826 0.0225448
R44294 vdd.n10826 vdd.n10825 0.0225448
R44295 vdd.n10841 vdd.n10840 0.0225448
R44296 vdd.n10842 vdd.n10841 0.0225448
R44297 vdd.n10838 vdd.n10837 0.0225448
R44298 vdd.n10834 vdd.n10833 0.0225448
R44299 vdd.n10835 vdd.n10834 0.0225448
R44300 vdd.n10844 vdd.n10843 0.0225448
R44301 vdd.n10843 vdd.n10842 0.0225448
R44302 vdd.n10824 vdd.n10800 0.0225448
R44303 vdd.n10825 vdd.n10824 0.0225448
R44304 vdd.n10822 vdd.n10821 0.0225448
R44305 vdd.n10866 vdd.n10864 0.0225448
R44306 vdd.n10866 vdd.n10865 0.0225448
R44307 vdd.n10877 vdd.n10876 0.0225448
R44308 vdd.n10876 vdd.n10875 0.0225448
R44309 vdd.n10891 vdd.n10890 0.0225448
R44310 vdd.n10892 vdd.n10891 0.0225448
R44311 vdd.n10888 vdd.n10887 0.0225448
R44312 vdd.n10884 vdd.n10883 0.0225448
R44313 vdd.n10885 vdd.n10884 0.0225448
R44314 vdd.n10894 vdd.n10893 0.0225448
R44315 vdd.n10893 vdd.n10892 0.0225448
R44316 vdd.n10874 vdd.n10850 0.0225448
R44317 vdd.n10875 vdd.n10874 0.0225448
R44318 vdd.n10872 vdd.n10871 0.0225448
R44319 vdd.n10914 vdd.n10912 0.0225448
R44320 vdd.n10914 vdd.n10913 0.0225448
R44321 vdd.n10925 vdd.n10924 0.0225448
R44322 vdd.n10924 vdd.n10923 0.0225448
R44323 vdd.n10939 vdd.n10938 0.0225448
R44324 vdd.n10940 vdd.n10939 0.0225448
R44325 vdd.n10936 vdd.n10935 0.0225448
R44326 vdd.n10932 vdd.n10931 0.0225448
R44327 vdd.n10933 vdd.n10932 0.0225448
R44328 vdd.n10942 vdd.n10941 0.0225448
R44329 vdd.n10941 vdd.n10940 0.0225448
R44330 vdd.n10922 vdd.n10898 0.0225448
R44331 vdd.n10923 vdd.n10922 0.0225448
R44332 vdd.n10920 vdd.n10919 0.0225448
R44333 vdd.n11012 vdd.n11010 0.0225448
R44334 vdd.n11012 vdd.n11011 0.0225448
R44335 vdd.n11023 vdd.n11022 0.0225448
R44336 vdd.n11022 vdd.n11021 0.0225448
R44337 vdd.n11037 vdd.n11036 0.0225448
R44338 vdd.n11038 vdd.n11037 0.0225448
R44339 vdd.n11034 vdd.n11033 0.0225448
R44340 vdd.n11030 vdd.n11029 0.0225448
R44341 vdd.n11031 vdd.n11030 0.0225448
R44342 vdd.n11040 vdd.n11039 0.0225448
R44343 vdd.n11039 vdd.n11038 0.0225448
R44344 vdd.n11020 vdd.n10996 0.0225448
R44345 vdd.n11021 vdd.n11020 0.0225448
R44346 vdd.n11018 vdd.n11017 0.0225448
R44347 vdd.n10964 vdd.n10962 0.0225448
R44348 vdd.n10964 vdd.n10963 0.0225448
R44349 vdd.n10975 vdd.n10974 0.0225448
R44350 vdd.n10974 vdd.n10973 0.0225448
R44351 vdd.n10989 vdd.n10988 0.0225448
R44352 vdd.n10990 vdd.n10989 0.0225448
R44353 vdd.n10986 vdd.n10985 0.0225448
R44354 vdd.n10982 vdd.n10981 0.0225448
R44355 vdd.n10983 vdd.n10982 0.0225448
R44356 vdd.n10992 vdd.n10991 0.0225448
R44357 vdd.n10991 vdd.n10990 0.0225448
R44358 vdd.n10972 vdd.n10948 0.0225448
R44359 vdd.n10973 vdd.n10972 0.0225448
R44360 vdd.n10970 vdd.n10969 0.0225448
R44361 vdd.n11061 vdd.n11059 0.0225448
R44362 vdd.n11061 vdd.n11060 0.0225448
R44363 vdd.n11072 vdd.n11071 0.0225448
R44364 vdd.n11071 vdd.n11070 0.0225448
R44365 vdd.n11086 vdd.n11085 0.0225448
R44366 vdd.n11087 vdd.n11086 0.0225448
R44367 vdd.n11083 vdd.n11082 0.0225448
R44368 vdd.n11079 vdd.n11078 0.0225448
R44369 vdd.n11080 vdd.n11079 0.0225448
R44370 vdd.n11089 vdd.n11088 0.0225448
R44371 vdd.n11088 vdd.n11087 0.0225448
R44372 vdd.n11069 vdd.n11045 0.0225448
R44373 vdd.n11070 vdd.n11069 0.0225448
R44374 vdd.n11067 vdd.n11066 0.0225448
R44375 vdd.n11111 vdd.n11109 0.0225448
R44376 vdd.n11111 vdd.n11110 0.0225448
R44377 vdd.n11122 vdd.n11121 0.0225448
R44378 vdd.n11121 vdd.n11120 0.0225448
R44379 vdd.n11136 vdd.n11135 0.0225448
R44380 vdd.n11137 vdd.n11136 0.0225448
R44381 vdd.n11133 vdd.n11132 0.0225448
R44382 vdd.n11129 vdd.n11128 0.0225448
R44383 vdd.n11130 vdd.n11129 0.0225448
R44384 vdd.n11139 vdd.n11138 0.0225448
R44385 vdd.n11138 vdd.n11137 0.0225448
R44386 vdd.n11119 vdd.n11095 0.0225448
R44387 vdd.n11120 vdd.n11119 0.0225448
R44388 vdd.n11117 vdd.n11116 0.0225448
R44389 vdd.n11159 vdd.n11157 0.0225448
R44390 vdd.n11159 vdd.n11158 0.0225448
R44391 vdd.n11170 vdd.n11169 0.0225448
R44392 vdd.n11169 vdd.n11168 0.0225448
R44393 vdd.n11184 vdd.n11183 0.0225448
R44394 vdd.n11185 vdd.n11184 0.0225448
R44395 vdd.n11181 vdd.n11180 0.0225448
R44396 vdd.n11177 vdd.n11176 0.0225448
R44397 vdd.n11178 vdd.n11177 0.0225448
R44398 vdd.n11187 vdd.n11186 0.0225448
R44399 vdd.n11186 vdd.n11185 0.0225448
R44400 vdd.n11167 vdd.n11143 0.0225448
R44401 vdd.n11168 vdd.n11167 0.0225448
R44402 vdd.n11165 vdd.n11164 0.0225448
R44403 vdd.n10178 vdd.n10177 0.0225448
R44404 vdd.n10179 vdd.n10178 0.0225448
R44405 vdd.n10175 vdd.n10168 0.0225448
R44406 vdd.n10186 vdd.n10168 0.0225448
R44407 vdd.n10188 vdd.n10187 0.0225448
R44408 vdd.n10189 vdd.n10188 0.0225448
R44409 vdd.n10203 vdd.n10202 0.0225448
R44410 vdd.n10199 vdd.n10158 0.0225448
R44411 vdd.n10200 vdd.n10199 0.0225448
R44412 vdd.n10194 vdd.n10163 0.0225448
R44413 vdd.n10189 vdd.n10163 0.0225448
R44414 vdd.n10185 vdd.n10184 0.0225448
R44415 vdd.n10186 vdd.n10185 0.0225448
R44416 vdd.n10182 vdd.n10181 0.0225448
R44417 vdd.n11258 vdd.n11256 0.0225448
R44418 vdd.n11258 vdd.n11257 0.0225448
R44419 vdd.n11269 vdd.n11268 0.0225448
R44420 vdd.n11268 vdd.n11267 0.0225448
R44421 vdd.n11283 vdd.n11282 0.0225448
R44422 vdd.n11284 vdd.n11283 0.0225448
R44423 vdd.n11280 vdd.n11279 0.0225448
R44424 vdd.n11276 vdd.n11275 0.0225448
R44425 vdd.n11277 vdd.n11276 0.0225448
R44426 vdd.n11286 vdd.n11285 0.0225448
R44427 vdd.n11285 vdd.n11284 0.0225448
R44428 vdd.n11266 vdd.n11242 0.0225448
R44429 vdd.n11267 vdd.n11266 0.0225448
R44430 vdd.n11264 vdd.n11263 0.0225448
R44431 vdd.n11210 vdd.n11208 0.0225448
R44432 vdd.n11210 vdd.n11209 0.0225448
R44433 vdd.n11221 vdd.n11220 0.0225448
R44434 vdd.n11220 vdd.n11219 0.0225448
R44435 vdd.n11235 vdd.n11234 0.0225448
R44436 vdd.n11236 vdd.n11235 0.0225448
R44437 vdd.n11232 vdd.n11231 0.0225448
R44438 vdd.n11228 vdd.n11227 0.0225448
R44439 vdd.n11229 vdd.n11228 0.0225448
R44440 vdd.n11238 vdd.n11237 0.0225448
R44441 vdd.n11237 vdd.n11236 0.0225448
R44442 vdd.n11218 vdd.n11194 0.0225448
R44443 vdd.n11219 vdd.n11218 0.0225448
R44444 vdd.n11216 vdd.n11215 0.0225448
R44445 vdd.n11307 vdd.n11305 0.0225448
R44446 vdd.n11307 vdd.n11306 0.0225448
R44447 vdd.n11318 vdd.n11317 0.0225448
R44448 vdd.n11317 vdd.n11316 0.0225448
R44449 vdd.n11332 vdd.n11331 0.0225448
R44450 vdd.n11333 vdd.n11332 0.0225448
R44451 vdd.n11329 vdd.n11328 0.0225448
R44452 vdd.n11325 vdd.n11324 0.0225448
R44453 vdd.n11326 vdd.n11325 0.0225448
R44454 vdd.n11335 vdd.n11334 0.0225448
R44455 vdd.n11334 vdd.n11333 0.0225448
R44456 vdd.n11315 vdd.n11291 0.0225448
R44457 vdd.n11316 vdd.n11315 0.0225448
R44458 vdd.n11313 vdd.n11312 0.0225448
R44459 vdd.n11357 vdd.n11355 0.0225448
R44460 vdd.n11357 vdd.n11356 0.0225448
R44461 vdd.n11368 vdd.n11367 0.0225448
R44462 vdd.n11367 vdd.n11366 0.0225448
R44463 vdd.n11382 vdd.n11381 0.0225448
R44464 vdd.n11383 vdd.n11382 0.0225448
R44465 vdd.n11379 vdd.n11378 0.0225448
R44466 vdd.n11375 vdd.n11374 0.0225448
R44467 vdd.n11376 vdd.n11375 0.0225448
R44468 vdd.n11385 vdd.n11384 0.0225448
R44469 vdd.n11384 vdd.n11383 0.0225448
R44470 vdd.n11365 vdd.n11341 0.0225448
R44471 vdd.n11366 vdd.n11365 0.0225448
R44472 vdd.n11363 vdd.n11362 0.0225448
R44473 vdd.n11405 vdd.n11403 0.0225448
R44474 vdd.n11405 vdd.n11404 0.0225448
R44475 vdd.n11416 vdd.n11415 0.0225448
R44476 vdd.n11415 vdd.n11414 0.0225448
R44477 vdd.n11430 vdd.n11429 0.0225448
R44478 vdd.n11431 vdd.n11430 0.0225448
R44479 vdd.n11427 vdd.n11426 0.0225448
R44480 vdd.n11423 vdd.n11422 0.0225448
R44481 vdd.n11424 vdd.n11423 0.0225448
R44482 vdd.n11433 vdd.n11432 0.0225448
R44483 vdd.n11432 vdd.n11431 0.0225448
R44484 vdd.n11413 vdd.n11389 0.0225448
R44485 vdd.n11414 vdd.n11413 0.0225448
R44486 vdd.n11411 vdd.n11410 0.0225448
R44487 vdd.n11459 vdd.n11458 0.0225448
R44488 vdd.n11467 vdd.n11466 0.0225448
R44489 vdd.n11466 vdd.n11465 0.0225448
R44490 vdd.n11481 vdd.n11480 0.0225448
R44491 vdd.n11482 vdd.n11481 0.0225448
R44492 vdd.n11478 vdd.n11477 0.0225448
R44493 vdd.n11477 vdd.n11476 0.0225448
R44494 vdd.n11474 vdd.n11473 0.0225448
R44495 vdd.n11484 vdd.n11483 0.0225448
R44496 vdd.n11483 vdd.n11482 0.0225448
R44497 vdd.n11464 vdd.n11440 0.0225448
R44498 vdd.n11465 vdd.n11464 0.0225448
R44499 vdd.n11462 vdd.n11456 0.0225448
R44500 vdd.n11462 vdd.n11461 0.0225448
R44501 vdd.n11506 vdd.n11505 0.0225448
R44502 vdd.n11514 vdd.n11513 0.0225448
R44503 vdd.n11513 vdd.n11512 0.0225448
R44504 vdd.n11528 vdd.n11527 0.0225448
R44505 vdd.n11529 vdd.n11528 0.0225448
R44506 vdd.n11525 vdd.n11524 0.0225448
R44507 vdd.n11524 vdd.n11523 0.0225448
R44508 vdd.n11521 vdd.n11520 0.0225448
R44509 vdd.n11531 vdd.n11530 0.0225448
R44510 vdd.n11530 vdd.n11529 0.0225448
R44511 vdd.n11511 vdd.n11487 0.0225448
R44512 vdd.n11512 vdd.n11511 0.0225448
R44513 vdd.n11509 vdd.n11503 0.0225448
R44514 vdd.n11509 vdd.n11508 0.0225448
R44515 vdd.n11556 vdd.n11555 0.0225448
R44516 vdd.n11564 vdd.n11563 0.0225448
R44517 vdd.n11563 vdd.n11562 0.0225448
R44518 vdd.n11578 vdd.n11577 0.0225448
R44519 vdd.n11579 vdd.n11578 0.0225448
R44520 vdd.n11575 vdd.n11574 0.0225448
R44521 vdd.n11574 vdd.n11573 0.0225448
R44522 vdd.n11571 vdd.n11570 0.0225448
R44523 vdd.n11581 vdd.n11580 0.0225448
R44524 vdd.n11580 vdd.n11579 0.0225448
R44525 vdd.n11561 vdd.n11537 0.0225448
R44526 vdd.n11562 vdd.n11561 0.0225448
R44527 vdd.n11559 vdd.n11553 0.0225448
R44528 vdd.n11559 vdd.n11558 0.0225448
R44529 vdd.n11606 vdd.n11605 0.0225448
R44530 vdd.n11614 vdd.n11613 0.0225448
R44531 vdd.n11613 vdd.n11612 0.0225448
R44532 vdd.n11628 vdd.n11627 0.0225448
R44533 vdd.n11629 vdd.n11628 0.0225448
R44534 vdd.n11625 vdd.n11624 0.0225448
R44535 vdd.n11624 vdd.n11623 0.0225448
R44536 vdd.n11621 vdd.n11620 0.0225448
R44537 vdd.n11631 vdd.n11630 0.0225448
R44538 vdd.n11630 vdd.n11629 0.0225448
R44539 vdd.n11611 vdd.n11587 0.0225448
R44540 vdd.n11612 vdd.n11611 0.0225448
R44541 vdd.n11609 vdd.n11603 0.0225448
R44542 vdd.n11609 vdd.n11608 0.0225448
R44543 vdd.n11654 vdd.n11653 0.0225448
R44544 vdd.n11662 vdd.n11661 0.0225448
R44545 vdd.n11661 vdd.n11660 0.0225448
R44546 vdd.n11676 vdd.n11675 0.0225448
R44547 vdd.n11677 vdd.n11676 0.0225448
R44548 vdd.n11673 vdd.n11672 0.0225448
R44549 vdd.n11672 vdd.n11671 0.0225448
R44550 vdd.n11669 vdd.n11668 0.0225448
R44551 vdd.n11679 vdd.n11678 0.0225448
R44552 vdd.n11678 vdd.n11677 0.0225448
R44553 vdd.n11659 vdd.n11635 0.0225448
R44554 vdd.n11660 vdd.n11659 0.0225448
R44555 vdd.n11657 vdd.n11651 0.0225448
R44556 vdd.n11657 vdd.n11656 0.0225448
R44557 vdd.n482 vdd.n481 0.0225448
R44558 vdd.n479 vdd.n478 0.0225448
R44559 vdd.n478 vdd.n477 0.0225448
R44560 vdd.n468 vdd.n467 0.0225448
R44561 vdd.n469 vdd.n468 0.0225448
R44562 vdd.n465 vdd.n464 0.0225448
R44563 vdd.n464 vdd.n463 0.0225448
R44564 vdd.n461 vdd.n460 0.0225448
R44565 vdd.n470 vdd.n452 0.0225448
R44566 vdd.n470 vdd.n469 0.0225448
R44567 vdd.n476 vdd.n475 0.0225448
R44568 vdd.n477 vdd.n476 0.0225448
R44569 vdd.n486 vdd.n485 0.0225448
R44570 vdd.n485 vdd.n484 0.0225448
R44571 vdd.n11705 vdd.n11704 0.0225448
R44572 vdd.n11713 vdd.n11712 0.0225448
R44573 vdd.n11712 vdd.n11711 0.0225448
R44574 vdd.n11727 vdd.n11726 0.0225448
R44575 vdd.n11728 vdd.n11727 0.0225448
R44576 vdd.n11724 vdd.n11723 0.0225448
R44577 vdd.n11723 vdd.n11722 0.0225448
R44578 vdd.n11720 vdd.n11719 0.0225448
R44579 vdd.n11730 vdd.n11729 0.0225448
R44580 vdd.n11729 vdd.n11728 0.0225448
R44581 vdd.n11710 vdd.n11686 0.0225448
R44582 vdd.n11711 vdd.n11710 0.0225448
R44583 vdd.n11708 vdd.n11702 0.0225448
R44584 vdd.n11708 vdd.n11707 0.0225448
R44585 vdd.n11752 vdd.n11751 0.0225448
R44586 vdd.n11760 vdd.n11759 0.0225448
R44587 vdd.n11759 vdd.n11758 0.0225448
R44588 vdd.n11774 vdd.n11773 0.0225448
R44589 vdd.n11775 vdd.n11774 0.0225448
R44590 vdd.n11771 vdd.n11770 0.0225448
R44591 vdd.n11770 vdd.n11769 0.0225448
R44592 vdd.n11767 vdd.n11766 0.0225448
R44593 vdd.n11777 vdd.n11776 0.0225448
R44594 vdd.n11776 vdd.n11775 0.0225448
R44595 vdd.n11757 vdd.n11733 0.0225448
R44596 vdd.n11758 vdd.n11757 0.0225448
R44597 vdd.n11755 vdd.n11749 0.0225448
R44598 vdd.n11755 vdd.n11754 0.0225448
R44599 vdd.n11800 vdd.n11799 0.0225448
R44600 vdd.n11808 vdd.n11807 0.0225448
R44601 vdd.n11807 vdd.n11806 0.0225448
R44602 vdd.n11822 vdd.n11821 0.0225448
R44603 vdd.n11823 vdd.n11822 0.0225448
R44604 vdd.n11819 vdd.n11818 0.0225448
R44605 vdd.n11818 vdd.n11817 0.0225448
R44606 vdd.n11815 vdd.n11814 0.0225448
R44607 vdd.n11825 vdd.n11824 0.0225448
R44608 vdd.n11824 vdd.n11823 0.0225448
R44609 vdd.n11805 vdd.n11781 0.0225448
R44610 vdd.n11806 vdd.n11805 0.0225448
R44611 vdd.n11803 vdd.n11797 0.0225448
R44612 vdd.n11803 vdd.n11802 0.0225448
R44613 vdd.n11851 vdd.n11850 0.0225448
R44614 vdd.n11859 vdd.n11858 0.0225448
R44615 vdd.n11858 vdd.n11857 0.0225448
R44616 vdd.n11873 vdd.n11872 0.0225448
R44617 vdd.n11874 vdd.n11873 0.0225448
R44618 vdd.n11870 vdd.n11869 0.0225448
R44619 vdd.n11869 vdd.n11868 0.0225448
R44620 vdd.n11866 vdd.n11865 0.0225448
R44621 vdd.n11876 vdd.n11875 0.0225448
R44622 vdd.n11875 vdd.n11874 0.0225448
R44623 vdd.n11856 vdd.n11832 0.0225448
R44624 vdd.n11857 vdd.n11856 0.0225448
R44625 vdd.n11854 vdd.n11848 0.0225448
R44626 vdd.n11854 vdd.n11853 0.0225448
R44627 vdd.n11901 vdd.n11900 0.0225448
R44628 vdd.n11909 vdd.n11908 0.0225448
R44629 vdd.n11908 vdd.n11907 0.0225448
R44630 vdd.n11923 vdd.n11922 0.0225448
R44631 vdd.n11924 vdd.n11923 0.0225448
R44632 vdd.n11920 vdd.n11919 0.0225448
R44633 vdd.n11919 vdd.n11918 0.0225448
R44634 vdd.n11916 vdd.n11915 0.0225448
R44635 vdd.n11926 vdd.n11925 0.0225448
R44636 vdd.n11925 vdd.n11924 0.0225448
R44637 vdd.n11906 vdd.n11882 0.0225448
R44638 vdd.n11907 vdd.n11906 0.0225448
R44639 vdd.n11904 vdd.n11898 0.0225448
R44640 vdd.n11904 vdd.n11903 0.0225448
R44641 vdd.n11949 vdd.n11948 0.0225448
R44642 vdd.n11957 vdd.n11956 0.0225448
R44643 vdd.n11956 vdd.n11955 0.0225448
R44644 vdd.n11971 vdd.n11970 0.0225448
R44645 vdd.n11972 vdd.n11971 0.0225448
R44646 vdd.n11968 vdd.n11967 0.0225448
R44647 vdd.n11967 vdd.n11966 0.0225448
R44648 vdd.n11964 vdd.n11963 0.0225448
R44649 vdd.n11974 vdd.n11973 0.0225448
R44650 vdd.n11973 vdd.n11972 0.0225448
R44651 vdd.n11954 vdd.n11930 0.0225448
R44652 vdd.n11955 vdd.n11954 0.0225448
R44653 vdd.n11952 vdd.n11946 0.0225448
R44654 vdd.n11952 vdd.n11951 0.0225448
R44655 vdd.n11999 vdd.n11998 0.0225448
R44656 vdd.n12007 vdd.n12006 0.0225448
R44657 vdd.n12006 vdd.n12005 0.0225448
R44658 vdd.n12021 vdd.n12020 0.0225448
R44659 vdd.n12022 vdd.n12021 0.0225448
R44660 vdd.n12018 vdd.n12017 0.0225448
R44661 vdd.n12017 vdd.n12016 0.0225448
R44662 vdd.n12014 vdd.n12013 0.0225448
R44663 vdd.n12024 vdd.n12023 0.0225448
R44664 vdd.n12023 vdd.n12022 0.0225448
R44665 vdd.n12004 vdd.n11980 0.0225448
R44666 vdd.n12005 vdd.n12004 0.0225448
R44667 vdd.n12002 vdd.n11996 0.0225448
R44668 vdd.n12002 vdd.n12001 0.0225448
R44669 vdd.n12046 vdd.n12045 0.0225448
R44670 vdd.n12054 vdd.n12053 0.0225448
R44671 vdd.n12053 vdd.n12052 0.0225448
R44672 vdd.n12068 vdd.n12067 0.0225448
R44673 vdd.n12069 vdd.n12068 0.0225448
R44674 vdd.n12065 vdd.n12064 0.0225448
R44675 vdd.n12064 vdd.n12063 0.0225448
R44676 vdd.n12061 vdd.n12060 0.0225448
R44677 vdd.n12071 vdd.n12070 0.0225448
R44678 vdd.n12070 vdd.n12069 0.0225448
R44679 vdd.n12051 vdd.n12027 0.0225448
R44680 vdd.n12052 vdd.n12051 0.0225448
R44681 vdd.n12049 vdd.n12043 0.0225448
R44682 vdd.n12049 vdd.n12048 0.0225448
R44683 vdd.n12096 vdd.n12095 0.0225448
R44684 vdd.n12104 vdd.n12103 0.0225448
R44685 vdd.n12103 vdd.n12102 0.0225448
R44686 vdd.n12118 vdd.n12117 0.0225448
R44687 vdd.n12119 vdd.n12118 0.0225448
R44688 vdd.n12115 vdd.n12114 0.0225448
R44689 vdd.n12114 vdd.n12113 0.0225448
R44690 vdd.n12111 vdd.n12110 0.0225448
R44691 vdd.n12121 vdd.n12120 0.0225448
R44692 vdd.n12120 vdd.n12119 0.0225448
R44693 vdd.n12101 vdd.n12077 0.0225448
R44694 vdd.n12102 vdd.n12101 0.0225448
R44695 vdd.n12099 vdd.n12093 0.0225448
R44696 vdd.n12099 vdd.n12098 0.0225448
R44697 vdd.n12146 vdd.n12145 0.0225448
R44698 vdd.n12154 vdd.n12153 0.0225448
R44699 vdd.n12153 vdd.n12152 0.0225448
R44700 vdd.n12168 vdd.n12167 0.0225448
R44701 vdd.n12169 vdd.n12168 0.0225448
R44702 vdd.n12165 vdd.n12164 0.0225448
R44703 vdd.n12164 vdd.n12163 0.0225448
R44704 vdd.n12161 vdd.n12160 0.0225448
R44705 vdd.n12171 vdd.n12170 0.0225448
R44706 vdd.n12170 vdd.n12169 0.0225448
R44707 vdd.n12151 vdd.n12127 0.0225448
R44708 vdd.n12152 vdd.n12151 0.0225448
R44709 vdd.n12149 vdd.n12143 0.0225448
R44710 vdd.n12149 vdd.n12148 0.0225448
R44711 vdd.n12194 vdd.n12193 0.0225448
R44712 vdd.n12202 vdd.n12201 0.0225448
R44713 vdd.n12201 vdd.n12200 0.0225448
R44714 vdd.n12216 vdd.n12215 0.0225448
R44715 vdd.n12217 vdd.n12216 0.0225448
R44716 vdd.n12213 vdd.n12212 0.0225448
R44717 vdd.n12212 vdd.n12211 0.0225448
R44718 vdd.n12209 vdd.n12208 0.0225448
R44719 vdd.n12219 vdd.n12218 0.0225448
R44720 vdd.n12218 vdd.n12217 0.0225448
R44721 vdd.n12199 vdd.n12175 0.0225448
R44722 vdd.n12200 vdd.n12199 0.0225448
R44723 vdd.n12197 vdd.n12191 0.0225448
R44724 vdd.n12197 vdd.n12196 0.0225448
R44725 vdd.n237 vdd.n236 0.0225448
R44726 vdd.n234 vdd.n233 0.0225448
R44727 vdd.n233 vdd.n232 0.0225448
R44728 vdd.n223 vdd.n222 0.0225448
R44729 vdd.n224 vdd.n223 0.0225448
R44730 vdd.n220 vdd.n219 0.0225448
R44731 vdd.n219 vdd.n218 0.0225448
R44732 vdd.n216 vdd.n215 0.0225448
R44733 vdd.n225 vdd.n207 0.0225448
R44734 vdd.n225 vdd.n224 0.0225448
R44735 vdd.n231 vdd.n230 0.0225448
R44736 vdd.n232 vdd.n231 0.0225448
R44737 vdd.n241 vdd.n240 0.0225448
R44738 vdd.n240 vdd.n239 0.0225448
R44739 vdd.n12245 vdd.n12244 0.0225448
R44740 vdd.n12253 vdd.n12252 0.0225448
R44741 vdd.n12252 vdd.n12251 0.0225448
R44742 vdd.n12267 vdd.n12266 0.0225448
R44743 vdd.n12268 vdd.n12267 0.0225448
R44744 vdd.n12264 vdd.n12263 0.0225448
R44745 vdd.n12263 vdd.n12262 0.0225448
R44746 vdd.n12260 vdd.n12259 0.0225448
R44747 vdd.n12270 vdd.n12269 0.0225448
R44748 vdd.n12269 vdd.n12268 0.0225448
R44749 vdd.n12250 vdd.n12226 0.0225448
R44750 vdd.n12251 vdd.n12250 0.0225448
R44751 vdd.n12248 vdd.n12242 0.0225448
R44752 vdd.n12248 vdd.n12247 0.0225448
R44753 vdd.n12292 vdd.n12291 0.0225448
R44754 vdd.n12300 vdd.n12299 0.0225448
R44755 vdd.n12299 vdd.n12298 0.0225448
R44756 vdd.n12314 vdd.n12313 0.0225448
R44757 vdd.n12315 vdd.n12314 0.0225448
R44758 vdd.n12311 vdd.n12310 0.0225448
R44759 vdd.n12310 vdd.n12309 0.0225448
R44760 vdd.n12307 vdd.n12306 0.0225448
R44761 vdd.n12317 vdd.n12316 0.0225448
R44762 vdd.n12316 vdd.n12315 0.0225448
R44763 vdd.n12297 vdd.n12273 0.0225448
R44764 vdd.n12298 vdd.n12297 0.0225448
R44765 vdd.n12295 vdd.n12289 0.0225448
R44766 vdd.n12295 vdd.n12294 0.0225448
R44767 vdd.n12342 vdd.n12341 0.0225448
R44768 vdd.n12350 vdd.n12349 0.0225448
R44769 vdd.n12349 vdd.n12348 0.0225448
R44770 vdd.n12364 vdd.n12363 0.0225448
R44771 vdd.n12365 vdd.n12364 0.0225448
R44772 vdd.n12361 vdd.n12360 0.0225448
R44773 vdd.n12360 vdd.n12359 0.0225448
R44774 vdd.n12357 vdd.n12356 0.0225448
R44775 vdd.n12367 vdd.n12366 0.0225448
R44776 vdd.n12366 vdd.n12365 0.0225448
R44777 vdd.n12347 vdd.n12323 0.0225448
R44778 vdd.n12348 vdd.n12347 0.0225448
R44779 vdd.n12345 vdd.n12339 0.0225448
R44780 vdd.n12345 vdd.n12344 0.0225448
R44781 vdd.n12392 vdd.n12391 0.0225448
R44782 vdd.n12400 vdd.n12399 0.0225448
R44783 vdd.n12399 vdd.n12398 0.0225448
R44784 vdd.n12414 vdd.n12413 0.0225448
R44785 vdd.n12415 vdd.n12414 0.0225448
R44786 vdd.n12411 vdd.n12410 0.0225448
R44787 vdd.n12410 vdd.n12409 0.0225448
R44788 vdd.n12407 vdd.n12406 0.0225448
R44789 vdd.n12417 vdd.n12416 0.0225448
R44790 vdd.n12416 vdd.n12415 0.0225448
R44791 vdd.n12397 vdd.n12373 0.0225448
R44792 vdd.n12398 vdd.n12397 0.0225448
R44793 vdd.n12395 vdd.n12389 0.0225448
R44794 vdd.n12395 vdd.n12394 0.0225448
R44795 vdd.n12440 vdd.n12439 0.0225448
R44796 vdd.n12448 vdd.n12447 0.0225448
R44797 vdd.n12447 vdd.n12446 0.0225448
R44798 vdd.n12462 vdd.n12461 0.0225448
R44799 vdd.n12463 vdd.n12462 0.0225448
R44800 vdd.n12459 vdd.n12458 0.0225448
R44801 vdd.n12458 vdd.n12457 0.0225448
R44802 vdd.n12455 vdd.n12454 0.0225448
R44803 vdd.n12465 vdd.n12464 0.0225448
R44804 vdd.n12464 vdd.n12463 0.0225448
R44805 vdd.n12445 vdd.n12421 0.0225448
R44806 vdd.n12446 vdd.n12445 0.0225448
R44807 vdd.n12443 vdd.n12437 0.0225448
R44808 vdd.n12443 vdd.n12442 0.0225448
R44809 vdd vdd 0.0218816
R44810 vdd vdd 0.0218816
R44811 vdd vdd 0.0218816
R44812 vdd vdd 0.0218816
R44813 vdd vdd 0.0218816
R44814 vdd vdd 0.0218816
R44815 vdd.n7802 vdd.n7752 0.0216765
R44816 vdd.n7802 vdd.n7801 0.0216765
R44817 vdd.n7557 vdd.n7507 0.0216765
R44818 vdd.n7557 vdd.n7556 0.0216765
R44819 vdd.n7359 vdd.n7309 0.0216765
R44820 vdd.n7359 vdd.n7358 0.0216765
R44821 vdd.n7113 vdd.n7063 0.0216765
R44822 vdd.n7113 vdd.n7112 0.0216765
R44823 vdd.n4660 vdd.n4610 0.0216765
R44824 vdd.n4660 vdd.n4659 0.0216765
R44825 vdd.n4415 vdd.n4365 0.0216765
R44826 vdd.n4415 vdd.n4414 0.0216765
R44827 vdd.n4217 vdd.n4167 0.0216765
R44828 vdd.n4217 vdd.n4216 0.0216765
R44829 vdd.n3971 vdd.n3921 0.0216765
R44830 vdd.n3971 vdd.n3970 0.0216765
R44831 vdd.n1518 vdd.n1468 0.0216765
R44832 vdd.n1518 vdd.n1517 0.0216765
R44833 vdd.n1273 vdd.n1223 0.0216765
R44834 vdd.n1273 vdd.n1272 0.0216765
R44835 vdd.n1075 vdd.n1025 0.0216765
R44836 vdd.n1075 vdd.n1074 0.0216765
R44837 vdd.n829 vdd.n779 0.0216765
R44838 vdd.n829 vdd.n828 0.0216765
R44839 vdd.n10452 vdd.n10402 0.0216765
R44840 vdd.n10452 vdd.n10451 0.0216765
R44841 vdd.n10206 vdd.n10156 0.0216765
R44842 vdd.n10206 vdd.n10205 0.0216765
R44843 vdd.n488 vdd.n438 0.0216765
R44844 vdd.n488 vdd.n487 0.0216765
R44845 vdd.n243 vdd.n193 0.0216765
R44846 vdd.n243 vdd.n242 0.0216765
R44847 vdd.n118 vdd.n117 0.0196536
R44848 vdd.n166 vdd.n165 0.0196536
R44849 vdd.n267 vdd.n266 0.0196536
R44850 vdd.n315 vdd.n314 0.0196536
R44851 vdd.n363 vdd.n362 0.0196536
R44852 vdd.n411 vdd.n410 0.0196536
R44853 vdd.n512 vdd.n511 0.0196536
R44854 vdd.n560 vdd.n559 0.0196536
R44855 vdd.n7432 vdd.n7431 0.0196536
R44856 vdd.n7480 vdd.n7479 0.0196536
R44857 vdd.n7581 vdd.n7580 0.0196536
R44858 vdd.n7629 vdd.n7628 0.0196536
R44859 vdd.n7677 vdd.n7676 0.0196536
R44860 vdd.n7725 vdd.n7724 0.0196536
R44861 vdd.n7826 vdd.n7825 0.0196536
R44862 vdd.n6939 vdd.n6938 0.0196536
R44863 vdd.n7874 vdd.n7873 0.0196536
R44864 vdd.n7921 vdd.n7920 0.0196536
R44865 vdd.n7971 vdd.n7970 0.0196536
R44866 vdd.n8021 vdd.n8020 0.0196536
R44867 vdd.n8069 vdd.n8068 0.0196536
R44868 vdd.n7797 vdd.n7796 0.0196536
R44869 vdd.n8120 vdd.n8119 0.0196536
R44870 vdd.n8167 vdd.n8166 0.0196536
R44871 vdd.n8215 vdd.n8214 0.0196536
R44872 vdd.n8266 vdd.n8265 0.0196536
R44873 vdd.n8316 vdd.n8315 0.0196536
R44874 vdd.n8364 vdd.n8363 0.0196536
R44875 vdd.n8414 vdd.n8413 0.0196536
R44876 vdd.n8461 vdd.n8460 0.0196536
R44877 vdd.n8511 vdd.n8510 0.0196536
R44878 vdd.n8561 vdd.n8560 0.0196536
R44879 vdd.n8609 vdd.n8608 0.0196536
R44880 vdd.n7552 vdd.n7551 0.0196536
R44881 vdd.n8660 vdd.n8659 0.0196536
R44882 vdd.n8707 vdd.n8706 0.0196536
R44883 vdd.n8757 vdd.n8756 0.0196536
R44884 vdd.n8807 vdd.n8806 0.0196536
R44885 vdd.n8855 vdd.n8854 0.0196536
R44886 vdd.n4290 vdd.n4289 0.0196536
R44887 vdd.n4338 vdd.n4337 0.0196536
R44888 vdd.n4439 vdd.n4438 0.0196536
R44889 vdd.n4487 vdd.n4486 0.0196536
R44890 vdd.n4535 vdd.n4534 0.0196536
R44891 vdd.n4583 vdd.n4582 0.0196536
R44892 vdd.n4684 vdd.n4683 0.0196536
R44893 vdd.n3797 vdd.n3796 0.0196536
R44894 vdd.n4732 vdd.n4731 0.0196536
R44895 vdd.n4779 vdd.n4778 0.0196536
R44896 vdd.n4829 vdd.n4828 0.0196536
R44897 vdd.n4879 vdd.n4878 0.0196536
R44898 vdd.n4927 vdd.n4926 0.0196536
R44899 vdd.n4655 vdd.n4654 0.0196536
R44900 vdd.n4978 vdd.n4977 0.0196536
R44901 vdd.n5025 vdd.n5024 0.0196536
R44902 vdd.n5073 vdd.n5072 0.0196536
R44903 vdd.n5124 vdd.n5123 0.0196536
R44904 vdd.n5174 vdd.n5173 0.0196536
R44905 vdd.n5222 vdd.n5221 0.0196536
R44906 vdd.n5272 vdd.n5271 0.0196536
R44907 vdd.n5319 vdd.n5318 0.0196536
R44908 vdd.n5369 vdd.n5368 0.0196536
R44909 vdd.n5419 vdd.n5418 0.0196536
R44910 vdd.n5467 vdd.n5466 0.0196536
R44911 vdd.n4410 vdd.n4409 0.0196536
R44912 vdd.n5518 vdd.n5517 0.0196536
R44913 vdd.n5565 vdd.n5564 0.0196536
R44914 vdd.n5615 vdd.n5614 0.0196536
R44915 vdd.n5665 vdd.n5664 0.0196536
R44916 vdd.n5713 vdd.n5712 0.0196536
R44917 vdd.n1148 vdd.n1147 0.0196536
R44918 vdd.n1196 vdd.n1195 0.0196536
R44919 vdd.n1297 vdd.n1296 0.0196536
R44920 vdd.n1345 vdd.n1344 0.0196536
R44921 vdd.n1393 vdd.n1392 0.0196536
R44922 vdd.n1441 vdd.n1440 0.0196536
R44923 vdd.n1542 vdd.n1541 0.0196536
R44924 vdd.n655 vdd.n654 0.0196536
R44925 vdd.n1590 vdd.n1589 0.0196536
R44926 vdd.n1637 vdd.n1636 0.0196536
R44927 vdd.n1687 vdd.n1686 0.0196536
R44928 vdd.n1737 vdd.n1736 0.0196536
R44929 vdd.n1785 vdd.n1784 0.0196536
R44930 vdd.n1513 vdd.n1512 0.0196536
R44931 vdd.n1836 vdd.n1835 0.0196536
R44932 vdd.n1883 vdd.n1882 0.0196536
R44933 vdd.n1931 vdd.n1930 0.0196536
R44934 vdd.n1982 vdd.n1981 0.0196536
R44935 vdd.n2032 vdd.n2031 0.0196536
R44936 vdd.n2080 vdd.n2079 0.0196536
R44937 vdd.n2130 vdd.n2129 0.0196536
R44938 vdd.n2177 vdd.n2176 0.0196536
R44939 vdd.n2227 vdd.n2226 0.0196536
R44940 vdd.n2277 vdd.n2276 0.0196536
R44941 vdd.n2325 vdd.n2324 0.0196536
R44942 vdd.n1268 vdd.n1267 0.0196536
R44943 vdd.n2376 vdd.n2375 0.0196536
R44944 vdd.n2423 vdd.n2422 0.0196536
R44945 vdd.n2473 vdd.n2472 0.0196536
R44946 vdd.n2523 vdd.n2522 0.0196536
R44947 vdd.n2571 vdd.n2570 0.0196536
R44948 vdd.n11460 vdd.n11459 0.0196536
R44949 vdd.n11507 vdd.n11506 0.0196536
R44950 vdd.n11557 vdd.n11556 0.0196536
R44951 vdd.n11607 vdd.n11606 0.0196536
R44952 vdd.n11655 vdd.n11654 0.0196536
R44953 vdd.n483 vdd.n482 0.0196536
R44954 vdd.n11706 vdd.n11705 0.0196536
R44955 vdd.n11753 vdd.n11752 0.0196536
R44956 vdd.n11801 vdd.n11800 0.0196536
R44957 vdd.n11852 vdd.n11851 0.0196536
R44958 vdd.n11902 vdd.n11901 0.0196536
R44959 vdd.n11950 vdd.n11949 0.0196536
R44960 vdd.n12000 vdd.n11999 0.0196536
R44961 vdd.n12047 vdd.n12046 0.0196536
R44962 vdd.n12097 vdd.n12096 0.0196536
R44963 vdd.n12147 vdd.n12146 0.0196536
R44964 vdd.n12195 vdd.n12194 0.0196536
R44965 vdd.n238 vdd.n237 0.0196536
R44966 vdd.n12246 vdd.n12245 0.0196536
R44967 vdd.n12293 vdd.n12292 0.0196536
R44968 vdd.n12343 vdd.n12342 0.0196536
R44969 vdd.n12393 vdd.n12392 0.0196536
R44970 vdd.n12441 vdd.n12440 0.0196536
R44971 vdd.n12482 vdd.n12481 0.0196151
R44972 vdd.n12503 vdd.n12502 0.0196151
R44973 vdd.n133 vdd.n132 0.0196151
R44974 vdd.n181 vdd.n180 0.0196151
R44975 vdd.n282 vdd.n281 0.0196151
R44976 vdd.n330 vdd.n329 0.0196151
R44977 vdd.n378 vdd.n377 0.0196151
R44978 vdd.n426 vdd.n425 0.0196151
R44979 vdd.n527 vdd.n526 0.0196151
R44980 vdd.n575 vdd.n574 0.0196151
R44981 vdd.n6990 vdd.n6981 0.0196151
R44982 vdd.n7005 vdd.n7004 0.0196151
R44983 vdd.n7038 vdd.n7029 0.0196151
R44984 vdd.n7053 vdd.n7052 0.0196151
R44985 vdd.n7140 vdd.n7131 0.0196151
R44986 vdd.n7155 vdd.n7154 0.0196151
R44987 vdd.n7188 vdd.n7179 0.0196151
R44988 vdd.n7203 vdd.n7202 0.0196151
R44989 vdd.n7236 vdd.n7227 0.0196151
R44990 vdd.n7251 vdd.n7250 0.0196151
R44991 vdd.n7284 vdd.n7275 0.0196151
R44992 vdd.n7299 vdd.n7298 0.0196151
R44993 vdd.n7386 vdd.n7377 0.0196151
R44994 vdd.n7401 vdd.n7400 0.0196151
R44995 vdd.n8906 vdd.n8897 0.0196151
R44996 vdd.n8921 vdd.n8920 0.0196151
R44997 vdd.n7447 vdd.n7446 0.0196151
R44998 vdd.n7495 vdd.n7494 0.0196151
R44999 vdd.n7596 vdd.n7595 0.0196151
R45000 vdd.n7644 vdd.n7643 0.0196151
R45001 vdd.n7692 vdd.n7691 0.0196151
R45002 vdd.n7740 vdd.n7739 0.0196151
R45003 vdd.n7841 vdd.n7840 0.0196151
R45004 vdd.n6954 vdd.n6953 0.0196151
R45005 vdd.n7889 vdd.n7888 0.0196151
R45006 vdd.n7936 vdd.n7935 0.0196151
R45007 vdd.n7986 vdd.n7985 0.0196151
R45008 vdd.n8036 vdd.n8035 0.0196151
R45009 vdd.n8084 vdd.n8083 0.0196151
R45010 vdd.n7776 vdd.n7775 0.0196151
R45011 vdd.n8135 vdd.n8134 0.0196151
R45012 vdd.n8182 vdd.n8181 0.0196151
R45013 vdd.n8230 vdd.n8229 0.0196151
R45014 vdd.n8281 vdd.n8280 0.0196151
R45015 vdd.n8331 vdd.n8330 0.0196151
R45016 vdd.n8379 vdd.n8378 0.0196151
R45017 vdd.n8429 vdd.n8428 0.0196151
R45018 vdd.n8476 vdd.n8475 0.0196151
R45019 vdd.n8526 vdd.n8525 0.0196151
R45020 vdd.n8576 vdd.n8575 0.0196151
R45021 vdd.n8624 vdd.n8623 0.0196151
R45022 vdd.n7531 vdd.n7530 0.0196151
R45023 vdd.n8675 vdd.n8674 0.0196151
R45024 vdd.n8722 vdd.n8721 0.0196151
R45025 vdd.n8772 vdd.n8771 0.0196151
R45026 vdd.n8822 vdd.n8821 0.0196151
R45027 vdd.n8870 vdd.n8869 0.0196151
R45028 vdd.n9003 vdd.n8994 0.0196151
R45029 vdd.n9018 vdd.n9017 0.0196151
R45030 vdd.n8955 vdd.n8946 0.0196151
R45031 vdd.n8970 vdd.n8969 0.0196151
R45032 vdd.n9052 vdd.n9043 0.0196151
R45033 vdd.n9067 vdd.n9066 0.0196151
R45034 vdd.n9102 vdd.n9093 0.0196151
R45035 vdd.n9117 vdd.n9116 0.0196151
R45036 vdd.n9150 vdd.n9141 0.0196151
R45037 vdd.n9165 vdd.n9164 0.0196151
R45038 vdd.n7334 vdd.n7333 0.0196151
R45039 vdd.n7355 vdd.n7354 0.0196151
R45040 vdd.n9298 vdd.n9289 0.0196151
R45041 vdd.n9313 vdd.n9312 0.0196151
R45042 vdd.n9249 vdd.n9240 0.0196151
R45043 vdd.n9264 vdd.n9263 0.0196151
R45044 vdd.n9201 vdd.n9192 0.0196151
R45045 vdd.n9216 vdd.n9215 0.0196151
R45046 vdd.n9347 vdd.n9338 0.0196151
R45047 vdd.n9362 vdd.n9361 0.0196151
R45048 vdd.n9397 vdd.n9388 0.0196151
R45049 vdd.n9412 vdd.n9411 0.0196151
R45050 vdd.n9445 vdd.n9436 0.0196151
R45051 vdd.n9460 vdd.n9459 0.0196151
R45052 vdd.n9543 vdd.n9534 0.0196151
R45053 vdd.n9558 vdd.n9557 0.0196151
R45054 vdd.n9495 vdd.n9486 0.0196151
R45055 vdd.n9510 vdd.n9509 0.0196151
R45056 vdd.n9592 vdd.n9583 0.0196151
R45057 vdd.n9607 vdd.n9606 0.0196151
R45058 vdd.n9642 vdd.n9633 0.0196151
R45059 vdd.n9657 vdd.n9656 0.0196151
R45060 vdd.n9690 vdd.n9681 0.0196151
R45061 vdd.n9705 vdd.n9704 0.0196151
R45062 vdd.n7088 vdd.n7087 0.0196151
R45063 vdd.n7109 vdd.n7108 0.0196151
R45064 vdd.n9789 vdd.n9780 0.0196151
R45065 vdd.n9804 vdd.n9803 0.0196151
R45066 vdd.n9741 vdd.n9732 0.0196151
R45067 vdd.n9756 vdd.n9755 0.0196151
R45068 vdd.n9838 vdd.n9829 0.0196151
R45069 vdd.n9853 vdd.n9852 0.0196151
R45070 vdd.n9888 vdd.n9879 0.0196151
R45071 vdd.n9903 vdd.n9902 0.0196151
R45072 vdd.n9936 vdd.n9927 0.0196151
R45073 vdd.n9951 vdd.n9950 0.0196151
R45074 vdd.n3848 vdd.n3839 0.0196151
R45075 vdd.n3863 vdd.n3862 0.0196151
R45076 vdd.n3896 vdd.n3887 0.0196151
R45077 vdd.n3911 vdd.n3910 0.0196151
R45078 vdd.n3998 vdd.n3989 0.0196151
R45079 vdd.n4013 vdd.n4012 0.0196151
R45080 vdd.n4046 vdd.n4037 0.0196151
R45081 vdd.n4061 vdd.n4060 0.0196151
R45082 vdd.n4094 vdd.n4085 0.0196151
R45083 vdd.n4109 vdd.n4108 0.0196151
R45084 vdd.n4142 vdd.n4133 0.0196151
R45085 vdd.n4157 vdd.n4156 0.0196151
R45086 vdd.n4244 vdd.n4235 0.0196151
R45087 vdd.n4259 vdd.n4258 0.0196151
R45088 vdd.n5764 vdd.n5755 0.0196151
R45089 vdd.n5779 vdd.n5778 0.0196151
R45090 vdd.n4305 vdd.n4304 0.0196151
R45091 vdd.n4353 vdd.n4352 0.0196151
R45092 vdd.n4454 vdd.n4453 0.0196151
R45093 vdd.n4502 vdd.n4501 0.0196151
R45094 vdd.n4550 vdd.n4549 0.0196151
R45095 vdd.n4598 vdd.n4597 0.0196151
R45096 vdd.n4699 vdd.n4698 0.0196151
R45097 vdd.n3812 vdd.n3811 0.0196151
R45098 vdd.n4747 vdd.n4746 0.0196151
R45099 vdd.n4794 vdd.n4793 0.0196151
R45100 vdd.n4844 vdd.n4843 0.0196151
R45101 vdd.n4894 vdd.n4893 0.0196151
R45102 vdd.n4942 vdd.n4941 0.0196151
R45103 vdd.n4634 vdd.n4633 0.0196151
R45104 vdd.n4993 vdd.n4992 0.0196151
R45105 vdd.n5040 vdd.n5039 0.0196151
R45106 vdd.n5088 vdd.n5087 0.0196151
R45107 vdd.n5139 vdd.n5138 0.0196151
R45108 vdd.n5189 vdd.n5188 0.0196151
R45109 vdd.n5237 vdd.n5236 0.0196151
R45110 vdd.n5287 vdd.n5286 0.0196151
R45111 vdd.n5334 vdd.n5333 0.0196151
R45112 vdd.n5384 vdd.n5383 0.0196151
R45113 vdd.n5434 vdd.n5433 0.0196151
R45114 vdd.n5482 vdd.n5481 0.0196151
R45115 vdd.n4389 vdd.n4388 0.0196151
R45116 vdd.n5533 vdd.n5532 0.0196151
R45117 vdd.n5580 vdd.n5579 0.0196151
R45118 vdd.n5630 vdd.n5629 0.0196151
R45119 vdd.n5680 vdd.n5679 0.0196151
R45120 vdd.n5728 vdd.n5727 0.0196151
R45121 vdd.n5861 vdd.n5852 0.0196151
R45122 vdd.n5876 vdd.n5875 0.0196151
R45123 vdd.n5813 vdd.n5804 0.0196151
R45124 vdd.n5828 vdd.n5827 0.0196151
R45125 vdd.n5910 vdd.n5901 0.0196151
R45126 vdd.n5925 vdd.n5924 0.0196151
R45127 vdd.n5960 vdd.n5951 0.0196151
R45128 vdd.n5975 vdd.n5974 0.0196151
R45129 vdd.n6008 vdd.n5999 0.0196151
R45130 vdd.n6023 vdd.n6022 0.0196151
R45131 vdd.n4192 vdd.n4191 0.0196151
R45132 vdd.n4213 vdd.n4212 0.0196151
R45133 vdd.n6156 vdd.n6147 0.0196151
R45134 vdd.n6171 vdd.n6170 0.0196151
R45135 vdd.n6107 vdd.n6098 0.0196151
R45136 vdd.n6122 vdd.n6121 0.0196151
R45137 vdd.n6059 vdd.n6050 0.0196151
R45138 vdd.n6074 vdd.n6073 0.0196151
R45139 vdd.n6205 vdd.n6196 0.0196151
R45140 vdd.n6220 vdd.n6219 0.0196151
R45141 vdd.n6255 vdd.n6246 0.0196151
R45142 vdd.n6270 vdd.n6269 0.0196151
R45143 vdd.n6303 vdd.n6294 0.0196151
R45144 vdd.n6318 vdd.n6317 0.0196151
R45145 vdd.n6401 vdd.n6392 0.0196151
R45146 vdd.n6416 vdd.n6415 0.0196151
R45147 vdd.n6353 vdd.n6344 0.0196151
R45148 vdd.n6368 vdd.n6367 0.0196151
R45149 vdd.n6450 vdd.n6441 0.0196151
R45150 vdd.n6465 vdd.n6464 0.0196151
R45151 vdd.n6500 vdd.n6491 0.0196151
R45152 vdd.n6515 vdd.n6514 0.0196151
R45153 vdd.n6548 vdd.n6539 0.0196151
R45154 vdd.n6563 vdd.n6562 0.0196151
R45155 vdd.n3946 vdd.n3945 0.0196151
R45156 vdd.n3967 vdd.n3966 0.0196151
R45157 vdd.n6647 vdd.n6638 0.0196151
R45158 vdd.n6662 vdd.n6661 0.0196151
R45159 vdd.n6599 vdd.n6590 0.0196151
R45160 vdd.n6614 vdd.n6613 0.0196151
R45161 vdd.n6696 vdd.n6687 0.0196151
R45162 vdd.n6711 vdd.n6710 0.0196151
R45163 vdd.n6746 vdd.n6737 0.0196151
R45164 vdd.n6761 vdd.n6760 0.0196151
R45165 vdd.n6794 vdd.n6785 0.0196151
R45166 vdd.n6809 vdd.n6808 0.0196151
R45167 vdd.n706 vdd.n697 0.0196151
R45168 vdd.n721 vdd.n720 0.0196151
R45169 vdd.n754 vdd.n745 0.0196151
R45170 vdd.n769 vdd.n768 0.0196151
R45171 vdd.n856 vdd.n847 0.0196151
R45172 vdd.n871 vdd.n870 0.0196151
R45173 vdd.n904 vdd.n895 0.0196151
R45174 vdd.n919 vdd.n918 0.0196151
R45175 vdd.n952 vdd.n943 0.0196151
R45176 vdd.n967 vdd.n966 0.0196151
R45177 vdd.n1000 vdd.n991 0.0196151
R45178 vdd.n1015 vdd.n1014 0.0196151
R45179 vdd.n1102 vdd.n1093 0.0196151
R45180 vdd.n1117 vdd.n1116 0.0196151
R45181 vdd.n2622 vdd.n2613 0.0196151
R45182 vdd.n2637 vdd.n2636 0.0196151
R45183 vdd.n1163 vdd.n1162 0.0196151
R45184 vdd.n1211 vdd.n1210 0.0196151
R45185 vdd.n1312 vdd.n1311 0.0196151
R45186 vdd.n1360 vdd.n1359 0.0196151
R45187 vdd.n1408 vdd.n1407 0.0196151
R45188 vdd.n1456 vdd.n1455 0.0196151
R45189 vdd.n1557 vdd.n1556 0.0196151
R45190 vdd.n670 vdd.n669 0.0196151
R45191 vdd.n1605 vdd.n1604 0.0196151
R45192 vdd.n1652 vdd.n1651 0.0196151
R45193 vdd.n1702 vdd.n1701 0.0196151
R45194 vdd.n1752 vdd.n1751 0.0196151
R45195 vdd.n1800 vdd.n1799 0.0196151
R45196 vdd.n1492 vdd.n1491 0.0196151
R45197 vdd.n1851 vdd.n1850 0.0196151
R45198 vdd.n1898 vdd.n1897 0.0196151
R45199 vdd.n1946 vdd.n1945 0.0196151
R45200 vdd.n1997 vdd.n1996 0.0196151
R45201 vdd.n2047 vdd.n2046 0.0196151
R45202 vdd.n2095 vdd.n2094 0.0196151
R45203 vdd.n2145 vdd.n2144 0.0196151
R45204 vdd.n2192 vdd.n2191 0.0196151
R45205 vdd.n2242 vdd.n2241 0.0196151
R45206 vdd.n2292 vdd.n2291 0.0196151
R45207 vdd.n2340 vdd.n2339 0.0196151
R45208 vdd.n1247 vdd.n1246 0.0196151
R45209 vdd.n2391 vdd.n2390 0.0196151
R45210 vdd.n2438 vdd.n2437 0.0196151
R45211 vdd.n2488 vdd.n2487 0.0196151
R45212 vdd.n2538 vdd.n2537 0.0196151
R45213 vdd.n2586 vdd.n2585 0.0196151
R45214 vdd.n2719 vdd.n2710 0.0196151
R45215 vdd.n2734 vdd.n2733 0.0196151
R45216 vdd.n2671 vdd.n2662 0.0196151
R45217 vdd.n2686 vdd.n2685 0.0196151
R45218 vdd.n2768 vdd.n2759 0.0196151
R45219 vdd.n2783 vdd.n2782 0.0196151
R45220 vdd.n2818 vdd.n2809 0.0196151
R45221 vdd.n2833 vdd.n2832 0.0196151
R45222 vdd.n2866 vdd.n2857 0.0196151
R45223 vdd.n2881 vdd.n2880 0.0196151
R45224 vdd.n1050 vdd.n1049 0.0196151
R45225 vdd.n1071 vdd.n1070 0.0196151
R45226 vdd.n3014 vdd.n3005 0.0196151
R45227 vdd.n3029 vdd.n3028 0.0196151
R45228 vdd.n2965 vdd.n2956 0.0196151
R45229 vdd.n2980 vdd.n2979 0.0196151
R45230 vdd.n2917 vdd.n2908 0.0196151
R45231 vdd.n2932 vdd.n2931 0.0196151
R45232 vdd.n3063 vdd.n3054 0.0196151
R45233 vdd.n3078 vdd.n3077 0.0196151
R45234 vdd.n3113 vdd.n3104 0.0196151
R45235 vdd.n3128 vdd.n3127 0.0196151
R45236 vdd.n3161 vdd.n3152 0.0196151
R45237 vdd.n3176 vdd.n3175 0.0196151
R45238 vdd.n3259 vdd.n3250 0.0196151
R45239 vdd.n3274 vdd.n3273 0.0196151
R45240 vdd.n3211 vdd.n3202 0.0196151
R45241 vdd.n3226 vdd.n3225 0.0196151
R45242 vdd.n3308 vdd.n3299 0.0196151
R45243 vdd.n3323 vdd.n3322 0.0196151
R45244 vdd.n3358 vdd.n3349 0.0196151
R45245 vdd.n3373 vdd.n3372 0.0196151
R45246 vdd.n3406 vdd.n3397 0.0196151
R45247 vdd.n3421 vdd.n3420 0.0196151
R45248 vdd.n804 vdd.n803 0.0196151
R45249 vdd.n825 vdd.n824 0.0196151
R45250 vdd.n3505 vdd.n3496 0.0196151
R45251 vdd.n3520 vdd.n3519 0.0196151
R45252 vdd.n3457 vdd.n3448 0.0196151
R45253 vdd.n3472 vdd.n3471 0.0196151
R45254 vdd.n3554 vdd.n3545 0.0196151
R45255 vdd.n3569 vdd.n3568 0.0196151
R45256 vdd.n3604 vdd.n3595 0.0196151
R45257 vdd.n3619 vdd.n3618 0.0196151
R45258 vdd.n3652 vdd.n3643 0.0196151
R45259 vdd.n3667 vdd.n3666 0.0196151
R45260 vdd.n610 vdd.n601 0.0196151
R45261 vdd.n625 vdd.n624 0.0196151
R45262 vdd.n3751 vdd.n3742 0.0196151
R45263 vdd.n3766 vdd.n3765 0.0196151
R45264 vdd.n3703 vdd.n3694 0.0196151
R45265 vdd.n3718 vdd.n3717 0.0196151
R45266 vdd.n6893 vdd.n6884 0.0196151
R45267 vdd.n6908 vdd.n6907 0.0196151
R45268 vdd.n6845 vdd.n6836 0.0196151
R45269 vdd.n6860 vdd.n6859 0.0196151
R45270 vdd.n10035 vdd.n10026 0.0196151
R45271 vdd.n10050 vdd.n10049 0.0196151
R45272 vdd.n9987 vdd.n9978 0.0196151
R45273 vdd.n10002 vdd.n10001 0.0196151
R45274 vdd.n10083 vdd.n10074 0.0196151
R45275 vdd.n10098 vdd.n10097 0.0196151
R45276 vdd.n10131 vdd.n10122 0.0196151
R45277 vdd.n10146 vdd.n10145 0.0196151
R45278 vdd.n10233 vdd.n10224 0.0196151
R45279 vdd.n10248 vdd.n10247 0.0196151
R45280 vdd.n10281 vdd.n10272 0.0196151
R45281 vdd.n10296 vdd.n10295 0.0196151
R45282 vdd.n10329 vdd.n10320 0.0196151
R45283 vdd.n10344 vdd.n10343 0.0196151
R45284 vdd.n10377 vdd.n10368 0.0196151
R45285 vdd.n10392 vdd.n10391 0.0196151
R45286 vdd.n10479 vdd.n10470 0.0196151
R45287 vdd.n10494 vdd.n10493 0.0196151
R45288 vdd.n71 vdd.n62 0.0196151
R45289 vdd.n86 vdd.n85 0.0196151
R45290 vdd.n23 vdd.n14 0.0196151
R45291 vdd.n38 vdd.n37 0.0196151
R45292 vdd.n10527 vdd.n10518 0.0196151
R45293 vdd.n10542 vdd.n10541 0.0196151
R45294 vdd.n10577 vdd.n10568 0.0196151
R45295 vdd.n10592 vdd.n10591 0.0196151
R45296 vdd.n10625 vdd.n10616 0.0196151
R45297 vdd.n10640 vdd.n10639 0.0196151
R45298 vdd.n10427 vdd.n10426 0.0196151
R45299 vdd.n10448 vdd.n10447 0.0196151
R45300 vdd.n10773 vdd.n10764 0.0196151
R45301 vdd.n10788 vdd.n10787 0.0196151
R45302 vdd.n10724 vdd.n10715 0.0196151
R45303 vdd.n10739 vdd.n10738 0.0196151
R45304 vdd.n10676 vdd.n10667 0.0196151
R45305 vdd.n10691 vdd.n10690 0.0196151
R45306 vdd.n10822 vdd.n10813 0.0196151
R45307 vdd.n10837 vdd.n10836 0.0196151
R45308 vdd.n10872 vdd.n10863 0.0196151
R45309 vdd.n10887 vdd.n10886 0.0196151
R45310 vdd.n10920 vdd.n10911 0.0196151
R45311 vdd.n10935 vdd.n10934 0.0196151
R45312 vdd.n11018 vdd.n11009 0.0196151
R45313 vdd.n11033 vdd.n11032 0.0196151
R45314 vdd.n10970 vdd.n10961 0.0196151
R45315 vdd.n10985 vdd.n10984 0.0196151
R45316 vdd.n11067 vdd.n11058 0.0196151
R45317 vdd.n11082 vdd.n11081 0.0196151
R45318 vdd.n11117 vdd.n11108 0.0196151
R45319 vdd.n11132 vdd.n11131 0.0196151
R45320 vdd.n11165 vdd.n11156 0.0196151
R45321 vdd.n11180 vdd.n11179 0.0196151
R45322 vdd.n10181 vdd.n10180 0.0196151
R45323 vdd.n10202 vdd.n10201 0.0196151
R45324 vdd.n11264 vdd.n11255 0.0196151
R45325 vdd.n11279 vdd.n11278 0.0196151
R45326 vdd.n11216 vdd.n11207 0.0196151
R45327 vdd.n11231 vdd.n11230 0.0196151
R45328 vdd.n11313 vdd.n11304 0.0196151
R45329 vdd.n11328 vdd.n11327 0.0196151
R45330 vdd.n11363 vdd.n11354 0.0196151
R45331 vdd.n11378 vdd.n11377 0.0196151
R45332 vdd.n11411 vdd.n11402 0.0196151
R45333 vdd.n11426 vdd.n11425 0.0196151
R45334 vdd.n11475 vdd.n11474 0.0196151
R45335 vdd.n11522 vdd.n11521 0.0196151
R45336 vdd.n11572 vdd.n11571 0.0196151
R45337 vdd.n11622 vdd.n11621 0.0196151
R45338 vdd.n11670 vdd.n11669 0.0196151
R45339 vdd.n462 vdd.n461 0.0196151
R45340 vdd.n11721 vdd.n11720 0.0196151
R45341 vdd.n11768 vdd.n11767 0.0196151
R45342 vdd.n11816 vdd.n11815 0.0196151
R45343 vdd.n11867 vdd.n11866 0.0196151
R45344 vdd.n11917 vdd.n11916 0.0196151
R45345 vdd.n11965 vdd.n11964 0.0196151
R45346 vdd.n12015 vdd.n12014 0.0196151
R45347 vdd.n12062 vdd.n12061 0.0196151
R45348 vdd.n12112 vdd.n12111 0.0196151
R45349 vdd.n12162 vdd.n12161 0.0196151
R45350 vdd.n12210 vdd.n12209 0.0196151
R45351 vdd.n217 vdd.n216 0.0196151
R45352 vdd.n12261 vdd.n12260 0.0196151
R45353 vdd.n12308 vdd.n12307 0.0196151
R45354 vdd.n12358 vdd.n12357 0.0196151
R45355 vdd.n12408 vdd.n12407 0.0196151
R45356 vdd.n12456 vdd.n12455 0.0196151
R45357 vdd.n7803 vdd.n7802 0.0185921
R45358 vdd.n7558 vdd.n7557 0.0185921
R45359 vdd.n7361 vdd.n7359 0.0185921
R45360 vdd.n7115 vdd.n7113 0.0185921
R45361 vdd.n4661 vdd.n4660 0.0185921
R45362 vdd.n4416 vdd.n4415 0.0185921
R45363 vdd.n4219 vdd.n4217 0.0185921
R45364 vdd.n3973 vdd.n3971 0.0185921
R45365 vdd.n1519 vdd.n1518 0.0185921
R45366 vdd.n1274 vdd.n1273 0.0185921
R45367 vdd.n1077 vdd.n1075 0.0185921
R45368 vdd.n831 vdd.n829 0.0185921
R45369 vdd.n10454 vdd.n10452 0.0185921
R45370 vdd.n10208 vdd.n10206 0.0185921
R45371 vdd.n489 vdd.n488 0.0185921
R45372 vdd.n244 vdd.n243 0.0185921
R45373 vdd vdd 0.0169474
R45374 vdd vdd 0.0169474
R45375 vdd vdd 0.0169474
R45376 vdd vdd 0.0169474
R45377 vdd vdd 0.0169474
R45378 vdd vdd 0.0169474
R45379 vdd vdd 0.0169474
R45380 vdd vdd 0.0169474
R45381 vdd.n7803 vdd 0.0136579
R45382 vdd.n7558 vdd 0.0136579
R45383 vdd.n4661 vdd 0.0136579
R45384 vdd.n4416 vdd 0.0136579
R45385 vdd vdd 0.0136579
R45386 vdd.n1519 vdd 0.0136579
R45387 vdd.n1274 vdd 0.0136579
R45388 vdd.n489 vdd 0.0136579
R45389 vdd.n244 vdd 0.0136579
R45390 vdd.n12472 vdd.n12471 0.0130799
R45391 vdd.n12471 vdd.n12470 0.0130799
R45392 vdd.n12475 vdd.n12474 0.0130799
R45393 vdd.n12474 vdd.n12473 0.0130799
R45394 vdd.n12498 vdd.n12497 0.0130799
R45395 vdd.n12497 vdd.n12496 0.0130799
R45396 vdd.n12500 vdd.n12499 0.0130799
R45397 vdd.n12477 vdd.n12476 0.0130799
R45398 vdd.n104 vdd.n97 0.0130799
R45399 vdd.n104 vdd.n102 0.0130799
R45400 vdd.n128 vdd.n127 0.0130799
R45401 vdd.n127 vdd.n103 0.0130799
R45402 vdd.n112 vdd.n110 0.0130799
R45403 vdd.n110 vdd.n109 0.0130799
R45404 vdd.n115 vdd.n111 0.0130799
R45405 vdd.n130 vdd.n129 0.0130799
R45406 vdd.n152 vdd.n145 0.0130799
R45407 vdd.n152 vdd.n150 0.0130799
R45408 vdd.n176 vdd.n175 0.0130799
R45409 vdd.n175 vdd.n151 0.0130799
R45410 vdd.n160 vdd.n158 0.0130799
R45411 vdd.n158 vdd.n157 0.0130799
R45412 vdd.n163 vdd.n159 0.0130799
R45413 vdd.n178 vdd.n177 0.0130799
R45414 vdd.n253 vdd.n246 0.0130799
R45415 vdd.n253 vdd.n251 0.0130799
R45416 vdd.n277 vdd.n276 0.0130799
R45417 vdd.n276 vdd.n252 0.0130799
R45418 vdd.n261 vdd.n259 0.0130799
R45419 vdd.n259 vdd.n258 0.0130799
R45420 vdd.n264 vdd.n260 0.0130799
R45421 vdd.n279 vdd.n278 0.0130799
R45422 vdd.n301 vdd.n294 0.0130799
R45423 vdd.n301 vdd.n299 0.0130799
R45424 vdd.n325 vdd.n324 0.0130799
R45425 vdd.n324 vdd.n300 0.0130799
R45426 vdd.n309 vdd.n307 0.0130799
R45427 vdd.n307 vdd.n306 0.0130799
R45428 vdd.n312 vdd.n308 0.0130799
R45429 vdd.n327 vdd.n326 0.0130799
R45430 vdd.n349 vdd.n342 0.0130799
R45431 vdd.n349 vdd.n347 0.0130799
R45432 vdd.n373 vdd.n372 0.0130799
R45433 vdd.n372 vdd.n348 0.0130799
R45434 vdd.n357 vdd.n355 0.0130799
R45435 vdd.n355 vdd.n354 0.0130799
R45436 vdd.n360 vdd.n356 0.0130799
R45437 vdd.n375 vdd.n374 0.0130799
R45438 vdd.n397 vdd.n390 0.0130799
R45439 vdd.n397 vdd.n395 0.0130799
R45440 vdd.n421 vdd.n420 0.0130799
R45441 vdd.n420 vdd.n396 0.0130799
R45442 vdd.n405 vdd.n403 0.0130799
R45443 vdd.n403 vdd.n402 0.0130799
R45444 vdd.n408 vdd.n404 0.0130799
R45445 vdd.n423 vdd.n422 0.0130799
R45446 vdd.n498 vdd.n491 0.0130799
R45447 vdd.n498 vdd.n496 0.0130799
R45448 vdd.n522 vdd.n521 0.0130799
R45449 vdd.n521 vdd.n497 0.0130799
R45450 vdd.n506 vdd.n504 0.0130799
R45451 vdd.n504 vdd.n503 0.0130799
R45452 vdd.n509 vdd.n505 0.0130799
R45453 vdd.n524 vdd.n523 0.0130799
R45454 vdd.n546 vdd.n539 0.0130799
R45455 vdd.n546 vdd.n544 0.0130799
R45456 vdd.n570 vdd.n569 0.0130799
R45457 vdd.n569 vdd.n545 0.0130799
R45458 vdd.n554 vdd.n552 0.0130799
R45459 vdd.n552 vdd.n551 0.0130799
R45460 vdd.n557 vdd.n553 0.0130799
R45461 vdd.n572 vdd.n571 0.0130799
R45462 vdd.n6974 vdd.n6967 0.0130799
R45463 vdd.n6974 vdd.n6972 0.0130799
R45464 vdd.n6987 vdd.n6980 0.0130799
R45465 vdd.n6980 vdd.n6979 0.0130799
R45466 vdd.n6998 vdd.n6997 0.0130799
R45467 vdd.n6997 vdd.n6973 0.0130799
R45468 vdd.n7000 vdd.n6999 0.0130799
R45469 vdd.n6986 vdd.n6985 0.0130799
R45470 vdd.n7022 vdd.n7015 0.0130799
R45471 vdd.n7022 vdd.n7020 0.0130799
R45472 vdd.n7035 vdd.n7028 0.0130799
R45473 vdd.n7028 vdd.n7027 0.0130799
R45474 vdd.n7046 vdd.n7045 0.0130799
R45475 vdd.n7045 vdd.n7021 0.0130799
R45476 vdd.n7048 vdd.n7047 0.0130799
R45477 vdd.n7034 vdd.n7033 0.0130799
R45478 vdd.n7124 vdd.n7117 0.0130799
R45479 vdd.n7124 vdd.n7122 0.0130799
R45480 vdd.n7137 vdd.n7130 0.0130799
R45481 vdd.n7130 vdd.n7129 0.0130799
R45482 vdd.n7148 vdd.n7147 0.0130799
R45483 vdd.n7147 vdd.n7123 0.0130799
R45484 vdd.n7150 vdd.n7149 0.0130799
R45485 vdd.n7136 vdd.n7135 0.0130799
R45486 vdd.n7172 vdd.n7165 0.0130799
R45487 vdd.n7172 vdd.n7170 0.0130799
R45488 vdd.n7185 vdd.n7178 0.0130799
R45489 vdd.n7178 vdd.n7177 0.0130799
R45490 vdd.n7196 vdd.n7195 0.0130799
R45491 vdd.n7195 vdd.n7171 0.0130799
R45492 vdd.n7198 vdd.n7197 0.0130799
R45493 vdd.n7184 vdd.n7183 0.0130799
R45494 vdd.n7220 vdd.n7213 0.0130799
R45495 vdd.n7220 vdd.n7218 0.0130799
R45496 vdd.n7233 vdd.n7226 0.0130799
R45497 vdd.n7226 vdd.n7225 0.0130799
R45498 vdd.n7244 vdd.n7243 0.0130799
R45499 vdd.n7243 vdd.n7219 0.0130799
R45500 vdd.n7246 vdd.n7245 0.0130799
R45501 vdd.n7232 vdd.n7231 0.0130799
R45502 vdd.n7268 vdd.n7261 0.0130799
R45503 vdd.n7268 vdd.n7266 0.0130799
R45504 vdd.n7281 vdd.n7274 0.0130799
R45505 vdd.n7274 vdd.n7273 0.0130799
R45506 vdd.n7292 vdd.n7291 0.0130799
R45507 vdd.n7291 vdd.n7267 0.0130799
R45508 vdd.n7294 vdd.n7293 0.0130799
R45509 vdd.n7280 vdd.n7279 0.0130799
R45510 vdd.n7370 vdd.n7363 0.0130799
R45511 vdd.n7370 vdd.n7368 0.0130799
R45512 vdd.n7383 vdd.n7376 0.0130799
R45513 vdd.n7376 vdd.n7375 0.0130799
R45514 vdd.n7394 vdd.n7393 0.0130799
R45515 vdd.n7393 vdd.n7369 0.0130799
R45516 vdd.n7396 vdd.n7395 0.0130799
R45517 vdd.n7382 vdd.n7381 0.0130799
R45518 vdd.n8890 vdd.n8883 0.0130799
R45519 vdd.n8890 vdd.n8888 0.0130799
R45520 vdd.n8903 vdd.n8896 0.0130799
R45521 vdd.n8896 vdd.n8895 0.0130799
R45522 vdd.n8914 vdd.n8913 0.0130799
R45523 vdd.n8913 vdd.n8889 0.0130799
R45524 vdd.n8916 vdd.n8915 0.0130799
R45525 vdd.n8902 vdd.n8901 0.0130799
R45526 vdd.n7418 vdd.n7411 0.0130799
R45527 vdd.n7418 vdd.n7416 0.0130799
R45528 vdd.n7442 vdd.n7441 0.0130799
R45529 vdd.n7441 vdd.n7417 0.0130799
R45530 vdd.n7426 vdd.n7424 0.0130799
R45531 vdd.n7424 vdd.n7423 0.0130799
R45532 vdd.n7429 vdd.n7425 0.0130799
R45533 vdd.n7444 vdd.n7443 0.0130799
R45534 vdd.n7466 vdd.n7459 0.0130799
R45535 vdd.n7466 vdd.n7464 0.0130799
R45536 vdd.n7490 vdd.n7489 0.0130799
R45537 vdd.n7489 vdd.n7465 0.0130799
R45538 vdd.n7474 vdd.n7472 0.0130799
R45539 vdd.n7472 vdd.n7471 0.0130799
R45540 vdd.n7477 vdd.n7473 0.0130799
R45541 vdd.n7492 vdd.n7491 0.0130799
R45542 vdd.n7567 vdd.n7560 0.0130799
R45543 vdd.n7567 vdd.n7565 0.0130799
R45544 vdd.n7591 vdd.n7590 0.0130799
R45545 vdd.n7590 vdd.n7566 0.0130799
R45546 vdd.n7575 vdd.n7573 0.0130799
R45547 vdd.n7573 vdd.n7572 0.0130799
R45548 vdd.n7578 vdd.n7574 0.0130799
R45549 vdd.n7593 vdd.n7592 0.0130799
R45550 vdd.n7615 vdd.n7608 0.0130799
R45551 vdd.n7615 vdd.n7613 0.0130799
R45552 vdd.n7639 vdd.n7638 0.0130799
R45553 vdd.n7638 vdd.n7614 0.0130799
R45554 vdd.n7623 vdd.n7621 0.0130799
R45555 vdd.n7621 vdd.n7620 0.0130799
R45556 vdd.n7626 vdd.n7622 0.0130799
R45557 vdd.n7641 vdd.n7640 0.0130799
R45558 vdd.n7663 vdd.n7656 0.0130799
R45559 vdd.n7663 vdd.n7661 0.0130799
R45560 vdd.n7687 vdd.n7686 0.0130799
R45561 vdd.n7686 vdd.n7662 0.0130799
R45562 vdd.n7671 vdd.n7669 0.0130799
R45563 vdd.n7669 vdd.n7668 0.0130799
R45564 vdd.n7674 vdd.n7670 0.0130799
R45565 vdd.n7689 vdd.n7688 0.0130799
R45566 vdd.n7711 vdd.n7704 0.0130799
R45567 vdd.n7711 vdd.n7709 0.0130799
R45568 vdd.n7735 vdd.n7734 0.0130799
R45569 vdd.n7734 vdd.n7710 0.0130799
R45570 vdd.n7719 vdd.n7717 0.0130799
R45571 vdd.n7717 vdd.n7716 0.0130799
R45572 vdd.n7722 vdd.n7718 0.0130799
R45573 vdd.n7737 vdd.n7736 0.0130799
R45574 vdd.n7812 vdd.n7805 0.0130799
R45575 vdd.n7812 vdd.n7810 0.0130799
R45576 vdd.n7836 vdd.n7835 0.0130799
R45577 vdd.n7835 vdd.n7811 0.0130799
R45578 vdd.n7820 vdd.n7818 0.0130799
R45579 vdd.n7818 vdd.n7817 0.0130799
R45580 vdd.n7823 vdd.n7819 0.0130799
R45581 vdd.n7838 vdd.n7837 0.0130799
R45582 vdd.n6925 vdd.n6918 0.0130799
R45583 vdd.n6925 vdd.n6923 0.0130799
R45584 vdd.n6949 vdd.n6948 0.0130799
R45585 vdd.n6948 vdd.n6924 0.0130799
R45586 vdd.n6933 vdd.n6931 0.0130799
R45587 vdd.n6931 vdd.n6930 0.0130799
R45588 vdd.n6936 vdd.n6932 0.0130799
R45589 vdd.n6951 vdd.n6950 0.0130799
R45590 vdd.n7860 vdd.n7853 0.0130799
R45591 vdd.n7860 vdd.n7858 0.0130799
R45592 vdd.n7884 vdd.n7883 0.0130799
R45593 vdd.n7883 vdd.n7859 0.0130799
R45594 vdd.n7868 vdd.n7866 0.0130799
R45595 vdd.n7866 vdd.n7865 0.0130799
R45596 vdd.n7871 vdd.n7867 0.0130799
R45597 vdd.n7886 vdd.n7885 0.0130799
R45598 vdd.n7907 vdd.n7900 0.0130799
R45599 vdd.n7907 vdd.n7905 0.0130799
R45600 vdd.n7931 vdd.n7930 0.0130799
R45601 vdd.n7930 vdd.n7906 0.0130799
R45602 vdd.n7915 vdd.n7913 0.0130799
R45603 vdd.n7913 vdd.n7912 0.0130799
R45604 vdd.n7918 vdd.n7914 0.0130799
R45605 vdd.n7933 vdd.n7932 0.0130799
R45606 vdd.n7957 vdd.n7950 0.0130799
R45607 vdd.n7957 vdd.n7955 0.0130799
R45608 vdd.n7981 vdd.n7980 0.0130799
R45609 vdd.n7980 vdd.n7956 0.0130799
R45610 vdd.n7965 vdd.n7963 0.0130799
R45611 vdd.n7963 vdd.n7962 0.0130799
R45612 vdd.n7968 vdd.n7964 0.0130799
R45613 vdd.n7983 vdd.n7982 0.0130799
R45614 vdd.n8007 vdd.n8000 0.0130799
R45615 vdd.n8007 vdd.n8005 0.0130799
R45616 vdd.n8031 vdd.n8030 0.0130799
R45617 vdd.n8030 vdd.n8006 0.0130799
R45618 vdd.n8015 vdd.n8013 0.0130799
R45619 vdd.n8013 vdd.n8012 0.0130799
R45620 vdd.n8018 vdd.n8014 0.0130799
R45621 vdd.n8033 vdd.n8032 0.0130799
R45622 vdd.n8055 vdd.n8048 0.0130799
R45623 vdd.n8055 vdd.n8053 0.0130799
R45624 vdd.n8079 vdd.n8078 0.0130799
R45625 vdd.n8078 vdd.n8054 0.0130799
R45626 vdd.n8063 vdd.n8061 0.0130799
R45627 vdd.n8061 vdd.n8060 0.0130799
R45628 vdd.n8066 vdd.n8062 0.0130799
R45629 vdd.n8081 vdd.n8080 0.0130799
R45630 vdd.n7787 vdd.n7786 0.0130799
R45631 vdd.n7786 vdd.n7764 0.0130799
R45632 vdd.n7770 vdd.n7769 0.0130799
R45633 vdd.n7769 vdd.n7767 0.0130799
R45634 vdd.n7761 vdd.n7760 0.0130799
R45635 vdd.n7760 vdd.n7758 0.0130799
R45636 vdd.n7756 vdd.n7754 0.0130799
R45637 vdd.n7772 vdd.n7771 0.0130799
R45638 vdd.n8106 vdd.n8099 0.0130799
R45639 vdd.n8106 vdd.n8104 0.0130799
R45640 vdd.n8130 vdd.n8129 0.0130799
R45641 vdd.n8129 vdd.n8105 0.0130799
R45642 vdd.n8114 vdd.n8112 0.0130799
R45643 vdd.n8112 vdd.n8111 0.0130799
R45644 vdd.n8117 vdd.n8113 0.0130799
R45645 vdd.n8132 vdd.n8131 0.0130799
R45646 vdd.n8153 vdd.n8146 0.0130799
R45647 vdd.n8153 vdd.n8151 0.0130799
R45648 vdd.n8177 vdd.n8176 0.0130799
R45649 vdd.n8176 vdd.n8152 0.0130799
R45650 vdd.n8161 vdd.n8159 0.0130799
R45651 vdd.n8159 vdd.n8158 0.0130799
R45652 vdd.n8164 vdd.n8160 0.0130799
R45653 vdd.n8179 vdd.n8178 0.0130799
R45654 vdd.n8201 vdd.n8194 0.0130799
R45655 vdd.n8201 vdd.n8199 0.0130799
R45656 vdd.n8225 vdd.n8224 0.0130799
R45657 vdd.n8224 vdd.n8200 0.0130799
R45658 vdd.n8209 vdd.n8207 0.0130799
R45659 vdd.n8207 vdd.n8206 0.0130799
R45660 vdd.n8212 vdd.n8208 0.0130799
R45661 vdd.n8227 vdd.n8226 0.0130799
R45662 vdd.n8252 vdd.n8245 0.0130799
R45663 vdd.n8252 vdd.n8250 0.0130799
R45664 vdd.n8276 vdd.n8275 0.0130799
R45665 vdd.n8275 vdd.n8251 0.0130799
R45666 vdd.n8260 vdd.n8258 0.0130799
R45667 vdd.n8258 vdd.n8257 0.0130799
R45668 vdd.n8263 vdd.n8259 0.0130799
R45669 vdd.n8278 vdd.n8277 0.0130799
R45670 vdd.n8302 vdd.n8295 0.0130799
R45671 vdd.n8302 vdd.n8300 0.0130799
R45672 vdd.n8326 vdd.n8325 0.0130799
R45673 vdd.n8325 vdd.n8301 0.0130799
R45674 vdd.n8310 vdd.n8308 0.0130799
R45675 vdd.n8308 vdd.n8307 0.0130799
R45676 vdd.n8313 vdd.n8309 0.0130799
R45677 vdd.n8328 vdd.n8327 0.0130799
R45678 vdd.n8350 vdd.n8343 0.0130799
R45679 vdd.n8350 vdd.n8348 0.0130799
R45680 vdd.n8374 vdd.n8373 0.0130799
R45681 vdd.n8373 vdd.n8349 0.0130799
R45682 vdd.n8358 vdd.n8356 0.0130799
R45683 vdd.n8356 vdd.n8355 0.0130799
R45684 vdd.n8361 vdd.n8357 0.0130799
R45685 vdd.n8376 vdd.n8375 0.0130799
R45686 vdd.n8400 vdd.n8393 0.0130799
R45687 vdd.n8400 vdd.n8398 0.0130799
R45688 vdd.n8424 vdd.n8423 0.0130799
R45689 vdd.n8423 vdd.n8399 0.0130799
R45690 vdd.n8408 vdd.n8406 0.0130799
R45691 vdd.n8406 vdd.n8405 0.0130799
R45692 vdd.n8411 vdd.n8407 0.0130799
R45693 vdd.n8426 vdd.n8425 0.0130799
R45694 vdd.n8447 vdd.n8440 0.0130799
R45695 vdd.n8447 vdd.n8445 0.0130799
R45696 vdd.n8471 vdd.n8470 0.0130799
R45697 vdd.n8470 vdd.n8446 0.0130799
R45698 vdd.n8455 vdd.n8453 0.0130799
R45699 vdd.n8453 vdd.n8452 0.0130799
R45700 vdd.n8458 vdd.n8454 0.0130799
R45701 vdd.n8473 vdd.n8472 0.0130799
R45702 vdd.n8497 vdd.n8490 0.0130799
R45703 vdd.n8497 vdd.n8495 0.0130799
R45704 vdd.n8521 vdd.n8520 0.0130799
R45705 vdd.n8520 vdd.n8496 0.0130799
R45706 vdd.n8505 vdd.n8503 0.0130799
R45707 vdd.n8503 vdd.n8502 0.0130799
R45708 vdd.n8508 vdd.n8504 0.0130799
R45709 vdd.n8523 vdd.n8522 0.0130799
R45710 vdd.n8547 vdd.n8540 0.0130799
R45711 vdd.n8547 vdd.n8545 0.0130799
R45712 vdd.n8571 vdd.n8570 0.0130799
R45713 vdd.n8570 vdd.n8546 0.0130799
R45714 vdd.n8555 vdd.n8553 0.0130799
R45715 vdd.n8553 vdd.n8552 0.0130799
R45716 vdd.n8558 vdd.n8554 0.0130799
R45717 vdd.n8573 vdd.n8572 0.0130799
R45718 vdd.n8595 vdd.n8588 0.0130799
R45719 vdd.n8595 vdd.n8593 0.0130799
R45720 vdd.n8619 vdd.n8618 0.0130799
R45721 vdd.n8618 vdd.n8594 0.0130799
R45722 vdd.n8603 vdd.n8601 0.0130799
R45723 vdd.n8601 vdd.n8600 0.0130799
R45724 vdd.n8606 vdd.n8602 0.0130799
R45725 vdd.n8621 vdd.n8620 0.0130799
R45726 vdd.n7542 vdd.n7541 0.0130799
R45727 vdd.n7541 vdd.n7519 0.0130799
R45728 vdd.n7525 vdd.n7524 0.0130799
R45729 vdd.n7524 vdd.n7522 0.0130799
R45730 vdd.n7516 vdd.n7515 0.0130799
R45731 vdd.n7515 vdd.n7513 0.0130799
R45732 vdd.n7511 vdd.n7509 0.0130799
R45733 vdd.n7527 vdd.n7526 0.0130799
R45734 vdd.n8646 vdd.n8639 0.0130799
R45735 vdd.n8646 vdd.n8644 0.0130799
R45736 vdd.n8670 vdd.n8669 0.0130799
R45737 vdd.n8669 vdd.n8645 0.0130799
R45738 vdd.n8654 vdd.n8652 0.0130799
R45739 vdd.n8652 vdd.n8651 0.0130799
R45740 vdd.n8657 vdd.n8653 0.0130799
R45741 vdd.n8672 vdd.n8671 0.0130799
R45742 vdd.n8693 vdd.n8686 0.0130799
R45743 vdd.n8693 vdd.n8691 0.0130799
R45744 vdd.n8717 vdd.n8716 0.0130799
R45745 vdd.n8716 vdd.n8692 0.0130799
R45746 vdd.n8701 vdd.n8699 0.0130799
R45747 vdd.n8699 vdd.n8698 0.0130799
R45748 vdd.n8704 vdd.n8700 0.0130799
R45749 vdd.n8719 vdd.n8718 0.0130799
R45750 vdd.n8743 vdd.n8736 0.0130799
R45751 vdd.n8743 vdd.n8741 0.0130799
R45752 vdd.n8767 vdd.n8766 0.0130799
R45753 vdd.n8766 vdd.n8742 0.0130799
R45754 vdd.n8751 vdd.n8749 0.0130799
R45755 vdd.n8749 vdd.n8748 0.0130799
R45756 vdd.n8754 vdd.n8750 0.0130799
R45757 vdd.n8769 vdd.n8768 0.0130799
R45758 vdd.n8793 vdd.n8786 0.0130799
R45759 vdd.n8793 vdd.n8791 0.0130799
R45760 vdd.n8817 vdd.n8816 0.0130799
R45761 vdd.n8816 vdd.n8792 0.0130799
R45762 vdd.n8801 vdd.n8799 0.0130799
R45763 vdd.n8799 vdd.n8798 0.0130799
R45764 vdd.n8804 vdd.n8800 0.0130799
R45765 vdd.n8819 vdd.n8818 0.0130799
R45766 vdd.n8841 vdd.n8834 0.0130799
R45767 vdd.n8841 vdd.n8839 0.0130799
R45768 vdd.n8865 vdd.n8864 0.0130799
R45769 vdd.n8864 vdd.n8840 0.0130799
R45770 vdd.n8849 vdd.n8847 0.0130799
R45771 vdd.n8847 vdd.n8846 0.0130799
R45772 vdd.n8852 vdd.n8848 0.0130799
R45773 vdd.n8867 vdd.n8866 0.0130799
R45774 vdd.n8987 vdd.n8980 0.0130799
R45775 vdd.n8987 vdd.n8985 0.0130799
R45776 vdd.n9000 vdd.n8993 0.0130799
R45777 vdd.n8993 vdd.n8992 0.0130799
R45778 vdd.n9011 vdd.n9010 0.0130799
R45779 vdd.n9010 vdd.n8986 0.0130799
R45780 vdd.n9013 vdd.n9012 0.0130799
R45781 vdd.n8999 vdd.n8998 0.0130799
R45782 vdd.n8939 vdd.n8932 0.0130799
R45783 vdd.n8939 vdd.n8937 0.0130799
R45784 vdd.n8952 vdd.n8945 0.0130799
R45785 vdd.n8945 vdd.n8944 0.0130799
R45786 vdd.n8963 vdd.n8962 0.0130799
R45787 vdd.n8962 vdd.n8938 0.0130799
R45788 vdd.n8965 vdd.n8964 0.0130799
R45789 vdd.n8951 vdd.n8950 0.0130799
R45790 vdd.n9036 vdd.n9029 0.0130799
R45791 vdd.n9036 vdd.n9034 0.0130799
R45792 vdd.n9049 vdd.n9042 0.0130799
R45793 vdd.n9042 vdd.n9041 0.0130799
R45794 vdd.n9060 vdd.n9059 0.0130799
R45795 vdd.n9059 vdd.n9035 0.0130799
R45796 vdd.n9062 vdd.n9061 0.0130799
R45797 vdd.n9048 vdd.n9047 0.0130799
R45798 vdd.n9086 vdd.n9079 0.0130799
R45799 vdd.n9086 vdd.n9084 0.0130799
R45800 vdd.n9099 vdd.n9092 0.0130799
R45801 vdd.n9092 vdd.n9091 0.0130799
R45802 vdd.n9110 vdd.n9109 0.0130799
R45803 vdd.n9109 vdd.n9085 0.0130799
R45804 vdd.n9112 vdd.n9111 0.0130799
R45805 vdd.n9098 vdd.n9097 0.0130799
R45806 vdd.n9134 vdd.n9127 0.0130799
R45807 vdd.n9134 vdd.n9132 0.0130799
R45808 vdd.n9147 vdd.n9140 0.0130799
R45809 vdd.n9140 vdd.n9139 0.0130799
R45810 vdd.n9158 vdd.n9157 0.0130799
R45811 vdd.n9157 vdd.n9133 0.0130799
R45812 vdd.n9160 vdd.n9159 0.0130799
R45813 vdd.n9146 vdd.n9145 0.0130799
R45814 vdd.n7345 vdd.n7344 0.0130799
R45815 vdd.n7344 vdd.n7343 0.0130799
R45816 vdd.n7326 vdd.n7323 0.0130799
R45817 vdd.n7326 vdd.n7320 0.0130799
R45818 vdd.n7350 vdd.n7349 0.0130799
R45819 vdd.n7350 vdd.n7315 0.0130799
R45820 vdd.n7357 vdd.n7312 0.0130799
R45821 vdd.n7325 vdd.n7324 0.0130799
R45822 vdd.n9282 vdd.n9275 0.0130799
R45823 vdd.n9282 vdd.n9280 0.0130799
R45824 vdd.n9295 vdd.n9288 0.0130799
R45825 vdd.n9288 vdd.n9287 0.0130799
R45826 vdd.n9306 vdd.n9305 0.0130799
R45827 vdd.n9305 vdd.n9281 0.0130799
R45828 vdd.n9308 vdd.n9307 0.0130799
R45829 vdd.n9294 vdd.n9293 0.0130799
R45830 vdd.n9233 vdd.n9226 0.0130799
R45831 vdd.n9233 vdd.n9231 0.0130799
R45832 vdd.n9246 vdd.n9239 0.0130799
R45833 vdd.n9239 vdd.n9238 0.0130799
R45834 vdd.n9257 vdd.n9256 0.0130799
R45835 vdd.n9256 vdd.n9232 0.0130799
R45836 vdd.n9259 vdd.n9258 0.0130799
R45837 vdd.n9245 vdd.n9244 0.0130799
R45838 vdd.n9185 vdd.n9178 0.0130799
R45839 vdd.n9185 vdd.n9183 0.0130799
R45840 vdd.n9198 vdd.n9191 0.0130799
R45841 vdd.n9191 vdd.n9190 0.0130799
R45842 vdd.n9209 vdd.n9208 0.0130799
R45843 vdd.n9208 vdd.n9184 0.0130799
R45844 vdd.n9211 vdd.n9210 0.0130799
R45845 vdd.n9197 vdd.n9196 0.0130799
R45846 vdd.n9331 vdd.n9324 0.0130799
R45847 vdd.n9331 vdd.n9329 0.0130799
R45848 vdd.n9344 vdd.n9337 0.0130799
R45849 vdd.n9337 vdd.n9336 0.0130799
R45850 vdd.n9355 vdd.n9354 0.0130799
R45851 vdd.n9354 vdd.n9330 0.0130799
R45852 vdd.n9357 vdd.n9356 0.0130799
R45853 vdd.n9343 vdd.n9342 0.0130799
R45854 vdd.n9381 vdd.n9374 0.0130799
R45855 vdd.n9381 vdd.n9379 0.0130799
R45856 vdd.n9394 vdd.n9387 0.0130799
R45857 vdd.n9387 vdd.n9386 0.0130799
R45858 vdd.n9405 vdd.n9404 0.0130799
R45859 vdd.n9404 vdd.n9380 0.0130799
R45860 vdd.n9407 vdd.n9406 0.0130799
R45861 vdd.n9393 vdd.n9392 0.0130799
R45862 vdd.n9429 vdd.n9422 0.0130799
R45863 vdd.n9429 vdd.n9427 0.0130799
R45864 vdd.n9442 vdd.n9435 0.0130799
R45865 vdd.n9435 vdd.n9434 0.0130799
R45866 vdd.n9453 vdd.n9452 0.0130799
R45867 vdd.n9452 vdd.n9428 0.0130799
R45868 vdd.n9455 vdd.n9454 0.0130799
R45869 vdd.n9441 vdd.n9440 0.0130799
R45870 vdd.n9527 vdd.n9520 0.0130799
R45871 vdd.n9527 vdd.n9525 0.0130799
R45872 vdd.n9540 vdd.n9533 0.0130799
R45873 vdd.n9533 vdd.n9532 0.0130799
R45874 vdd.n9551 vdd.n9550 0.0130799
R45875 vdd.n9550 vdd.n9526 0.0130799
R45876 vdd.n9553 vdd.n9552 0.0130799
R45877 vdd.n9539 vdd.n9538 0.0130799
R45878 vdd.n9479 vdd.n9472 0.0130799
R45879 vdd.n9479 vdd.n9477 0.0130799
R45880 vdd.n9492 vdd.n9485 0.0130799
R45881 vdd.n9485 vdd.n9484 0.0130799
R45882 vdd.n9503 vdd.n9502 0.0130799
R45883 vdd.n9502 vdd.n9478 0.0130799
R45884 vdd.n9505 vdd.n9504 0.0130799
R45885 vdd.n9491 vdd.n9490 0.0130799
R45886 vdd.n9576 vdd.n9569 0.0130799
R45887 vdd.n9576 vdd.n9574 0.0130799
R45888 vdd.n9589 vdd.n9582 0.0130799
R45889 vdd.n9582 vdd.n9581 0.0130799
R45890 vdd.n9600 vdd.n9599 0.0130799
R45891 vdd.n9599 vdd.n9575 0.0130799
R45892 vdd.n9602 vdd.n9601 0.0130799
R45893 vdd.n9588 vdd.n9587 0.0130799
R45894 vdd.n9626 vdd.n9619 0.0130799
R45895 vdd.n9626 vdd.n9624 0.0130799
R45896 vdd.n9639 vdd.n9632 0.0130799
R45897 vdd.n9632 vdd.n9631 0.0130799
R45898 vdd.n9650 vdd.n9649 0.0130799
R45899 vdd.n9649 vdd.n9625 0.0130799
R45900 vdd.n9652 vdd.n9651 0.0130799
R45901 vdd.n9638 vdd.n9637 0.0130799
R45902 vdd.n9674 vdd.n9667 0.0130799
R45903 vdd.n9674 vdd.n9672 0.0130799
R45904 vdd.n9687 vdd.n9680 0.0130799
R45905 vdd.n9680 vdd.n9679 0.0130799
R45906 vdd.n9698 vdd.n9697 0.0130799
R45907 vdd.n9697 vdd.n9673 0.0130799
R45908 vdd.n9700 vdd.n9699 0.0130799
R45909 vdd.n9686 vdd.n9685 0.0130799
R45910 vdd.n7099 vdd.n7098 0.0130799
R45911 vdd.n7098 vdd.n7097 0.0130799
R45912 vdd.n7080 vdd.n7077 0.0130799
R45913 vdd.n7080 vdd.n7074 0.0130799
R45914 vdd.n7104 vdd.n7103 0.0130799
R45915 vdd.n7104 vdd.n7069 0.0130799
R45916 vdd.n7111 vdd.n7066 0.0130799
R45917 vdd.n7079 vdd.n7078 0.0130799
R45918 vdd.n9773 vdd.n9766 0.0130799
R45919 vdd.n9773 vdd.n9771 0.0130799
R45920 vdd.n9786 vdd.n9779 0.0130799
R45921 vdd.n9779 vdd.n9778 0.0130799
R45922 vdd.n9797 vdd.n9796 0.0130799
R45923 vdd.n9796 vdd.n9772 0.0130799
R45924 vdd.n9799 vdd.n9798 0.0130799
R45925 vdd.n9785 vdd.n9784 0.0130799
R45926 vdd.n9725 vdd.n9718 0.0130799
R45927 vdd.n9725 vdd.n9723 0.0130799
R45928 vdd.n9738 vdd.n9731 0.0130799
R45929 vdd.n9731 vdd.n9730 0.0130799
R45930 vdd.n9749 vdd.n9748 0.0130799
R45931 vdd.n9748 vdd.n9724 0.0130799
R45932 vdd.n9751 vdd.n9750 0.0130799
R45933 vdd.n9737 vdd.n9736 0.0130799
R45934 vdd.n9822 vdd.n9815 0.0130799
R45935 vdd.n9822 vdd.n9820 0.0130799
R45936 vdd.n9835 vdd.n9828 0.0130799
R45937 vdd.n9828 vdd.n9827 0.0130799
R45938 vdd.n9846 vdd.n9845 0.0130799
R45939 vdd.n9845 vdd.n9821 0.0130799
R45940 vdd.n9848 vdd.n9847 0.0130799
R45941 vdd.n9834 vdd.n9833 0.0130799
R45942 vdd.n9872 vdd.n9865 0.0130799
R45943 vdd.n9872 vdd.n9870 0.0130799
R45944 vdd.n9885 vdd.n9878 0.0130799
R45945 vdd.n9878 vdd.n9877 0.0130799
R45946 vdd.n9896 vdd.n9895 0.0130799
R45947 vdd.n9895 vdd.n9871 0.0130799
R45948 vdd.n9898 vdd.n9897 0.0130799
R45949 vdd.n9884 vdd.n9883 0.0130799
R45950 vdd.n9920 vdd.n9913 0.0130799
R45951 vdd.n9920 vdd.n9918 0.0130799
R45952 vdd.n9933 vdd.n9926 0.0130799
R45953 vdd.n9926 vdd.n9925 0.0130799
R45954 vdd.n9944 vdd.n9943 0.0130799
R45955 vdd.n9943 vdd.n9919 0.0130799
R45956 vdd.n9946 vdd.n9945 0.0130799
R45957 vdd.n9932 vdd.n9931 0.0130799
R45958 vdd.n3832 vdd.n3825 0.0130799
R45959 vdd.n3832 vdd.n3830 0.0130799
R45960 vdd.n3845 vdd.n3838 0.0130799
R45961 vdd.n3838 vdd.n3837 0.0130799
R45962 vdd.n3856 vdd.n3855 0.0130799
R45963 vdd.n3855 vdd.n3831 0.0130799
R45964 vdd.n3858 vdd.n3857 0.0130799
R45965 vdd.n3844 vdd.n3843 0.0130799
R45966 vdd.n3880 vdd.n3873 0.0130799
R45967 vdd.n3880 vdd.n3878 0.0130799
R45968 vdd.n3893 vdd.n3886 0.0130799
R45969 vdd.n3886 vdd.n3885 0.0130799
R45970 vdd.n3904 vdd.n3903 0.0130799
R45971 vdd.n3903 vdd.n3879 0.0130799
R45972 vdd.n3906 vdd.n3905 0.0130799
R45973 vdd.n3892 vdd.n3891 0.0130799
R45974 vdd.n3982 vdd.n3975 0.0130799
R45975 vdd.n3982 vdd.n3980 0.0130799
R45976 vdd.n3995 vdd.n3988 0.0130799
R45977 vdd.n3988 vdd.n3987 0.0130799
R45978 vdd.n4006 vdd.n4005 0.0130799
R45979 vdd.n4005 vdd.n3981 0.0130799
R45980 vdd.n4008 vdd.n4007 0.0130799
R45981 vdd.n3994 vdd.n3993 0.0130799
R45982 vdd.n4030 vdd.n4023 0.0130799
R45983 vdd.n4030 vdd.n4028 0.0130799
R45984 vdd.n4043 vdd.n4036 0.0130799
R45985 vdd.n4036 vdd.n4035 0.0130799
R45986 vdd.n4054 vdd.n4053 0.0130799
R45987 vdd.n4053 vdd.n4029 0.0130799
R45988 vdd.n4056 vdd.n4055 0.0130799
R45989 vdd.n4042 vdd.n4041 0.0130799
R45990 vdd.n4078 vdd.n4071 0.0130799
R45991 vdd.n4078 vdd.n4076 0.0130799
R45992 vdd.n4091 vdd.n4084 0.0130799
R45993 vdd.n4084 vdd.n4083 0.0130799
R45994 vdd.n4102 vdd.n4101 0.0130799
R45995 vdd.n4101 vdd.n4077 0.0130799
R45996 vdd.n4104 vdd.n4103 0.0130799
R45997 vdd.n4090 vdd.n4089 0.0130799
R45998 vdd.n4126 vdd.n4119 0.0130799
R45999 vdd.n4126 vdd.n4124 0.0130799
R46000 vdd.n4139 vdd.n4132 0.0130799
R46001 vdd.n4132 vdd.n4131 0.0130799
R46002 vdd.n4150 vdd.n4149 0.0130799
R46003 vdd.n4149 vdd.n4125 0.0130799
R46004 vdd.n4152 vdd.n4151 0.0130799
R46005 vdd.n4138 vdd.n4137 0.0130799
R46006 vdd.n4228 vdd.n4221 0.0130799
R46007 vdd.n4228 vdd.n4226 0.0130799
R46008 vdd.n4241 vdd.n4234 0.0130799
R46009 vdd.n4234 vdd.n4233 0.0130799
R46010 vdd.n4252 vdd.n4251 0.0130799
R46011 vdd.n4251 vdd.n4227 0.0130799
R46012 vdd.n4254 vdd.n4253 0.0130799
R46013 vdd.n4240 vdd.n4239 0.0130799
R46014 vdd.n5748 vdd.n5741 0.0130799
R46015 vdd.n5748 vdd.n5746 0.0130799
R46016 vdd.n5761 vdd.n5754 0.0130799
R46017 vdd.n5754 vdd.n5753 0.0130799
R46018 vdd.n5772 vdd.n5771 0.0130799
R46019 vdd.n5771 vdd.n5747 0.0130799
R46020 vdd.n5774 vdd.n5773 0.0130799
R46021 vdd.n5760 vdd.n5759 0.0130799
R46022 vdd.n4276 vdd.n4269 0.0130799
R46023 vdd.n4276 vdd.n4274 0.0130799
R46024 vdd.n4300 vdd.n4299 0.0130799
R46025 vdd.n4299 vdd.n4275 0.0130799
R46026 vdd.n4284 vdd.n4282 0.0130799
R46027 vdd.n4282 vdd.n4281 0.0130799
R46028 vdd.n4287 vdd.n4283 0.0130799
R46029 vdd.n4302 vdd.n4301 0.0130799
R46030 vdd.n4324 vdd.n4317 0.0130799
R46031 vdd.n4324 vdd.n4322 0.0130799
R46032 vdd.n4348 vdd.n4347 0.0130799
R46033 vdd.n4347 vdd.n4323 0.0130799
R46034 vdd.n4332 vdd.n4330 0.0130799
R46035 vdd.n4330 vdd.n4329 0.0130799
R46036 vdd.n4335 vdd.n4331 0.0130799
R46037 vdd.n4350 vdd.n4349 0.0130799
R46038 vdd.n4425 vdd.n4418 0.0130799
R46039 vdd.n4425 vdd.n4423 0.0130799
R46040 vdd.n4449 vdd.n4448 0.0130799
R46041 vdd.n4448 vdd.n4424 0.0130799
R46042 vdd.n4433 vdd.n4431 0.0130799
R46043 vdd.n4431 vdd.n4430 0.0130799
R46044 vdd.n4436 vdd.n4432 0.0130799
R46045 vdd.n4451 vdd.n4450 0.0130799
R46046 vdd.n4473 vdd.n4466 0.0130799
R46047 vdd.n4473 vdd.n4471 0.0130799
R46048 vdd.n4497 vdd.n4496 0.0130799
R46049 vdd.n4496 vdd.n4472 0.0130799
R46050 vdd.n4481 vdd.n4479 0.0130799
R46051 vdd.n4479 vdd.n4478 0.0130799
R46052 vdd.n4484 vdd.n4480 0.0130799
R46053 vdd.n4499 vdd.n4498 0.0130799
R46054 vdd.n4521 vdd.n4514 0.0130799
R46055 vdd.n4521 vdd.n4519 0.0130799
R46056 vdd.n4545 vdd.n4544 0.0130799
R46057 vdd.n4544 vdd.n4520 0.0130799
R46058 vdd.n4529 vdd.n4527 0.0130799
R46059 vdd.n4527 vdd.n4526 0.0130799
R46060 vdd.n4532 vdd.n4528 0.0130799
R46061 vdd.n4547 vdd.n4546 0.0130799
R46062 vdd.n4569 vdd.n4562 0.0130799
R46063 vdd.n4569 vdd.n4567 0.0130799
R46064 vdd.n4593 vdd.n4592 0.0130799
R46065 vdd.n4592 vdd.n4568 0.0130799
R46066 vdd.n4577 vdd.n4575 0.0130799
R46067 vdd.n4575 vdd.n4574 0.0130799
R46068 vdd.n4580 vdd.n4576 0.0130799
R46069 vdd.n4595 vdd.n4594 0.0130799
R46070 vdd.n4670 vdd.n4663 0.0130799
R46071 vdd.n4670 vdd.n4668 0.0130799
R46072 vdd.n4694 vdd.n4693 0.0130799
R46073 vdd.n4693 vdd.n4669 0.0130799
R46074 vdd.n4678 vdd.n4676 0.0130799
R46075 vdd.n4676 vdd.n4675 0.0130799
R46076 vdd.n4681 vdd.n4677 0.0130799
R46077 vdd.n4696 vdd.n4695 0.0130799
R46078 vdd.n3783 vdd.n3776 0.0130799
R46079 vdd.n3783 vdd.n3781 0.0130799
R46080 vdd.n3807 vdd.n3806 0.0130799
R46081 vdd.n3806 vdd.n3782 0.0130799
R46082 vdd.n3791 vdd.n3789 0.0130799
R46083 vdd.n3789 vdd.n3788 0.0130799
R46084 vdd.n3794 vdd.n3790 0.0130799
R46085 vdd.n3809 vdd.n3808 0.0130799
R46086 vdd.n4718 vdd.n4711 0.0130799
R46087 vdd.n4718 vdd.n4716 0.0130799
R46088 vdd.n4742 vdd.n4741 0.0130799
R46089 vdd.n4741 vdd.n4717 0.0130799
R46090 vdd.n4726 vdd.n4724 0.0130799
R46091 vdd.n4724 vdd.n4723 0.0130799
R46092 vdd.n4729 vdd.n4725 0.0130799
R46093 vdd.n4744 vdd.n4743 0.0130799
R46094 vdd.n4765 vdd.n4758 0.0130799
R46095 vdd.n4765 vdd.n4763 0.0130799
R46096 vdd.n4789 vdd.n4788 0.0130799
R46097 vdd.n4788 vdd.n4764 0.0130799
R46098 vdd.n4773 vdd.n4771 0.0130799
R46099 vdd.n4771 vdd.n4770 0.0130799
R46100 vdd.n4776 vdd.n4772 0.0130799
R46101 vdd.n4791 vdd.n4790 0.0130799
R46102 vdd.n4815 vdd.n4808 0.0130799
R46103 vdd.n4815 vdd.n4813 0.0130799
R46104 vdd.n4839 vdd.n4838 0.0130799
R46105 vdd.n4838 vdd.n4814 0.0130799
R46106 vdd.n4823 vdd.n4821 0.0130799
R46107 vdd.n4821 vdd.n4820 0.0130799
R46108 vdd.n4826 vdd.n4822 0.0130799
R46109 vdd.n4841 vdd.n4840 0.0130799
R46110 vdd.n4865 vdd.n4858 0.0130799
R46111 vdd.n4865 vdd.n4863 0.0130799
R46112 vdd.n4889 vdd.n4888 0.0130799
R46113 vdd.n4888 vdd.n4864 0.0130799
R46114 vdd.n4873 vdd.n4871 0.0130799
R46115 vdd.n4871 vdd.n4870 0.0130799
R46116 vdd.n4876 vdd.n4872 0.0130799
R46117 vdd.n4891 vdd.n4890 0.0130799
R46118 vdd.n4913 vdd.n4906 0.0130799
R46119 vdd.n4913 vdd.n4911 0.0130799
R46120 vdd.n4937 vdd.n4936 0.0130799
R46121 vdd.n4936 vdd.n4912 0.0130799
R46122 vdd.n4921 vdd.n4919 0.0130799
R46123 vdd.n4919 vdd.n4918 0.0130799
R46124 vdd.n4924 vdd.n4920 0.0130799
R46125 vdd.n4939 vdd.n4938 0.0130799
R46126 vdd.n4645 vdd.n4644 0.0130799
R46127 vdd.n4644 vdd.n4622 0.0130799
R46128 vdd.n4628 vdd.n4627 0.0130799
R46129 vdd.n4627 vdd.n4625 0.0130799
R46130 vdd.n4619 vdd.n4618 0.0130799
R46131 vdd.n4618 vdd.n4616 0.0130799
R46132 vdd.n4614 vdd.n4612 0.0130799
R46133 vdd.n4630 vdd.n4629 0.0130799
R46134 vdd.n4964 vdd.n4957 0.0130799
R46135 vdd.n4964 vdd.n4962 0.0130799
R46136 vdd.n4988 vdd.n4987 0.0130799
R46137 vdd.n4987 vdd.n4963 0.0130799
R46138 vdd.n4972 vdd.n4970 0.0130799
R46139 vdd.n4970 vdd.n4969 0.0130799
R46140 vdd.n4975 vdd.n4971 0.0130799
R46141 vdd.n4990 vdd.n4989 0.0130799
R46142 vdd.n5011 vdd.n5004 0.0130799
R46143 vdd.n5011 vdd.n5009 0.0130799
R46144 vdd.n5035 vdd.n5034 0.0130799
R46145 vdd.n5034 vdd.n5010 0.0130799
R46146 vdd.n5019 vdd.n5017 0.0130799
R46147 vdd.n5017 vdd.n5016 0.0130799
R46148 vdd.n5022 vdd.n5018 0.0130799
R46149 vdd.n5037 vdd.n5036 0.0130799
R46150 vdd.n5059 vdd.n5052 0.0130799
R46151 vdd.n5059 vdd.n5057 0.0130799
R46152 vdd.n5083 vdd.n5082 0.0130799
R46153 vdd.n5082 vdd.n5058 0.0130799
R46154 vdd.n5067 vdd.n5065 0.0130799
R46155 vdd.n5065 vdd.n5064 0.0130799
R46156 vdd.n5070 vdd.n5066 0.0130799
R46157 vdd.n5085 vdd.n5084 0.0130799
R46158 vdd.n5110 vdd.n5103 0.0130799
R46159 vdd.n5110 vdd.n5108 0.0130799
R46160 vdd.n5134 vdd.n5133 0.0130799
R46161 vdd.n5133 vdd.n5109 0.0130799
R46162 vdd.n5118 vdd.n5116 0.0130799
R46163 vdd.n5116 vdd.n5115 0.0130799
R46164 vdd.n5121 vdd.n5117 0.0130799
R46165 vdd.n5136 vdd.n5135 0.0130799
R46166 vdd.n5160 vdd.n5153 0.0130799
R46167 vdd.n5160 vdd.n5158 0.0130799
R46168 vdd.n5184 vdd.n5183 0.0130799
R46169 vdd.n5183 vdd.n5159 0.0130799
R46170 vdd.n5168 vdd.n5166 0.0130799
R46171 vdd.n5166 vdd.n5165 0.0130799
R46172 vdd.n5171 vdd.n5167 0.0130799
R46173 vdd.n5186 vdd.n5185 0.0130799
R46174 vdd.n5208 vdd.n5201 0.0130799
R46175 vdd.n5208 vdd.n5206 0.0130799
R46176 vdd.n5232 vdd.n5231 0.0130799
R46177 vdd.n5231 vdd.n5207 0.0130799
R46178 vdd.n5216 vdd.n5214 0.0130799
R46179 vdd.n5214 vdd.n5213 0.0130799
R46180 vdd.n5219 vdd.n5215 0.0130799
R46181 vdd.n5234 vdd.n5233 0.0130799
R46182 vdd.n5258 vdd.n5251 0.0130799
R46183 vdd.n5258 vdd.n5256 0.0130799
R46184 vdd.n5282 vdd.n5281 0.0130799
R46185 vdd.n5281 vdd.n5257 0.0130799
R46186 vdd.n5266 vdd.n5264 0.0130799
R46187 vdd.n5264 vdd.n5263 0.0130799
R46188 vdd.n5269 vdd.n5265 0.0130799
R46189 vdd.n5284 vdd.n5283 0.0130799
R46190 vdd.n5305 vdd.n5298 0.0130799
R46191 vdd.n5305 vdd.n5303 0.0130799
R46192 vdd.n5329 vdd.n5328 0.0130799
R46193 vdd.n5328 vdd.n5304 0.0130799
R46194 vdd.n5313 vdd.n5311 0.0130799
R46195 vdd.n5311 vdd.n5310 0.0130799
R46196 vdd.n5316 vdd.n5312 0.0130799
R46197 vdd.n5331 vdd.n5330 0.0130799
R46198 vdd.n5355 vdd.n5348 0.0130799
R46199 vdd.n5355 vdd.n5353 0.0130799
R46200 vdd.n5379 vdd.n5378 0.0130799
R46201 vdd.n5378 vdd.n5354 0.0130799
R46202 vdd.n5363 vdd.n5361 0.0130799
R46203 vdd.n5361 vdd.n5360 0.0130799
R46204 vdd.n5366 vdd.n5362 0.0130799
R46205 vdd.n5381 vdd.n5380 0.0130799
R46206 vdd.n5405 vdd.n5398 0.0130799
R46207 vdd.n5405 vdd.n5403 0.0130799
R46208 vdd.n5429 vdd.n5428 0.0130799
R46209 vdd.n5428 vdd.n5404 0.0130799
R46210 vdd.n5413 vdd.n5411 0.0130799
R46211 vdd.n5411 vdd.n5410 0.0130799
R46212 vdd.n5416 vdd.n5412 0.0130799
R46213 vdd.n5431 vdd.n5430 0.0130799
R46214 vdd.n5453 vdd.n5446 0.0130799
R46215 vdd.n5453 vdd.n5451 0.0130799
R46216 vdd.n5477 vdd.n5476 0.0130799
R46217 vdd.n5476 vdd.n5452 0.0130799
R46218 vdd.n5461 vdd.n5459 0.0130799
R46219 vdd.n5459 vdd.n5458 0.0130799
R46220 vdd.n5464 vdd.n5460 0.0130799
R46221 vdd.n5479 vdd.n5478 0.0130799
R46222 vdd.n4400 vdd.n4399 0.0130799
R46223 vdd.n4399 vdd.n4377 0.0130799
R46224 vdd.n4383 vdd.n4382 0.0130799
R46225 vdd.n4382 vdd.n4380 0.0130799
R46226 vdd.n4374 vdd.n4373 0.0130799
R46227 vdd.n4373 vdd.n4371 0.0130799
R46228 vdd.n4369 vdd.n4367 0.0130799
R46229 vdd.n4385 vdd.n4384 0.0130799
R46230 vdd.n5504 vdd.n5497 0.0130799
R46231 vdd.n5504 vdd.n5502 0.0130799
R46232 vdd.n5528 vdd.n5527 0.0130799
R46233 vdd.n5527 vdd.n5503 0.0130799
R46234 vdd.n5512 vdd.n5510 0.0130799
R46235 vdd.n5510 vdd.n5509 0.0130799
R46236 vdd.n5515 vdd.n5511 0.0130799
R46237 vdd.n5530 vdd.n5529 0.0130799
R46238 vdd.n5551 vdd.n5544 0.0130799
R46239 vdd.n5551 vdd.n5549 0.0130799
R46240 vdd.n5575 vdd.n5574 0.0130799
R46241 vdd.n5574 vdd.n5550 0.0130799
R46242 vdd.n5559 vdd.n5557 0.0130799
R46243 vdd.n5557 vdd.n5556 0.0130799
R46244 vdd.n5562 vdd.n5558 0.0130799
R46245 vdd.n5577 vdd.n5576 0.0130799
R46246 vdd.n5601 vdd.n5594 0.0130799
R46247 vdd.n5601 vdd.n5599 0.0130799
R46248 vdd.n5625 vdd.n5624 0.0130799
R46249 vdd.n5624 vdd.n5600 0.0130799
R46250 vdd.n5609 vdd.n5607 0.0130799
R46251 vdd.n5607 vdd.n5606 0.0130799
R46252 vdd.n5612 vdd.n5608 0.0130799
R46253 vdd.n5627 vdd.n5626 0.0130799
R46254 vdd.n5651 vdd.n5644 0.0130799
R46255 vdd.n5651 vdd.n5649 0.0130799
R46256 vdd.n5675 vdd.n5674 0.0130799
R46257 vdd.n5674 vdd.n5650 0.0130799
R46258 vdd.n5659 vdd.n5657 0.0130799
R46259 vdd.n5657 vdd.n5656 0.0130799
R46260 vdd.n5662 vdd.n5658 0.0130799
R46261 vdd.n5677 vdd.n5676 0.0130799
R46262 vdd.n5699 vdd.n5692 0.0130799
R46263 vdd.n5699 vdd.n5697 0.0130799
R46264 vdd.n5723 vdd.n5722 0.0130799
R46265 vdd.n5722 vdd.n5698 0.0130799
R46266 vdd.n5707 vdd.n5705 0.0130799
R46267 vdd.n5705 vdd.n5704 0.0130799
R46268 vdd.n5710 vdd.n5706 0.0130799
R46269 vdd.n5725 vdd.n5724 0.0130799
R46270 vdd.n5845 vdd.n5838 0.0130799
R46271 vdd.n5845 vdd.n5843 0.0130799
R46272 vdd.n5858 vdd.n5851 0.0130799
R46273 vdd.n5851 vdd.n5850 0.0130799
R46274 vdd.n5869 vdd.n5868 0.0130799
R46275 vdd.n5868 vdd.n5844 0.0130799
R46276 vdd.n5871 vdd.n5870 0.0130799
R46277 vdd.n5857 vdd.n5856 0.0130799
R46278 vdd.n5797 vdd.n5790 0.0130799
R46279 vdd.n5797 vdd.n5795 0.0130799
R46280 vdd.n5810 vdd.n5803 0.0130799
R46281 vdd.n5803 vdd.n5802 0.0130799
R46282 vdd.n5821 vdd.n5820 0.0130799
R46283 vdd.n5820 vdd.n5796 0.0130799
R46284 vdd.n5823 vdd.n5822 0.0130799
R46285 vdd.n5809 vdd.n5808 0.0130799
R46286 vdd.n5894 vdd.n5887 0.0130799
R46287 vdd.n5894 vdd.n5892 0.0130799
R46288 vdd.n5907 vdd.n5900 0.0130799
R46289 vdd.n5900 vdd.n5899 0.0130799
R46290 vdd.n5918 vdd.n5917 0.0130799
R46291 vdd.n5917 vdd.n5893 0.0130799
R46292 vdd.n5920 vdd.n5919 0.0130799
R46293 vdd.n5906 vdd.n5905 0.0130799
R46294 vdd.n5944 vdd.n5937 0.0130799
R46295 vdd.n5944 vdd.n5942 0.0130799
R46296 vdd.n5957 vdd.n5950 0.0130799
R46297 vdd.n5950 vdd.n5949 0.0130799
R46298 vdd.n5968 vdd.n5967 0.0130799
R46299 vdd.n5967 vdd.n5943 0.0130799
R46300 vdd.n5970 vdd.n5969 0.0130799
R46301 vdd.n5956 vdd.n5955 0.0130799
R46302 vdd.n5992 vdd.n5985 0.0130799
R46303 vdd.n5992 vdd.n5990 0.0130799
R46304 vdd.n6005 vdd.n5998 0.0130799
R46305 vdd.n5998 vdd.n5997 0.0130799
R46306 vdd.n6016 vdd.n6015 0.0130799
R46307 vdd.n6015 vdd.n5991 0.0130799
R46308 vdd.n6018 vdd.n6017 0.0130799
R46309 vdd.n6004 vdd.n6003 0.0130799
R46310 vdd.n4203 vdd.n4202 0.0130799
R46311 vdd.n4202 vdd.n4201 0.0130799
R46312 vdd.n4184 vdd.n4181 0.0130799
R46313 vdd.n4184 vdd.n4178 0.0130799
R46314 vdd.n4208 vdd.n4207 0.0130799
R46315 vdd.n4208 vdd.n4173 0.0130799
R46316 vdd.n4215 vdd.n4170 0.0130799
R46317 vdd.n4183 vdd.n4182 0.0130799
R46318 vdd.n6140 vdd.n6133 0.0130799
R46319 vdd.n6140 vdd.n6138 0.0130799
R46320 vdd.n6153 vdd.n6146 0.0130799
R46321 vdd.n6146 vdd.n6145 0.0130799
R46322 vdd.n6164 vdd.n6163 0.0130799
R46323 vdd.n6163 vdd.n6139 0.0130799
R46324 vdd.n6166 vdd.n6165 0.0130799
R46325 vdd.n6152 vdd.n6151 0.0130799
R46326 vdd.n6091 vdd.n6084 0.0130799
R46327 vdd.n6091 vdd.n6089 0.0130799
R46328 vdd.n6104 vdd.n6097 0.0130799
R46329 vdd.n6097 vdd.n6096 0.0130799
R46330 vdd.n6115 vdd.n6114 0.0130799
R46331 vdd.n6114 vdd.n6090 0.0130799
R46332 vdd.n6117 vdd.n6116 0.0130799
R46333 vdd.n6103 vdd.n6102 0.0130799
R46334 vdd.n6043 vdd.n6036 0.0130799
R46335 vdd.n6043 vdd.n6041 0.0130799
R46336 vdd.n6056 vdd.n6049 0.0130799
R46337 vdd.n6049 vdd.n6048 0.0130799
R46338 vdd.n6067 vdd.n6066 0.0130799
R46339 vdd.n6066 vdd.n6042 0.0130799
R46340 vdd.n6069 vdd.n6068 0.0130799
R46341 vdd.n6055 vdd.n6054 0.0130799
R46342 vdd.n6189 vdd.n6182 0.0130799
R46343 vdd.n6189 vdd.n6187 0.0130799
R46344 vdd.n6202 vdd.n6195 0.0130799
R46345 vdd.n6195 vdd.n6194 0.0130799
R46346 vdd.n6213 vdd.n6212 0.0130799
R46347 vdd.n6212 vdd.n6188 0.0130799
R46348 vdd.n6215 vdd.n6214 0.0130799
R46349 vdd.n6201 vdd.n6200 0.0130799
R46350 vdd.n6239 vdd.n6232 0.0130799
R46351 vdd.n6239 vdd.n6237 0.0130799
R46352 vdd.n6252 vdd.n6245 0.0130799
R46353 vdd.n6245 vdd.n6244 0.0130799
R46354 vdd.n6263 vdd.n6262 0.0130799
R46355 vdd.n6262 vdd.n6238 0.0130799
R46356 vdd.n6265 vdd.n6264 0.0130799
R46357 vdd.n6251 vdd.n6250 0.0130799
R46358 vdd.n6287 vdd.n6280 0.0130799
R46359 vdd.n6287 vdd.n6285 0.0130799
R46360 vdd.n6300 vdd.n6293 0.0130799
R46361 vdd.n6293 vdd.n6292 0.0130799
R46362 vdd.n6311 vdd.n6310 0.0130799
R46363 vdd.n6310 vdd.n6286 0.0130799
R46364 vdd.n6313 vdd.n6312 0.0130799
R46365 vdd.n6299 vdd.n6298 0.0130799
R46366 vdd.n6385 vdd.n6378 0.0130799
R46367 vdd.n6385 vdd.n6383 0.0130799
R46368 vdd.n6398 vdd.n6391 0.0130799
R46369 vdd.n6391 vdd.n6390 0.0130799
R46370 vdd.n6409 vdd.n6408 0.0130799
R46371 vdd.n6408 vdd.n6384 0.0130799
R46372 vdd.n6411 vdd.n6410 0.0130799
R46373 vdd.n6397 vdd.n6396 0.0130799
R46374 vdd.n6337 vdd.n6330 0.0130799
R46375 vdd.n6337 vdd.n6335 0.0130799
R46376 vdd.n6350 vdd.n6343 0.0130799
R46377 vdd.n6343 vdd.n6342 0.0130799
R46378 vdd.n6361 vdd.n6360 0.0130799
R46379 vdd.n6360 vdd.n6336 0.0130799
R46380 vdd.n6363 vdd.n6362 0.0130799
R46381 vdd.n6349 vdd.n6348 0.0130799
R46382 vdd.n6434 vdd.n6427 0.0130799
R46383 vdd.n6434 vdd.n6432 0.0130799
R46384 vdd.n6447 vdd.n6440 0.0130799
R46385 vdd.n6440 vdd.n6439 0.0130799
R46386 vdd.n6458 vdd.n6457 0.0130799
R46387 vdd.n6457 vdd.n6433 0.0130799
R46388 vdd.n6460 vdd.n6459 0.0130799
R46389 vdd.n6446 vdd.n6445 0.0130799
R46390 vdd.n6484 vdd.n6477 0.0130799
R46391 vdd.n6484 vdd.n6482 0.0130799
R46392 vdd.n6497 vdd.n6490 0.0130799
R46393 vdd.n6490 vdd.n6489 0.0130799
R46394 vdd.n6508 vdd.n6507 0.0130799
R46395 vdd.n6507 vdd.n6483 0.0130799
R46396 vdd.n6510 vdd.n6509 0.0130799
R46397 vdd.n6496 vdd.n6495 0.0130799
R46398 vdd.n6532 vdd.n6525 0.0130799
R46399 vdd.n6532 vdd.n6530 0.0130799
R46400 vdd.n6545 vdd.n6538 0.0130799
R46401 vdd.n6538 vdd.n6537 0.0130799
R46402 vdd.n6556 vdd.n6555 0.0130799
R46403 vdd.n6555 vdd.n6531 0.0130799
R46404 vdd.n6558 vdd.n6557 0.0130799
R46405 vdd.n6544 vdd.n6543 0.0130799
R46406 vdd.n3957 vdd.n3956 0.0130799
R46407 vdd.n3956 vdd.n3955 0.0130799
R46408 vdd.n3938 vdd.n3935 0.0130799
R46409 vdd.n3938 vdd.n3932 0.0130799
R46410 vdd.n3962 vdd.n3961 0.0130799
R46411 vdd.n3962 vdd.n3927 0.0130799
R46412 vdd.n3969 vdd.n3924 0.0130799
R46413 vdd.n3937 vdd.n3936 0.0130799
R46414 vdd.n6631 vdd.n6624 0.0130799
R46415 vdd.n6631 vdd.n6629 0.0130799
R46416 vdd.n6644 vdd.n6637 0.0130799
R46417 vdd.n6637 vdd.n6636 0.0130799
R46418 vdd.n6655 vdd.n6654 0.0130799
R46419 vdd.n6654 vdd.n6630 0.0130799
R46420 vdd.n6657 vdd.n6656 0.0130799
R46421 vdd.n6643 vdd.n6642 0.0130799
R46422 vdd.n6583 vdd.n6576 0.0130799
R46423 vdd.n6583 vdd.n6581 0.0130799
R46424 vdd.n6596 vdd.n6589 0.0130799
R46425 vdd.n6589 vdd.n6588 0.0130799
R46426 vdd.n6607 vdd.n6606 0.0130799
R46427 vdd.n6606 vdd.n6582 0.0130799
R46428 vdd.n6609 vdd.n6608 0.0130799
R46429 vdd.n6595 vdd.n6594 0.0130799
R46430 vdd.n6680 vdd.n6673 0.0130799
R46431 vdd.n6680 vdd.n6678 0.0130799
R46432 vdd.n6693 vdd.n6686 0.0130799
R46433 vdd.n6686 vdd.n6685 0.0130799
R46434 vdd.n6704 vdd.n6703 0.0130799
R46435 vdd.n6703 vdd.n6679 0.0130799
R46436 vdd.n6706 vdd.n6705 0.0130799
R46437 vdd.n6692 vdd.n6691 0.0130799
R46438 vdd.n6730 vdd.n6723 0.0130799
R46439 vdd.n6730 vdd.n6728 0.0130799
R46440 vdd.n6743 vdd.n6736 0.0130799
R46441 vdd.n6736 vdd.n6735 0.0130799
R46442 vdd.n6754 vdd.n6753 0.0130799
R46443 vdd.n6753 vdd.n6729 0.0130799
R46444 vdd.n6756 vdd.n6755 0.0130799
R46445 vdd.n6742 vdd.n6741 0.0130799
R46446 vdd.n6778 vdd.n6771 0.0130799
R46447 vdd.n6778 vdd.n6776 0.0130799
R46448 vdd.n6791 vdd.n6784 0.0130799
R46449 vdd.n6784 vdd.n6783 0.0130799
R46450 vdd.n6802 vdd.n6801 0.0130799
R46451 vdd.n6801 vdd.n6777 0.0130799
R46452 vdd.n6804 vdd.n6803 0.0130799
R46453 vdd.n6790 vdd.n6789 0.0130799
R46454 vdd.n690 vdd.n683 0.0130799
R46455 vdd.n690 vdd.n688 0.0130799
R46456 vdd.n703 vdd.n696 0.0130799
R46457 vdd.n696 vdd.n695 0.0130799
R46458 vdd.n714 vdd.n713 0.0130799
R46459 vdd.n713 vdd.n689 0.0130799
R46460 vdd.n716 vdd.n715 0.0130799
R46461 vdd.n702 vdd.n701 0.0130799
R46462 vdd.n738 vdd.n731 0.0130799
R46463 vdd.n738 vdd.n736 0.0130799
R46464 vdd.n751 vdd.n744 0.0130799
R46465 vdd.n744 vdd.n743 0.0130799
R46466 vdd.n762 vdd.n761 0.0130799
R46467 vdd.n761 vdd.n737 0.0130799
R46468 vdd.n764 vdd.n763 0.0130799
R46469 vdd.n750 vdd.n749 0.0130799
R46470 vdd.n840 vdd.n833 0.0130799
R46471 vdd.n840 vdd.n838 0.0130799
R46472 vdd.n853 vdd.n846 0.0130799
R46473 vdd.n846 vdd.n845 0.0130799
R46474 vdd.n864 vdd.n863 0.0130799
R46475 vdd.n863 vdd.n839 0.0130799
R46476 vdd.n866 vdd.n865 0.0130799
R46477 vdd.n852 vdd.n851 0.0130799
R46478 vdd.n888 vdd.n881 0.0130799
R46479 vdd.n888 vdd.n886 0.0130799
R46480 vdd.n901 vdd.n894 0.0130799
R46481 vdd.n894 vdd.n893 0.0130799
R46482 vdd.n912 vdd.n911 0.0130799
R46483 vdd.n911 vdd.n887 0.0130799
R46484 vdd.n914 vdd.n913 0.0130799
R46485 vdd.n900 vdd.n899 0.0130799
R46486 vdd.n936 vdd.n929 0.0130799
R46487 vdd.n936 vdd.n934 0.0130799
R46488 vdd.n949 vdd.n942 0.0130799
R46489 vdd.n942 vdd.n941 0.0130799
R46490 vdd.n960 vdd.n959 0.0130799
R46491 vdd.n959 vdd.n935 0.0130799
R46492 vdd.n962 vdd.n961 0.0130799
R46493 vdd.n948 vdd.n947 0.0130799
R46494 vdd.n984 vdd.n977 0.0130799
R46495 vdd.n984 vdd.n982 0.0130799
R46496 vdd.n997 vdd.n990 0.0130799
R46497 vdd.n990 vdd.n989 0.0130799
R46498 vdd.n1008 vdd.n1007 0.0130799
R46499 vdd.n1007 vdd.n983 0.0130799
R46500 vdd.n1010 vdd.n1009 0.0130799
R46501 vdd.n996 vdd.n995 0.0130799
R46502 vdd.n1086 vdd.n1079 0.0130799
R46503 vdd.n1086 vdd.n1084 0.0130799
R46504 vdd.n1099 vdd.n1092 0.0130799
R46505 vdd.n1092 vdd.n1091 0.0130799
R46506 vdd.n1110 vdd.n1109 0.0130799
R46507 vdd.n1109 vdd.n1085 0.0130799
R46508 vdd.n1112 vdd.n1111 0.0130799
R46509 vdd.n1098 vdd.n1097 0.0130799
R46510 vdd.n2606 vdd.n2599 0.0130799
R46511 vdd.n2606 vdd.n2604 0.0130799
R46512 vdd.n2619 vdd.n2612 0.0130799
R46513 vdd.n2612 vdd.n2611 0.0130799
R46514 vdd.n2630 vdd.n2629 0.0130799
R46515 vdd.n2629 vdd.n2605 0.0130799
R46516 vdd.n2632 vdd.n2631 0.0130799
R46517 vdd.n2618 vdd.n2617 0.0130799
R46518 vdd.n1134 vdd.n1127 0.0130799
R46519 vdd.n1134 vdd.n1132 0.0130799
R46520 vdd.n1158 vdd.n1157 0.0130799
R46521 vdd.n1157 vdd.n1133 0.0130799
R46522 vdd.n1142 vdd.n1140 0.0130799
R46523 vdd.n1140 vdd.n1139 0.0130799
R46524 vdd.n1145 vdd.n1141 0.0130799
R46525 vdd.n1160 vdd.n1159 0.0130799
R46526 vdd.n1182 vdd.n1175 0.0130799
R46527 vdd.n1182 vdd.n1180 0.0130799
R46528 vdd.n1206 vdd.n1205 0.0130799
R46529 vdd.n1205 vdd.n1181 0.0130799
R46530 vdd.n1190 vdd.n1188 0.0130799
R46531 vdd.n1188 vdd.n1187 0.0130799
R46532 vdd.n1193 vdd.n1189 0.0130799
R46533 vdd.n1208 vdd.n1207 0.0130799
R46534 vdd.n1283 vdd.n1276 0.0130799
R46535 vdd.n1283 vdd.n1281 0.0130799
R46536 vdd.n1307 vdd.n1306 0.0130799
R46537 vdd.n1306 vdd.n1282 0.0130799
R46538 vdd.n1291 vdd.n1289 0.0130799
R46539 vdd.n1289 vdd.n1288 0.0130799
R46540 vdd.n1294 vdd.n1290 0.0130799
R46541 vdd.n1309 vdd.n1308 0.0130799
R46542 vdd.n1331 vdd.n1324 0.0130799
R46543 vdd.n1331 vdd.n1329 0.0130799
R46544 vdd.n1355 vdd.n1354 0.0130799
R46545 vdd.n1354 vdd.n1330 0.0130799
R46546 vdd.n1339 vdd.n1337 0.0130799
R46547 vdd.n1337 vdd.n1336 0.0130799
R46548 vdd.n1342 vdd.n1338 0.0130799
R46549 vdd.n1357 vdd.n1356 0.0130799
R46550 vdd.n1379 vdd.n1372 0.0130799
R46551 vdd.n1379 vdd.n1377 0.0130799
R46552 vdd.n1403 vdd.n1402 0.0130799
R46553 vdd.n1402 vdd.n1378 0.0130799
R46554 vdd.n1387 vdd.n1385 0.0130799
R46555 vdd.n1385 vdd.n1384 0.0130799
R46556 vdd.n1390 vdd.n1386 0.0130799
R46557 vdd.n1405 vdd.n1404 0.0130799
R46558 vdd.n1427 vdd.n1420 0.0130799
R46559 vdd.n1427 vdd.n1425 0.0130799
R46560 vdd.n1451 vdd.n1450 0.0130799
R46561 vdd.n1450 vdd.n1426 0.0130799
R46562 vdd.n1435 vdd.n1433 0.0130799
R46563 vdd.n1433 vdd.n1432 0.0130799
R46564 vdd.n1438 vdd.n1434 0.0130799
R46565 vdd.n1453 vdd.n1452 0.0130799
R46566 vdd.n1528 vdd.n1521 0.0130799
R46567 vdd.n1528 vdd.n1526 0.0130799
R46568 vdd.n1552 vdd.n1551 0.0130799
R46569 vdd.n1551 vdd.n1527 0.0130799
R46570 vdd.n1536 vdd.n1534 0.0130799
R46571 vdd.n1534 vdd.n1533 0.0130799
R46572 vdd.n1539 vdd.n1535 0.0130799
R46573 vdd.n1554 vdd.n1553 0.0130799
R46574 vdd.n641 vdd.n634 0.0130799
R46575 vdd.n641 vdd.n639 0.0130799
R46576 vdd.n665 vdd.n664 0.0130799
R46577 vdd.n664 vdd.n640 0.0130799
R46578 vdd.n649 vdd.n647 0.0130799
R46579 vdd.n647 vdd.n646 0.0130799
R46580 vdd.n652 vdd.n648 0.0130799
R46581 vdd.n667 vdd.n666 0.0130799
R46582 vdd.n1576 vdd.n1569 0.0130799
R46583 vdd.n1576 vdd.n1574 0.0130799
R46584 vdd.n1600 vdd.n1599 0.0130799
R46585 vdd.n1599 vdd.n1575 0.0130799
R46586 vdd.n1584 vdd.n1582 0.0130799
R46587 vdd.n1582 vdd.n1581 0.0130799
R46588 vdd.n1587 vdd.n1583 0.0130799
R46589 vdd.n1602 vdd.n1601 0.0130799
R46590 vdd.n1623 vdd.n1616 0.0130799
R46591 vdd.n1623 vdd.n1621 0.0130799
R46592 vdd.n1647 vdd.n1646 0.0130799
R46593 vdd.n1646 vdd.n1622 0.0130799
R46594 vdd.n1631 vdd.n1629 0.0130799
R46595 vdd.n1629 vdd.n1628 0.0130799
R46596 vdd.n1634 vdd.n1630 0.0130799
R46597 vdd.n1649 vdd.n1648 0.0130799
R46598 vdd.n1673 vdd.n1666 0.0130799
R46599 vdd.n1673 vdd.n1671 0.0130799
R46600 vdd.n1697 vdd.n1696 0.0130799
R46601 vdd.n1696 vdd.n1672 0.0130799
R46602 vdd.n1681 vdd.n1679 0.0130799
R46603 vdd.n1679 vdd.n1678 0.0130799
R46604 vdd.n1684 vdd.n1680 0.0130799
R46605 vdd.n1699 vdd.n1698 0.0130799
R46606 vdd.n1723 vdd.n1716 0.0130799
R46607 vdd.n1723 vdd.n1721 0.0130799
R46608 vdd.n1747 vdd.n1746 0.0130799
R46609 vdd.n1746 vdd.n1722 0.0130799
R46610 vdd.n1731 vdd.n1729 0.0130799
R46611 vdd.n1729 vdd.n1728 0.0130799
R46612 vdd.n1734 vdd.n1730 0.0130799
R46613 vdd.n1749 vdd.n1748 0.0130799
R46614 vdd.n1771 vdd.n1764 0.0130799
R46615 vdd.n1771 vdd.n1769 0.0130799
R46616 vdd.n1795 vdd.n1794 0.0130799
R46617 vdd.n1794 vdd.n1770 0.0130799
R46618 vdd.n1779 vdd.n1777 0.0130799
R46619 vdd.n1777 vdd.n1776 0.0130799
R46620 vdd.n1782 vdd.n1778 0.0130799
R46621 vdd.n1797 vdd.n1796 0.0130799
R46622 vdd.n1503 vdd.n1502 0.0130799
R46623 vdd.n1502 vdd.n1480 0.0130799
R46624 vdd.n1486 vdd.n1485 0.0130799
R46625 vdd.n1485 vdd.n1483 0.0130799
R46626 vdd.n1477 vdd.n1476 0.0130799
R46627 vdd.n1476 vdd.n1474 0.0130799
R46628 vdd.n1472 vdd.n1470 0.0130799
R46629 vdd.n1488 vdd.n1487 0.0130799
R46630 vdd.n1822 vdd.n1815 0.0130799
R46631 vdd.n1822 vdd.n1820 0.0130799
R46632 vdd.n1846 vdd.n1845 0.0130799
R46633 vdd.n1845 vdd.n1821 0.0130799
R46634 vdd.n1830 vdd.n1828 0.0130799
R46635 vdd.n1828 vdd.n1827 0.0130799
R46636 vdd.n1833 vdd.n1829 0.0130799
R46637 vdd.n1848 vdd.n1847 0.0130799
R46638 vdd.n1869 vdd.n1862 0.0130799
R46639 vdd.n1869 vdd.n1867 0.0130799
R46640 vdd.n1893 vdd.n1892 0.0130799
R46641 vdd.n1892 vdd.n1868 0.0130799
R46642 vdd.n1877 vdd.n1875 0.0130799
R46643 vdd.n1875 vdd.n1874 0.0130799
R46644 vdd.n1880 vdd.n1876 0.0130799
R46645 vdd.n1895 vdd.n1894 0.0130799
R46646 vdd.n1917 vdd.n1910 0.0130799
R46647 vdd.n1917 vdd.n1915 0.0130799
R46648 vdd.n1941 vdd.n1940 0.0130799
R46649 vdd.n1940 vdd.n1916 0.0130799
R46650 vdd.n1925 vdd.n1923 0.0130799
R46651 vdd.n1923 vdd.n1922 0.0130799
R46652 vdd.n1928 vdd.n1924 0.0130799
R46653 vdd.n1943 vdd.n1942 0.0130799
R46654 vdd.n1968 vdd.n1961 0.0130799
R46655 vdd.n1968 vdd.n1966 0.0130799
R46656 vdd.n1992 vdd.n1991 0.0130799
R46657 vdd.n1991 vdd.n1967 0.0130799
R46658 vdd.n1976 vdd.n1974 0.0130799
R46659 vdd.n1974 vdd.n1973 0.0130799
R46660 vdd.n1979 vdd.n1975 0.0130799
R46661 vdd.n1994 vdd.n1993 0.0130799
R46662 vdd.n2018 vdd.n2011 0.0130799
R46663 vdd.n2018 vdd.n2016 0.0130799
R46664 vdd.n2042 vdd.n2041 0.0130799
R46665 vdd.n2041 vdd.n2017 0.0130799
R46666 vdd.n2026 vdd.n2024 0.0130799
R46667 vdd.n2024 vdd.n2023 0.0130799
R46668 vdd.n2029 vdd.n2025 0.0130799
R46669 vdd.n2044 vdd.n2043 0.0130799
R46670 vdd.n2066 vdd.n2059 0.0130799
R46671 vdd.n2066 vdd.n2064 0.0130799
R46672 vdd.n2090 vdd.n2089 0.0130799
R46673 vdd.n2089 vdd.n2065 0.0130799
R46674 vdd.n2074 vdd.n2072 0.0130799
R46675 vdd.n2072 vdd.n2071 0.0130799
R46676 vdd.n2077 vdd.n2073 0.0130799
R46677 vdd.n2092 vdd.n2091 0.0130799
R46678 vdd.n2116 vdd.n2109 0.0130799
R46679 vdd.n2116 vdd.n2114 0.0130799
R46680 vdd.n2140 vdd.n2139 0.0130799
R46681 vdd.n2139 vdd.n2115 0.0130799
R46682 vdd.n2124 vdd.n2122 0.0130799
R46683 vdd.n2122 vdd.n2121 0.0130799
R46684 vdd.n2127 vdd.n2123 0.0130799
R46685 vdd.n2142 vdd.n2141 0.0130799
R46686 vdd.n2163 vdd.n2156 0.0130799
R46687 vdd.n2163 vdd.n2161 0.0130799
R46688 vdd.n2187 vdd.n2186 0.0130799
R46689 vdd.n2186 vdd.n2162 0.0130799
R46690 vdd.n2171 vdd.n2169 0.0130799
R46691 vdd.n2169 vdd.n2168 0.0130799
R46692 vdd.n2174 vdd.n2170 0.0130799
R46693 vdd.n2189 vdd.n2188 0.0130799
R46694 vdd.n2213 vdd.n2206 0.0130799
R46695 vdd.n2213 vdd.n2211 0.0130799
R46696 vdd.n2237 vdd.n2236 0.0130799
R46697 vdd.n2236 vdd.n2212 0.0130799
R46698 vdd.n2221 vdd.n2219 0.0130799
R46699 vdd.n2219 vdd.n2218 0.0130799
R46700 vdd.n2224 vdd.n2220 0.0130799
R46701 vdd.n2239 vdd.n2238 0.0130799
R46702 vdd.n2263 vdd.n2256 0.0130799
R46703 vdd.n2263 vdd.n2261 0.0130799
R46704 vdd.n2287 vdd.n2286 0.0130799
R46705 vdd.n2286 vdd.n2262 0.0130799
R46706 vdd.n2271 vdd.n2269 0.0130799
R46707 vdd.n2269 vdd.n2268 0.0130799
R46708 vdd.n2274 vdd.n2270 0.0130799
R46709 vdd.n2289 vdd.n2288 0.0130799
R46710 vdd.n2311 vdd.n2304 0.0130799
R46711 vdd.n2311 vdd.n2309 0.0130799
R46712 vdd.n2335 vdd.n2334 0.0130799
R46713 vdd.n2334 vdd.n2310 0.0130799
R46714 vdd.n2319 vdd.n2317 0.0130799
R46715 vdd.n2317 vdd.n2316 0.0130799
R46716 vdd.n2322 vdd.n2318 0.0130799
R46717 vdd.n2337 vdd.n2336 0.0130799
R46718 vdd.n1258 vdd.n1257 0.0130799
R46719 vdd.n1257 vdd.n1235 0.0130799
R46720 vdd.n1241 vdd.n1240 0.0130799
R46721 vdd.n1240 vdd.n1238 0.0130799
R46722 vdd.n1232 vdd.n1231 0.0130799
R46723 vdd.n1231 vdd.n1229 0.0130799
R46724 vdd.n1227 vdd.n1225 0.0130799
R46725 vdd.n1243 vdd.n1242 0.0130799
R46726 vdd.n2362 vdd.n2355 0.0130799
R46727 vdd.n2362 vdd.n2360 0.0130799
R46728 vdd.n2386 vdd.n2385 0.0130799
R46729 vdd.n2385 vdd.n2361 0.0130799
R46730 vdd.n2370 vdd.n2368 0.0130799
R46731 vdd.n2368 vdd.n2367 0.0130799
R46732 vdd.n2373 vdd.n2369 0.0130799
R46733 vdd.n2388 vdd.n2387 0.0130799
R46734 vdd.n2409 vdd.n2402 0.0130799
R46735 vdd.n2409 vdd.n2407 0.0130799
R46736 vdd.n2433 vdd.n2432 0.0130799
R46737 vdd.n2432 vdd.n2408 0.0130799
R46738 vdd.n2417 vdd.n2415 0.0130799
R46739 vdd.n2415 vdd.n2414 0.0130799
R46740 vdd.n2420 vdd.n2416 0.0130799
R46741 vdd.n2435 vdd.n2434 0.0130799
R46742 vdd.n2459 vdd.n2452 0.0130799
R46743 vdd.n2459 vdd.n2457 0.0130799
R46744 vdd.n2483 vdd.n2482 0.0130799
R46745 vdd.n2482 vdd.n2458 0.0130799
R46746 vdd.n2467 vdd.n2465 0.0130799
R46747 vdd.n2465 vdd.n2464 0.0130799
R46748 vdd.n2470 vdd.n2466 0.0130799
R46749 vdd.n2485 vdd.n2484 0.0130799
R46750 vdd.n2509 vdd.n2502 0.0130799
R46751 vdd.n2509 vdd.n2507 0.0130799
R46752 vdd.n2533 vdd.n2532 0.0130799
R46753 vdd.n2532 vdd.n2508 0.0130799
R46754 vdd.n2517 vdd.n2515 0.0130799
R46755 vdd.n2515 vdd.n2514 0.0130799
R46756 vdd.n2520 vdd.n2516 0.0130799
R46757 vdd.n2535 vdd.n2534 0.0130799
R46758 vdd.n2557 vdd.n2550 0.0130799
R46759 vdd.n2557 vdd.n2555 0.0130799
R46760 vdd.n2581 vdd.n2580 0.0130799
R46761 vdd.n2580 vdd.n2556 0.0130799
R46762 vdd.n2565 vdd.n2563 0.0130799
R46763 vdd.n2563 vdd.n2562 0.0130799
R46764 vdd.n2568 vdd.n2564 0.0130799
R46765 vdd.n2583 vdd.n2582 0.0130799
R46766 vdd.n2703 vdd.n2696 0.0130799
R46767 vdd.n2703 vdd.n2701 0.0130799
R46768 vdd.n2716 vdd.n2709 0.0130799
R46769 vdd.n2709 vdd.n2708 0.0130799
R46770 vdd.n2727 vdd.n2726 0.0130799
R46771 vdd.n2726 vdd.n2702 0.0130799
R46772 vdd.n2729 vdd.n2728 0.0130799
R46773 vdd.n2715 vdd.n2714 0.0130799
R46774 vdd.n2655 vdd.n2648 0.0130799
R46775 vdd.n2655 vdd.n2653 0.0130799
R46776 vdd.n2668 vdd.n2661 0.0130799
R46777 vdd.n2661 vdd.n2660 0.0130799
R46778 vdd.n2679 vdd.n2678 0.0130799
R46779 vdd.n2678 vdd.n2654 0.0130799
R46780 vdd.n2681 vdd.n2680 0.0130799
R46781 vdd.n2667 vdd.n2666 0.0130799
R46782 vdd.n2752 vdd.n2745 0.0130799
R46783 vdd.n2752 vdd.n2750 0.0130799
R46784 vdd.n2765 vdd.n2758 0.0130799
R46785 vdd.n2758 vdd.n2757 0.0130799
R46786 vdd.n2776 vdd.n2775 0.0130799
R46787 vdd.n2775 vdd.n2751 0.0130799
R46788 vdd.n2778 vdd.n2777 0.0130799
R46789 vdd.n2764 vdd.n2763 0.0130799
R46790 vdd.n2802 vdd.n2795 0.0130799
R46791 vdd.n2802 vdd.n2800 0.0130799
R46792 vdd.n2815 vdd.n2808 0.0130799
R46793 vdd.n2808 vdd.n2807 0.0130799
R46794 vdd.n2826 vdd.n2825 0.0130799
R46795 vdd.n2825 vdd.n2801 0.0130799
R46796 vdd.n2828 vdd.n2827 0.0130799
R46797 vdd.n2814 vdd.n2813 0.0130799
R46798 vdd.n2850 vdd.n2843 0.0130799
R46799 vdd.n2850 vdd.n2848 0.0130799
R46800 vdd.n2863 vdd.n2856 0.0130799
R46801 vdd.n2856 vdd.n2855 0.0130799
R46802 vdd.n2874 vdd.n2873 0.0130799
R46803 vdd.n2873 vdd.n2849 0.0130799
R46804 vdd.n2876 vdd.n2875 0.0130799
R46805 vdd.n2862 vdd.n2861 0.0130799
R46806 vdd.n1061 vdd.n1060 0.0130799
R46807 vdd.n1060 vdd.n1059 0.0130799
R46808 vdd.n1042 vdd.n1039 0.0130799
R46809 vdd.n1042 vdd.n1036 0.0130799
R46810 vdd.n1066 vdd.n1065 0.0130799
R46811 vdd.n1066 vdd.n1031 0.0130799
R46812 vdd.n1073 vdd.n1028 0.0130799
R46813 vdd.n1041 vdd.n1040 0.0130799
R46814 vdd.n2998 vdd.n2991 0.0130799
R46815 vdd.n2998 vdd.n2996 0.0130799
R46816 vdd.n3011 vdd.n3004 0.0130799
R46817 vdd.n3004 vdd.n3003 0.0130799
R46818 vdd.n3022 vdd.n3021 0.0130799
R46819 vdd.n3021 vdd.n2997 0.0130799
R46820 vdd.n3024 vdd.n3023 0.0130799
R46821 vdd.n3010 vdd.n3009 0.0130799
R46822 vdd.n2949 vdd.n2942 0.0130799
R46823 vdd.n2949 vdd.n2947 0.0130799
R46824 vdd.n2962 vdd.n2955 0.0130799
R46825 vdd.n2955 vdd.n2954 0.0130799
R46826 vdd.n2973 vdd.n2972 0.0130799
R46827 vdd.n2972 vdd.n2948 0.0130799
R46828 vdd.n2975 vdd.n2974 0.0130799
R46829 vdd.n2961 vdd.n2960 0.0130799
R46830 vdd.n2901 vdd.n2894 0.0130799
R46831 vdd.n2901 vdd.n2899 0.0130799
R46832 vdd.n2914 vdd.n2907 0.0130799
R46833 vdd.n2907 vdd.n2906 0.0130799
R46834 vdd.n2925 vdd.n2924 0.0130799
R46835 vdd.n2924 vdd.n2900 0.0130799
R46836 vdd.n2927 vdd.n2926 0.0130799
R46837 vdd.n2913 vdd.n2912 0.0130799
R46838 vdd.n3047 vdd.n3040 0.0130799
R46839 vdd.n3047 vdd.n3045 0.0130799
R46840 vdd.n3060 vdd.n3053 0.0130799
R46841 vdd.n3053 vdd.n3052 0.0130799
R46842 vdd.n3071 vdd.n3070 0.0130799
R46843 vdd.n3070 vdd.n3046 0.0130799
R46844 vdd.n3073 vdd.n3072 0.0130799
R46845 vdd.n3059 vdd.n3058 0.0130799
R46846 vdd.n3097 vdd.n3090 0.0130799
R46847 vdd.n3097 vdd.n3095 0.0130799
R46848 vdd.n3110 vdd.n3103 0.0130799
R46849 vdd.n3103 vdd.n3102 0.0130799
R46850 vdd.n3121 vdd.n3120 0.0130799
R46851 vdd.n3120 vdd.n3096 0.0130799
R46852 vdd.n3123 vdd.n3122 0.0130799
R46853 vdd.n3109 vdd.n3108 0.0130799
R46854 vdd.n3145 vdd.n3138 0.0130799
R46855 vdd.n3145 vdd.n3143 0.0130799
R46856 vdd.n3158 vdd.n3151 0.0130799
R46857 vdd.n3151 vdd.n3150 0.0130799
R46858 vdd.n3169 vdd.n3168 0.0130799
R46859 vdd.n3168 vdd.n3144 0.0130799
R46860 vdd.n3171 vdd.n3170 0.0130799
R46861 vdd.n3157 vdd.n3156 0.0130799
R46862 vdd.n3243 vdd.n3236 0.0130799
R46863 vdd.n3243 vdd.n3241 0.0130799
R46864 vdd.n3256 vdd.n3249 0.0130799
R46865 vdd.n3249 vdd.n3248 0.0130799
R46866 vdd.n3267 vdd.n3266 0.0130799
R46867 vdd.n3266 vdd.n3242 0.0130799
R46868 vdd.n3269 vdd.n3268 0.0130799
R46869 vdd.n3255 vdd.n3254 0.0130799
R46870 vdd.n3195 vdd.n3188 0.0130799
R46871 vdd.n3195 vdd.n3193 0.0130799
R46872 vdd.n3208 vdd.n3201 0.0130799
R46873 vdd.n3201 vdd.n3200 0.0130799
R46874 vdd.n3219 vdd.n3218 0.0130799
R46875 vdd.n3218 vdd.n3194 0.0130799
R46876 vdd.n3221 vdd.n3220 0.0130799
R46877 vdd.n3207 vdd.n3206 0.0130799
R46878 vdd.n3292 vdd.n3285 0.0130799
R46879 vdd.n3292 vdd.n3290 0.0130799
R46880 vdd.n3305 vdd.n3298 0.0130799
R46881 vdd.n3298 vdd.n3297 0.0130799
R46882 vdd.n3316 vdd.n3315 0.0130799
R46883 vdd.n3315 vdd.n3291 0.0130799
R46884 vdd.n3318 vdd.n3317 0.0130799
R46885 vdd.n3304 vdd.n3303 0.0130799
R46886 vdd.n3342 vdd.n3335 0.0130799
R46887 vdd.n3342 vdd.n3340 0.0130799
R46888 vdd.n3355 vdd.n3348 0.0130799
R46889 vdd.n3348 vdd.n3347 0.0130799
R46890 vdd.n3366 vdd.n3365 0.0130799
R46891 vdd.n3365 vdd.n3341 0.0130799
R46892 vdd.n3368 vdd.n3367 0.0130799
R46893 vdd.n3354 vdd.n3353 0.0130799
R46894 vdd.n3390 vdd.n3383 0.0130799
R46895 vdd.n3390 vdd.n3388 0.0130799
R46896 vdd.n3403 vdd.n3396 0.0130799
R46897 vdd.n3396 vdd.n3395 0.0130799
R46898 vdd.n3414 vdd.n3413 0.0130799
R46899 vdd.n3413 vdd.n3389 0.0130799
R46900 vdd.n3416 vdd.n3415 0.0130799
R46901 vdd.n3402 vdd.n3401 0.0130799
R46902 vdd.n815 vdd.n814 0.0130799
R46903 vdd.n814 vdd.n813 0.0130799
R46904 vdd.n796 vdd.n793 0.0130799
R46905 vdd.n796 vdd.n790 0.0130799
R46906 vdd.n820 vdd.n819 0.0130799
R46907 vdd.n820 vdd.n785 0.0130799
R46908 vdd.n827 vdd.n782 0.0130799
R46909 vdd.n795 vdd.n794 0.0130799
R46910 vdd.n3489 vdd.n3482 0.0130799
R46911 vdd.n3489 vdd.n3487 0.0130799
R46912 vdd.n3502 vdd.n3495 0.0130799
R46913 vdd.n3495 vdd.n3494 0.0130799
R46914 vdd.n3513 vdd.n3512 0.0130799
R46915 vdd.n3512 vdd.n3488 0.0130799
R46916 vdd.n3515 vdd.n3514 0.0130799
R46917 vdd.n3501 vdd.n3500 0.0130799
R46918 vdd.n3441 vdd.n3434 0.0130799
R46919 vdd.n3441 vdd.n3439 0.0130799
R46920 vdd.n3454 vdd.n3447 0.0130799
R46921 vdd.n3447 vdd.n3446 0.0130799
R46922 vdd.n3465 vdd.n3464 0.0130799
R46923 vdd.n3464 vdd.n3440 0.0130799
R46924 vdd.n3467 vdd.n3466 0.0130799
R46925 vdd.n3453 vdd.n3452 0.0130799
R46926 vdd.n3538 vdd.n3531 0.0130799
R46927 vdd.n3538 vdd.n3536 0.0130799
R46928 vdd.n3551 vdd.n3544 0.0130799
R46929 vdd.n3544 vdd.n3543 0.0130799
R46930 vdd.n3562 vdd.n3561 0.0130799
R46931 vdd.n3561 vdd.n3537 0.0130799
R46932 vdd.n3564 vdd.n3563 0.0130799
R46933 vdd.n3550 vdd.n3549 0.0130799
R46934 vdd.n3588 vdd.n3581 0.0130799
R46935 vdd.n3588 vdd.n3586 0.0130799
R46936 vdd.n3601 vdd.n3594 0.0130799
R46937 vdd.n3594 vdd.n3593 0.0130799
R46938 vdd.n3612 vdd.n3611 0.0130799
R46939 vdd.n3611 vdd.n3587 0.0130799
R46940 vdd.n3614 vdd.n3613 0.0130799
R46941 vdd.n3600 vdd.n3599 0.0130799
R46942 vdd.n3636 vdd.n3629 0.0130799
R46943 vdd.n3636 vdd.n3634 0.0130799
R46944 vdd.n3649 vdd.n3642 0.0130799
R46945 vdd.n3642 vdd.n3641 0.0130799
R46946 vdd.n3660 vdd.n3659 0.0130799
R46947 vdd.n3659 vdd.n3635 0.0130799
R46948 vdd.n3662 vdd.n3661 0.0130799
R46949 vdd.n3648 vdd.n3647 0.0130799
R46950 vdd.n594 vdd.n587 0.0130799
R46951 vdd.n594 vdd.n592 0.0130799
R46952 vdd.n607 vdd.n600 0.0130799
R46953 vdd.n600 vdd.n599 0.0130799
R46954 vdd.n618 vdd.n617 0.0130799
R46955 vdd.n617 vdd.n593 0.0130799
R46956 vdd.n620 vdd.n619 0.0130799
R46957 vdd.n606 vdd.n605 0.0130799
R46958 vdd.n3735 vdd.n3728 0.0130799
R46959 vdd.n3735 vdd.n3733 0.0130799
R46960 vdd.n3748 vdd.n3741 0.0130799
R46961 vdd.n3741 vdd.n3740 0.0130799
R46962 vdd.n3759 vdd.n3758 0.0130799
R46963 vdd.n3758 vdd.n3734 0.0130799
R46964 vdd.n3761 vdd.n3760 0.0130799
R46965 vdd.n3747 vdd.n3746 0.0130799
R46966 vdd.n3687 vdd.n3680 0.0130799
R46967 vdd.n3687 vdd.n3685 0.0130799
R46968 vdd.n3700 vdd.n3693 0.0130799
R46969 vdd.n3693 vdd.n3692 0.0130799
R46970 vdd.n3711 vdd.n3710 0.0130799
R46971 vdd.n3710 vdd.n3686 0.0130799
R46972 vdd.n3713 vdd.n3712 0.0130799
R46973 vdd.n3699 vdd.n3698 0.0130799
R46974 vdd.n6877 vdd.n6870 0.0130799
R46975 vdd.n6877 vdd.n6875 0.0130799
R46976 vdd.n6890 vdd.n6883 0.0130799
R46977 vdd.n6883 vdd.n6882 0.0130799
R46978 vdd.n6901 vdd.n6900 0.0130799
R46979 vdd.n6900 vdd.n6876 0.0130799
R46980 vdd.n6903 vdd.n6902 0.0130799
R46981 vdd.n6889 vdd.n6888 0.0130799
R46982 vdd.n6829 vdd.n6822 0.0130799
R46983 vdd.n6829 vdd.n6827 0.0130799
R46984 vdd.n6842 vdd.n6835 0.0130799
R46985 vdd.n6835 vdd.n6834 0.0130799
R46986 vdd.n6853 vdd.n6852 0.0130799
R46987 vdd.n6852 vdd.n6828 0.0130799
R46988 vdd.n6855 vdd.n6854 0.0130799
R46989 vdd.n6841 vdd.n6840 0.0130799
R46990 vdd.n10019 vdd.n10012 0.0130799
R46991 vdd.n10019 vdd.n10017 0.0130799
R46992 vdd.n10032 vdd.n10025 0.0130799
R46993 vdd.n10025 vdd.n10024 0.0130799
R46994 vdd.n10043 vdd.n10042 0.0130799
R46995 vdd.n10042 vdd.n10018 0.0130799
R46996 vdd.n10045 vdd.n10044 0.0130799
R46997 vdd.n10031 vdd.n10030 0.0130799
R46998 vdd.n9971 vdd.n9964 0.0130799
R46999 vdd.n9971 vdd.n9969 0.0130799
R47000 vdd.n9984 vdd.n9977 0.0130799
R47001 vdd.n9977 vdd.n9976 0.0130799
R47002 vdd.n9995 vdd.n9994 0.0130799
R47003 vdd.n9994 vdd.n9970 0.0130799
R47004 vdd.n9997 vdd.n9996 0.0130799
R47005 vdd.n9983 vdd.n9982 0.0130799
R47006 vdd.n10067 vdd.n10060 0.0130799
R47007 vdd.n10067 vdd.n10065 0.0130799
R47008 vdd.n10080 vdd.n10073 0.0130799
R47009 vdd.n10073 vdd.n10072 0.0130799
R47010 vdd.n10091 vdd.n10090 0.0130799
R47011 vdd.n10090 vdd.n10066 0.0130799
R47012 vdd.n10093 vdd.n10092 0.0130799
R47013 vdd.n10079 vdd.n10078 0.0130799
R47014 vdd.n10115 vdd.n10108 0.0130799
R47015 vdd.n10115 vdd.n10113 0.0130799
R47016 vdd.n10128 vdd.n10121 0.0130799
R47017 vdd.n10121 vdd.n10120 0.0130799
R47018 vdd.n10139 vdd.n10138 0.0130799
R47019 vdd.n10138 vdd.n10114 0.0130799
R47020 vdd.n10141 vdd.n10140 0.0130799
R47021 vdd.n10127 vdd.n10126 0.0130799
R47022 vdd.n10217 vdd.n10210 0.0130799
R47023 vdd.n10217 vdd.n10215 0.0130799
R47024 vdd.n10230 vdd.n10223 0.0130799
R47025 vdd.n10223 vdd.n10222 0.0130799
R47026 vdd.n10241 vdd.n10240 0.0130799
R47027 vdd.n10240 vdd.n10216 0.0130799
R47028 vdd.n10243 vdd.n10242 0.0130799
R47029 vdd.n10229 vdd.n10228 0.0130799
R47030 vdd.n10265 vdd.n10258 0.0130799
R47031 vdd.n10265 vdd.n10263 0.0130799
R47032 vdd.n10278 vdd.n10271 0.0130799
R47033 vdd.n10271 vdd.n10270 0.0130799
R47034 vdd.n10289 vdd.n10288 0.0130799
R47035 vdd.n10288 vdd.n10264 0.0130799
R47036 vdd.n10291 vdd.n10290 0.0130799
R47037 vdd.n10277 vdd.n10276 0.0130799
R47038 vdd.n10313 vdd.n10306 0.0130799
R47039 vdd.n10313 vdd.n10311 0.0130799
R47040 vdd.n10326 vdd.n10319 0.0130799
R47041 vdd.n10319 vdd.n10318 0.0130799
R47042 vdd.n10337 vdd.n10336 0.0130799
R47043 vdd.n10336 vdd.n10312 0.0130799
R47044 vdd.n10339 vdd.n10338 0.0130799
R47045 vdd.n10325 vdd.n10324 0.0130799
R47046 vdd.n10361 vdd.n10354 0.0130799
R47047 vdd.n10361 vdd.n10359 0.0130799
R47048 vdd.n10374 vdd.n10367 0.0130799
R47049 vdd.n10367 vdd.n10366 0.0130799
R47050 vdd.n10385 vdd.n10384 0.0130799
R47051 vdd.n10384 vdd.n10360 0.0130799
R47052 vdd.n10387 vdd.n10386 0.0130799
R47053 vdd.n10373 vdd.n10372 0.0130799
R47054 vdd.n10463 vdd.n10456 0.0130799
R47055 vdd.n10463 vdd.n10461 0.0130799
R47056 vdd.n10476 vdd.n10469 0.0130799
R47057 vdd.n10469 vdd.n10468 0.0130799
R47058 vdd.n10487 vdd.n10486 0.0130799
R47059 vdd.n10486 vdd.n10462 0.0130799
R47060 vdd.n10489 vdd.n10488 0.0130799
R47061 vdd.n10475 vdd.n10474 0.0130799
R47062 vdd.n55 vdd.n48 0.0130799
R47063 vdd.n55 vdd.n53 0.0130799
R47064 vdd.n68 vdd.n61 0.0130799
R47065 vdd.n61 vdd.n60 0.0130799
R47066 vdd.n79 vdd.n78 0.0130799
R47067 vdd.n78 vdd.n54 0.0130799
R47068 vdd.n81 vdd.n80 0.0130799
R47069 vdd.n67 vdd.n66 0.0130799
R47070 vdd.n7 vdd.n0 0.0130799
R47071 vdd.n7 vdd.n5 0.0130799
R47072 vdd.n20 vdd.n13 0.0130799
R47073 vdd.n13 vdd.n12 0.0130799
R47074 vdd.n31 vdd.n30 0.0130799
R47075 vdd.n30 vdd.n6 0.0130799
R47076 vdd.n33 vdd.n32 0.0130799
R47077 vdd.n19 vdd.n18 0.0130799
R47078 vdd.n10511 vdd.n10504 0.0130799
R47079 vdd.n10511 vdd.n10509 0.0130799
R47080 vdd.n10524 vdd.n10517 0.0130799
R47081 vdd.n10517 vdd.n10516 0.0130799
R47082 vdd.n10535 vdd.n10534 0.0130799
R47083 vdd.n10534 vdd.n10510 0.0130799
R47084 vdd.n10537 vdd.n10536 0.0130799
R47085 vdd.n10523 vdd.n10522 0.0130799
R47086 vdd.n10561 vdd.n10554 0.0130799
R47087 vdd.n10561 vdd.n10559 0.0130799
R47088 vdd.n10574 vdd.n10567 0.0130799
R47089 vdd.n10567 vdd.n10566 0.0130799
R47090 vdd.n10585 vdd.n10584 0.0130799
R47091 vdd.n10584 vdd.n10560 0.0130799
R47092 vdd.n10587 vdd.n10586 0.0130799
R47093 vdd.n10573 vdd.n10572 0.0130799
R47094 vdd.n10609 vdd.n10602 0.0130799
R47095 vdd.n10609 vdd.n10607 0.0130799
R47096 vdd.n10622 vdd.n10615 0.0130799
R47097 vdd.n10615 vdd.n10614 0.0130799
R47098 vdd.n10633 vdd.n10632 0.0130799
R47099 vdd.n10632 vdd.n10608 0.0130799
R47100 vdd.n10635 vdd.n10634 0.0130799
R47101 vdd.n10621 vdd.n10620 0.0130799
R47102 vdd.n10438 vdd.n10437 0.0130799
R47103 vdd.n10437 vdd.n10436 0.0130799
R47104 vdd.n10419 vdd.n10416 0.0130799
R47105 vdd.n10419 vdd.n10413 0.0130799
R47106 vdd.n10443 vdd.n10442 0.0130799
R47107 vdd.n10443 vdd.n10408 0.0130799
R47108 vdd.n10450 vdd.n10405 0.0130799
R47109 vdd.n10418 vdd.n10417 0.0130799
R47110 vdd.n10757 vdd.n10750 0.0130799
R47111 vdd.n10757 vdd.n10755 0.0130799
R47112 vdd.n10770 vdd.n10763 0.0130799
R47113 vdd.n10763 vdd.n10762 0.0130799
R47114 vdd.n10781 vdd.n10780 0.0130799
R47115 vdd.n10780 vdd.n10756 0.0130799
R47116 vdd.n10783 vdd.n10782 0.0130799
R47117 vdd.n10769 vdd.n10768 0.0130799
R47118 vdd.n10708 vdd.n10701 0.0130799
R47119 vdd.n10708 vdd.n10706 0.0130799
R47120 vdd.n10721 vdd.n10714 0.0130799
R47121 vdd.n10714 vdd.n10713 0.0130799
R47122 vdd.n10732 vdd.n10731 0.0130799
R47123 vdd.n10731 vdd.n10707 0.0130799
R47124 vdd.n10734 vdd.n10733 0.0130799
R47125 vdd.n10720 vdd.n10719 0.0130799
R47126 vdd.n10660 vdd.n10653 0.0130799
R47127 vdd.n10660 vdd.n10658 0.0130799
R47128 vdd.n10673 vdd.n10666 0.0130799
R47129 vdd.n10666 vdd.n10665 0.0130799
R47130 vdd.n10684 vdd.n10683 0.0130799
R47131 vdd.n10683 vdd.n10659 0.0130799
R47132 vdd.n10686 vdd.n10685 0.0130799
R47133 vdd.n10672 vdd.n10671 0.0130799
R47134 vdd.n10806 vdd.n10799 0.0130799
R47135 vdd.n10806 vdd.n10804 0.0130799
R47136 vdd.n10819 vdd.n10812 0.0130799
R47137 vdd.n10812 vdd.n10811 0.0130799
R47138 vdd.n10830 vdd.n10829 0.0130799
R47139 vdd.n10829 vdd.n10805 0.0130799
R47140 vdd.n10832 vdd.n10831 0.0130799
R47141 vdd.n10818 vdd.n10817 0.0130799
R47142 vdd.n10856 vdd.n10849 0.0130799
R47143 vdd.n10856 vdd.n10854 0.0130799
R47144 vdd.n10869 vdd.n10862 0.0130799
R47145 vdd.n10862 vdd.n10861 0.0130799
R47146 vdd.n10880 vdd.n10879 0.0130799
R47147 vdd.n10879 vdd.n10855 0.0130799
R47148 vdd.n10882 vdd.n10881 0.0130799
R47149 vdd.n10868 vdd.n10867 0.0130799
R47150 vdd.n10904 vdd.n10897 0.0130799
R47151 vdd.n10904 vdd.n10902 0.0130799
R47152 vdd.n10917 vdd.n10910 0.0130799
R47153 vdd.n10910 vdd.n10909 0.0130799
R47154 vdd.n10928 vdd.n10927 0.0130799
R47155 vdd.n10927 vdd.n10903 0.0130799
R47156 vdd.n10930 vdd.n10929 0.0130799
R47157 vdd.n10916 vdd.n10915 0.0130799
R47158 vdd.n11002 vdd.n10995 0.0130799
R47159 vdd.n11002 vdd.n11000 0.0130799
R47160 vdd.n11015 vdd.n11008 0.0130799
R47161 vdd.n11008 vdd.n11007 0.0130799
R47162 vdd.n11026 vdd.n11025 0.0130799
R47163 vdd.n11025 vdd.n11001 0.0130799
R47164 vdd.n11028 vdd.n11027 0.0130799
R47165 vdd.n11014 vdd.n11013 0.0130799
R47166 vdd.n10954 vdd.n10947 0.0130799
R47167 vdd.n10954 vdd.n10952 0.0130799
R47168 vdd.n10967 vdd.n10960 0.0130799
R47169 vdd.n10960 vdd.n10959 0.0130799
R47170 vdd.n10978 vdd.n10977 0.0130799
R47171 vdd.n10977 vdd.n10953 0.0130799
R47172 vdd.n10980 vdd.n10979 0.0130799
R47173 vdd.n10966 vdd.n10965 0.0130799
R47174 vdd.n11051 vdd.n11044 0.0130799
R47175 vdd.n11051 vdd.n11049 0.0130799
R47176 vdd.n11064 vdd.n11057 0.0130799
R47177 vdd.n11057 vdd.n11056 0.0130799
R47178 vdd.n11075 vdd.n11074 0.0130799
R47179 vdd.n11074 vdd.n11050 0.0130799
R47180 vdd.n11077 vdd.n11076 0.0130799
R47181 vdd.n11063 vdd.n11062 0.0130799
R47182 vdd.n11101 vdd.n11094 0.0130799
R47183 vdd.n11101 vdd.n11099 0.0130799
R47184 vdd.n11114 vdd.n11107 0.0130799
R47185 vdd.n11107 vdd.n11106 0.0130799
R47186 vdd.n11125 vdd.n11124 0.0130799
R47187 vdd.n11124 vdd.n11100 0.0130799
R47188 vdd.n11127 vdd.n11126 0.0130799
R47189 vdd.n11113 vdd.n11112 0.0130799
R47190 vdd.n11149 vdd.n11142 0.0130799
R47191 vdd.n11149 vdd.n11147 0.0130799
R47192 vdd.n11162 vdd.n11155 0.0130799
R47193 vdd.n11155 vdd.n11154 0.0130799
R47194 vdd.n11173 vdd.n11172 0.0130799
R47195 vdd.n11172 vdd.n11148 0.0130799
R47196 vdd.n11175 vdd.n11174 0.0130799
R47197 vdd.n11161 vdd.n11160 0.0130799
R47198 vdd.n10192 vdd.n10191 0.0130799
R47199 vdd.n10191 vdd.n10190 0.0130799
R47200 vdd.n10173 vdd.n10170 0.0130799
R47201 vdd.n10173 vdd.n10167 0.0130799
R47202 vdd.n10197 vdd.n10196 0.0130799
R47203 vdd.n10197 vdd.n10162 0.0130799
R47204 vdd.n10204 vdd.n10159 0.0130799
R47205 vdd.n10172 vdd.n10171 0.0130799
R47206 vdd.n11248 vdd.n11241 0.0130799
R47207 vdd.n11248 vdd.n11246 0.0130799
R47208 vdd.n11261 vdd.n11254 0.0130799
R47209 vdd.n11254 vdd.n11253 0.0130799
R47210 vdd.n11272 vdd.n11271 0.0130799
R47211 vdd.n11271 vdd.n11247 0.0130799
R47212 vdd.n11274 vdd.n11273 0.0130799
R47213 vdd.n11260 vdd.n11259 0.0130799
R47214 vdd.n11200 vdd.n11193 0.0130799
R47215 vdd.n11200 vdd.n11198 0.0130799
R47216 vdd.n11213 vdd.n11206 0.0130799
R47217 vdd.n11206 vdd.n11205 0.0130799
R47218 vdd.n11224 vdd.n11223 0.0130799
R47219 vdd.n11223 vdd.n11199 0.0130799
R47220 vdd.n11226 vdd.n11225 0.0130799
R47221 vdd.n11212 vdd.n11211 0.0130799
R47222 vdd.n11297 vdd.n11290 0.0130799
R47223 vdd.n11297 vdd.n11295 0.0130799
R47224 vdd.n11310 vdd.n11303 0.0130799
R47225 vdd.n11303 vdd.n11302 0.0130799
R47226 vdd.n11321 vdd.n11320 0.0130799
R47227 vdd.n11320 vdd.n11296 0.0130799
R47228 vdd.n11323 vdd.n11322 0.0130799
R47229 vdd.n11309 vdd.n11308 0.0130799
R47230 vdd.n11347 vdd.n11340 0.0130799
R47231 vdd.n11347 vdd.n11345 0.0130799
R47232 vdd.n11360 vdd.n11353 0.0130799
R47233 vdd.n11353 vdd.n11352 0.0130799
R47234 vdd.n11371 vdd.n11370 0.0130799
R47235 vdd.n11370 vdd.n11346 0.0130799
R47236 vdd.n11373 vdd.n11372 0.0130799
R47237 vdd.n11359 vdd.n11358 0.0130799
R47238 vdd.n11395 vdd.n11388 0.0130799
R47239 vdd.n11395 vdd.n11393 0.0130799
R47240 vdd.n11408 vdd.n11401 0.0130799
R47241 vdd.n11401 vdd.n11400 0.0130799
R47242 vdd.n11419 vdd.n11418 0.0130799
R47243 vdd.n11418 vdd.n11394 0.0130799
R47244 vdd.n11421 vdd.n11420 0.0130799
R47245 vdd.n11407 vdd.n11406 0.0130799
R47246 vdd.n11446 vdd.n11439 0.0130799
R47247 vdd.n11446 vdd.n11444 0.0130799
R47248 vdd.n11470 vdd.n11469 0.0130799
R47249 vdd.n11469 vdd.n11445 0.0130799
R47250 vdd.n11454 vdd.n11452 0.0130799
R47251 vdd.n11452 vdd.n11451 0.0130799
R47252 vdd.n11457 vdd.n11453 0.0130799
R47253 vdd.n11472 vdd.n11471 0.0130799
R47254 vdd.n11493 vdd.n11486 0.0130799
R47255 vdd.n11493 vdd.n11491 0.0130799
R47256 vdd.n11517 vdd.n11516 0.0130799
R47257 vdd.n11516 vdd.n11492 0.0130799
R47258 vdd.n11501 vdd.n11499 0.0130799
R47259 vdd.n11499 vdd.n11498 0.0130799
R47260 vdd.n11504 vdd.n11500 0.0130799
R47261 vdd.n11519 vdd.n11518 0.0130799
R47262 vdd.n11543 vdd.n11536 0.0130799
R47263 vdd.n11543 vdd.n11541 0.0130799
R47264 vdd.n11567 vdd.n11566 0.0130799
R47265 vdd.n11566 vdd.n11542 0.0130799
R47266 vdd.n11551 vdd.n11549 0.0130799
R47267 vdd.n11549 vdd.n11548 0.0130799
R47268 vdd.n11554 vdd.n11550 0.0130799
R47269 vdd.n11569 vdd.n11568 0.0130799
R47270 vdd.n11593 vdd.n11586 0.0130799
R47271 vdd.n11593 vdd.n11591 0.0130799
R47272 vdd.n11617 vdd.n11616 0.0130799
R47273 vdd.n11616 vdd.n11592 0.0130799
R47274 vdd.n11601 vdd.n11599 0.0130799
R47275 vdd.n11599 vdd.n11598 0.0130799
R47276 vdd.n11604 vdd.n11600 0.0130799
R47277 vdd.n11619 vdd.n11618 0.0130799
R47278 vdd.n11641 vdd.n11634 0.0130799
R47279 vdd.n11641 vdd.n11639 0.0130799
R47280 vdd.n11665 vdd.n11664 0.0130799
R47281 vdd.n11664 vdd.n11640 0.0130799
R47282 vdd.n11649 vdd.n11647 0.0130799
R47283 vdd.n11647 vdd.n11646 0.0130799
R47284 vdd.n11652 vdd.n11648 0.0130799
R47285 vdd.n11667 vdd.n11666 0.0130799
R47286 vdd.n473 vdd.n472 0.0130799
R47287 vdd.n472 vdd.n450 0.0130799
R47288 vdd.n456 vdd.n455 0.0130799
R47289 vdd.n455 vdd.n453 0.0130799
R47290 vdd.n447 vdd.n446 0.0130799
R47291 vdd.n446 vdd.n444 0.0130799
R47292 vdd.n442 vdd.n440 0.0130799
R47293 vdd.n458 vdd.n457 0.0130799
R47294 vdd.n11692 vdd.n11685 0.0130799
R47295 vdd.n11692 vdd.n11690 0.0130799
R47296 vdd.n11716 vdd.n11715 0.0130799
R47297 vdd.n11715 vdd.n11691 0.0130799
R47298 vdd.n11700 vdd.n11698 0.0130799
R47299 vdd.n11698 vdd.n11697 0.0130799
R47300 vdd.n11703 vdd.n11699 0.0130799
R47301 vdd.n11718 vdd.n11717 0.0130799
R47302 vdd.n11739 vdd.n11732 0.0130799
R47303 vdd.n11739 vdd.n11737 0.0130799
R47304 vdd.n11763 vdd.n11762 0.0130799
R47305 vdd.n11762 vdd.n11738 0.0130799
R47306 vdd.n11747 vdd.n11745 0.0130799
R47307 vdd.n11745 vdd.n11744 0.0130799
R47308 vdd.n11750 vdd.n11746 0.0130799
R47309 vdd.n11765 vdd.n11764 0.0130799
R47310 vdd.n11787 vdd.n11780 0.0130799
R47311 vdd.n11787 vdd.n11785 0.0130799
R47312 vdd.n11811 vdd.n11810 0.0130799
R47313 vdd.n11810 vdd.n11786 0.0130799
R47314 vdd.n11795 vdd.n11793 0.0130799
R47315 vdd.n11793 vdd.n11792 0.0130799
R47316 vdd.n11798 vdd.n11794 0.0130799
R47317 vdd.n11813 vdd.n11812 0.0130799
R47318 vdd.n11838 vdd.n11831 0.0130799
R47319 vdd.n11838 vdd.n11836 0.0130799
R47320 vdd.n11862 vdd.n11861 0.0130799
R47321 vdd.n11861 vdd.n11837 0.0130799
R47322 vdd.n11846 vdd.n11844 0.0130799
R47323 vdd.n11844 vdd.n11843 0.0130799
R47324 vdd.n11849 vdd.n11845 0.0130799
R47325 vdd.n11864 vdd.n11863 0.0130799
R47326 vdd.n11888 vdd.n11881 0.0130799
R47327 vdd.n11888 vdd.n11886 0.0130799
R47328 vdd.n11912 vdd.n11911 0.0130799
R47329 vdd.n11911 vdd.n11887 0.0130799
R47330 vdd.n11896 vdd.n11894 0.0130799
R47331 vdd.n11894 vdd.n11893 0.0130799
R47332 vdd.n11899 vdd.n11895 0.0130799
R47333 vdd.n11914 vdd.n11913 0.0130799
R47334 vdd.n11936 vdd.n11929 0.0130799
R47335 vdd.n11936 vdd.n11934 0.0130799
R47336 vdd.n11960 vdd.n11959 0.0130799
R47337 vdd.n11959 vdd.n11935 0.0130799
R47338 vdd.n11944 vdd.n11942 0.0130799
R47339 vdd.n11942 vdd.n11941 0.0130799
R47340 vdd.n11947 vdd.n11943 0.0130799
R47341 vdd.n11962 vdd.n11961 0.0130799
R47342 vdd.n11986 vdd.n11979 0.0130799
R47343 vdd.n11986 vdd.n11984 0.0130799
R47344 vdd.n12010 vdd.n12009 0.0130799
R47345 vdd.n12009 vdd.n11985 0.0130799
R47346 vdd.n11994 vdd.n11992 0.0130799
R47347 vdd.n11992 vdd.n11991 0.0130799
R47348 vdd.n11997 vdd.n11993 0.0130799
R47349 vdd.n12012 vdd.n12011 0.0130799
R47350 vdd.n12033 vdd.n12026 0.0130799
R47351 vdd.n12033 vdd.n12031 0.0130799
R47352 vdd.n12057 vdd.n12056 0.0130799
R47353 vdd.n12056 vdd.n12032 0.0130799
R47354 vdd.n12041 vdd.n12039 0.0130799
R47355 vdd.n12039 vdd.n12038 0.0130799
R47356 vdd.n12044 vdd.n12040 0.0130799
R47357 vdd.n12059 vdd.n12058 0.0130799
R47358 vdd.n12083 vdd.n12076 0.0130799
R47359 vdd.n12083 vdd.n12081 0.0130799
R47360 vdd.n12107 vdd.n12106 0.0130799
R47361 vdd.n12106 vdd.n12082 0.0130799
R47362 vdd.n12091 vdd.n12089 0.0130799
R47363 vdd.n12089 vdd.n12088 0.0130799
R47364 vdd.n12094 vdd.n12090 0.0130799
R47365 vdd.n12109 vdd.n12108 0.0130799
R47366 vdd.n12133 vdd.n12126 0.0130799
R47367 vdd.n12133 vdd.n12131 0.0130799
R47368 vdd.n12157 vdd.n12156 0.0130799
R47369 vdd.n12156 vdd.n12132 0.0130799
R47370 vdd.n12141 vdd.n12139 0.0130799
R47371 vdd.n12139 vdd.n12138 0.0130799
R47372 vdd.n12144 vdd.n12140 0.0130799
R47373 vdd.n12159 vdd.n12158 0.0130799
R47374 vdd.n12181 vdd.n12174 0.0130799
R47375 vdd.n12181 vdd.n12179 0.0130799
R47376 vdd.n12205 vdd.n12204 0.0130799
R47377 vdd.n12204 vdd.n12180 0.0130799
R47378 vdd.n12189 vdd.n12187 0.0130799
R47379 vdd.n12187 vdd.n12186 0.0130799
R47380 vdd.n12192 vdd.n12188 0.0130799
R47381 vdd.n12207 vdd.n12206 0.0130799
R47382 vdd.n228 vdd.n227 0.0130799
R47383 vdd.n227 vdd.n205 0.0130799
R47384 vdd.n211 vdd.n210 0.0130799
R47385 vdd.n210 vdd.n208 0.0130799
R47386 vdd.n202 vdd.n201 0.0130799
R47387 vdd.n201 vdd.n199 0.0130799
R47388 vdd.n197 vdd.n195 0.0130799
R47389 vdd.n213 vdd.n212 0.0130799
R47390 vdd.n12232 vdd.n12225 0.0130799
R47391 vdd.n12232 vdd.n12230 0.0130799
R47392 vdd.n12256 vdd.n12255 0.0130799
R47393 vdd.n12255 vdd.n12231 0.0130799
R47394 vdd.n12240 vdd.n12238 0.0130799
R47395 vdd.n12238 vdd.n12237 0.0130799
R47396 vdd.n12243 vdd.n12239 0.0130799
R47397 vdd.n12258 vdd.n12257 0.0130799
R47398 vdd.n12279 vdd.n12272 0.0130799
R47399 vdd.n12279 vdd.n12277 0.0130799
R47400 vdd.n12303 vdd.n12302 0.0130799
R47401 vdd.n12302 vdd.n12278 0.0130799
R47402 vdd.n12287 vdd.n12285 0.0130799
R47403 vdd.n12285 vdd.n12284 0.0130799
R47404 vdd.n12290 vdd.n12286 0.0130799
R47405 vdd.n12305 vdd.n12304 0.0130799
R47406 vdd.n12329 vdd.n12322 0.0130799
R47407 vdd.n12329 vdd.n12327 0.0130799
R47408 vdd.n12353 vdd.n12352 0.0130799
R47409 vdd.n12352 vdd.n12328 0.0130799
R47410 vdd.n12337 vdd.n12335 0.0130799
R47411 vdd.n12335 vdd.n12334 0.0130799
R47412 vdd.n12340 vdd.n12336 0.0130799
R47413 vdd.n12355 vdd.n12354 0.0130799
R47414 vdd.n12379 vdd.n12372 0.0130799
R47415 vdd.n12379 vdd.n12377 0.0130799
R47416 vdd.n12403 vdd.n12402 0.0130799
R47417 vdd.n12402 vdd.n12378 0.0130799
R47418 vdd.n12387 vdd.n12385 0.0130799
R47419 vdd.n12385 vdd.n12384 0.0130799
R47420 vdd.n12390 vdd.n12386 0.0130799
R47421 vdd.n12405 vdd.n12404 0.0130799
R47422 vdd.n12427 vdd.n12420 0.0130799
R47423 vdd.n12427 vdd.n12425 0.0130799
R47424 vdd.n12451 vdd.n12450 0.0130799
R47425 vdd.n12450 vdd.n12426 0.0130799
R47426 vdd.n12435 vdd.n12433 0.0130799
R47427 vdd.n12433 vdd.n12432 0.0130799
R47428 vdd.n12438 vdd.n12434 0.0130799
R47429 vdd.n12453 vdd.n12452 0.0130799
R47430 vdd vdd 0.0120132
R47431 vdd vdd 0.0120132
R47432 vdd vdd 0.0120132
R47433 vdd vdd 0.0120132
R47434 vdd vdd 0.0120132
R47435 vdd vdd 0.0120132
R47436 vdd vdd 0.0120132
R47437 vdd vdd 0.0120132
R47438 vdd vdd 0.00872368
R47439 vdd vdd 0.00872368
R47440 vdd.n119 vdd.n118 0.00463816
R47441 vdd.n167 vdd.n166 0.00463816
R47442 vdd.n268 vdd.n267 0.00463816
R47443 vdd.n316 vdd.n315 0.00463816
R47444 vdd.n364 vdd.n363 0.00463816
R47445 vdd.n412 vdd.n411 0.00463816
R47446 vdd.n513 vdd.n512 0.00463816
R47447 vdd.n561 vdd.n560 0.00463816
R47448 vdd.n7433 vdd.n7432 0.00463816
R47449 vdd.n7481 vdd.n7480 0.00463816
R47450 vdd.n7582 vdd.n7581 0.00463816
R47451 vdd.n7630 vdd.n7629 0.00463816
R47452 vdd.n7678 vdd.n7677 0.00463816
R47453 vdd.n7726 vdd.n7725 0.00463816
R47454 vdd.n7827 vdd.n7826 0.00463816
R47455 vdd.n6940 vdd.n6939 0.00463816
R47456 vdd.n7875 vdd.n7874 0.00463816
R47457 vdd.n7922 vdd.n7921 0.00463816
R47458 vdd.n7972 vdd.n7971 0.00463816
R47459 vdd.n8022 vdd.n8021 0.00463816
R47460 vdd.n8070 vdd.n8069 0.00463816
R47461 vdd.n7798 vdd.n7797 0.00463816
R47462 vdd.n8121 vdd.n8120 0.00463816
R47463 vdd.n8168 vdd.n8167 0.00463816
R47464 vdd.n8216 vdd.n8215 0.00463816
R47465 vdd.n8267 vdd.n8266 0.00463816
R47466 vdd.n8317 vdd.n8316 0.00463816
R47467 vdd.n8365 vdd.n8364 0.00463816
R47468 vdd.n8415 vdd.n8414 0.00463816
R47469 vdd.n8462 vdd.n8461 0.00463816
R47470 vdd.n8512 vdd.n8511 0.00463816
R47471 vdd.n8562 vdd.n8561 0.00463816
R47472 vdd.n8610 vdd.n8609 0.00463816
R47473 vdd.n7553 vdd.n7552 0.00463816
R47474 vdd.n8661 vdd.n8660 0.00463816
R47475 vdd.n8708 vdd.n8707 0.00463816
R47476 vdd.n8758 vdd.n8757 0.00463816
R47477 vdd.n8808 vdd.n8807 0.00463816
R47478 vdd.n8856 vdd.n8855 0.00463816
R47479 vdd.n4291 vdd.n4290 0.00463816
R47480 vdd.n4339 vdd.n4338 0.00463816
R47481 vdd.n4440 vdd.n4439 0.00463816
R47482 vdd.n4488 vdd.n4487 0.00463816
R47483 vdd.n4536 vdd.n4535 0.00463816
R47484 vdd.n4584 vdd.n4583 0.00463816
R47485 vdd.n4685 vdd.n4684 0.00463816
R47486 vdd.n3798 vdd.n3797 0.00463816
R47487 vdd.n4733 vdd.n4732 0.00463816
R47488 vdd.n4780 vdd.n4779 0.00463816
R47489 vdd.n4830 vdd.n4829 0.00463816
R47490 vdd.n4880 vdd.n4879 0.00463816
R47491 vdd.n4928 vdd.n4927 0.00463816
R47492 vdd.n4656 vdd.n4655 0.00463816
R47493 vdd.n4979 vdd.n4978 0.00463816
R47494 vdd.n5026 vdd.n5025 0.00463816
R47495 vdd.n5074 vdd.n5073 0.00463816
R47496 vdd.n5125 vdd.n5124 0.00463816
R47497 vdd.n5175 vdd.n5174 0.00463816
R47498 vdd.n5223 vdd.n5222 0.00463816
R47499 vdd.n5273 vdd.n5272 0.00463816
R47500 vdd.n5320 vdd.n5319 0.00463816
R47501 vdd.n5370 vdd.n5369 0.00463816
R47502 vdd.n5420 vdd.n5419 0.00463816
R47503 vdd.n5468 vdd.n5467 0.00463816
R47504 vdd.n4411 vdd.n4410 0.00463816
R47505 vdd.n5519 vdd.n5518 0.00463816
R47506 vdd.n5566 vdd.n5565 0.00463816
R47507 vdd.n5616 vdd.n5615 0.00463816
R47508 vdd.n5666 vdd.n5665 0.00463816
R47509 vdd.n5714 vdd.n5713 0.00463816
R47510 vdd.n1149 vdd.n1148 0.00463816
R47511 vdd.n1197 vdd.n1196 0.00463816
R47512 vdd.n1298 vdd.n1297 0.00463816
R47513 vdd.n1346 vdd.n1345 0.00463816
R47514 vdd.n1394 vdd.n1393 0.00463816
R47515 vdd.n1442 vdd.n1441 0.00463816
R47516 vdd.n1543 vdd.n1542 0.00463816
R47517 vdd.n656 vdd.n655 0.00463816
R47518 vdd.n1591 vdd.n1590 0.00463816
R47519 vdd.n1638 vdd.n1637 0.00463816
R47520 vdd.n1688 vdd.n1687 0.00463816
R47521 vdd.n1738 vdd.n1737 0.00463816
R47522 vdd.n1786 vdd.n1785 0.00463816
R47523 vdd.n1514 vdd.n1513 0.00463816
R47524 vdd.n1837 vdd.n1836 0.00463816
R47525 vdd.n1884 vdd.n1883 0.00463816
R47526 vdd.n1932 vdd.n1931 0.00463816
R47527 vdd.n1983 vdd.n1982 0.00463816
R47528 vdd.n2033 vdd.n2032 0.00463816
R47529 vdd.n2081 vdd.n2080 0.00463816
R47530 vdd.n2131 vdd.n2130 0.00463816
R47531 vdd.n2178 vdd.n2177 0.00463816
R47532 vdd.n2228 vdd.n2227 0.00463816
R47533 vdd.n2278 vdd.n2277 0.00463816
R47534 vdd.n2326 vdd.n2325 0.00463816
R47535 vdd.n1269 vdd.n1268 0.00463816
R47536 vdd.n2377 vdd.n2376 0.00463816
R47537 vdd.n2424 vdd.n2423 0.00463816
R47538 vdd.n2474 vdd.n2473 0.00463816
R47539 vdd.n2524 vdd.n2523 0.00463816
R47540 vdd.n2572 vdd.n2571 0.00463816
R47541 vdd.n11461 vdd.n11460 0.00463816
R47542 vdd.n11508 vdd.n11507 0.00463816
R47543 vdd.n11558 vdd.n11557 0.00463816
R47544 vdd.n11608 vdd.n11607 0.00463816
R47545 vdd.n11656 vdd.n11655 0.00463816
R47546 vdd.n484 vdd.n483 0.00463816
R47547 vdd.n11707 vdd.n11706 0.00463816
R47548 vdd.n11754 vdd.n11753 0.00463816
R47549 vdd.n11802 vdd.n11801 0.00463816
R47550 vdd.n11853 vdd.n11852 0.00463816
R47551 vdd.n11903 vdd.n11902 0.00463816
R47552 vdd.n11951 vdd.n11950 0.00463816
R47553 vdd.n12001 vdd.n12000 0.00463816
R47554 vdd.n12048 vdd.n12047 0.00463816
R47555 vdd.n12098 vdd.n12097 0.00463816
R47556 vdd.n12148 vdd.n12147 0.00463816
R47557 vdd.n12196 vdd.n12195 0.00463816
R47558 vdd.n239 vdd.n238 0.00463816
R47559 vdd.n12247 vdd.n12246 0.00463816
R47560 vdd.n12294 vdd.n12293 0.00463816
R47561 vdd.n12344 vdd.n12343 0.00463816
R47562 vdd.n12394 vdd.n12393 0.00463816
R47563 vdd.n12442 vdd.n12441 0.00463816
R47564 vdd.n12504 vdd.n12503 0.00442942
R47565 vdd.n12481 vdd.n12480 0.00442942
R47566 vdd.n134 vdd.n133 0.00442942
R47567 vdd.n182 vdd.n181 0.00442942
R47568 vdd.n283 vdd.n282 0.00442942
R47569 vdd.n331 vdd.n330 0.00442942
R47570 vdd.n379 vdd.n378 0.00442942
R47571 vdd.n427 vdd.n426 0.00442942
R47572 vdd.n528 vdd.n527 0.00442942
R47573 vdd.n576 vdd.n575 0.00442942
R47574 vdd.n7004 vdd.n7003 0.00442942
R47575 vdd.n6983 vdd.n6981 0.00442942
R47576 vdd.n7052 vdd.n7051 0.00442942
R47577 vdd.n7031 vdd.n7029 0.00442942
R47578 vdd.n7154 vdd.n7153 0.00442942
R47579 vdd.n7133 vdd.n7131 0.00442942
R47580 vdd.n7202 vdd.n7201 0.00442942
R47581 vdd.n7181 vdd.n7179 0.00442942
R47582 vdd.n7250 vdd.n7249 0.00442942
R47583 vdd.n7229 vdd.n7227 0.00442942
R47584 vdd.n7298 vdd.n7297 0.00442942
R47585 vdd.n7277 vdd.n7275 0.00442942
R47586 vdd.n7400 vdd.n7399 0.00442942
R47587 vdd.n7379 vdd.n7377 0.00442942
R47588 vdd.n8920 vdd.n8919 0.00442942
R47589 vdd.n8899 vdd.n8897 0.00442942
R47590 vdd.n7448 vdd.n7447 0.00442942
R47591 vdd.n7496 vdd.n7495 0.00442942
R47592 vdd.n7597 vdd.n7596 0.00442942
R47593 vdd.n7645 vdd.n7644 0.00442942
R47594 vdd.n7693 vdd.n7692 0.00442942
R47595 vdd.n7741 vdd.n7740 0.00442942
R47596 vdd.n7842 vdd.n7841 0.00442942
R47597 vdd.n6955 vdd.n6954 0.00442942
R47598 vdd.n7890 vdd.n7889 0.00442942
R47599 vdd.n7937 vdd.n7936 0.00442942
R47600 vdd.n7987 vdd.n7986 0.00442942
R47601 vdd.n8037 vdd.n8036 0.00442942
R47602 vdd.n8085 vdd.n8084 0.00442942
R47603 vdd.n7777 vdd.n7776 0.00442942
R47604 vdd.n8136 vdd.n8135 0.00442942
R47605 vdd.n8183 vdd.n8182 0.00442942
R47606 vdd.n8231 vdd.n8230 0.00442942
R47607 vdd.n8282 vdd.n8281 0.00442942
R47608 vdd.n8332 vdd.n8331 0.00442942
R47609 vdd.n8380 vdd.n8379 0.00442942
R47610 vdd.n8430 vdd.n8429 0.00442942
R47611 vdd.n8477 vdd.n8476 0.00442942
R47612 vdd.n8527 vdd.n8526 0.00442942
R47613 vdd.n8577 vdd.n8576 0.00442942
R47614 vdd.n8625 vdd.n8624 0.00442942
R47615 vdd.n7532 vdd.n7531 0.00442942
R47616 vdd.n8676 vdd.n8675 0.00442942
R47617 vdd.n8723 vdd.n8722 0.00442942
R47618 vdd.n8773 vdd.n8772 0.00442942
R47619 vdd.n8823 vdd.n8822 0.00442942
R47620 vdd.n8871 vdd.n8870 0.00442942
R47621 vdd.n9017 vdd.n9016 0.00442942
R47622 vdd.n8996 vdd.n8994 0.00442942
R47623 vdd.n8969 vdd.n8968 0.00442942
R47624 vdd.n8948 vdd.n8946 0.00442942
R47625 vdd.n9066 vdd.n9065 0.00442942
R47626 vdd.n9045 vdd.n9043 0.00442942
R47627 vdd.n9116 vdd.n9115 0.00442942
R47628 vdd.n9095 vdd.n9093 0.00442942
R47629 vdd.n9164 vdd.n9163 0.00442942
R47630 vdd.n9143 vdd.n9141 0.00442942
R47631 vdd.n7354 vdd.n7353 0.00442942
R47632 vdd.n7333 vdd.n7332 0.00442942
R47633 vdd.n9312 vdd.n9311 0.00442942
R47634 vdd.n9291 vdd.n9289 0.00442942
R47635 vdd.n9263 vdd.n9262 0.00442942
R47636 vdd.n9242 vdd.n9240 0.00442942
R47637 vdd.n9215 vdd.n9214 0.00442942
R47638 vdd.n9194 vdd.n9192 0.00442942
R47639 vdd.n9361 vdd.n9360 0.00442942
R47640 vdd.n9340 vdd.n9338 0.00442942
R47641 vdd.n9411 vdd.n9410 0.00442942
R47642 vdd.n9390 vdd.n9388 0.00442942
R47643 vdd.n9459 vdd.n9458 0.00442942
R47644 vdd.n9438 vdd.n9436 0.00442942
R47645 vdd.n9557 vdd.n9556 0.00442942
R47646 vdd.n9536 vdd.n9534 0.00442942
R47647 vdd.n9509 vdd.n9508 0.00442942
R47648 vdd.n9488 vdd.n9486 0.00442942
R47649 vdd.n9606 vdd.n9605 0.00442942
R47650 vdd.n9585 vdd.n9583 0.00442942
R47651 vdd.n9656 vdd.n9655 0.00442942
R47652 vdd.n9635 vdd.n9633 0.00442942
R47653 vdd.n9704 vdd.n9703 0.00442942
R47654 vdd.n9683 vdd.n9681 0.00442942
R47655 vdd.n7108 vdd.n7107 0.00442942
R47656 vdd.n7087 vdd.n7086 0.00442942
R47657 vdd.n9803 vdd.n9802 0.00442942
R47658 vdd.n9782 vdd.n9780 0.00442942
R47659 vdd.n9755 vdd.n9754 0.00442942
R47660 vdd.n9734 vdd.n9732 0.00442942
R47661 vdd.n9852 vdd.n9851 0.00442942
R47662 vdd.n9831 vdd.n9829 0.00442942
R47663 vdd.n9902 vdd.n9901 0.00442942
R47664 vdd.n9881 vdd.n9879 0.00442942
R47665 vdd.n9950 vdd.n9949 0.00442942
R47666 vdd.n9929 vdd.n9927 0.00442942
R47667 vdd.n3862 vdd.n3861 0.00442942
R47668 vdd.n3841 vdd.n3839 0.00442942
R47669 vdd.n3910 vdd.n3909 0.00442942
R47670 vdd.n3889 vdd.n3887 0.00442942
R47671 vdd.n4012 vdd.n4011 0.00442942
R47672 vdd.n3991 vdd.n3989 0.00442942
R47673 vdd.n4060 vdd.n4059 0.00442942
R47674 vdd.n4039 vdd.n4037 0.00442942
R47675 vdd.n4108 vdd.n4107 0.00442942
R47676 vdd.n4087 vdd.n4085 0.00442942
R47677 vdd.n4156 vdd.n4155 0.00442942
R47678 vdd.n4135 vdd.n4133 0.00442942
R47679 vdd.n4258 vdd.n4257 0.00442942
R47680 vdd.n4237 vdd.n4235 0.00442942
R47681 vdd.n5778 vdd.n5777 0.00442942
R47682 vdd.n5757 vdd.n5755 0.00442942
R47683 vdd.n4306 vdd.n4305 0.00442942
R47684 vdd.n4354 vdd.n4353 0.00442942
R47685 vdd.n4455 vdd.n4454 0.00442942
R47686 vdd.n4503 vdd.n4502 0.00442942
R47687 vdd.n4551 vdd.n4550 0.00442942
R47688 vdd.n4599 vdd.n4598 0.00442942
R47689 vdd.n4700 vdd.n4699 0.00442942
R47690 vdd.n3813 vdd.n3812 0.00442942
R47691 vdd.n4748 vdd.n4747 0.00442942
R47692 vdd.n4795 vdd.n4794 0.00442942
R47693 vdd.n4845 vdd.n4844 0.00442942
R47694 vdd.n4895 vdd.n4894 0.00442942
R47695 vdd.n4943 vdd.n4942 0.00442942
R47696 vdd.n4635 vdd.n4634 0.00442942
R47697 vdd.n4994 vdd.n4993 0.00442942
R47698 vdd.n5041 vdd.n5040 0.00442942
R47699 vdd.n5089 vdd.n5088 0.00442942
R47700 vdd.n5140 vdd.n5139 0.00442942
R47701 vdd.n5190 vdd.n5189 0.00442942
R47702 vdd.n5238 vdd.n5237 0.00442942
R47703 vdd.n5288 vdd.n5287 0.00442942
R47704 vdd.n5335 vdd.n5334 0.00442942
R47705 vdd.n5385 vdd.n5384 0.00442942
R47706 vdd.n5435 vdd.n5434 0.00442942
R47707 vdd.n5483 vdd.n5482 0.00442942
R47708 vdd.n4390 vdd.n4389 0.00442942
R47709 vdd.n5534 vdd.n5533 0.00442942
R47710 vdd.n5581 vdd.n5580 0.00442942
R47711 vdd.n5631 vdd.n5630 0.00442942
R47712 vdd.n5681 vdd.n5680 0.00442942
R47713 vdd.n5729 vdd.n5728 0.00442942
R47714 vdd.n5875 vdd.n5874 0.00442942
R47715 vdd.n5854 vdd.n5852 0.00442942
R47716 vdd.n5827 vdd.n5826 0.00442942
R47717 vdd.n5806 vdd.n5804 0.00442942
R47718 vdd.n5924 vdd.n5923 0.00442942
R47719 vdd.n5903 vdd.n5901 0.00442942
R47720 vdd.n5974 vdd.n5973 0.00442942
R47721 vdd.n5953 vdd.n5951 0.00442942
R47722 vdd.n6022 vdd.n6021 0.00442942
R47723 vdd.n6001 vdd.n5999 0.00442942
R47724 vdd.n4212 vdd.n4211 0.00442942
R47725 vdd.n4191 vdd.n4190 0.00442942
R47726 vdd.n6170 vdd.n6169 0.00442942
R47727 vdd.n6149 vdd.n6147 0.00442942
R47728 vdd.n6121 vdd.n6120 0.00442942
R47729 vdd.n6100 vdd.n6098 0.00442942
R47730 vdd.n6073 vdd.n6072 0.00442942
R47731 vdd.n6052 vdd.n6050 0.00442942
R47732 vdd.n6219 vdd.n6218 0.00442942
R47733 vdd.n6198 vdd.n6196 0.00442942
R47734 vdd.n6269 vdd.n6268 0.00442942
R47735 vdd.n6248 vdd.n6246 0.00442942
R47736 vdd.n6317 vdd.n6316 0.00442942
R47737 vdd.n6296 vdd.n6294 0.00442942
R47738 vdd.n6415 vdd.n6414 0.00442942
R47739 vdd.n6394 vdd.n6392 0.00442942
R47740 vdd.n6367 vdd.n6366 0.00442942
R47741 vdd.n6346 vdd.n6344 0.00442942
R47742 vdd.n6464 vdd.n6463 0.00442942
R47743 vdd.n6443 vdd.n6441 0.00442942
R47744 vdd.n6514 vdd.n6513 0.00442942
R47745 vdd.n6493 vdd.n6491 0.00442942
R47746 vdd.n6562 vdd.n6561 0.00442942
R47747 vdd.n6541 vdd.n6539 0.00442942
R47748 vdd.n3966 vdd.n3965 0.00442942
R47749 vdd.n3945 vdd.n3944 0.00442942
R47750 vdd.n6661 vdd.n6660 0.00442942
R47751 vdd.n6640 vdd.n6638 0.00442942
R47752 vdd.n6613 vdd.n6612 0.00442942
R47753 vdd.n6592 vdd.n6590 0.00442942
R47754 vdd.n6710 vdd.n6709 0.00442942
R47755 vdd.n6689 vdd.n6687 0.00442942
R47756 vdd.n6760 vdd.n6759 0.00442942
R47757 vdd.n6739 vdd.n6737 0.00442942
R47758 vdd.n6808 vdd.n6807 0.00442942
R47759 vdd.n6787 vdd.n6785 0.00442942
R47760 vdd.n720 vdd.n719 0.00442942
R47761 vdd.n699 vdd.n697 0.00442942
R47762 vdd.n768 vdd.n767 0.00442942
R47763 vdd.n747 vdd.n745 0.00442942
R47764 vdd.n870 vdd.n869 0.00442942
R47765 vdd.n849 vdd.n847 0.00442942
R47766 vdd.n918 vdd.n917 0.00442942
R47767 vdd.n897 vdd.n895 0.00442942
R47768 vdd.n966 vdd.n965 0.00442942
R47769 vdd.n945 vdd.n943 0.00442942
R47770 vdd.n1014 vdd.n1013 0.00442942
R47771 vdd.n993 vdd.n991 0.00442942
R47772 vdd.n1116 vdd.n1115 0.00442942
R47773 vdd.n1095 vdd.n1093 0.00442942
R47774 vdd.n2636 vdd.n2635 0.00442942
R47775 vdd.n2615 vdd.n2613 0.00442942
R47776 vdd.n1164 vdd.n1163 0.00442942
R47777 vdd.n1212 vdd.n1211 0.00442942
R47778 vdd.n1313 vdd.n1312 0.00442942
R47779 vdd.n1361 vdd.n1360 0.00442942
R47780 vdd.n1409 vdd.n1408 0.00442942
R47781 vdd.n1457 vdd.n1456 0.00442942
R47782 vdd.n1558 vdd.n1557 0.00442942
R47783 vdd.n671 vdd.n670 0.00442942
R47784 vdd.n1606 vdd.n1605 0.00442942
R47785 vdd.n1653 vdd.n1652 0.00442942
R47786 vdd.n1703 vdd.n1702 0.00442942
R47787 vdd.n1753 vdd.n1752 0.00442942
R47788 vdd.n1801 vdd.n1800 0.00442942
R47789 vdd.n1493 vdd.n1492 0.00442942
R47790 vdd.n1852 vdd.n1851 0.00442942
R47791 vdd.n1899 vdd.n1898 0.00442942
R47792 vdd.n1947 vdd.n1946 0.00442942
R47793 vdd.n1998 vdd.n1997 0.00442942
R47794 vdd.n2048 vdd.n2047 0.00442942
R47795 vdd.n2096 vdd.n2095 0.00442942
R47796 vdd.n2146 vdd.n2145 0.00442942
R47797 vdd.n2193 vdd.n2192 0.00442942
R47798 vdd.n2243 vdd.n2242 0.00442942
R47799 vdd.n2293 vdd.n2292 0.00442942
R47800 vdd.n2341 vdd.n2340 0.00442942
R47801 vdd.n1248 vdd.n1247 0.00442942
R47802 vdd.n2392 vdd.n2391 0.00442942
R47803 vdd.n2439 vdd.n2438 0.00442942
R47804 vdd.n2489 vdd.n2488 0.00442942
R47805 vdd.n2539 vdd.n2538 0.00442942
R47806 vdd.n2587 vdd.n2586 0.00442942
R47807 vdd.n2733 vdd.n2732 0.00442942
R47808 vdd.n2712 vdd.n2710 0.00442942
R47809 vdd.n2685 vdd.n2684 0.00442942
R47810 vdd.n2664 vdd.n2662 0.00442942
R47811 vdd.n2782 vdd.n2781 0.00442942
R47812 vdd.n2761 vdd.n2759 0.00442942
R47813 vdd.n2832 vdd.n2831 0.00442942
R47814 vdd.n2811 vdd.n2809 0.00442942
R47815 vdd.n2880 vdd.n2879 0.00442942
R47816 vdd.n2859 vdd.n2857 0.00442942
R47817 vdd.n1070 vdd.n1069 0.00442942
R47818 vdd.n1049 vdd.n1048 0.00442942
R47819 vdd.n3028 vdd.n3027 0.00442942
R47820 vdd.n3007 vdd.n3005 0.00442942
R47821 vdd.n2979 vdd.n2978 0.00442942
R47822 vdd.n2958 vdd.n2956 0.00442942
R47823 vdd.n2931 vdd.n2930 0.00442942
R47824 vdd.n2910 vdd.n2908 0.00442942
R47825 vdd.n3077 vdd.n3076 0.00442942
R47826 vdd.n3056 vdd.n3054 0.00442942
R47827 vdd.n3127 vdd.n3126 0.00442942
R47828 vdd.n3106 vdd.n3104 0.00442942
R47829 vdd.n3175 vdd.n3174 0.00442942
R47830 vdd.n3154 vdd.n3152 0.00442942
R47831 vdd.n3273 vdd.n3272 0.00442942
R47832 vdd.n3252 vdd.n3250 0.00442942
R47833 vdd.n3225 vdd.n3224 0.00442942
R47834 vdd.n3204 vdd.n3202 0.00442942
R47835 vdd.n3322 vdd.n3321 0.00442942
R47836 vdd.n3301 vdd.n3299 0.00442942
R47837 vdd.n3372 vdd.n3371 0.00442942
R47838 vdd.n3351 vdd.n3349 0.00442942
R47839 vdd.n3420 vdd.n3419 0.00442942
R47840 vdd.n3399 vdd.n3397 0.00442942
R47841 vdd.n824 vdd.n823 0.00442942
R47842 vdd.n803 vdd.n802 0.00442942
R47843 vdd.n3519 vdd.n3518 0.00442942
R47844 vdd.n3498 vdd.n3496 0.00442942
R47845 vdd.n3471 vdd.n3470 0.00442942
R47846 vdd.n3450 vdd.n3448 0.00442942
R47847 vdd.n3568 vdd.n3567 0.00442942
R47848 vdd.n3547 vdd.n3545 0.00442942
R47849 vdd.n3618 vdd.n3617 0.00442942
R47850 vdd.n3597 vdd.n3595 0.00442942
R47851 vdd.n3666 vdd.n3665 0.00442942
R47852 vdd.n3645 vdd.n3643 0.00442942
R47853 vdd.n624 vdd.n623 0.00442942
R47854 vdd.n603 vdd.n601 0.00442942
R47855 vdd.n3765 vdd.n3764 0.00442942
R47856 vdd.n3744 vdd.n3742 0.00442942
R47857 vdd.n3717 vdd.n3716 0.00442942
R47858 vdd.n3696 vdd.n3694 0.00442942
R47859 vdd.n6907 vdd.n6906 0.00442942
R47860 vdd.n6886 vdd.n6884 0.00442942
R47861 vdd.n6859 vdd.n6858 0.00442942
R47862 vdd.n6838 vdd.n6836 0.00442942
R47863 vdd.n10049 vdd.n10048 0.00442942
R47864 vdd.n10028 vdd.n10026 0.00442942
R47865 vdd.n10001 vdd.n10000 0.00442942
R47866 vdd.n9980 vdd.n9978 0.00442942
R47867 vdd.n10097 vdd.n10096 0.00442942
R47868 vdd.n10076 vdd.n10074 0.00442942
R47869 vdd.n10145 vdd.n10144 0.00442942
R47870 vdd.n10124 vdd.n10122 0.00442942
R47871 vdd.n10247 vdd.n10246 0.00442942
R47872 vdd.n10226 vdd.n10224 0.00442942
R47873 vdd.n10295 vdd.n10294 0.00442942
R47874 vdd.n10274 vdd.n10272 0.00442942
R47875 vdd.n10343 vdd.n10342 0.00442942
R47876 vdd.n10322 vdd.n10320 0.00442942
R47877 vdd.n10391 vdd.n10390 0.00442942
R47878 vdd.n10370 vdd.n10368 0.00442942
R47879 vdd.n10493 vdd.n10492 0.00442942
R47880 vdd.n10472 vdd.n10470 0.00442942
R47881 vdd.n85 vdd.n84 0.00442942
R47882 vdd.n64 vdd.n62 0.00442942
R47883 vdd.n37 vdd.n36 0.00442942
R47884 vdd.n16 vdd.n14 0.00442942
R47885 vdd.n10541 vdd.n10540 0.00442942
R47886 vdd.n10520 vdd.n10518 0.00442942
R47887 vdd.n10591 vdd.n10590 0.00442942
R47888 vdd.n10570 vdd.n10568 0.00442942
R47889 vdd.n10639 vdd.n10638 0.00442942
R47890 vdd.n10618 vdd.n10616 0.00442942
R47891 vdd.n10447 vdd.n10446 0.00442942
R47892 vdd.n10426 vdd.n10425 0.00442942
R47893 vdd.n10787 vdd.n10786 0.00442942
R47894 vdd.n10766 vdd.n10764 0.00442942
R47895 vdd.n10738 vdd.n10737 0.00442942
R47896 vdd.n10717 vdd.n10715 0.00442942
R47897 vdd.n10690 vdd.n10689 0.00442942
R47898 vdd.n10669 vdd.n10667 0.00442942
R47899 vdd.n10836 vdd.n10835 0.00442942
R47900 vdd.n10815 vdd.n10813 0.00442942
R47901 vdd.n10886 vdd.n10885 0.00442942
R47902 vdd.n10865 vdd.n10863 0.00442942
R47903 vdd.n10934 vdd.n10933 0.00442942
R47904 vdd.n10913 vdd.n10911 0.00442942
R47905 vdd.n11032 vdd.n11031 0.00442942
R47906 vdd.n11011 vdd.n11009 0.00442942
R47907 vdd.n10984 vdd.n10983 0.00442942
R47908 vdd.n10963 vdd.n10961 0.00442942
R47909 vdd.n11081 vdd.n11080 0.00442942
R47910 vdd.n11060 vdd.n11058 0.00442942
R47911 vdd.n11131 vdd.n11130 0.00442942
R47912 vdd.n11110 vdd.n11108 0.00442942
R47913 vdd.n11179 vdd.n11178 0.00442942
R47914 vdd.n11158 vdd.n11156 0.00442942
R47915 vdd.n10201 vdd.n10200 0.00442942
R47916 vdd.n10180 vdd.n10179 0.00442942
R47917 vdd.n11278 vdd.n11277 0.00442942
R47918 vdd.n11257 vdd.n11255 0.00442942
R47919 vdd.n11230 vdd.n11229 0.00442942
R47920 vdd.n11209 vdd.n11207 0.00442942
R47921 vdd.n11327 vdd.n11326 0.00442942
R47922 vdd.n11306 vdd.n11304 0.00442942
R47923 vdd.n11377 vdd.n11376 0.00442942
R47924 vdd.n11356 vdd.n11354 0.00442942
R47925 vdd.n11425 vdd.n11424 0.00442942
R47926 vdd.n11404 vdd.n11402 0.00442942
R47927 vdd.n11476 vdd.n11475 0.00442942
R47928 vdd.n11523 vdd.n11522 0.00442942
R47929 vdd.n11573 vdd.n11572 0.00442942
R47930 vdd.n11623 vdd.n11622 0.00442942
R47931 vdd.n11671 vdd.n11670 0.00442942
R47932 vdd.n463 vdd.n462 0.00442942
R47933 vdd.n11722 vdd.n11721 0.00442942
R47934 vdd.n11769 vdd.n11768 0.00442942
R47935 vdd.n11817 vdd.n11816 0.00442942
R47936 vdd.n11868 vdd.n11867 0.00442942
R47937 vdd.n11918 vdd.n11917 0.00442942
R47938 vdd.n11966 vdd.n11965 0.00442942
R47939 vdd.n12016 vdd.n12015 0.00442942
R47940 vdd.n12063 vdd.n12062 0.00442942
R47941 vdd.n12113 vdd.n12112 0.00442942
R47942 vdd.n12163 vdd.n12162 0.00442942
R47943 vdd.n12211 vdd.n12210 0.00442942
R47944 vdd.n218 vdd.n217 0.00442942
R47945 vdd.n12262 vdd.n12261 0.00442942
R47946 vdd.n12309 vdd.n12308 0.00442942
R47947 vdd.n12359 vdd.n12358 0.00442942
R47948 vdd.n12409 vdd.n12408 0.00442942
R47949 vdd.n12457 vdd.n12456 0.00442942
R47950 vdd vdd 0.00214474
R47951 vdd.n7346 vdd.n7310 0.00100279
R47952 vdd.n7100 vdd.n7064 0.00100279
R47953 vdd.n4204 vdd.n4168 0.00100279
R47954 vdd.n3958 vdd.n3922 0.00100279
R47955 vdd.n1062 vdd.n1026 0.00100279
R47956 vdd.n816 vdd.n780 0.00100279
R47957 vdd.n10439 vdd.n10403 0.00100279
R47958 vdd.n10193 vdd.n10157 0.00100279
R47959 vdd.n7788 vdd.n7753 0.00100279
R47960 vdd.n7543 vdd.n7508 0.00100279
R47961 vdd.n4646 vdd.n4611 0.00100279
R47962 vdd.n4401 vdd.n4366 0.00100279
R47963 vdd.n1504 vdd.n1469 0.00100279
R47964 vdd.n1259 vdd.n1224 0.00100279
R47965 vdd.n474 vdd.n439 0.00100279
R47966 vdd.n229 vdd.n194 0.00100279
R47967 vdd.n7804 vdd.n7803 0.00100001
R47968 vdd.n7559 vdd.n7558 0.00100001
R47969 vdd.n7362 vdd.n7361 0.00100001
R47970 vdd.n7116 vdd.n7115 0.00100001
R47971 vdd.n4662 vdd.n4661 0.00100001
R47972 vdd.n4417 vdd.n4416 0.00100001
R47973 vdd.n4220 vdd.n4219 0.00100001
R47974 vdd.n3974 vdd.n3973 0.00100001
R47975 vdd.n1520 vdd.n1519 0.00100001
R47976 vdd.n1275 vdd.n1274 0.00100001
R47977 vdd.n1078 vdd.n1077 0.00100001
R47978 vdd.n832 vdd.n831 0.00100001
R47979 vdd.n10455 vdd.n10454 0.00100001
R47980 vdd.n10209 vdd.n10208 0.00100001
R47981 vdd.n490 vdd.n489 0.00100001
R47982 vdd.n245 vdd.n244 0.00100001
R47983 vdd.n6965 vdd.n6964 0.000501408
R47984 vdd.n7947 vdd.n7946 0.000501408
R47985 vdd.n7948 vdd.n7899 0.000501408
R47986 vdd.n7997 vdd.n7996 0.000501408
R47987 vdd.n7852 vdd.n7851 0.000501408
R47988 vdd.n8095 vdd.n8094 0.000501408
R47989 vdd.n7751 vdd.n7750 0.000501408
R47990 vdd.n8241 vdd.n8240 0.000501408
R47991 vdd.n8193 vdd.n8192 0.000501408
R47992 vdd.n8243 vdd.n8145 0.000501408
R47993 vdd.n8292 vdd.n8291 0.000501408
R47994 vdd.n7703 vdd.n7702 0.000501408
R47995 vdd.n8390 vdd.n8389 0.000501408
R47996 vdd.n7655 vdd.n7654 0.000501408
R47997 vdd.n8487 vdd.n8486 0.000501408
R47998 vdd.n8488 vdd.n8439 0.000501408
R47999 vdd.n8537 vdd.n8536 0.000501408
R48000 vdd.n7607 vdd.n7606 0.000501408
R48001 vdd.n8635 vdd.n8634 0.000501408
R48002 vdd.n7506 vdd.n7505 0.000501408
R48003 vdd.n8733 vdd.n8732 0.000501408
R48004 vdd.n8734 vdd.n8685 0.000501408
R48005 vdd.n8783 vdd.n8782 0.000501408
R48006 vdd.n7458 vdd.n7457 0.000501408
R48007 vdd.n8881 vdd.n8880 0.000501408
R48008 vdd.n8930 vdd.n8929 0.000501408
R48009 vdd.n8979 vdd.n8978 0.000501408
R48010 vdd.n9027 vdd.n9026 0.000501408
R48011 vdd.n9076 vdd.n9075 0.000501408
R48012 vdd.n7410 vdd.n7409 0.000501408
R48013 vdd.n9174 vdd.n9173 0.000501408
R48014 vdd.n7308 vdd.n7307 0.000501408
R48015 vdd.n9225 vdd.n9224 0.000501408
R48016 vdd.n9273 vdd.n9272 0.000501408
R48017 vdd.n9322 vdd.n9321 0.000501408
R48018 vdd.n9371 vdd.n9370 0.000501408
R48019 vdd.n7260 vdd.n7259 0.000501408
R48020 vdd.n9469 vdd.n9468 0.000501408
R48021 vdd.n7212 vdd.n7211 0.000501408
R48022 vdd.n9519 vdd.n9518 0.000501408
R48023 vdd.n9567 vdd.n9566 0.000501408
R48024 vdd.n9616 vdd.n9615 0.000501408
R48025 vdd.n7164 vdd.n7163 0.000501408
R48026 vdd.n9714 vdd.n9713 0.000501408
R48027 vdd.n7062 vdd.n7061 0.000501408
R48028 vdd.n9765 vdd.n9764 0.000501408
R48029 vdd.n9813 vdd.n9812 0.000501408
R48030 vdd.n9862 vdd.n9861 0.000501408
R48031 vdd.n7014 vdd.n7013 0.000501408
R48032 vdd.n9960 vdd.n9959 0.000501408
R48033 vdd.n3823 vdd.n3822 0.000501408
R48034 vdd.n4805 vdd.n4804 0.000501408
R48035 vdd.n4806 vdd.n4757 0.000501408
R48036 vdd.n4855 vdd.n4854 0.000501408
R48037 vdd.n4710 vdd.n4709 0.000501408
R48038 vdd.n4953 vdd.n4952 0.000501408
R48039 vdd.n4609 vdd.n4608 0.000501408
R48040 vdd.n5099 vdd.n5098 0.000501408
R48041 vdd.n5051 vdd.n5050 0.000501408
R48042 vdd.n5101 vdd.n5003 0.000501408
R48043 vdd.n5150 vdd.n5149 0.000501408
R48044 vdd.n4561 vdd.n4560 0.000501408
R48045 vdd.n5248 vdd.n5247 0.000501408
R48046 vdd.n4513 vdd.n4512 0.000501408
R48047 vdd.n5345 vdd.n5344 0.000501408
R48048 vdd.n5346 vdd.n5297 0.000501408
R48049 vdd.n5395 vdd.n5394 0.000501408
R48050 vdd.n4465 vdd.n4464 0.000501408
R48051 vdd.n5493 vdd.n5492 0.000501408
R48052 vdd.n4364 vdd.n4363 0.000501408
R48053 vdd.n5591 vdd.n5590 0.000501408
R48054 vdd.n5592 vdd.n5543 0.000501408
R48055 vdd.n5641 vdd.n5640 0.000501408
R48056 vdd.n4316 vdd.n4315 0.000501408
R48057 vdd.n5739 vdd.n5738 0.000501408
R48058 vdd.n5788 vdd.n5787 0.000501408
R48059 vdd.n5837 vdd.n5836 0.000501408
R48060 vdd.n5885 vdd.n5884 0.000501408
R48061 vdd.n5934 vdd.n5933 0.000501408
R48062 vdd.n4268 vdd.n4267 0.000501408
R48063 vdd.n6032 vdd.n6031 0.000501408
R48064 vdd.n4166 vdd.n4165 0.000501408
R48065 vdd.n6083 vdd.n6082 0.000501408
R48066 vdd.n6131 vdd.n6130 0.000501408
R48067 vdd.n6180 vdd.n6179 0.000501408
R48068 vdd.n6229 vdd.n6228 0.000501408
R48069 vdd.n4118 vdd.n4117 0.000501408
R48070 vdd.n6327 vdd.n6326 0.000501408
R48071 vdd.n4070 vdd.n4069 0.000501408
R48072 vdd.n6377 vdd.n6376 0.000501408
R48073 vdd.n6425 vdd.n6424 0.000501408
R48074 vdd.n6474 vdd.n6473 0.000501408
R48075 vdd.n4022 vdd.n4021 0.000501408
R48076 vdd.n6572 vdd.n6571 0.000501408
R48077 vdd.n3920 vdd.n3919 0.000501408
R48078 vdd.n6623 vdd.n6622 0.000501408
R48079 vdd.n6671 vdd.n6670 0.000501408
R48080 vdd.n6720 vdd.n6719 0.000501408
R48081 vdd.n3872 vdd.n3871 0.000501408
R48082 vdd.n6818 vdd.n6817 0.000501408
R48083 vdd.n681 vdd.n680 0.000501408
R48084 vdd.n1663 vdd.n1662 0.000501408
R48085 vdd.n1664 vdd.n1615 0.000501408
R48086 vdd.n1713 vdd.n1712 0.000501408
R48087 vdd.n1568 vdd.n1567 0.000501408
R48088 vdd.n1811 vdd.n1810 0.000501408
R48089 vdd.n1467 vdd.n1466 0.000501408
R48090 vdd.n1957 vdd.n1956 0.000501408
R48091 vdd.n1909 vdd.n1908 0.000501408
R48092 vdd.n1959 vdd.n1861 0.000501408
R48093 vdd.n2008 vdd.n2007 0.000501408
R48094 vdd.n1419 vdd.n1418 0.000501408
R48095 vdd.n2106 vdd.n2105 0.000501408
R48096 vdd.n1371 vdd.n1370 0.000501408
R48097 vdd.n2203 vdd.n2202 0.000501408
R48098 vdd.n2204 vdd.n2155 0.000501408
R48099 vdd.n2253 vdd.n2252 0.000501408
R48100 vdd.n1323 vdd.n1322 0.000501408
R48101 vdd.n2351 vdd.n2350 0.000501408
R48102 vdd.n1222 vdd.n1221 0.000501408
R48103 vdd.n2449 vdd.n2448 0.000501408
R48104 vdd.n2450 vdd.n2401 0.000501408
R48105 vdd.n2499 vdd.n2498 0.000501408
R48106 vdd.n1174 vdd.n1173 0.000501408
R48107 vdd.n2597 vdd.n2596 0.000501408
R48108 vdd.n2646 vdd.n2645 0.000501408
R48109 vdd.n2695 vdd.n2694 0.000501408
R48110 vdd.n2743 vdd.n2742 0.000501408
R48111 vdd.n2792 vdd.n2791 0.000501408
R48112 vdd.n1126 vdd.n1125 0.000501408
R48113 vdd.n2890 vdd.n2889 0.000501408
R48114 vdd.n1024 vdd.n1023 0.000501408
R48115 vdd.n2941 vdd.n2940 0.000501408
R48116 vdd.n2989 vdd.n2988 0.000501408
R48117 vdd.n3038 vdd.n3037 0.000501408
R48118 vdd.n3087 vdd.n3086 0.000501408
R48119 vdd.n976 vdd.n975 0.000501408
R48120 vdd.n3185 vdd.n3184 0.000501408
R48121 vdd.n928 vdd.n927 0.000501408
R48122 vdd.n3235 vdd.n3234 0.000501408
R48123 vdd.n3283 vdd.n3282 0.000501408
R48124 vdd.n3332 vdd.n3331 0.000501408
R48125 vdd.n880 vdd.n879 0.000501408
R48126 vdd.n3430 vdd.n3429 0.000501408
R48127 vdd.n778 vdd.n777 0.000501408
R48128 vdd.n3481 vdd.n3480 0.000501408
R48129 vdd.n3529 vdd.n3528 0.000501408
R48130 vdd.n3578 vdd.n3577 0.000501408
R48131 vdd.n730 vdd.n729 0.000501408
R48132 vdd.n3676 vdd.n3675 0.000501408
R48133 vdd.n10011 vdd.n10010 0.000501408
R48134 vdd.n10059 vdd.n10058 0.000501408
R48135 vdd.n6869 vdd.n6868 0.000501408
R48136 vdd.n6917 vdd.n6916 0.000501408
R48137 vdd.n3727 vdd.n3726 0.000501408
R48138 vdd.n3775 vdd.n3774 0.000501408
R48139 vdd.n47 vdd.n46 0.000501408
R48140 vdd.n95 vdd.n94 0.000501408
R48141 vdd.n10551 vdd.n10550 0.000501408
R48142 vdd.n10503 vdd.n10502 0.000501408
R48143 vdd.n10649 vdd.n10648 0.000501408
R48144 vdd.n10401 vdd.n10400 0.000501408
R48145 vdd.n10700 vdd.n10699 0.000501408
R48146 vdd.n10748 vdd.n10747 0.000501408
R48147 vdd.n10797 vdd.n10796 0.000501408
R48148 vdd.n10846 vdd.n10845 0.000501408
R48149 vdd.n10353 vdd.n10352 0.000501408
R48150 vdd.n10944 vdd.n10943 0.000501408
R48151 vdd.n10305 vdd.n10304 0.000501408
R48152 vdd.n10994 vdd.n10993 0.000501408
R48153 vdd.n11042 vdd.n11041 0.000501408
R48154 vdd.n11091 vdd.n11090 0.000501408
R48155 vdd.n10257 vdd.n10256 0.000501408
R48156 vdd.n11189 vdd.n11188 0.000501408
R48157 vdd.n10155 vdd.n10154 0.000501408
R48158 vdd.n11240 vdd.n11239 0.000501408
R48159 vdd.n11288 vdd.n11287 0.000501408
R48160 vdd.n11337 vdd.n11336 0.000501408
R48161 vdd.n10107 vdd.n10106 0.000501408
R48162 vdd.n11435 vdd.n11434 0.000501408
R48163 vdd.n586 vdd.n585 0.000501408
R48164 vdd.n11533 vdd.n11532 0.000501408
R48165 vdd.n11534 vdd.n11485 0.000501408
R48166 vdd.n11583 vdd.n11582 0.000501408
R48167 vdd.n538 vdd.n537 0.000501408
R48168 vdd.n11681 vdd.n11680 0.000501408
R48169 vdd.n437 vdd.n436 0.000501408
R48170 vdd.n11827 vdd.n11826 0.000501408
R48171 vdd.n11779 vdd.n11778 0.000501408
R48172 vdd.n11829 vdd.n11731 0.000501408
R48173 vdd.n11878 vdd.n11877 0.000501408
R48174 vdd.n389 vdd.n388 0.000501408
R48175 vdd.n11976 vdd.n11975 0.000501408
R48176 vdd.n341 vdd.n340 0.000501408
R48177 vdd.n12073 vdd.n12072 0.000501408
R48178 vdd.n12074 vdd.n12025 0.000501408
R48179 vdd.n12123 vdd.n12122 0.000501408
R48180 vdd.n293 vdd.n292 0.000501408
R48181 vdd.n12221 vdd.n12220 0.000501408
R48182 vdd.n192 vdd.n191 0.000501408
R48183 vdd.n12319 vdd.n12318 0.000501408
R48184 vdd.n12320 vdd.n12271 0.000501408
R48185 vdd.n12369 vdd.n12368 0.000501408
R48186 vdd.n144 vdd.n143 0.000501408
R48187 vdd.n12467 vdd.n12466 0.000501408
R48188 vdd.n12517 vdd.n12516 0.000501408
R48189 d1.n1 d1.t0 40.0866
R48190 d1.n13 d1.t14 40.0866
R48191 d1.n11 d1.t12 40.0866
R48192 d1.n109 d1.t62 40.0866
R48193 d1.n110 d1.t60 40.0866
R48194 d1.n112 d1.t58 40.0866
R48195 d1.n114 d1.t56 40.0866
R48196 d1.n116 d1.t54 40.0866
R48197 d1.n118 d1.t52 40.0866
R48198 d1.n120 d1.t50 40.0866
R48199 d1.n122 d1.t48 40.0866
R48200 d1.n124 d1.t32 40.0866
R48201 d1.n126 d1.t34 40.0866
R48202 d1.n129 d1.t36 40.0866
R48203 d1.n132 d1.t38 40.0866
R48204 d1.n135 d1.t40 40.0866
R48205 d1.n138 d1.t42 40.0866
R48206 d1.n141 d1.t44 40.0866
R48207 d1.n144 d1.t46 40.0866
R48208 d1.n69 d1.t94 40.0866
R48209 d1.n70 d1.t92 40.0866
R48210 d1.n72 d1.t90 40.0866
R48211 d1.n74 d1.t88 40.0866
R48212 d1.n76 d1.t86 40.0866
R48213 d1.n78 d1.t84 40.0866
R48214 d1.n80 d1.t82 40.0866
R48215 d1.n82 d1.t80 40.0866
R48216 d1.n84 d1.t64 40.0866
R48217 d1.n86 d1.t66 40.0866
R48218 d1.n89 d1.t68 40.0866
R48219 d1.n92 d1.t70 40.0866
R48220 d1.n95 d1.t72 40.0866
R48221 d1.n98 d1.t74 40.0866
R48222 d1.n101 d1.t76 40.0866
R48223 d1.n104 d1.t78 40.0866
R48224 d1.n30 d1.t126 40.0866
R48225 d1.n31 d1.t124 40.0866
R48226 d1.n33 d1.t122 40.0866
R48227 d1.n35 d1.t120 40.0866
R48228 d1.n37 d1.t118 40.0866
R48229 d1.n39 d1.t116 40.0866
R48230 d1.n41 d1.t114 40.0866
R48231 d1.n43 d1.t112 40.0866
R48232 d1.n45 d1.t96 40.0866
R48233 d1.n47 d1.t98 40.0866
R48234 d1.n50 d1.t100 40.0866
R48235 d1.n53 d1.t102 40.0866
R48236 d1.n56 d1.t104 40.0866
R48237 d1.n59 d1.t106 40.0866
R48238 d1.n62 d1.t108 40.0866
R48239 d1.n65 d1.t110 40.0866
R48240 d1.n15 d1.t30 40.0866
R48241 d1.n16 d1.t28 40.0866
R48242 d1.n18 d1.t26 40.0866
R48243 d1.n20 d1.t24 40.0866
R48244 d1.n22 d1.t22 40.0866
R48245 d1.n24 d1.t20 40.0866
R48246 d1.n26 d1.t18 40.0866
R48247 d1.n28 d1.t16 40.0866
R48248 d1.n9 d1.t10 40.0866
R48249 d1.n7 d1.t8 40.0866
R48250 d1.n5 d1.t6 40.0866
R48251 d1.n3 d1.t4 40.0866
R48252 d1.n0 d1.t2 40.0866
R48253 d1.n108 d1.n68 25.9475
R48254 d1.n149 d1.n148 25.9475
R48255 d1.n13 d1.t15 23.8528
R48256 d1.n11 d1.t13 23.8528
R48257 d1.n109 d1.t63 23.8528
R48258 d1.n110 d1.t61 23.8528
R48259 d1.n112 d1.t59 23.8528
R48260 d1.n114 d1.t57 23.8528
R48261 d1.n116 d1.t55 23.8528
R48262 d1.n118 d1.t53 23.8528
R48263 d1.n120 d1.t51 23.8528
R48264 d1.n122 d1.t49 23.8528
R48265 d1.n124 d1.t33 23.8528
R48266 d1.n126 d1.t35 23.8528
R48267 d1.n129 d1.t37 23.8528
R48268 d1.n132 d1.t39 23.8528
R48269 d1.n135 d1.t41 23.8528
R48270 d1.n138 d1.t43 23.8528
R48271 d1.n141 d1.t45 23.8528
R48272 d1.n144 d1.t47 23.8528
R48273 d1.n69 d1.t95 23.8528
R48274 d1.n70 d1.t93 23.8528
R48275 d1.n72 d1.t91 23.8528
R48276 d1.n74 d1.t89 23.8528
R48277 d1.n76 d1.t87 23.8528
R48278 d1.n78 d1.t85 23.8528
R48279 d1.n80 d1.t83 23.8528
R48280 d1.n82 d1.t81 23.8528
R48281 d1.n84 d1.t65 23.8528
R48282 d1.n86 d1.t67 23.8528
R48283 d1.n89 d1.t69 23.8528
R48284 d1.n92 d1.t71 23.8528
R48285 d1.n95 d1.t73 23.8528
R48286 d1.n98 d1.t75 23.8528
R48287 d1.n101 d1.t77 23.8528
R48288 d1.n104 d1.t79 23.8528
R48289 d1.n30 d1.t127 23.8528
R48290 d1.n31 d1.t125 23.8528
R48291 d1.n33 d1.t123 23.8528
R48292 d1.n35 d1.t121 23.8528
R48293 d1.n37 d1.t119 23.8528
R48294 d1.n39 d1.t117 23.8528
R48295 d1.n41 d1.t115 23.8528
R48296 d1.n43 d1.t113 23.8528
R48297 d1.n45 d1.t97 23.8528
R48298 d1.n47 d1.t99 23.8528
R48299 d1.n50 d1.t101 23.8528
R48300 d1.n53 d1.t103 23.8528
R48301 d1.n56 d1.t105 23.8528
R48302 d1.n59 d1.t107 23.8528
R48303 d1.n62 d1.t109 23.8528
R48304 d1.n65 d1.t111 23.8528
R48305 d1.n15 d1.t31 23.8528
R48306 d1.n16 d1.t29 23.8528
R48307 d1.n18 d1.t27 23.8528
R48308 d1.n20 d1.t25 23.8528
R48309 d1.n22 d1.t23 23.8528
R48310 d1.n24 d1.t21 23.8528
R48311 d1.n26 d1.t19 23.8528
R48312 d1.n28 d1.t17 23.8528
R48313 d1.n9 d1.t11 23.8528
R48314 d1.n7 d1.t9 23.8528
R48315 d1.n5 d1.t7 23.8528
R48316 d1.n3 d1.t5 23.8528
R48317 d1.n0 d1.t3 23.8528
R48318 d1.n1 d1.t1 23.8528
R48319 d1.n148 d1.n108 22.8755
R48320 d1.n147 d1.n146 10.6976
R48321 d1.n107 d1.n106 10.6976
R48322 d1.n68 d1.n67 10.6976
R48323 d1.n150 d1.n149 10.6976
R48324 d1.n111 d1 5.95687
R48325 d1.n128 d1.n125 5.95687
R48326 d1.n71 d1 5.95687
R48327 d1.n88 d1.n85 5.95687
R48328 d1.n32 d1 5.95687
R48329 d1.n49 d1.n46 5.95687
R48330 d1.n17 d1 5.95687
R48331 d1.n156 d1.n2 5.95687
R48332 d1.n115 d1.n113 5.95675
R48333 d1.n117 d1.n115 5.95675
R48334 d1.n119 d1.n117 5.95675
R48335 d1.n134 d1.n131 5.95675
R48336 d1.n137 d1.n134 5.95675
R48337 d1.n140 d1.n137 5.95675
R48338 d1.n146 d1.n143 5.95675
R48339 d1.n123 d1.n121 5.95675
R48340 d1.n75 d1.n73 5.95675
R48341 d1.n77 d1.n75 5.95675
R48342 d1.n79 d1.n77 5.95675
R48343 d1.n94 d1.n91 5.95675
R48344 d1.n97 d1.n94 5.95675
R48345 d1.n100 d1.n97 5.95675
R48346 d1.n106 d1.n103 5.95675
R48347 d1.n83 d1.n81 5.95675
R48348 d1.n36 d1.n34 5.95675
R48349 d1.n38 d1.n36 5.95675
R48350 d1.n40 d1.n38 5.95675
R48351 d1.n55 d1.n52 5.95675
R48352 d1.n58 d1.n55 5.95675
R48353 d1.n61 d1.n58 5.95675
R48354 d1.n67 d1.n64 5.95675
R48355 d1.n44 d1.n42 5.95675
R48356 d1.n21 d1.n19 5.95675
R48357 d1.n23 d1.n21 5.95675
R48358 d1.n25 d1.n23 5.95675
R48359 d1.n29 d1.n27 5.95675
R48360 d1.n151 d1.n150 5.95675
R48361 d1.n155 d1.n154 5.95675
R48362 d1.n154 d1.n153 5.95675
R48363 d1.n153 d1.n152 5.95675
R48364 d1.n113 d1.n111 5.36034
R48365 d1.n121 d1.n119 5.36034
R48366 d1.n73 d1.n71 5.36034
R48367 d1.n81 d1.n79 5.36034
R48368 d1.n34 d1.n32 5.36034
R48369 d1.n42 d1.n40 5.36034
R48370 d1.n19 d1.n17 5.36034
R48371 d1.n27 d1.n25 5.36034
R48372 d1.n152 d1.n151 5.36034
R48373 d1.n156 d1.n155 5.36034
R48374 d1.n131 d1.n128 5.36034
R48375 d1.n143 d1.n140 5.36034
R48376 d1.n91 d1.n88 5.36034
R48377 d1.n103 d1.n100 5.36034
R48378 d1.n52 d1.n49 5.36034
R48379 d1.n64 d1.n61 5.36034
R48380 d1.n148 d1.n147 3.07249
R48381 d1.n108 d1.n107 3.07249
R48382 d1.n147 d1.n123 1.82237
R48383 d1.n107 d1.n83 1.82237
R48384 d1.n68 d1.n44 1.82237
R48385 d1.n149 d1.n29 1.82237
R48386 d1.n14 d1.n13 0.2505
R48387 d1.n12 d1.n11 0.2505
R48388 d1 d1.n109 0.2505
R48389 d1 d1.n112 0.2505
R48390 d1 d1.n116 0.2505
R48391 d1 d1.n120 0.2505
R48392 d1.n125 d1.n124 0.2505
R48393 d1.n127 d1.n126 0.2505
R48394 d1.n130 d1.n129 0.2505
R48395 d1.n133 d1.n132 0.2505
R48396 d1.n136 d1.n135 0.2505
R48397 d1.n139 d1.n138 0.2505
R48398 d1.n142 d1.n141 0.2505
R48399 d1.n145 d1.n144 0.2505
R48400 d1 d1.n69 0.2505
R48401 d1 d1.n72 0.2505
R48402 d1 d1.n76 0.2505
R48403 d1 d1.n80 0.2505
R48404 d1.n85 d1.n84 0.2505
R48405 d1.n87 d1.n86 0.2505
R48406 d1.n90 d1.n89 0.2505
R48407 d1.n93 d1.n92 0.2505
R48408 d1.n96 d1.n95 0.2505
R48409 d1.n99 d1.n98 0.2505
R48410 d1.n102 d1.n101 0.2505
R48411 d1.n105 d1.n104 0.2505
R48412 d1 d1.n30 0.2505
R48413 d1 d1.n33 0.2505
R48414 d1 d1.n37 0.2505
R48415 d1 d1.n41 0.2505
R48416 d1.n46 d1.n45 0.2505
R48417 d1.n48 d1.n47 0.2505
R48418 d1.n51 d1.n50 0.2505
R48419 d1.n54 d1.n53 0.2505
R48420 d1.n57 d1.n56 0.2505
R48421 d1.n60 d1.n59 0.2505
R48422 d1.n63 d1.n62 0.2505
R48423 d1.n66 d1.n65 0.2505
R48424 d1 d1.n15 0.2505
R48425 d1 d1.n18 0.2505
R48426 d1 d1.n22 0.2505
R48427 d1 d1.n26 0.2505
R48428 d1.n10 d1.n9 0.2505
R48429 d1.n8 d1.n7 0.2505
R48430 d1.n6 d1.n5 0.2505
R48431 d1.n4 d1.n3 0.2505
R48432 d1.n157 d1.n0 0.2505
R48433 d1.n2 d1.n1 0.2505
R48434 d1 d1.n110 0.188
R48435 d1 d1.n114 0.188
R48436 d1 d1.n118 0.188
R48437 d1 d1.n122 0.188
R48438 d1 d1.n70 0.188
R48439 d1 d1.n74 0.188
R48440 d1 d1.n78 0.188
R48441 d1 d1.n82 0.188
R48442 d1 d1.n31 0.188
R48443 d1 d1.n35 0.188
R48444 d1 d1.n39 0.188
R48445 d1 d1.n43 0.188
R48446 d1 d1.n16 0.188
R48447 d1 d1.n20 0.188
R48448 d1 d1.n24 0.188
R48449 d1 d1.n28 0.188
R48450 d1.n14 d1 0.063
R48451 d1.n12 d1 0.063
R48452 d1 d1 0.063
R48453 d1 d1 0.063
R48454 d1 d1 0.063
R48455 d1 d1 0.063
R48456 d1.n125 d1 0.063
R48457 d1.n127 d1 0.063
R48458 d1.n130 d1 0.063
R48459 d1.n133 d1 0.063
R48460 d1.n136 d1 0.063
R48461 d1.n139 d1 0.063
R48462 d1.n142 d1 0.063
R48463 d1.n145 d1 0.063
R48464 d1 d1 0.063
R48465 d1 d1 0.063
R48466 d1 d1 0.063
R48467 d1 d1 0.063
R48468 d1.n85 d1 0.063
R48469 d1.n87 d1 0.063
R48470 d1.n90 d1 0.063
R48471 d1.n93 d1 0.063
R48472 d1.n96 d1 0.063
R48473 d1.n99 d1 0.063
R48474 d1.n102 d1 0.063
R48475 d1.n105 d1 0.063
R48476 d1 d1 0.063
R48477 d1 d1 0.063
R48478 d1 d1 0.063
R48479 d1 d1 0.063
R48480 d1.n46 d1 0.063
R48481 d1.n48 d1 0.063
R48482 d1.n51 d1 0.063
R48483 d1.n54 d1 0.063
R48484 d1.n57 d1 0.063
R48485 d1.n60 d1 0.063
R48486 d1.n63 d1 0.063
R48487 d1.n66 d1 0.063
R48488 d1 d1 0.063
R48489 d1 d1 0.063
R48490 d1 d1 0.063
R48491 d1 d1 0.063
R48492 d1.n10 d1 0.063
R48493 d1.n8 d1 0.063
R48494 d1.n6 d1 0.063
R48495 d1.n4 d1 0.063
R48496 d1 d1.n157 0.063
R48497 d1.n2 d1 0.063
R48498 d1.n111 d1 0.000617139
R48499 d1.n119 d1 0.000617139
R48500 d1.n117 d1 0.000617139
R48501 d1.n115 d1 0.000617139
R48502 d1.n113 d1 0.000617139
R48503 d1.n128 d1.n127 0.000617139
R48504 d1.n140 d1.n139 0.000617139
R48505 d1.n137 d1.n136 0.000617139
R48506 d1.n134 d1.n133 0.000617139
R48507 d1.n131 d1.n130 0.000617139
R48508 d1.n146 d1.n145 0.000617139
R48509 d1.n143 d1.n142 0.000617139
R48510 d1.n123 d1 0.000617139
R48511 d1.n121 d1 0.000617139
R48512 d1.n71 d1 0.000617139
R48513 d1.n79 d1 0.000617139
R48514 d1.n77 d1 0.000617139
R48515 d1.n75 d1 0.000617139
R48516 d1.n73 d1 0.000617139
R48517 d1.n88 d1.n87 0.000617139
R48518 d1.n100 d1.n99 0.000617139
R48519 d1.n97 d1.n96 0.000617139
R48520 d1.n94 d1.n93 0.000617139
R48521 d1.n91 d1.n90 0.000617139
R48522 d1.n106 d1.n105 0.000617139
R48523 d1.n103 d1.n102 0.000617139
R48524 d1.n83 d1 0.000617139
R48525 d1.n81 d1 0.000617139
R48526 d1.n32 d1 0.000617139
R48527 d1.n40 d1 0.000617139
R48528 d1.n38 d1 0.000617139
R48529 d1.n36 d1 0.000617139
R48530 d1.n34 d1 0.000617139
R48531 d1.n49 d1.n48 0.000617139
R48532 d1.n61 d1.n60 0.000617139
R48533 d1.n58 d1.n57 0.000617139
R48534 d1.n55 d1.n54 0.000617139
R48535 d1.n52 d1.n51 0.000617139
R48536 d1.n67 d1.n66 0.000617139
R48537 d1.n64 d1.n63 0.000617139
R48538 d1.n44 d1 0.000617139
R48539 d1.n42 d1 0.000617139
R48540 d1.n17 d1 0.000617139
R48541 d1.n25 d1 0.000617139
R48542 d1.n23 d1 0.000617139
R48543 d1.n21 d1 0.000617139
R48544 d1.n19 d1 0.000617139
R48545 d1.n29 d1 0.000617139
R48546 d1.n27 d1 0.000617139
R48547 d1.n151 d1.n12 0.000617139
R48548 d1.n150 d1.n14 0.000617139
R48549 d1.n155 d1.n4 0.000617139
R48550 d1.n154 d1.n6 0.000617139
R48551 d1.n153 d1.n8 0.000617139
R48552 d1.n152 d1.n10 0.000617139
R48553 d1.n157 d1.n156 0.000617139
R48554 d2.n66 d2.t0 40.0866
R48555 d2.n55 d2.t16 40.0866
R48556 d2.n56 d2.t22 40.0866
R48557 d2.n53 d2.t30 40.0866
R48558 d2.n47 d2.t28 40.0866
R48559 d2.n48 d2.t26 40.0866
R48560 d2.n49 d2.t24 40.0866
R48561 d2.n58 d2.t20 40.0866
R48562 d2.n60 d2.t18 40.0866
R48563 d2.n37 d2.t32 40.0866
R48564 d2.n38 d2.t38 40.0866
R48565 d2.n35 d2.t46 40.0866
R48566 d2.n29 d2.t44 40.0866
R48567 d2.n30 d2.t42 40.0866
R48568 d2.n31 d2.t40 40.0866
R48569 d2.n40 d2.t36 40.0866
R48570 d2.n42 d2.t34 40.0866
R48571 d2.n20 d2.t48 40.0866
R48572 d2.n21 d2.t54 40.0866
R48573 d2.n18 d2.t62 40.0866
R48574 d2.n12 d2.t60 40.0866
R48575 d2.n13 d2.t58 40.0866
R48576 d2.n14 d2.t56 40.0866
R48577 d2.n23 d2.t52 40.0866
R48578 d2.n25 d2.t50 40.0866
R48579 d2.n2 d2.t6 40.0866
R48580 d2.n10 d2.t14 40.0866
R48581 d2.n6 d2.t12 40.0866
R48582 d2.n7 d2.t10 40.0866
R48583 d2.n0 d2.t8 40.0866
R48584 d2.n4 d2.t4 40.0866
R48585 d2.n69 d2.t2 40.0866
R48586 d2.n65 d2.n64 25.7145
R48587 d2.n46 d2.n28 25.7131
R48588 d2.n55 d2.t17 23.8528
R48589 d2.n56 d2.t23 23.8528
R48590 d2.n53 d2.t31 23.8528
R48591 d2.n47 d2.t29 23.8528
R48592 d2.n48 d2.t27 23.8528
R48593 d2.n49 d2.t25 23.8528
R48594 d2.n58 d2.t21 23.8528
R48595 d2.n60 d2.t19 23.8528
R48596 d2.n37 d2.t33 23.8528
R48597 d2.n38 d2.t39 23.8528
R48598 d2.n35 d2.t47 23.8528
R48599 d2.n29 d2.t45 23.8528
R48600 d2.n30 d2.t43 23.8528
R48601 d2.n31 d2.t41 23.8528
R48602 d2.n40 d2.t37 23.8528
R48603 d2.n42 d2.t35 23.8528
R48604 d2.n20 d2.t49 23.8528
R48605 d2.n21 d2.t55 23.8528
R48606 d2.n18 d2.t63 23.8528
R48607 d2.n12 d2.t61 23.8528
R48608 d2.n13 d2.t59 23.8528
R48609 d2.n14 d2.t57 23.8528
R48610 d2.n23 d2.t53 23.8528
R48611 d2.n25 d2.t51 23.8528
R48612 d2.n2 d2.t7 23.8528
R48613 d2.n10 d2.t15 23.8528
R48614 d2.n6 d2.t13 23.8528
R48615 d2.n7 d2.t11 23.8528
R48616 d2.n0 d2.t9 23.8528
R48617 d2.n4 d2.t5 23.8528
R48618 d2.n69 d2.t3 23.8528
R48619 d2.n66 d2.t1 23.8528
R48620 d2.n64 d2.n46 20.7519
R48621 d2.n59 d2.n57 9.35243
R48622 d2.n41 d2.n39 9.35243
R48623 d2.n24 d2.n22 9.35243
R48624 d2.n5 d2.n3 9.35243
R48625 d2.n62 d2.n61 9.35243
R48626 d2.n44 d2.n43 9.35243
R48627 d2.n27 d2.n26 9.35243
R48628 d2.n68 d2.n67 9.35243
R48629 d2.n54 d2.n52 9.33579
R48630 d2.n36 d2.n34 9.33579
R48631 d2.n19 d2.n17 9.33579
R48632 d2.n11 d2.n9 9.33579
R48633 d2.n51 d2.n50 9.32359
R48634 d2.n33 d2.n32 9.32359
R48635 d2.n16 d2.n15 9.32359
R48636 d2.n52 d2.n51 9.24786
R48637 d2.n61 d2.n59 9.24786
R48638 d2.n34 d2.n33 9.24786
R48639 d2.n43 d2.n41 9.24786
R48640 d2.n17 d2.n16 9.24786
R48641 d2.n26 d2.n24 9.24786
R48642 d2.n9 d2.n8 9.24786
R48643 d2.n68 d2.n5 9.24786
R48644 d2.n46 d2.n45 5.79918
R48645 d2.n64 d2.n63 5.7978
R48646 d2.n3 d2.n1 2.79465
R48647 d2.n45 d2.n44 1.51198
R48648 d2.n67 d2.n65 1.51198
R48649 d2.n63 d2.n54 1.39016
R48650 d2.n28 d2.n19 1.39016
R48651 d2.n63 d2.n62 1.35282
R48652 d2.n28 d2.n27 1.35282
R48653 d2.n45 d2.n36 1.231
R48654 d2.n65 d2.n11 1.231
R48655 d2.n52 d2.n47 0.624393
R48656 d2.n51 d2.n48 0.624393
R48657 d2.n59 d2.n58 0.624393
R48658 d2.n61 d2.n60 0.624393
R48659 d2.n34 d2.n29 0.624393
R48660 d2.n33 d2.n30 0.624393
R48661 d2.n41 d2.n40 0.624393
R48662 d2.n43 d2.n42 0.624393
R48663 d2.n17 d2.n12 0.624393
R48664 d2.n16 d2.n13 0.624393
R48665 d2.n24 d2.n23 0.624393
R48666 d2.n26 d2.n25 0.624393
R48667 d2.n9 d2.n6 0.624393
R48668 d2.n8 d2.n7 0.624393
R48669 d2.n5 d2.n4 0.624393
R48670 d2.n69 d2.n68 0.624393
R48671 d2.n55 d2 0.313
R48672 d2.n56 d2 0.313
R48673 d2.n58 d2 0.313
R48674 d2.n60 d2 0.313
R48675 d2.n37 d2 0.313
R48676 d2.n38 d2 0.313
R48677 d2.n40 d2 0.313
R48678 d2.n42 d2 0.313
R48679 d2.n20 d2 0.313
R48680 d2.n21 d2 0.313
R48681 d2.n23 d2 0.313
R48682 d2.n25 d2 0.313
R48683 d2.n2 d2 0.313
R48684 d2.n4 d2 0.313
R48685 d2 d2.n69 0.313
R48686 d2.n66 d2 0.313
R48687 d2.n62 d2.n55 0.301802
R48688 d2.n57 d2.n56 0.301802
R48689 d2.n54 d2.n53 0.301802
R48690 d2.n50 d2.n49 0.301802
R48691 d2.n44 d2.n37 0.301802
R48692 d2.n39 d2.n38 0.301802
R48693 d2.n36 d2.n35 0.301802
R48694 d2.n32 d2.n31 0.301802
R48695 d2.n27 d2.n20 0.301802
R48696 d2.n22 d2.n21 0.301802
R48697 d2.n19 d2.n18 0.301802
R48698 d2.n15 d2.n14 0.301802
R48699 d2.n3 d2.n2 0.301802
R48700 d2.n11 d2.n10 0.301802
R48701 d2.n1 d2.n0 0.301802
R48702 d2.n67 d2.n66 0.301802
R48703 d2.n53 d2 0.188
R48704 d2.n47 d2 0.188
R48705 d2.n48 d2 0.188
R48706 d2.n49 d2 0.188
R48707 d2.n35 d2 0.188
R48708 d2.n29 d2 0.188
R48709 d2.n30 d2 0.188
R48710 d2.n31 d2 0.188
R48711 d2.n18 d2 0.188
R48712 d2.n12 d2 0.188
R48713 d2.n13 d2 0.188
R48714 d2.n14 d2 0.188
R48715 d2.n10 d2 0.188
R48716 d2.n6 d2 0.188
R48717 d2.n7 d2 0.188
R48718 d2.n0 d2 0.188
R48719 d2 d2 0.063
R48720 d2 d2 0.063
R48721 d2 d2 0.063
R48722 d2 d2 0.063
R48723 d2 d2 0.063
R48724 d2 d2 0.063
R48725 d2 d2 0.063
R48726 d2 d2 0.063
R48727 d2 d2 0.063
R48728 d2 d2 0.063
R48729 d2 d2 0.063
R48730 d2 d2 0.063
R48731 d2 d2 0.063
R48732 d2 d2 0.063
R48733 d2 d2 0.063
R48734 d2 d2 0.063
R48735 d3.n64 d3.t0 40.0866
R48736 d3.n51 d3.t12 40.0866
R48737 d3.n41 d3.t8 40.0866
R48738 d3.n15 d3.t30 40.0866
R48739 d3.n1 d3.t26 40.0866
R48740 d3.n10 d3.t28 40.0866
R48741 d3.n0 d3.t24 40.0866
R48742 d3.n20 d3.t22 40.0866
R48743 d3.n35 d3.t16 40.0866
R48744 d3.n30 d3.t18 40.0866
R48745 d3.n21 d3.t20 40.0866
R48746 d3.n56 d3.t14 40.0795
R48747 d3.n42 d3.t10 40.0795
R48748 d3.n62 d3.t6 40.0795
R48749 d3.n81 d3.t4 40.0322
R48750 d3.n74 d3.t2 40.0251
R48751 d3.n40 d3.n19 31.476
R48752 d3.n63 d3.n61 31.4135
R48753 d3.n56 d3.t15 23.8528
R48754 d3.n42 d3.t11 23.8528
R48755 d3.n51 d3.t13 23.8528
R48756 d3.n15 d3.t31 23.8528
R48757 d3.n1 d3.t27 23.8528
R48758 d3.n10 d3.t29 23.8528
R48759 d3.n0 d3.t25 23.8528
R48760 d3.n20 d3.t23 23.8528
R48761 d3.n30 d3.t19 23.8528
R48762 d3.n21 d3.t21 23.8528
R48763 d3.n62 d3.t7 23.8528
R48764 d3.n41 d3.t9 23.8457
R48765 d3.n35 d3.t17 23.8457
R48766 d3.n64 d3.t1 23.8457
R48767 d3.n81 d3.t5 23.7914
R48768 d3.n74 d3.t3 23.7914
R48769 d3.n61 d3.n40 21.8199
R48770 d3.n61 d3.n60 12.6287
R48771 d3.n40 d3.n39 12.5662
R48772 d3.n58 d3.n50 6.088
R48773 d3.n59 d3.n46 6.088
R48774 d3.n57 d3.n55 6.088
R48775 d3.n17 d3.n9 6.088
R48776 d3.n18 d3.n5 6.088
R48777 d3.n16 d3.n14 6.088
R48778 d3.n37 d3.n29 6.088
R48779 d3.n36 d3.n34 6.088
R48780 d3.n38 d3.n25 6.088
R48781 d3.n68 d3.n67 6.088
R48782 d3.n54 d3.n53 5.88488
R48783 d3.n45 d3.n44 5.88488
R48784 d3.n49 d3.n48 5.88488
R48785 d3.n13 d3.n12 5.88488
R48786 d3.n4 d3.n3 5.88488
R48787 d3.n8 d3.n7 5.88488
R48788 d3.n24 d3.n23 5.88488
R48789 d3.n33 d3.n32 5.88488
R48790 d3.n28 d3.n27 5.88488
R48791 d3.n70 d3.n69 5.88488
R48792 d3.n77 d3.n76 5.88488
R48793 d3.n73 d3.n72 5.88488
R48794 d3.n53 d3.n52 5.65675
R48795 d3.n48 d3.n47 5.65675
R48796 d3.n44 d3.n43 5.65675
R48797 d3.n12 d3.n11 5.65675
R48798 d3.n7 d3.n6 5.65675
R48799 d3.n3 d3.n2 5.65675
R48800 d3.n23 d3.n22 5.65675
R48801 d3.n27 d3.n26 5.65675
R48802 d3.n32 d3.n31 5.65675
R48803 d3.n80 d3.n70 5.65675
R48804 d3.n79 d3.n73 5.65675
R48805 d3.n78 d3.n77 5.65675
R48806 d3.n55 d3.n54 5.51612
R48807 d3.n50 d3.n49 5.51612
R48808 d3.n46 d3.n45 5.51612
R48809 d3.n14 d3.n13 5.51612
R48810 d3.n9 d3.n8 5.51612
R48811 d3.n5 d3.n4 5.51612
R48812 d3.n25 d3.n24 5.51612
R48813 d3.n29 d3.n28 5.51612
R48814 d3.n34 d3.n33 5.51612
R48815 d3.n69 d3.n68 5.51612
R48816 d3.n72 d3.n71 5.51612
R48817 d3.n76 d3.n75 5.51612
R48818 d3.n52 d3.n51 1.59714
R48819 d3.n11 d3.n10 1.59714
R48820 d3.n36 d3.n35 1.59714
R48821 d3.n22 d3.n21 1.59714
R48822 d3.n81 d3.n80 1.59714
R48823 d3.n65 d3.n64 1.59714
R48824 d3.n60 d3.n41 1.59703
R48825 d3.n19 d3.n0 1.59703
R48826 d3.n57 d3.n56 1.45966
R48827 d3.n43 d3.n42 1.45966
R48828 d3.n16 d3.n15 1.45966
R48829 d3.n2 d3.n1 1.45966
R48830 d3.n31 d3.n30 1.45966
R48831 d3.n78 d3.n74 1.45966
R48832 d3.n39 d3.n20 1.27758
R48833 d3.n63 d3.n62 1.27758
R48834 d3.n74 d3 0.384875
R48835 d3.n58 d3.n57 0.332778
R48836 d3.n59 d3.n58 0.332778
R48837 d3.n17 d3.n16 0.332778
R48838 d3.n18 d3.n17 0.332778
R48839 d3.n38 d3.n37 0.332778
R48840 d3.n37 d3.n36 0.332778
R48841 d3.n80 d3.n79 0.332778
R48842 d3.n79 d3.n78 0.332778
R48843 d3.n67 d3.n66 0.332778
R48844 d3.n66 d3.n65 0.332778
R48845 d3.n42 d3 0.313
R48846 d3.n41 d3 0.313
R48847 d3.n1 d3 0.313
R48848 d3.n0 d3 0.313
R48849 d3.n35 d3 0.313
R48850 d3.n30 d3 0.313
R48851 d3.n64 d3 0.313
R48852 d3 d3.n81 0.259875
R48853 d3.n56 d3 0.2505
R48854 d3.n15 d3 0.2505
R48855 d3.n20 d3 0.2505
R48856 d3.n62 d3 0.2505
R48857 d3.n51 d3 0.188
R48858 d3.n10 d3 0.188
R48859 d3.n21 d3 0.188
R48860 d3.n39 d3.n38 0.182579
R48861 d3.n67 d3.n63 0.182579
R48862 d3 d3 0.063
R48863 d3 d3 0.063
R48864 d3 d3 0.063
R48865 d3 d3 0.063
R48866 d3.n60 d3.n59 0.000617139
R48867 d3.n19 d3.n18 0.000617139
R48868 d4.n8 d4.n3 45.8392
R48869 d4.n15 d4.n13 45.8392
R48870 d4.n14 d4.t0 40.0866
R48871 d4.n11 d4.t4 40.0866
R48872 d4.n6 d4.t8 40.0866
R48873 d4.n2 d4.t12 40.0866
R48874 d4.n10 d4.t6 40.0322
R48875 d4.n5 d4.t10 40.0322
R48876 d4.n1 d4.t14 40.0322
R48877 d4.n16 d4.t2 40.0322
R48878 d4.n13 d4.n12 24.8948
R48879 d4.n8 d4.n7 24.8948
R48880 d4.n9 d4.t7 23.8528
R48881 d4.n11 d4.t5 23.8528
R48882 d4.n4 d4.t11 23.8528
R48883 d4.n6 d4.t9 23.8528
R48884 d4.n0 d4.t15 23.8528
R48885 d4.n2 d4.t13 23.8528
R48886 d4.n17 d4.t3 23.8528
R48887 d4.n14 d4.t1 23.8528
R48888 d4.n13 d4.n8 19.7227
R48889 d4.n12 d4.n11 1.76105
R48890 d4.n3 d4.n2 1.76105
R48891 d4.n7 d4.n5 1.74408
R48892 d4.n16 d4.n15 1.74408
R48893 d4.n15 d4.n14 1.51486
R48894 d4.n7 d4.n6 1.51486
R48895 d4.n12 d4.n10 1.49789
R48896 d4.n3 d4.n1 1.49789
R48897 d4.n11 d4 0.313
R48898 d4.n6 d4 0.313
R48899 d4.n2 d4 0.313
R48900 d4.n14 d4 0.313
R48901 d4.n9 d4 0.188
R48902 d4.n4 d4 0.188
R48903 d4.n0 d4 0.188
R48904 d4 d4.n17 0.188
R48905 d4 d4 0.063
R48906 d4 d4 0.063
R48907 d4 d4 0.063
R48908 d4 d4 0.063
R48909 d4.n10 d4.n9 0.0548478
R48910 d4.n5 d4.n4 0.0548478
R48911 d4.n1 d4.n0 0.0548478
R48912 d4.n17 d4.n16 0.0548478
R48913 d5.n4 d5.t0 40.0866
R48914 d5.n2 d5.t4 40.0866
R48915 d5.n1 d5.t6 40.0866
R48916 d5.n0 d5.t2 40.0866
R48917 d5.n3 d5 24.7257
R48918 d5.n5 d5 24.4414
R48919 d5.n2 d5.t5 23.8528
R48920 d5.n1 d5.t7 23.8528
R48921 d5.n0 d5.t3 23.8528
R48922 d5.n4 d5.t1 23.8528
R48923 d5.n5 d5.n3 23.1567
R48924 d5 d5.n5 2.13198
R48925 d5.n3 d5 1.84761
R48926 d5 d5.n2 0.313
R48927 d5 d5.n1 0.313
R48928 d5 d5.n0 0.313
R48929 d5 d5.n4 0.313
R48930 d6 d6 48.8947
R48931 d6.n1 d6.t0 40.0866
R48932 d6.n0 d6.t2 40.0866
R48933 d6.n0 d6.t3 23.8528
R48934 d6.n1 d6.t1 23.8528
R48935 d6 d6.n0 0.313
R48936 d6 d6.n1 0.313
R48937 vrefl.n0 vrefl 3.74286
R48938 vrefl vrefl.n0 0.0363796
R48939 vrefl.n0 vrefl 0.016125
R48940 vrefl vrefl 0.00223611
R48941 vrefl vrefl 0.00165741
R48942 vrefl vrefl 0.0010787
R48943 vrefl vrefl 0.0010787
R48944 d7.n0 d7.t0 40.0866
R48945 d7.n0 d7.t1 23.8528
R48946 d7 d7.n0 0.313
R48947 vout vout 0.00354878
C0 d6 d7 5.23e-19
C1 d2 X1/X2/X1/X1/X1/X1/X1/vin1 -0.0257f
C2 X1/X2/X2/X1/X1/X2/X2/vin1 X2/X1/X1/X2/X2/X1/X1/vin2 0.00232f
C3 X2/X1/X1/X1/X1/X2/vrefh X2/X1/X1/X1/X1/X2/X1/vin1 7.11e-33
C4 X1/X2/X2/X1/X2/vrefh X2/X1/X1/X2/X2/X1/X1/vin2 0.0128f
C5 X1/X2/X2/X2/X2/X2/X1/vin1 X2/X1/X1/X1/X1/X2/vrefh 0.00437f
C6 X2/X1/X3/vin2 d5 -0.00244f
C7 d0 X1/X2/X2/X1/X1/X2/vrefh 0.00385f
C8 d0 X3/vin1 0.0184f
C9 d0 X2/X1/X3/vin1 -0.00274f
C10 d4 X2/X1/X1/X1/X1/X1/X1/vin2 8.21e-20
C11 d1 X1/X2/X3/vin1 -0.00249f
C12 X1/X3/vin1 X1/X3/vin2 -1.23e-20
C13 X1/X2/X2/X1/X1/X1/X2/vin1 X2/X1/X1/X2/X2/X2/X1/vin2 0.00232f
C14 X1/X2/X2/X1/X1/X2/X1/vin2 X2/X1/X1/X2/X2/X1/X2/vin1 0.00232f
C15 d1 X3/vin1 0.0325f
C16 d1 X2/X1/X3/vin1 0.0416f
C17 d2 d3 4.92f
C18 X2/X1/X3/m1_994_178# d6 0.00105f
C19 X1/X2/X2/X1/X2/X2/vrefh X2/X1/X1/X2/X1/X2/X1/vin2 0.0128f
C20 X2/X3/vin1 d1 0.0144f
C21 d4 X2/vrefh 0.00449f
C22 X1/X2/X2/X1/X1/X1/X1/vin1 X2/X1/X2/vrefh 0.00437f
C23 X1/X2/X2/X2/vrefh X2/X1/X1/X2/X1/X1/X1/vin2 0.0128f
C24 X1/X2/X2/X1/X2/vrefh X2/X1/X1/X2/X2/vrefh 0.117f
C25 d2 X2/X1/X1/X1/X1/X1/X1/m1_688_n494# 1.95e-19
C26 X1/X2/X2/X2/X2/X1/X1/vin1 X2/X1/X1/X1/X2/vrefh 0.00437f
C27 X2/X3/m1_994_178# d6 0.0045f
C28 X1/X2/X2/X2/X1/X2/X2/vin1 X2/X1/X1/X1/X2/X1/X1/vin2 0.00232f
C29 X1/X2/X2/X2/X2/X1/X1/vin2 X2/X1/X1/X1/X1/X2/X2/vin1 0.00232f
C30 X1/X2/X2/X2/X2/X2/X2/vin1 X2/X1/X1/X1/X1/X1/X1/vin2 0.00232f
C31 X1/X2/X2/X2/X1/X1/X1/vin2 X2/X1/X1/X1/X2/X2/X2/vin1 0.00232f
C32 X1/X2/X3/vin1 d5 0.0463f
C33 d5 X3/vin1 0.0663f
C34 d5 X2/X1/X3/vin1 -0.00244f
C35 X2/X3/vin2 X2/X3/m1_688_n494# -0.0081f
C36 d4 X1/X2/X2/X2/X2/X2/X2/m1_688_n494# 8.99e-20
C37 d0 d1 3.64f
C38 X1/X2/X2/X2/X2/X1/X2/vin1 X2/X1/X1/X1/X1/X2/X1/vin2 0.00232f
C39 X1/X2/X2/X2/X2/X2/X1/vin2 X2/X1/X1/X1/X1/X1/X2/vin1 0.00232f
C40 d0 X2/X1/X1/X2/vrefh 0.00385f
C41 d2 X1/X2/vrefh -0.157f
C42 X1/X2/X2/vrefh X3/m1_994_178# 4.63e-19
C43 d0 X1/X2/X2/X2/vrefh 0.00385f
C44 X1/X2/X2/X1/X2/X2/vrefh X2/X1/X1/X2/X1/X2/vrefh 0.117f
C45 X1/X2/X2/X2/X1/X2/X1/vin2 X2/X1/X1/X1/X2/X2/vrefh 0.0128f
C46 d2 X2/X1/X1/X1/X1/X1/X3/vin1 0.00301f
C47 X1/X2/X3/vin2 X3/vin1 0.00523f
C48 X2/X3/m1_688_n494# d6 0.0249f
C49 X1/X2/X2/X2/vrefh X2/X1/X1/X2/vrefh 0.117f
C50 X1/X2/X2/X1/X1/X1/X1/vin2 X2/X1/X2/vrefh 0.0128f
C51 d4 d0 1.8e-19
C52 d3 X2/X1/X1/X1/X1/X1/X1/m1_688_n494# 1.28e-19
C53 X1/X2/X2/X2/X2/X1/X1/vin2 X2/X1/X1/X1/X2/vrefh 0.0128f
C54 X2/X3/vin2 X3/vin2 0.142f
C55 d0 d5 -0.525f
C56 d4 X1/X2/X2/X2/X2/X2/X3/vin2 1.57e-19
C57 d1 d5 4.52f
C58 X1/X3/m1_994_178# d6 0.00555f
C59 d1 X1/X2/X2/X1/X1/X1/X1/m1_688_n494# 1.39e-20
C60 d1 X2/X1/X1/X2/X2/X2/X2/m1_994_178# 2.78e-20
C61 X1/X2/X2/X1/X1/X2/vrefh X2/X1/X1/X2/X2/X2/vrefh 0.117f
C62 X1/X2/X2/vrefh d7 3.76e-19
C63 d2 X2/X1/X1/X1/X1/X1/X1/vin1 0.00798f
C64 X3/vin2 d6 3.1f
C65 d4 X2/X1/X1/X1/X1/X1/X1/m1_994_178# 1.8e-19
C66 X1/X2/X3/m1_994_178# d6 0.00105f
C67 d1 X1/X2/X3/vin2 -0.00873f
C68 d6 X3/m1_688_n494# 0.00114f
C69 X1/X2/X2/X1/X2/X2/vrefh X2/X1/X1/X2/X1/X2/X1/vin1 0.00437f
C70 d0 X2/X1/X1/X1/X2/X2/vrefh 0.00385f
C71 X1/X3/vin1 X1/X3/m1_994_178# -0.00136f
C72 X2/X1/X3/vin2 d6 0.013f
C73 X1/X2/X2/X2/X1/X2/X1/vin2 X2/X1/X1/X1/X2/X1/X2/vin1 0.00232f
C74 X1/X3/m1_688_n494# d6 0.026f
C75 X1/X2/X2/X1/X2/X2/X2/vin1 X2/X1/X1/X2/X1/X1/X1/vin2 0.00232f
C76 d0 X2/X1/X1/X2/X1/X2/vrefh 0.00385f
C77 X2/X1/X3/m1_688_n494# d6 0.00114f
C78 X1/X2/X2/X1/X1/X2/X1/vin2 X2/X1/X1/X2/X2/X2/vrefh 0.0128f
C79 X1/X2/X2/X1/X2/X2/X1/vin2 X2/X1/X1/X2/X1/X2/vrefh 0.0128f
C80 d0 X2/X1/X1/X1/X2/vrefh 0.00385f
C81 X1/X2/X3/vin2 d5 0.0348f
C82 d0 X2/X1/X1/X2/X2/X2/vrefh 0.00385f
C83 X2/X3/vin1 X2/X3/vin2 -1.23e-20
C84 d2 X2/X1/X1/X1/X1/X1/X1/vin2 1.68e-19
C85 X1/X3/vin1 X1/X3/m1_688_n494# -0.0135f
C86 d3 X2/X1/X1/X1/X1/X1/X1/vin1 0.00492f
C87 X2/X3/m1_994_178# X2/X3/m1_688_n494# 2.84e-32
C88 d0 X1/X2/X2/X1/X2/vrefh 0.00385f
C89 d2 X2/vrefh 0.0108f
C90 X1/X3/vin2 X1/X3/m1_688_n494# -0.0081f
C91 X1/X2/X3/m1_688_n494# X3/vin1 5.96e-19
C92 X1/X2/X2/X2/X1/X2/X1/vin1 X2/X1/X1/X1/X2/X2/vrefh 0.00437f
C93 X3/vin1 d6 2.49f
C94 X1/X2/X2/vrefh X2/X1/X2/vrefh 0.0959f
C95 X3/vin1 X3/m1_994_178# 0.0255f
C96 X2/X3/vin1 d6 0.013f
C97 X2/X1/X3/m1_994_178# X3/vin2 4.87e-19
C98 X1/X2/X2/X1/X1/X1/X1/vin2 X2/X1/X1/X2/X2/X2/X2/vin1 0.00232f
C99 X1/X2/X2/X1/X2/X1/X1/vin2 X2/X1/X1/X2/X1/X2/X2/vin1 0.00232f
C100 d1 X1/X2/X2/X1/X1/X1/X1/vin1 0.00124f
C101 d2 X1/X2/X2/X2/X2/X2/X2/m1_688_n494# 1.95e-19
C102 X1/X3/vin1 X3/vin1 0.0385f
C103 d0 X1/X2/X2/X2/X1/X2/vrefh 0.00385f
C104 X2/X3/m1_994_178# X3/vin2 0.021f
C105 X1/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X2/X1/X1/vin2 0.0128f
C106 X1/X2/X2/X2/X1/X2/vrefh X2/X1/X1/X1/X2/X2/X1/vin2 0.0128f
C107 X1/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X2/X1/X1/vin1 0.00437f
C108 X1/X3/vin2 X3/vin1 0.173f
C109 d3 X2/X1/X1/X1/X1/X1/X1/vin2 1.14e-19
C110 d2 X2/X2/vrefh -0.157f
C111 d0 X3/m1_994_178# 2.73e-19
C112 X3/vin1 d7 0.0158f
C113 d2 d0 3.9e-19
C114 d3 X2/vrefh 0.00665f
C115 X1/X2/X2/X1/X2/X1/X2/vin1 X2/X1/X1/X2/X1/X2/X1/vin2 0.00232f
C116 d4 X1/X2/X2/X2/X2/X2/X2/m1_994_178# 1.8e-19
C117 d1 X3/m1_994_178# 4.67e-19
C118 X2/X1/X2/vrefh X3/vin2 3.04e-19
C119 d2 d1 1.48e-20
C120 X1/X2/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X1/X2/vrefh 0.117f
C121 d2 X1/X2/X2/X2/X2/X2/X3/vin2 0.00369f
C122 X2/X3/m1_688_n494# X3/vin2 0.0725f
C123 d4 d2 -0.0245f
C124 X1/X2/X3/m1_688_n494# d5 0.00103f
C125 d3 X1/X2/X2/X2/X2/X2/X2/m1_688_n494# 1.28e-19
C126 d5 d6 0.0012f
C127 d0 X1/X2/X2/X2/X2/vrefh 0.00385f
C128 d5 X3/m1_994_178# 9.9e-19
C129 d2 X2/X1/X1/X1/X1/X1/X1/m1_994_178# 3.9e-19
C130 d0 d7 1.37e-19
C131 X1/X2/X2/X1/X1/X2/X1/vin1 X2/X1/X1/X2/X2/X2/vrefh 0.00437f
C132 d1 d7 2.34e-19
C133 X1/X2/X2/X1/X2/X2/X1/vin1 X2/X1/X1/X2/X1/X2/vrefh 0.00437f
C134 X2/X3/vin1 X2/X3/m1_994_178# -0.00136f
C135 X1/X2/X2/X2/X1/X2/vrefh X2/X1/X1/X1/X2/X2/vrefh 0.117f
C136 X1/X2/X3/vin2 d6 0.013f
C137 d2 X2/X1/X1/X1/X1/X1/X3/m1_994_178# 2.97e-20
C138 d0 d3 2.56e-19
C139 X1/X2/X2/X1/X1/X2/vrefh X2/X1/X1/X2/X2/X2/X1/vin2 0.0128f
C140 d2 X2/X2/X1/X1/X1/X1/X1/vin1 -0.0257f
C141 X1/X2/X2/vrefh X3/vin1 0.0274f
C142 X1/X2/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X1/X2/X1/vin2 0.0128f
C143 X1/X3/m1_994_178# X1/X3/m1_688_n494# 5.68e-32
C144 d1 X2/X1/X3/m1_994_178# 4.67e-19
C145 X1/X3/vin2 d5 0.00217f
C146 d3 X1/X2/X2/X2/X2/X2/X3/vin2 0.0028f
C147 X2/X1/X3/vin2 X3/vin2 0.00486f
C148 X1/X2/X2/X1/X2/X1/X1/vin1 X2/X1/X1/X2/X2/vrefh 0.00437f
C149 d5 d7 4.95e-19
C150 d4 d3 5f
C151 X1/X2/X2/X2/X1/X1/X2/vin1 X2/X1/X1/X1/X2/X2/X1/vin2 0.00232f
C152 X2/X1/X3/m1_688_n494# X3/vin2 5.64e-19
C153 X2/X3/vin1 X2/X3/m1_688_n494# -0.0135f
C154 X1/X2/X2/X2/X2/X2/X1/vin2 X2/X1/X1/X1/X1/X2/vrefh 0.0128f
C155 d3 X2/X1/X1/X1/X1/X1/X1/m1_994_178# 2.56e-19
C156 X2/vrefh X2/X1/X1/X1/X1/X1/X1/vin1 0.0048f
C157 d4 X2/X1/X1/X1/X1/X1/X1/m1_688_n494# 8.99e-20
C158 X1/X2/X2/X2/X1/X1/X1/vin1 X2/X1/X1/X2/vrefh 0.00437f
C159 X1/X3/m1_994_178# X3/vin1 0.0205f
C160 d0 X1/X2/X2/vrefh 0.0571f
C161 d0 X2/X1/X2/vrefh 0.0562f
C162 X1/X2/X2/X2/X1/X2/vrefh X2/X1/X1/X1/X2/X2/X1/vin1 0.00437f
C163 d1 X1/X2/X2/X1/X1/X1/X1/m1_994_178# 2.78e-20
C164 d1 X2/X1/X2/vrefh 0.00168f
C165 X1/X2/X3/m1_994_178# X3/vin1 5.17e-19
C166 X2/X3/vin1 X3/vin2 0.0407f
C167 d0 X2/X1/X1/X2/X2/vrefh 0.00385f
C168 X3/vin1 X3/m1_688_n494# 0.035f
C169 d0 X1/X2/X2/X2/X2/X2/vrefh 0.00385f
C170 X1/X2/X2/X1/X2/X1/X1/vin2 X2/X1/X1/X2/X2/vrefh 0.0128f
C171 X1/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X2/vrefh 0.117f
C172 X2/X3/vin2 d6 0.00829f
C173 X1/X3/m1_688_n494# X3/vin1 0.0725f
C174 X2/vrefh X2/X1/X1/X1/X1/X1/X1/vin2 0.0128f
C175 d1 X2/X1/X1/X2/X2/X2/X2/m1_688_n494# 1.39e-20
C176 X1/X2/X2/X2/X1/X1/X1/vin2 X2/X1/X1/X2/vrefh 0.0128f
C177 d2 X1/X2/X2/X2/X2/X2/X2/m1_994_178# 3.9e-19
C178 d0 X2/X1/X1/X1/X1/X2/vrefh 0.00385f
C179 X1/X2/X3/m1_688_n494# d6 0.00114f
C180 d0 X3/vin2 1.31e-19
C181 X3/m1_994_178# d6 0.00105f
C182 d1 X3/vin2 3.83e-19
C183 X1/X2/X2/X1/X2/vrefh X2/X1/X1/X2/X2/X1/X1/vin1 0.00437f
C184 d0 X3/m1_688_n494# 1.37e-19
C185 d2 X2/X1/X1/X1/X1/X1/X3/m1_688_n494# 1.48e-20
C186 d1 X3/m1_688_n494# 2.34e-19
C187 X1/X2/X2/X1/X2/X2/X1/vin2 X2/X1/X1/X2/X1/X1/X2/vin1 0.00232f
C188 d4 X2/X1/X1/X1/X1/X1/X1/vin1 0.00332f
C189 X2/X1/X3/vin2 d0 -0.00274f
C190 X1/X2/X2/X1/X1/X2/vrefh X2/X1/X1/X2/X2/X2/X1/vin1 0.00437f
C191 X2/X1/X3/vin2 d1 0.0344f
C192 X1/X3/vin1 d6 0.00739f
C193 X1/X2/X2/X2/vrefh X2/X1/X1/X2/X1/X1/X1/vin1 0.00437f
C194 X1/X2/X2/X2/X2/X2/vrefh X2/X1/X1/X1/X1/X2/X1/vin1 0.00437f
C195 d0 X1/X2/X2/X1/X2/X2/vrefh 0.00385f
C196 X2/X1/X3/m1_688_n494# d1 5.18e-19
C197 X1/X3/vin2 d6 0.0889f
C198 d5 X3/vin2 0.00102f
C199 X1/X2/X3/m1_994_178# d5 9.9e-19
C200 d3 X1/X2/X2/X2/X2/X2/X2/m1_994_178# 2.56e-19
C201 d5 X3/m1_688_n494# 4.95e-19
C202 d6.t2 vss 0.0335f
C203 d6.t3 vss 0.0205f
C204 d6.n0 vss 0.257f
C205 d6.t0 vss 0.0335f
C206 d6.t1 vss 0.0205f
C207 d6.n1 vss 0.257f
C208 d5.t2 vss 0.083f
C209 d5.t3 vss 0.0509f
C210 d5.n0 vss 0.638f
C211 d5.t6 vss 0.083f
C212 d5.t7 vss 0.0509f
C213 d5.n1 vss 0.638f
C214 d5.t4 vss 0.083f
C215 d5.t5 vss 0.0509f
C216 d5.n2 vss 0.638f
C217 d5.n3 vss 6.2f
C218 d5.t0 vss 0.083f
C219 d5.t1 vss 0.0509f
C220 d5.n4 vss 0.638f
C221 d5.n5 vss 6.2f
C222 d4.t3 vss 0.0229f
C223 d4.t2 vss 0.0372f
C224 d4.t15 vss 0.0229f
C225 d4.n0 vss 0.135f
C226 d4.t14 vss 0.0372f
C227 d4.n1 vss 0.329f
C228 d4.t12 vss 0.0373f
C229 d4.t13 vss 0.0229f
C230 d4.n2 vss 0.507f
C231 d4.n3 vss 3.23f
C232 d4.t11 vss 0.0229f
C233 d4.n4 vss 0.135f
C234 d4.t10 vss 0.0372f
C235 d4.n5 vss 0.368f
C236 d4.t8 vss 0.0373f
C237 d4.t9 vss 0.0229f
C238 d4.n6 vss 0.468f
C239 d4.n7 vss 1.91f
C240 d4.n8 vss 5.84f
C241 d4.t7 vss 0.0229f
C242 d4.n9 vss 0.135f
C243 d4.t6 vss 0.0372f
C244 d4.n10 vss 0.329f
C245 d4.t4 vss 0.0373f
C246 d4.t5 vss 0.0229f
C247 d4.n11 vss 0.507f
C248 d4.n12 vss 1.91f
C249 d4.n13 vss 5.84f
C250 d4.t0 vss 0.0373f
C251 d4.t1 vss 0.0229f
C252 d4.n14 vss 0.468f
C253 d4.n15 vss 3.23f
C254 d4.n16 vss 0.368f
C255 d4.n17 vss 0.135f
C256 d3.t4 vss 0.0303f
C257 d3.t5 vss 0.0186f
C258 d3.t24 vss 0.0304f
C259 d3.t25 vss 0.0187f
C260 d3.n0 vss 0.417f
C261 d3.t26 vss 0.0304f
C262 d3.t27 vss 0.0187f
C263 d3.n1 vss 0.407f
C264 d3.n2 vss 0.539f
C265 d3.n3 vss 0.562f
C266 d3.n4 vss 0.556f
C267 d3.n5 vss 0.565f
C268 d3.n6 vss 0.375f
C269 d3.n7 vss 0.588f
C270 d3.n8 vss 0.581f
C271 d3.n9 vss 0.591f
C272 d3.t29 vss 0.0187f
C273 d3.t28 vss 0.0304f
C274 d3.n10 vss 0.411f
C275 d3.n11 vss 0.5f
C276 d3.n12 vss 0.562f
C277 d3.n13 vss 0.556f
C278 d3.n14 vss 0.565f
C279 d3.t31 vss 0.0187f
C280 d3.t30 vss 0.0304f
C281 d3.n15 vss 0.404f
C282 d3.n16 vss 0.558f
C283 d3.n17 vss 0.395f
C284 d3.n18 vss 0.347f
C285 d3.n19 vss 1.75f
C286 d3.t23 vss 0.0187f
C287 d3.t22 vss 0.0304f
C288 d3.n20 vss 0.377f
C289 d3.t21 vss 0.0187f
C290 d3.t20 vss 0.0304f
C291 d3.n21 vss 0.411f
C292 d3.n22 vss 0.5f
C293 d3.n23 vss 0.562f
C294 d3.n24 vss 0.556f
C295 d3.n25 vss 0.565f
C296 d3.n26 vss 0.375f
C297 d3.n27 vss 0.588f
C298 d3.n28 vss 0.581f
C299 d3.n29 vss 0.591f
C300 d3.t18 vss 0.0304f
C301 d3.t19 vss 0.0187f
C302 d3.n30 vss 0.407f
C303 d3.n31 vss 0.539f
C304 d3.n32 vss 0.562f
C305 d3.n33 vss 0.556f
C306 d3.n34 vss 0.565f
C307 d3.t16 vss 0.0304f
C308 d3.t17 vss 0.0188f
C309 d3.n35 vss 0.424f
C310 d3.n36 vss 0.519f
C311 d3.n37 vss 0.395f
C312 d3.n38 vss 0.368f
C313 d3.n39 vss 0.789f
C314 d3.n40 vss 3.59f
C315 d3.t8 vss 0.0304f
C316 d3.t9 vss 0.0188f
C317 d3.n41 vss 0.424f
C318 d3.t10 vss 0.0306f
C319 d3.t11 vss 0.0187f
C320 d3.n42 vss 0.414f
C321 d3.n43 vss 0.539f
C322 d3.n44 vss 0.562f
C323 d3.n45 vss 0.556f
C324 d3.n46 vss 0.565f
C325 d3.n47 vss 0.375f
C326 d3.n48 vss 0.588f
C327 d3.n49 vss 0.581f
C328 d3.n50 vss 0.591f
C329 d3.t13 vss 0.0187f
C330 d3.t12 vss 0.0304f
C331 d3.n51 vss 0.411f
C332 d3.n52 vss 0.5f
C333 d3.n53 vss 0.562f
C334 d3.n54 vss 0.556f
C335 d3.n55 vss 0.565f
C336 d3.t15 vss 0.0187f
C337 d3.t14 vss 0.0306f
C338 d3.n56 vss 0.411f
C339 d3.n57 vss 0.558f
C340 d3.n58 vss 0.395f
C341 d3.n59 vss 0.347f
C342 d3.n60 vss 0.747f
C343 d3.n61 vss 3.59f
C344 d3.t7 vss 0.0187f
C345 d3.t6 vss 0.0306f
C346 d3.n62 vss 0.384f
C347 d3.n63 vss 1.79f
C348 d3.t0 vss 0.0304f
C349 d3.t1 vss 0.0188f
C350 d3.n64 vss 0.424f
C351 d3.n65 vss 0.519f
C352 d3.n66 vss 0.395f
C353 d3.n67 vss 0.368f
C354 d3.n68 vss 0.565f
C355 d3.n69 vss 0.556f
C356 d3.n70 vss 0.562f
C357 d3.n71 vss 0.591f
C358 d3.n72 vss 0.581f
C359 d3.n73 vss 0.588f
C360 d3.t3 vss 0.0186f
C361 d3.t2 vss 0.0304f
C362 d3.n74 vss 0.418f
C363 d3.n75 vss 0.565f
C364 d3.n76 vss 0.556f
C365 d3.n77 vss 0.562f
C366 d3.n78 vss 0.539f
C367 d3.n79 vss 0.375f
C368 d3.n80 vss 0.5f
C369 d3.n81 vss 0.415f
C370 d2.t2 vss 0.0587f
C371 d2.t3 vss 0.036f
C372 d2.t9 vss 0.036f
C373 d2.t8 vss 0.0587f
C374 d2.n0 vss 0.486f
C375 d2.n1 vss 2.12f
C376 d2.t6 vss 0.0587f
C377 d2.t7 vss 0.036f
C378 d2.n2 vss 0.497f
C379 d2.n3 vss 2.13f
C380 d2.t4 vss 0.0587f
C381 d2.t5 vss 0.036f
C382 d2.n4 vss 0.575f
C383 d2.n5 vss 2.46f
C384 d2.t13 vss 0.036f
C385 d2.t12 vss 0.0587f
C386 d2.n6 vss 0.564f
C387 d2.t11 vss 0.036f
C388 d2.t10 vss 0.0587f
C389 d2.n7 vss 0.563f
C390 d2.n8 vss 2.45f
C391 d2.n9 vss 2.46f
C392 d2.t15 vss 0.036f
C393 d2.t14 vss 0.0587f
C394 d2.n10 vss 0.486f
C395 d2.n11 vss 1.75f
C396 d2.t61 vss 0.036f
C397 d2.t60 vss 0.0587f
C398 d2.n12 vss 0.564f
C399 d2.t59 vss 0.036f
C400 d2.t58 vss 0.0587f
C401 d2.n13 vss 0.563f
C402 d2.t57 vss 0.036f
C403 d2.t56 vss 0.0587f
C404 d2.n14 vss 0.486f
C405 d2.n15 vss 2.12f
C406 d2.n16 vss 2.45f
C407 d2.n17 vss 2.46f
C408 d2.t63 vss 0.036f
C409 d2.t62 vss 0.0587f
C410 d2.n18 vss 0.486f
C411 d2.n19 vss 1.79f
C412 d2.t48 vss 0.0587f
C413 d2.t49 vss 0.036f
C414 d2.n20 vss 0.497f
C415 d2.t54 vss 0.0587f
C416 d2.t55 vss 0.036f
C417 d2.n21 vss 0.497f
C418 d2.n22 vss 2.13f
C419 d2.t52 vss 0.0587f
C420 d2.t53 vss 0.036f
C421 d2.n23 vss 0.575f
C422 d2.n24 vss 2.46f
C423 d2.t50 vss 0.0587f
C424 d2.t51 vss 0.036f
C425 d2.n25 vss 0.574f
C426 d2.n26 vss 2.46f
C427 d2.n27 vss 1.68f
C428 d2.n28 vss 3.67f
C429 d2.t45 vss 0.036f
C430 d2.t44 vss 0.0587f
C431 d2.n29 vss 0.564f
C432 d2.t43 vss 0.036f
C433 d2.t42 vss 0.0587f
C434 d2.n30 vss 0.563f
C435 d2.t41 vss 0.036f
C436 d2.t40 vss 0.0587f
C437 d2.n31 vss 0.486f
C438 d2.n32 vss 2.12f
C439 d2.n33 vss 2.45f
C440 d2.n34 vss 2.46f
C441 d2.t47 vss 0.036f
C442 d2.t46 vss 0.0587f
C443 d2.n35 vss 0.486f
C444 d2.n36 vss 1.75f
C445 d2.t32 vss 0.0587f
C446 d2.t33 vss 0.036f
C447 d2.n37 vss 0.497f
C448 d2.t38 vss 0.0587f
C449 d2.t39 vss 0.036f
C450 d2.n38 vss 0.497f
C451 d2.n39 vss 2.13f
C452 d2.t36 vss 0.0587f
C453 d2.t37 vss 0.036f
C454 d2.n40 vss 0.575f
C455 d2.n41 vss 2.46f
C456 d2.t34 vss 0.0587f
C457 d2.t35 vss 0.036f
C458 d2.n42 vss 0.574f
C459 d2.n43 vss 2.46f
C460 d2.n44 vss 1.73f
C461 d2.n45 vss 1.43f
C462 d2.n46 vss 5.83f
C463 d2.t29 vss 0.036f
C464 d2.t28 vss 0.0587f
C465 d2.n47 vss 0.564f
C466 d2.t27 vss 0.036f
C467 d2.t26 vss 0.0587f
C468 d2.n48 vss 0.563f
C469 d2.t25 vss 0.036f
C470 d2.t24 vss 0.0587f
C471 d2.n49 vss 0.486f
C472 d2.n50 vss 2.12f
C473 d2.n51 vss 2.45f
C474 d2.n52 vss 2.46f
C475 d2.t31 vss 0.036f
C476 d2.t30 vss 0.0587f
C477 d2.n53 vss 0.486f
C478 d2.n54 vss 1.79f
C479 d2.t16 vss 0.0587f
C480 d2.t17 vss 0.036f
C481 d2.n55 vss 0.497f
C482 d2.t22 vss 0.0587f
C483 d2.t23 vss 0.036f
C484 d2.n56 vss 0.497f
C485 d2.n57 vss 2.13f
C486 d2.t20 vss 0.0587f
C487 d2.t21 vss 0.036f
C488 d2.n58 vss 0.575f
C489 d2.n59 vss 2.46f
C490 d2.t18 vss 0.0587f
C491 d2.t19 vss 0.036f
C492 d2.n60 vss 0.574f
C493 d2.n61 vss 2.46f
C494 d2.n62 vss 1.68f
C495 d2.n63 vss 1.43f
C496 d2.n64 vss 5.83f
C497 d2.n65 vss 3.67f
C498 d2.t0 vss 0.0587f
C499 d2.t1 vss 0.036f
C500 d2.n66 vss 0.497f
C501 d2.n67 vss 1.73f
C502 d2.n68 vss 2.46f
C503 d2.n69 vss 0.574f
C504 d1.t2 vss 0.056f
C505 d1.t3 vss 0.0343f
C506 d1.n0 vss 0.425f
C507 d1.t0 vss 0.056f
C508 d1.t1 vss 0.0343f
C509 d1.n1 vss 0.425f
C510 d1.n2 vss 0.535f
C511 d1.t4 vss 0.056f
C512 d1.t5 vss 0.0343f
C513 d1.n3 vss 0.425f
C514 d1.n4 vss 0.0262f
C515 d1.t6 vss 0.056f
C516 d1.t7 vss 0.0343f
C517 d1.n5 vss 0.425f
C518 d1.n6 vss 0.0262f
C519 d1.t8 vss 0.056f
C520 d1.t9 vss 0.0343f
C521 d1.n7 vss 0.425f
C522 d1.n8 vss 0.0262f
C523 d1.t10 vss 0.056f
C524 d1.t11 vss 0.0343f
C525 d1.n9 vss 0.425f
C526 d1.n10 vss 0.0262f
C527 d1.t12 vss 0.056f
C528 d1.t13 vss 0.0343f
C529 d1.n11 vss 0.425f
C530 d1.n12 vss 0.0262f
C531 d1.t14 vss 0.056f
C532 d1.t15 vss 0.0343f
C533 d1.n13 vss 0.425f
C534 d1.n14 vss 0.0262f
C535 d1.t31 vss 0.0343f
C536 d1.t30 vss 0.056f
C537 d1.n15 vss 0.425f
C538 d1.t29 vss 0.0343f
C539 d1.t28 vss 0.056f
C540 d1.n16 vss 0.42f
C541 d1.n17 vss 1.01f
C542 d1.t27 vss 0.0343f
C543 d1.t26 vss 0.056f
C544 d1.n18 vss 0.425f
C545 d1.n19 vss 1.07f
C546 d1.t25 vss 0.0343f
C547 d1.t24 vss 0.056f
C548 d1.n20 vss 0.42f
C549 d1.n21 vss 0.997f
C550 d1.t23 vss 0.0343f
C551 d1.t22 vss 0.056f
C552 d1.n22 vss 0.425f
C553 d1.n23 vss 0.997f
C554 d1.t21 vss 0.0343f
C555 d1.t20 vss 0.056f
C556 d1.n24 vss 0.42f
C557 d1.n25 vss 1.01f
C558 d1.t19 vss 0.0343f
C559 d1.t18 vss 0.056f
C560 d1.n26 vss 0.425f
C561 d1.n27 vss 1.07f
C562 d1.t17 vss 0.0343f
C563 d1.t16 vss 0.056f
C564 d1.n28 vss 0.42f
C565 d1.n29 vss 0.651f
C566 d1.t127 vss 0.0343f
C567 d1.t126 vss 0.056f
C568 d1.n30 vss 0.425f
C569 d1.t125 vss 0.0343f
C570 d1.t124 vss 0.056f
C571 d1.n31 vss 0.42f
C572 d1.n32 vss 1.01f
C573 d1.t123 vss 0.0343f
C574 d1.t122 vss 0.056f
C575 d1.n33 vss 0.425f
C576 d1.n34 vss 1.07f
C577 d1.t121 vss 0.0343f
C578 d1.t120 vss 0.056f
C579 d1.n35 vss 0.42f
C580 d1.n36 vss 0.997f
C581 d1.t119 vss 0.0343f
C582 d1.t118 vss 0.056f
C583 d1.n37 vss 0.425f
C584 d1.n38 vss 0.997f
C585 d1.t117 vss 0.0343f
C586 d1.t116 vss 0.056f
C587 d1.n39 vss 0.42f
C588 d1.n40 vss 1.01f
C589 d1.t115 vss 0.0343f
C590 d1.t114 vss 0.056f
C591 d1.n41 vss 0.425f
C592 d1.n42 vss 1.07f
C593 d1.t113 vss 0.0343f
C594 d1.t112 vss 0.056f
C595 d1.n43 vss 0.42f
C596 d1.n44 vss 0.651f
C597 d1.t96 vss 0.056f
C598 d1.t97 vss 0.0343f
C599 d1.n45 vss 0.425f
C600 d1.n46 vss 0.535f
C601 d1.t98 vss 0.056f
C602 d1.t99 vss 0.0343f
C603 d1.n47 vss 0.425f
C604 d1.n48 vss 0.0262f
C605 d1.n49 vss 1.07f
C606 d1.t100 vss 0.056f
C607 d1.t101 vss 0.0343f
C608 d1.n50 vss 0.425f
C609 d1.n51 vss 0.0262f
C610 d1.n52 vss 1.01f
C611 d1.t102 vss 0.056f
C612 d1.t103 vss 0.0343f
C613 d1.n53 vss 0.425f
C614 d1.n54 vss 0.0262f
C615 d1.n55 vss 0.997f
C616 d1.t104 vss 0.056f
C617 d1.t105 vss 0.0343f
C618 d1.n56 vss 0.425f
C619 d1.n57 vss 0.0262f
C620 d1.n58 vss 0.997f
C621 d1.t106 vss 0.056f
C622 d1.t107 vss 0.0343f
C623 d1.n59 vss 0.425f
C624 d1.n60 vss 0.0262f
C625 d1.n61 vss 1.07f
C626 d1.t108 vss 0.056f
C627 d1.t109 vss 0.0343f
C628 d1.n62 vss 0.425f
C629 d1.n63 vss 0.0262f
C630 d1.n64 vss 1.01f
C631 d1.t110 vss 0.056f
C632 d1.t111 vss 0.0343f
C633 d1.n65 vss 0.425f
C634 d1.n66 vss 0.0262f
C635 d1.n67 vss 1.42f
C636 d1.n68 vss 3.26f
C637 d1.t95 vss 0.0343f
C638 d1.t94 vss 0.056f
C639 d1.n69 vss 0.425f
C640 d1.t93 vss 0.0343f
C641 d1.t92 vss 0.056f
C642 d1.n70 vss 0.42f
C643 d1.n71 vss 1.01f
C644 d1.t91 vss 0.0343f
C645 d1.t90 vss 0.056f
C646 d1.n72 vss 0.425f
C647 d1.n73 vss 1.07f
C648 d1.t89 vss 0.0343f
C649 d1.t88 vss 0.056f
C650 d1.n74 vss 0.42f
C651 d1.n75 vss 0.997f
C652 d1.t87 vss 0.0343f
C653 d1.t86 vss 0.056f
C654 d1.n76 vss 0.425f
C655 d1.n77 vss 0.997f
C656 d1.t85 vss 0.0343f
C657 d1.t84 vss 0.056f
C658 d1.n78 vss 0.42f
C659 d1.n79 vss 1.01f
C660 d1.t83 vss 0.0343f
C661 d1.t82 vss 0.056f
C662 d1.n80 vss 0.425f
C663 d1.n81 vss 1.07f
C664 d1.t81 vss 0.0343f
C665 d1.t80 vss 0.056f
C666 d1.n82 vss 0.42f
C667 d1.n83 vss 0.651f
C668 d1.t64 vss 0.056f
C669 d1.t65 vss 0.0343f
C670 d1.n84 vss 0.425f
C671 d1.n85 vss 0.535f
C672 d1.t66 vss 0.056f
C673 d1.t67 vss 0.0343f
C674 d1.n86 vss 0.425f
C675 d1.n87 vss 0.0262f
C676 d1.n88 vss 1.07f
C677 d1.t68 vss 0.056f
C678 d1.t69 vss 0.0343f
C679 d1.n89 vss 0.425f
C680 d1.n90 vss 0.0262f
C681 d1.n91 vss 1.01f
C682 d1.t70 vss 0.056f
C683 d1.t71 vss 0.0343f
C684 d1.n92 vss 0.425f
C685 d1.n93 vss 0.0262f
C686 d1.n94 vss 0.997f
C687 d1.t72 vss 0.056f
C688 d1.t73 vss 0.0343f
C689 d1.n95 vss 0.425f
C690 d1.n96 vss 0.0262f
C691 d1.n97 vss 0.997f
C692 d1.t74 vss 0.056f
C693 d1.t75 vss 0.0343f
C694 d1.n98 vss 0.425f
C695 d1.n99 vss 0.0262f
C696 d1.n100 vss 1.07f
C697 d1.t76 vss 0.056f
C698 d1.t77 vss 0.0343f
C699 d1.n101 vss 0.425f
C700 d1.n102 vss 0.0262f
C701 d1.n103 vss 1.01f
C702 d1.t78 vss 0.056f
C703 d1.t79 vss 0.0343f
C704 d1.n104 vss 0.425f
C705 d1.n105 vss 0.0262f
C706 d1.n106 vss 1.42f
C707 d1.n107 vss 1.32f
C708 d1.n108 vss 4.36f
C709 d1.t63 vss 0.0343f
C710 d1.t62 vss 0.056f
C711 d1.n109 vss 0.425f
C712 d1.t61 vss 0.0343f
C713 d1.t60 vss 0.056f
C714 d1.n110 vss 0.42f
C715 d1.n111 vss 1.01f
C716 d1.t59 vss 0.0343f
C717 d1.t58 vss 0.056f
C718 d1.n112 vss 0.425f
C719 d1.n113 vss 1.07f
C720 d1.t57 vss 0.0343f
C721 d1.t56 vss 0.056f
C722 d1.n114 vss 0.42f
C723 d1.n115 vss 0.997f
C724 d1.t55 vss 0.0343f
C725 d1.t54 vss 0.056f
C726 d1.n116 vss 0.425f
C727 d1.n117 vss 0.997f
C728 d1.t53 vss 0.0343f
C729 d1.t52 vss 0.056f
C730 d1.n118 vss 0.42f
C731 d1.n119 vss 1.01f
C732 d1.t51 vss 0.0343f
C733 d1.t50 vss 0.056f
C734 d1.n120 vss 0.425f
C735 d1.n121 vss 1.07f
C736 d1.t49 vss 0.0343f
C737 d1.t48 vss 0.056f
C738 d1.n122 vss 0.42f
C739 d1.n123 vss 0.651f
C740 d1.t32 vss 0.056f
C741 d1.t33 vss 0.0343f
C742 d1.n124 vss 0.425f
C743 d1.n125 vss 0.535f
C744 d1.t34 vss 0.056f
C745 d1.t35 vss 0.0343f
C746 d1.n126 vss 0.425f
C747 d1.n127 vss 0.0262f
C748 d1.n128 vss 1.07f
C749 d1.t36 vss 0.056f
C750 d1.t37 vss 0.0343f
C751 d1.n129 vss 0.425f
C752 d1.n130 vss 0.0262f
C753 d1.n131 vss 1.01f
C754 d1.t38 vss 0.056f
C755 d1.t39 vss 0.0343f
C756 d1.n132 vss 0.425f
C757 d1.n133 vss 0.0262f
C758 d1.n134 vss 0.997f
C759 d1.t40 vss 0.056f
C760 d1.t41 vss 0.0343f
C761 d1.n135 vss 0.425f
C762 d1.n136 vss 0.0262f
C763 d1.n137 vss 0.997f
C764 d1.t42 vss 0.056f
C765 d1.t43 vss 0.0343f
C766 d1.n138 vss 0.425f
C767 d1.n139 vss 0.0262f
C768 d1.n140 vss 1.07f
C769 d1.t44 vss 0.056f
C770 d1.t45 vss 0.0343f
C771 d1.n141 vss 0.425f
C772 d1.n142 vss 0.0262f
C773 d1.n143 vss 1.01f
C774 d1.t46 vss 0.056f
C775 d1.t47 vss 0.0343f
C776 d1.n144 vss 0.425f
C777 d1.n145 vss 0.0262f
C778 d1.n146 vss 1.42f
C779 d1.n147 vss 1.32f
C780 d1.n148 vss 4.36f
C781 d1.n149 vss 3.26f
C782 d1.n150 vss 1.42f
C783 d1.n151 vss 1.01f
C784 d1.n152 vss 1.07f
C785 d1.n153 vss 0.997f
C786 d1.n154 vss 0.997f
C787 d1.n155 vss 1.01f
C788 d1.n156 vss 1.07f
C789 d1.n157 vss 0.0262f
C790 vdd.n0 vss 0.00324f
C791 vdd.n1 vss 0.0112f
C792 vdd.n2 vss 0.0128f
C793 vdd.n3 vss 0.00413f
C794 vdd.n4 vss 0.00413f
C795 vdd.n5 vss 0.0471f
C796 vdd.n6 vss 0.0471f
C797 vdd.n7 vss 0.00324f
C798 vdd.n8 vss 0.00413f
C799 vdd.n9 vss 0.00413f
C800 vdd.n10 vss 0.00679f
C801 vdd.n11 vss 0.00413f
C802 vdd.n12 vss 0.0471f
C803 vdd.n13 vss 0.00324f
C804 vdd.n15 vss 0.00925f
C805 vdd.n16 vss 0.0471f
C806 vdd.n17 vss 0.00425f
C807 vdd.n18 vss 0.0424f
C808 vdd.n19 vss 0.0132f
C809 vdd.n20 vss 0.00324f
C810 vdd.n21 vss 0.0128f
C811 vdd.n22 vss 0.02f
C812 vdd.n23 vss 0.00425f
C813 vdd.n24 vss 0.00413f
C814 vdd.n25 vss 0.00251f
C815 vdd.n26 vss 0.0471f
C816 vdd.n27 vss 0.00251f
C817 vdd.n28 vss 0.00517f
C818 vdd.n29 vss 0.00679f
C819 vdd.n30 vss 0.00324f
C820 vdd.n31 vss 0.00324f
C821 vdd.n32 vss 0.0132f
C822 vdd.n33 vss 0.0424f
C823 vdd.n34 vss 0.02f
C824 vdd.n35 vss 0.00425f
C825 vdd.n36 vss 0.0471f
C826 vdd.n38 vss 0.00425f
C827 vdd.n39 vss 0.00925f
C828 vdd.n40 vss 0.00679f
C829 vdd.n41 vss 0.00517f
C830 vdd.n42 vss 0.00251f
C831 vdd.n43 vss 0.0471f
C832 vdd.n44 vss 0.00251f
C833 vdd.n45 vss 0.0112f
C834 vdd.n46 vss 0.0128f
C835 vdd.n47 vss 0.146f
C836 vdd.n48 vss 0.00324f
C837 vdd.n49 vss 0.0112f
C838 vdd.n50 vss 0.0128f
C839 vdd.n51 vss 0.00413f
C840 vdd.n52 vss 0.00413f
C841 vdd.n53 vss 0.0471f
C842 vdd.n54 vss 0.0471f
C843 vdd.n55 vss 0.00324f
C844 vdd.n56 vss 0.00413f
C845 vdd.n57 vss 0.00413f
C846 vdd.n58 vss 0.00679f
C847 vdd.n59 vss 0.00413f
C848 vdd.n60 vss 0.0471f
C849 vdd.n61 vss 0.00324f
C850 vdd.n63 vss 0.00925f
C851 vdd.n64 vss 0.0471f
C852 vdd.n65 vss 0.00425f
C853 vdd.n66 vss 0.0424f
C854 vdd.n67 vss 0.0132f
C855 vdd.n68 vss 0.00324f
C856 vdd.n69 vss 0.0128f
C857 vdd.n70 vss 0.02f
C858 vdd.n71 vss 0.00425f
C859 vdd.n72 vss 0.00413f
C860 vdd.n73 vss 0.00251f
C861 vdd.n74 vss 0.0471f
C862 vdd.n75 vss 0.00251f
C863 vdd.n76 vss 0.00517f
C864 vdd.n77 vss 0.00679f
C865 vdd.n78 vss 0.00324f
C866 vdd.n79 vss 0.00324f
C867 vdd.n80 vss 0.0132f
C868 vdd.n81 vss 0.0424f
C869 vdd.n82 vss 0.02f
C870 vdd.n83 vss 0.00425f
C871 vdd.n84 vss 0.0471f
C872 vdd.n86 vss 0.00425f
C873 vdd.n87 vss 0.00925f
C874 vdd.n88 vss 0.00679f
C875 vdd.n89 vss 0.00517f
C876 vdd.n90 vss 0.00251f
C877 vdd.n91 vss 0.0471f
C878 vdd.n92 vss 0.00251f
C879 vdd.n93 vss 0.0112f
C880 vdd.n94 vss 0.0128f
C881 vdd.n95 vss 0.146f
C882 vdd.n96 vss 0.0596f
C883 vdd.n97 vss 0.00324f
C884 vdd.n98 vss 0.0112f
C885 vdd.n99 vss 0.0128f
C886 vdd.n100 vss 0.00413f
C887 vdd.n101 vss 0.00413f
C888 vdd.n102 vss 0.0471f
C889 vdd.n103 vss 0.0471f
C890 vdd.n104 vss 0.00324f
C891 vdd.n105 vss 0.00413f
C892 vdd.n106 vss 0.00413f
C893 vdd.n107 vss 0.00679f
C894 vdd.n108 vss 0.00413f
C895 vdd.n109 vss 0.0471f
C896 vdd.n110 vss 0.00324f
C897 vdd.n111 vss 0.0424f
C898 vdd.n112 vss 0.00324f
C899 vdd.n113 vss 0.0128f
C900 vdd.n114 vss 0.02f
C901 vdd.n115 vss 0.0132f
C902 vdd.n116 vss 0.00925f
C903 vdd.n117 vss 0.00425f
C904 vdd.n119 vss 0.0471f
C905 vdd.n120 vss 0.00425f
C906 vdd.n121 vss 0.00413f
C907 vdd.n122 vss 0.00251f
C908 vdd.n123 vss 0.0471f
C909 vdd.n124 vss 0.00251f
C910 vdd.n125 vss 0.00517f
C911 vdd.n126 vss 0.00679f
C912 vdd.n127 vss 0.00324f
C913 vdd.n128 vss 0.00324f
C914 vdd.n129 vss 0.0132f
C915 vdd.n130 vss 0.0424f
C916 vdd.n131 vss 0.02f
C917 vdd.n132 vss 0.00425f
C918 vdd.n134 vss 0.0471f
C919 vdd.n135 vss 0.00425f
C920 vdd.n136 vss 0.00925f
C921 vdd.n137 vss 0.00679f
C922 vdd.n138 vss 0.00517f
C923 vdd.n139 vss 0.00251f
C924 vdd.n140 vss 0.0471f
C925 vdd.n141 vss 0.00251f
C926 vdd.n142 vss 0.0112f
C927 vdd.n143 vss 0.0128f
C928 vdd.n144 vss 0.0666f
C929 vdd.n145 vss 0.00324f
C930 vdd.n146 vss 0.0112f
C931 vdd.n147 vss 0.0128f
C932 vdd.n148 vss 0.00413f
C933 vdd.n149 vss 0.00413f
C934 vdd.n150 vss 0.0471f
C935 vdd.n151 vss 0.0471f
C936 vdd.n152 vss 0.00324f
C937 vdd.n153 vss 0.00413f
C938 vdd.n154 vss 0.00413f
C939 vdd.n155 vss 0.00679f
C940 vdd.n156 vss 0.00413f
C941 vdd.n157 vss 0.0471f
C942 vdd.n158 vss 0.00324f
C943 vdd.n159 vss 0.0424f
C944 vdd.n160 vss 0.00324f
C945 vdd.n161 vss 0.0128f
C946 vdd.n162 vss 0.02f
C947 vdd.n163 vss 0.0132f
C948 vdd.n164 vss 0.00925f
C949 vdd.n165 vss 0.00425f
C950 vdd.n167 vss 0.0471f
C951 vdd.n168 vss 0.00425f
C952 vdd.n169 vss 0.00413f
C953 vdd.n170 vss 0.00251f
C954 vdd.n171 vss 0.0471f
C955 vdd.n172 vss 0.00251f
C956 vdd.n173 vss 0.00517f
C957 vdd.n174 vss 0.00679f
C958 vdd.n175 vss 0.00324f
C959 vdd.n176 vss 0.00324f
C960 vdd.n177 vss 0.0132f
C961 vdd.n178 vss 0.0424f
C962 vdd.n179 vss 0.02f
C963 vdd.n180 vss 0.00425f
C964 vdd.n182 vss 0.0471f
C965 vdd.n183 vss 0.00425f
C966 vdd.n184 vss 0.00925f
C967 vdd.n185 vss 0.00679f
C968 vdd.n186 vss 0.00517f
C969 vdd.n187 vss 0.00251f
C970 vdd.n188 vss 0.0471f
C971 vdd.n189 vss 0.00251f
C972 vdd.n190 vss 0.0112f
C973 vdd.n191 vss 0.0128f
C974 vdd.n192 vss 0.0617f
C975 vdd.n193 vss 0.00335f
C976 vdd.n194 vss 0.0855f
C977 vdd.n195 vss 0.0107f
C978 vdd.n196 vss 0.0128f
C979 vdd.n197 vss 0.0424f
C980 vdd.n198 vss 0.00413f
C981 vdd.n199 vss 0.0471f
C982 vdd.n200 vss 0.00413f
C983 vdd.n201 vss 0.00324f
C984 vdd.n202 vss 0.00324f
C985 vdd.n203 vss 0.00679f
C986 vdd.n204 vss 0.00413f
C987 vdd.n205 vss 0.0471f
C988 vdd.n206 vss 0.00413f
C989 vdd.n207 vss 0.0105f
C990 vdd.n208 vss 0.0471f
C991 vdd.n209 vss 0.00413f
C992 vdd.n210 vss 0.00324f
C993 vdd.n211 vss 0.00324f
C994 vdd.n212 vss 0.0132f
C995 vdd.n213 vss 0.0424f
C996 vdd.n214 vss 0.0128f
C997 vdd.n215 vss 0.02f
C998 vdd.n216 vss 0.00425f
C999 vdd.n218 vss 0.0471f
C1000 vdd.n219 vss 0.00425f
C1001 vdd.n220 vss 0.00925f
C1002 vdd.n221 vss 0.00679f
C1003 vdd.n222 vss 0.00517f
C1004 vdd.n223 vss 0.00251f
C1005 vdd.n224 vss 0.0471f
C1006 vdd.n225 vss 0.00251f
C1007 vdd.n226 vss 0.00413f
C1008 vdd.n227 vss 0.00324f
C1009 vdd.n228 vss 0.00324f
C1010 vdd.n229 vss 0.00805f
C1011 vdd.n230 vss 0.0112f
C1012 vdd.n231 vss 0.00251f
C1013 vdd.n232 vss 0.0471f
C1014 vdd.n233 vss 0.00251f
C1015 vdd.n234 vss 0.00517f
C1016 vdd.n235 vss 0.00679f
C1017 vdd.n236 vss 0.00925f
C1018 vdd.n237 vss 0.00425f
C1019 vdd.n239 vss 0.0471f
C1020 vdd.n240 vss 0.00425f
C1021 vdd.n241 vss 0.00991f
C1022 vdd.n242 vss 0.0126f
C1023 vdd.n243 vss 0.0516f
C1024 vdd.n244 vss 0.0011f
C1025 vdd.n245 vss 0.0271f
C1026 vdd.n246 vss 0.00324f
C1027 vdd.n247 vss 0.0112f
C1028 vdd.n248 vss 0.0128f
C1029 vdd.n249 vss 0.00413f
C1030 vdd.n250 vss 0.00413f
C1031 vdd.n251 vss 0.0471f
C1032 vdd.n252 vss 0.0471f
C1033 vdd.n253 vss 0.00324f
C1034 vdd.n254 vss 0.00413f
C1035 vdd.n255 vss 0.00413f
C1036 vdd.n256 vss 0.00679f
C1037 vdd.n257 vss 0.00413f
C1038 vdd.n258 vss 0.0471f
C1039 vdd.n259 vss 0.00324f
C1040 vdd.n260 vss 0.0424f
C1041 vdd.n261 vss 0.00324f
C1042 vdd.n262 vss 0.0128f
C1043 vdd.n263 vss 0.02f
C1044 vdd.n264 vss 0.0132f
C1045 vdd.n265 vss 0.00925f
C1046 vdd.n266 vss 0.00425f
C1047 vdd.n268 vss 0.0471f
C1048 vdd.n269 vss 0.00425f
C1049 vdd.n270 vss 0.00413f
C1050 vdd.n271 vss 0.00251f
C1051 vdd.n272 vss 0.0471f
C1052 vdd.n273 vss 0.00251f
C1053 vdd.n274 vss 0.00517f
C1054 vdd.n275 vss 0.00679f
C1055 vdd.n276 vss 0.00324f
C1056 vdd.n277 vss 0.00324f
C1057 vdd.n278 vss 0.0132f
C1058 vdd.n279 vss 0.0424f
C1059 vdd.n280 vss 0.02f
C1060 vdd.n281 vss 0.00425f
C1061 vdd.n283 vss 0.0471f
C1062 vdd.n284 vss 0.00425f
C1063 vdd.n285 vss 0.00925f
C1064 vdd.n286 vss 0.00679f
C1065 vdd.n287 vss 0.00517f
C1066 vdd.n288 vss 0.00251f
C1067 vdd.n289 vss 0.0471f
C1068 vdd.n290 vss 0.00251f
C1069 vdd.n291 vss 0.0112f
C1070 vdd.n292 vss 0.0128f
C1071 vdd.n293 vss 0.0666f
C1072 vdd.n294 vss 0.00324f
C1073 vdd.n295 vss 0.0112f
C1074 vdd.n296 vss 0.0128f
C1075 vdd.n297 vss 0.00413f
C1076 vdd.n298 vss 0.00413f
C1077 vdd.n299 vss 0.0471f
C1078 vdd.n300 vss 0.0471f
C1079 vdd.n301 vss 0.00324f
C1080 vdd.n302 vss 0.00413f
C1081 vdd.n303 vss 0.00413f
C1082 vdd.n304 vss 0.00679f
C1083 vdd.n305 vss 0.00413f
C1084 vdd.n306 vss 0.0471f
C1085 vdd.n307 vss 0.00324f
C1086 vdd.n308 vss 0.0424f
C1087 vdd.n309 vss 0.00324f
C1088 vdd.n310 vss 0.0128f
C1089 vdd.n311 vss 0.02f
C1090 vdd.n312 vss 0.0132f
C1091 vdd.n313 vss 0.00925f
C1092 vdd.n314 vss 0.00425f
C1093 vdd.n316 vss 0.0471f
C1094 vdd.n317 vss 0.00425f
C1095 vdd.n318 vss 0.00413f
C1096 vdd.n319 vss 0.00251f
C1097 vdd.n320 vss 0.0471f
C1098 vdd.n321 vss 0.00251f
C1099 vdd.n322 vss 0.00517f
C1100 vdd.n323 vss 0.00679f
C1101 vdd.n324 vss 0.00324f
C1102 vdd.n325 vss 0.00324f
C1103 vdd.n326 vss 0.0132f
C1104 vdd.n327 vss 0.0424f
C1105 vdd.n328 vss 0.02f
C1106 vdd.n329 vss 0.00425f
C1107 vdd.n331 vss 0.0471f
C1108 vdd.n332 vss 0.00425f
C1109 vdd.n333 vss 0.00925f
C1110 vdd.n334 vss 0.00679f
C1111 vdd.n335 vss 0.00517f
C1112 vdd.n336 vss 0.00251f
C1113 vdd.n337 vss 0.0471f
C1114 vdd.n338 vss 0.00251f
C1115 vdd.n339 vss 0.0112f
C1116 vdd.n340 vss 0.0128f
C1117 vdd.n341 vss 0.0613f
C1118 vdd.n342 vss 0.00324f
C1119 vdd.n343 vss 0.0112f
C1120 vdd.n344 vss 0.0128f
C1121 vdd.n345 vss 0.00413f
C1122 vdd.n346 vss 0.00413f
C1123 vdd.n347 vss 0.0471f
C1124 vdd.n348 vss 0.0471f
C1125 vdd.n349 vss 0.00324f
C1126 vdd.n350 vss 0.00413f
C1127 vdd.n351 vss 0.00413f
C1128 vdd.n352 vss 0.00679f
C1129 vdd.n353 vss 0.00413f
C1130 vdd.n354 vss 0.0471f
C1131 vdd.n355 vss 0.00324f
C1132 vdd.n356 vss 0.0424f
C1133 vdd.n357 vss 0.00324f
C1134 vdd.n358 vss 0.0128f
C1135 vdd.n359 vss 0.02f
C1136 vdd.n360 vss 0.0132f
C1137 vdd.n361 vss 0.00925f
C1138 vdd.n362 vss 0.00425f
C1139 vdd.n364 vss 0.0471f
C1140 vdd.n365 vss 0.00425f
C1141 vdd.n366 vss 0.00413f
C1142 vdd.n367 vss 0.00251f
C1143 vdd.n368 vss 0.0471f
C1144 vdd.n369 vss 0.00251f
C1145 vdd.n370 vss 0.00517f
C1146 vdd.n371 vss 0.00679f
C1147 vdd.n372 vss 0.00324f
C1148 vdd.n373 vss 0.00324f
C1149 vdd.n374 vss 0.0132f
C1150 vdd.n375 vss 0.0424f
C1151 vdd.n376 vss 0.02f
C1152 vdd.n377 vss 0.00425f
C1153 vdd.n379 vss 0.0471f
C1154 vdd.n380 vss 0.00425f
C1155 vdd.n381 vss 0.00925f
C1156 vdd.n382 vss 0.00679f
C1157 vdd.n383 vss 0.00517f
C1158 vdd.n384 vss 0.00251f
C1159 vdd.n385 vss 0.0471f
C1160 vdd.n386 vss 0.00251f
C1161 vdd.n387 vss 0.0112f
C1162 vdd.n388 vss 0.0128f
C1163 vdd.n389 vss 0.0666f
C1164 vdd.n390 vss 0.00324f
C1165 vdd.n391 vss 0.0112f
C1166 vdd.n392 vss 0.0128f
C1167 vdd.n393 vss 0.00413f
C1168 vdd.n394 vss 0.00413f
C1169 vdd.n395 vss 0.0471f
C1170 vdd.n396 vss 0.0471f
C1171 vdd.n397 vss 0.00324f
C1172 vdd.n398 vss 0.00413f
C1173 vdd.n399 vss 0.00413f
C1174 vdd.n400 vss 0.00679f
C1175 vdd.n401 vss 0.00413f
C1176 vdd.n402 vss 0.0471f
C1177 vdd.n403 vss 0.00324f
C1178 vdd.n404 vss 0.0424f
C1179 vdd.n405 vss 0.00324f
C1180 vdd.n406 vss 0.0128f
C1181 vdd.n407 vss 0.02f
C1182 vdd.n408 vss 0.0132f
C1183 vdd.n409 vss 0.00925f
C1184 vdd.n410 vss 0.00425f
C1185 vdd.n412 vss 0.0471f
C1186 vdd.n413 vss 0.00425f
C1187 vdd.n414 vss 0.00413f
C1188 vdd.n415 vss 0.00251f
C1189 vdd.n416 vss 0.0471f
C1190 vdd.n417 vss 0.00251f
C1191 vdd.n418 vss 0.00517f
C1192 vdd.n419 vss 0.00679f
C1193 vdd.n420 vss 0.00324f
C1194 vdd.n421 vss 0.00324f
C1195 vdd.n422 vss 0.0132f
C1196 vdd.n423 vss 0.0424f
C1197 vdd.n424 vss 0.02f
C1198 vdd.n425 vss 0.00425f
C1199 vdd.n427 vss 0.0471f
C1200 vdd.n428 vss 0.00425f
C1201 vdd.n429 vss 0.00925f
C1202 vdd.n430 vss 0.00679f
C1203 vdd.n431 vss 0.00517f
C1204 vdd.n432 vss 0.00251f
C1205 vdd.n433 vss 0.0471f
C1206 vdd.n434 vss 0.00251f
C1207 vdd.n435 vss 0.0112f
C1208 vdd.n436 vss 0.0128f
C1209 vdd.n437 vss 0.0617f
C1210 vdd.n438 vss 0.00335f
C1211 vdd.n439 vss 0.0855f
C1212 vdd.n440 vss 0.0107f
C1213 vdd.n441 vss 0.0128f
C1214 vdd.n442 vss 0.0424f
C1215 vdd.n443 vss 0.00413f
C1216 vdd.n444 vss 0.0471f
C1217 vdd.n445 vss 0.00413f
C1218 vdd.n446 vss 0.00324f
C1219 vdd.n447 vss 0.00324f
C1220 vdd.n448 vss 0.00679f
C1221 vdd.n449 vss 0.00413f
C1222 vdd.n450 vss 0.0471f
C1223 vdd.n451 vss 0.00413f
C1224 vdd.n452 vss 0.0105f
C1225 vdd.n453 vss 0.0471f
C1226 vdd.n454 vss 0.00413f
C1227 vdd.n455 vss 0.00324f
C1228 vdd.n456 vss 0.00324f
C1229 vdd.n457 vss 0.0132f
C1230 vdd.n458 vss 0.0424f
C1231 vdd.n459 vss 0.0128f
C1232 vdd.n460 vss 0.02f
C1233 vdd.n461 vss 0.00425f
C1234 vdd.n463 vss 0.0471f
C1235 vdd.n464 vss 0.00425f
C1236 vdd.n465 vss 0.00925f
C1237 vdd.n466 vss 0.00679f
C1238 vdd.n467 vss 0.00517f
C1239 vdd.n468 vss 0.00251f
C1240 vdd.n469 vss 0.0471f
C1241 vdd.n470 vss 0.00251f
C1242 vdd.n471 vss 0.00413f
C1243 vdd.n472 vss 0.00324f
C1244 vdd.n473 vss 0.00324f
C1245 vdd.n474 vss 0.00805f
C1246 vdd.n475 vss 0.0112f
C1247 vdd.n476 vss 0.00251f
C1248 vdd.n477 vss 0.0471f
C1249 vdd.n478 vss 0.00251f
C1250 vdd.n479 vss 0.00517f
C1251 vdd.n480 vss 0.00679f
C1252 vdd.n481 vss 0.00925f
C1253 vdd.n482 vss 0.00425f
C1254 vdd.n484 vss 0.0471f
C1255 vdd.n485 vss 0.00425f
C1256 vdd.n486 vss 0.00991f
C1257 vdd.n487 vss 0.0126f
C1258 vdd.n488 vss 0.0516f
C1259 vdd.n489 vss 0.0011f
C1260 vdd.n490 vss 0.0271f
C1261 vdd.n491 vss 0.00324f
C1262 vdd.n492 vss 0.0112f
C1263 vdd.n493 vss 0.0128f
C1264 vdd.n494 vss 0.00413f
C1265 vdd.n495 vss 0.00413f
C1266 vdd.n496 vss 0.0471f
C1267 vdd.n497 vss 0.0471f
C1268 vdd.n498 vss 0.00324f
C1269 vdd.n499 vss 0.00413f
C1270 vdd.n500 vss 0.00413f
C1271 vdd.n501 vss 0.00679f
C1272 vdd.n502 vss 0.00413f
C1273 vdd.n503 vss 0.0471f
C1274 vdd.n504 vss 0.00324f
C1275 vdd.n505 vss 0.0424f
C1276 vdd.n506 vss 0.00324f
C1277 vdd.n507 vss 0.0128f
C1278 vdd.n508 vss 0.02f
C1279 vdd.n509 vss 0.0132f
C1280 vdd.n510 vss 0.00925f
C1281 vdd.n511 vss 0.00425f
C1282 vdd.n513 vss 0.0471f
C1283 vdd.n514 vss 0.00425f
C1284 vdd.n515 vss 0.00413f
C1285 vdd.n516 vss 0.00251f
C1286 vdd.n517 vss 0.0471f
C1287 vdd.n518 vss 0.00251f
C1288 vdd.n519 vss 0.00517f
C1289 vdd.n520 vss 0.00679f
C1290 vdd.n521 vss 0.00324f
C1291 vdd.n522 vss 0.00324f
C1292 vdd.n523 vss 0.0132f
C1293 vdd.n524 vss 0.0424f
C1294 vdd.n525 vss 0.02f
C1295 vdd.n526 vss 0.00425f
C1296 vdd.n528 vss 0.0471f
C1297 vdd.n529 vss 0.00425f
C1298 vdd.n530 vss 0.00925f
C1299 vdd.n531 vss 0.00679f
C1300 vdd.n532 vss 0.00517f
C1301 vdd.n533 vss 0.00251f
C1302 vdd.n534 vss 0.0471f
C1303 vdd.n535 vss 0.00251f
C1304 vdd.n536 vss 0.0112f
C1305 vdd.n537 vss 0.0128f
C1306 vdd.n538 vss 0.0666f
C1307 vdd.n539 vss 0.00324f
C1308 vdd.n540 vss 0.0112f
C1309 vdd.n541 vss 0.0128f
C1310 vdd.n542 vss 0.00413f
C1311 vdd.n543 vss 0.00413f
C1312 vdd.n544 vss 0.0471f
C1313 vdd.n545 vss 0.0471f
C1314 vdd.n546 vss 0.00324f
C1315 vdd.n547 vss 0.00413f
C1316 vdd.n548 vss 0.00413f
C1317 vdd.n549 vss 0.00679f
C1318 vdd.n550 vss 0.00413f
C1319 vdd.n551 vss 0.0471f
C1320 vdd.n552 vss 0.00324f
C1321 vdd.n553 vss 0.0424f
C1322 vdd.n554 vss 0.00324f
C1323 vdd.n555 vss 0.0128f
C1324 vdd.n556 vss 0.02f
C1325 vdd.n557 vss 0.0132f
C1326 vdd.n558 vss 0.00925f
C1327 vdd.n559 vss 0.00425f
C1328 vdd.n561 vss 0.0471f
C1329 vdd.n562 vss 0.00425f
C1330 vdd.n563 vss 0.00413f
C1331 vdd.n564 vss 0.00251f
C1332 vdd.n565 vss 0.0471f
C1333 vdd.n566 vss 0.00251f
C1334 vdd.n567 vss 0.00517f
C1335 vdd.n568 vss 0.00679f
C1336 vdd.n569 vss 0.00324f
C1337 vdd.n570 vss 0.00324f
C1338 vdd.n571 vss 0.0132f
C1339 vdd.n572 vss 0.0424f
C1340 vdd.n573 vss 0.02f
C1341 vdd.n574 vss 0.00425f
C1342 vdd.n576 vss 0.0471f
C1343 vdd.n577 vss 0.00425f
C1344 vdd.n578 vss 0.00925f
C1345 vdd.n579 vss 0.00679f
C1346 vdd.n580 vss 0.00517f
C1347 vdd.n581 vss 0.00251f
C1348 vdd.n582 vss 0.0471f
C1349 vdd.n583 vss 0.00251f
C1350 vdd.n584 vss 0.0112f
C1351 vdd.n585 vss 0.0128f
C1352 vdd.n586 vss 0.0599f
C1353 vdd.n587 vss 0.00324f
C1354 vdd.n588 vss 0.0112f
C1355 vdd.n589 vss 0.0128f
C1356 vdd.n590 vss 0.00413f
C1357 vdd.n591 vss 0.00413f
C1358 vdd.n592 vss 0.0471f
C1359 vdd.n593 vss 0.0471f
C1360 vdd.n594 vss 0.00324f
C1361 vdd.n595 vss 0.00413f
C1362 vdd.n596 vss 0.00413f
C1363 vdd.n597 vss 0.00679f
C1364 vdd.n598 vss 0.00413f
C1365 vdd.n599 vss 0.0471f
C1366 vdd.n600 vss 0.00324f
C1367 vdd.n602 vss 0.00925f
C1368 vdd.n603 vss 0.0471f
C1369 vdd.n604 vss 0.00425f
C1370 vdd.n605 vss 0.0424f
C1371 vdd.n606 vss 0.0132f
C1372 vdd.n607 vss 0.00324f
C1373 vdd.n608 vss 0.0128f
C1374 vdd.n609 vss 0.02f
C1375 vdd.n610 vss 0.00425f
C1376 vdd.n611 vss 0.00413f
C1377 vdd.n612 vss 0.00251f
C1378 vdd.n613 vss 0.0471f
C1379 vdd.n614 vss 0.00251f
C1380 vdd.n615 vss 0.00517f
C1381 vdd.n616 vss 0.00679f
C1382 vdd.n617 vss 0.00324f
C1383 vdd.n618 vss 0.00324f
C1384 vdd.n619 vss 0.0132f
C1385 vdd.n620 vss 0.0424f
C1386 vdd.n621 vss 0.02f
C1387 vdd.n622 vss 0.00425f
C1388 vdd.n623 vss 0.0471f
C1389 vdd.n625 vss 0.00425f
C1390 vdd.n626 vss 0.00925f
C1391 vdd.n627 vss 0.00679f
C1392 vdd.n628 vss 0.00517f
C1393 vdd.n629 vss 0.00251f
C1394 vdd.n630 vss 0.0471f
C1395 vdd.n631 vss 0.00251f
C1396 vdd.n632 vss 0.0112f
C1397 vdd.n633 vss 0.098f
C1398 vdd.n634 vss 0.00324f
C1399 vdd.n635 vss 0.0112f
C1400 vdd.n636 vss 0.0128f
C1401 vdd.n637 vss 0.00413f
C1402 vdd.n638 vss 0.00413f
C1403 vdd.n639 vss 0.0471f
C1404 vdd.n640 vss 0.0471f
C1405 vdd.n641 vss 0.00324f
C1406 vdd.n642 vss 0.00413f
C1407 vdd.n643 vss 0.00413f
C1408 vdd.n644 vss 0.00679f
C1409 vdd.n645 vss 0.00413f
C1410 vdd.n646 vss 0.0471f
C1411 vdd.n647 vss 0.00324f
C1412 vdd.n648 vss 0.0424f
C1413 vdd.n649 vss 0.00324f
C1414 vdd.n650 vss 0.0128f
C1415 vdd.n651 vss 0.02f
C1416 vdd.n652 vss 0.0132f
C1417 vdd.n653 vss 0.00925f
C1418 vdd.n654 vss 0.00425f
C1419 vdd.n656 vss 0.0471f
C1420 vdd.n657 vss 0.00425f
C1421 vdd.n658 vss 0.00413f
C1422 vdd.n659 vss 0.00251f
C1423 vdd.n660 vss 0.0471f
C1424 vdd.n661 vss 0.00251f
C1425 vdd.n662 vss 0.00517f
C1426 vdd.n663 vss 0.00679f
C1427 vdd.n664 vss 0.00324f
C1428 vdd.n665 vss 0.00324f
C1429 vdd.n666 vss 0.0132f
C1430 vdd.n667 vss 0.0424f
C1431 vdd.n668 vss 0.02f
C1432 vdd.n669 vss 0.00425f
C1433 vdd.n671 vss 0.0471f
C1434 vdd.n672 vss 0.00425f
C1435 vdd.n673 vss 0.00925f
C1436 vdd.n674 vss 0.00679f
C1437 vdd.n675 vss 0.00517f
C1438 vdd.n676 vss 0.00251f
C1439 vdd.n677 vss 0.0471f
C1440 vdd.n678 vss 0.00251f
C1441 vdd.n679 vss 0.0112f
C1442 vdd.n680 vss 0.0128f
C1443 vdd.n681 vss 0.0599f
C1444 vdd.n682 vss 0.202f
C1445 vdd.n683 vss 0.00324f
C1446 vdd.n684 vss 0.0112f
C1447 vdd.n685 vss 0.0128f
C1448 vdd.n686 vss 0.00413f
C1449 vdd.n687 vss 0.00413f
C1450 vdd.n688 vss 0.0471f
C1451 vdd.n689 vss 0.0471f
C1452 vdd.n690 vss 0.00324f
C1453 vdd.n691 vss 0.00413f
C1454 vdd.n692 vss 0.00413f
C1455 vdd.n693 vss 0.00679f
C1456 vdd.n694 vss 0.00413f
C1457 vdd.n695 vss 0.0471f
C1458 vdd.n696 vss 0.00324f
C1459 vdd.n698 vss 0.00925f
C1460 vdd.n699 vss 0.0471f
C1461 vdd.n700 vss 0.00425f
C1462 vdd.n701 vss 0.0424f
C1463 vdd.n702 vss 0.0132f
C1464 vdd.n703 vss 0.00324f
C1465 vdd.n704 vss 0.0128f
C1466 vdd.n705 vss 0.02f
C1467 vdd.n706 vss 0.00425f
C1468 vdd.n707 vss 0.00413f
C1469 vdd.n708 vss 0.00251f
C1470 vdd.n709 vss 0.0471f
C1471 vdd.n710 vss 0.00251f
C1472 vdd.n711 vss 0.00517f
C1473 vdd.n712 vss 0.00679f
C1474 vdd.n713 vss 0.00324f
C1475 vdd.n714 vss 0.00324f
C1476 vdd.n715 vss 0.0132f
C1477 vdd.n716 vss 0.0424f
C1478 vdd.n717 vss 0.02f
C1479 vdd.n718 vss 0.00425f
C1480 vdd.n719 vss 0.0471f
C1481 vdd.n721 vss 0.00425f
C1482 vdd.n722 vss 0.00925f
C1483 vdd.n723 vss 0.00679f
C1484 vdd.n724 vss 0.00517f
C1485 vdd.n725 vss 0.00251f
C1486 vdd.n726 vss 0.0471f
C1487 vdd.n727 vss 0.00251f
C1488 vdd.n728 vss 0.0112f
C1489 vdd.n729 vss 0.0128f
C1490 vdd.n730 vss 0.0692f
C1491 vdd.n731 vss 0.00324f
C1492 vdd.n732 vss 0.0112f
C1493 vdd.n733 vss 0.0128f
C1494 vdd.n734 vss 0.00413f
C1495 vdd.n735 vss 0.00413f
C1496 vdd.n736 vss 0.0471f
C1497 vdd.n737 vss 0.0471f
C1498 vdd.n738 vss 0.00324f
C1499 vdd.n739 vss 0.00413f
C1500 vdd.n740 vss 0.00413f
C1501 vdd.n741 vss 0.00679f
C1502 vdd.n742 vss 0.00413f
C1503 vdd.n743 vss 0.0471f
C1504 vdd.n744 vss 0.00324f
C1505 vdd.n746 vss 0.00925f
C1506 vdd.n747 vss 0.0471f
C1507 vdd.n748 vss 0.00425f
C1508 vdd.n749 vss 0.0424f
C1509 vdd.n750 vss 0.0132f
C1510 vdd.n751 vss 0.00324f
C1511 vdd.n752 vss 0.0128f
C1512 vdd.n753 vss 0.02f
C1513 vdd.n754 vss 0.00425f
C1514 vdd.n755 vss 0.00413f
C1515 vdd.n756 vss 0.00251f
C1516 vdd.n757 vss 0.0471f
C1517 vdd.n758 vss 0.00251f
C1518 vdd.n759 vss 0.00517f
C1519 vdd.n760 vss 0.00679f
C1520 vdd.n761 vss 0.00324f
C1521 vdd.n762 vss 0.00324f
C1522 vdd.n763 vss 0.0132f
C1523 vdd.n764 vss 0.0424f
C1524 vdd.n765 vss 0.02f
C1525 vdd.n766 vss 0.00425f
C1526 vdd.n767 vss 0.0471f
C1527 vdd.n769 vss 0.00425f
C1528 vdd.n770 vss 0.00925f
C1529 vdd.n771 vss 0.00679f
C1530 vdd.n772 vss 0.00517f
C1531 vdd.n773 vss 0.00251f
C1532 vdd.n774 vss 0.0471f
C1533 vdd.n775 vss 0.00251f
C1534 vdd.n776 vss 0.0112f
C1535 vdd.n777 vss 0.0128f
C1536 vdd.n778 vss 0.0619f
C1537 vdd.n779 vss 0.00335f
C1538 vdd.n780 vss 0.0855f
C1539 vdd.n781 vss 0.00991f
C1540 vdd.n782 vss 0.0424f
C1541 vdd.n783 vss 0.00679f
C1542 vdd.n784 vss 0.00413f
C1543 vdd.n785 vss 0.0471f
C1544 vdd.n786 vss 0.00251f
C1545 vdd.n787 vss 0.00679f
C1546 vdd.n788 vss 0.00413f
C1547 vdd.n789 vss 0.00413f
C1548 vdd.n790 vss 0.0471f
C1549 vdd.n791 vss 0.00251f
C1550 vdd.n792 vss 0.00413f
C1551 vdd.n793 vss 0.00324f
C1552 vdd.n794 vss 0.0132f
C1553 vdd.n795 vss 0.0424f
C1554 vdd.n796 vss 0.00324f
C1555 vdd.n797 vss 0.00413f
C1556 vdd.n798 vss 0.00517f
C1557 vdd.n799 vss 0.00679f
C1558 vdd.n800 vss 0.00925f
C1559 vdd.n801 vss 0.00425f
C1560 vdd.n802 vss 0.0471f
C1561 vdd.n804 vss 0.00425f
C1562 vdd.n805 vss 0.02f
C1563 vdd.n806 vss 0.0128f
C1564 vdd.n807 vss 0.0105f
C1565 vdd.n808 vss 0.00251f
C1566 vdd.n809 vss 0.0471f
C1567 vdd.n810 vss 0.00517f
C1568 vdd.n811 vss 0.00251f
C1569 vdd.n812 vss 0.0471f
C1570 vdd.n813 vss 0.0471f
C1571 vdd.n814 vss 0.00324f
C1572 vdd.n815 vss 0.00324f
C1573 vdd.n816 vss 0.00805f
C1574 vdd.n817 vss 0.0112f
C1575 vdd.n818 vss 0.0128f
C1576 vdd.n819 vss 0.00324f
C1577 vdd.n820 vss 0.00324f
C1578 vdd.n821 vss 0.00413f
C1579 vdd.n822 vss 0.00425f
C1580 vdd.n823 vss 0.0471f
C1581 vdd.n825 vss 0.00425f
C1582 vdd.n826 vss 0.00925f
C1583 vdd.n827 vss 0.0107f
C1584 vdd.n828 vss 0.0126f
C1585 vdd.n829 vss 0.0516f
C1586 vdd.n830 vss 0.00163f
C1587 vdd.n831 vss 0.00145f
C1588 vdd.n832 vss 0.0271f
C1589 vdd.n833 vss 0.00324f
C1590 vdd.n834 vss 0.0112f
C1591 vdd.n835 vss 0.0128f
C1592 vdd.n836 vss 0.00413f
C1593 vdd.n837 vss 0.00413f
C1594 vdd.n838 vss 0.0471f
C1595 vdd.n839 vss 0.0471f
C1596 vdd.n840 vss 0.00324f
C1597 vdd.n841 vss 0.00413f
C1598 vdd.n842 vss 0.00413f
C1599 vdd.n843 vss 0.00679f
C1600 vdd.n844 vss 0.00413f
C1601 vdd.n845 vss 0.0471f
C1602 vdd.n846 vss 0.00324f
C1603 vdd.n848 vss 0.00925f
C1604 vdd.n849 vss 0.0471f
C1605 vdd.n850 vss 0.00425f
C1606 vdd.n851 vss 0.0424f
C1607 vdd.n852 vss 0.0132f
C1608 vdd.n853 vss 0.00324f
C1609 vdd.n854 vss 0.0128f
C1610 vdd.n855 vss 0.02f
C1611 vdd.n856 vss 0.00425f
C1612 vdd.n857 vss 0.00413f
C1613 vdd.n858 vss 0.00251f
C1614 vdd.n859 vss 0.0471f
C1615 vdd.n860 vss 0.00251f
C1616 vdd.n861 vss 0.00517f
C1617 vdd.n862 vss 0.00679f
C1618 vdd.n863 vss 0.00324f
C1619 vdd.n864 vss 0.00324f
C1620 vdd.n865 vss 0.0132f
C1621 vdd.n866 vss 0.0424f
C1622 vdd.n867 vss 0.02f
C1623 vdd.n868 vss 0.00425f
C1624 vdd.n869 vss 0.0471f
C1625 vdd.n871 vss 0.00425f
C1626 vdd.n872 vss 0.00925f
C1627 vdd.n873 vss 0.00679f
C1628 vdd.n874 vss 0.00517f
C1629 vdd.n875 vss 0.00251f
C1630 vdd.n876 vss 0.0471f
C1631 vdd.n877 vss 0.00251f
C1632 vdd.n878 vss 0.0112f
C1633 vdd.n879 vss 0.0128f
C1634 vdd.n880 vss 0.0692f
C1635 vdd.n881 vss 0.00324f
C1636 vdd.n882 vss 0.0112f
C1637 vdd.n883 vss 0.0128f
C1638 vdd.n884 vss 0.00413f
C1639 vdd.n885 vss 0.00413f
C1640 vdd.n886 vss 0.0471f
C1641 vdd.n887 vss 0.0471f
C1642 vdd.n888 vss 0.00324f
C1643 vdd.n889 vss 0.00413f
C1644 vdd.n890 vss 0.00413f
C1645 vdd.n891 vss 0.00679f
C1646 vdd.n892 vss 0.00413f
C1647 vdd.n893 vss 0.0471f
C1648 vdd.n894 vss 0.00324f
C1649 vdd.n896 vss 0.00925f
C1650 vdd.n897 vss 0.0471f
C1651 vdd.n898 vss 0.00425f
C1652 vdd.n899 vss 0.0424f
C1653 vdd.n900 vss 0.0132f
C1654 vdd.n901 vss 0.00324f
C1655 vdd.n902 vss 0.0128f
C1656 vdd.n903 vss 0.02f
C1657 vdd.n904 vss 0.00425f
C1658 vdd.n905 vss 0.00413f
C1659 vdd.n906 vss 0.00251f
C1660 vdd.n907 vss 0.0471f
C1661 vdd.n908 vss 0.00251f
C1662 vdd.n909 vss 0.00517f
C1663 vdd.n910 vss 0.00679f
C1664 vdd.n911 vss 0.00324f
C1665 vdd.n912 vss 0.00324f
C1666 vdd.n913 vss 0.0132f
C1667 vdd.n914 vss 0.0424f
C1668 vdd.n915 vss 0.02f
C1669 vdd.n916 vss 0.00425f
C1670 vdd.n917 vss 0.0471f
C1671 vdd.n919 vss 0.00425f
C1672 vdd.n920 vss 0.00925f
C1673 vdd.n921 vss 0.00679f
C1674 vdd.n922 vss 0.00517f
C1675 vdd.n923 vss 0.00251f
C1676 vdd.n924 vss 0.0471f
C1677 vdd.n925 vss 0.00251f
C1678 vdd.n926 vss 0.0112f
C1679 vdd.n927 vss 0.0128f
C1680 vdd.n928 vss 0.0619f
C1681 vdd.n929 vss 0.00324f
C1682 vdd.n930 vss 0.0112f
C1683 vdd.n931 vss 0.0128f
C1684 vdd.n932 vss 0.00413f
C1685 vdd.n933 vss 0.00413f
C1686 vdd.n934 vss 0.0471f
C1687 vdd.n935 vss 0.0471f
C1688 vdd.n936 vss 0.00324f
C1689 vdd.n937 vss 0.00413f
C1690 vdd.n938 vss 0.00413f
C1691 vdd.n939 vss 0.00679f
C1692 vdd.n940 vss 0.00413f
C1693 vdd.n941 vss 0.0471f
C1694 vdd.n942 vss 0.00324f
C1695 vdd.n944 vss 0.00925f
C1696 vdd.n945 vss 0.0471f
C1697 vdd.n946 vss 0.00425f
C1698 vdd.n947 vss 0.0424f
C1699 vdd.n948 vss 0.0132f
C1700 vdd.n949 vss 0.00324f
C1701 vdd.n950 vss 0.0128f
C1702 vdd.n951 vss 0.02f
C1703 vdd.n952 vss 0.00425f
C1704 vdd.n953 vss 0.00413f
C1705 vdd.n954 vss 0.00251f
C1706 vdd.n955 vss 0.0471f
C1707 vdd.n956 vss 0.00251f
C1708 vdd.n957 vss 0.00517f
C1709 vdd.n958 vss 0.00679f
C1710 vdd.n959 vss 0.00324f
C1711 vdd.n960 vss 0.00324f
C1712 vdd.n961 vss 0.0132f
C1713 vdd.n962 vss 0.0424f
C1714 vdd.n963 vss 0.02f
C1715 vdd.n964 vss 0.00425f
C1716 vdd.n965 vss 0.0471f
C1717 vdd.n967 vss 0.00425f
C1718 vdd.n968 vss 0.00925f
C1719 vdd.n969 vss 0.00679f
C1720 vdd.n970 vss 0.00517f
C1721 vdd.n971 vss 0.00251f
C1722 vdd.n972 vss 0.0471f
C1723 vdd.n973 vss 0.00251f
C1724 vdd.n974 vss 0.0112f
C1725 vdd.n975 vss 0.0128f
C1726 vdd.n976 vss 0.0692f
C1727 vdd.n977 vss 0.00324f
C1728 vdd.n978 vss 0.0112f
C1729 vdd.n979 vss 0.0128f
C1730 vdd.n980 vss 0.00413f
C1731 vdd.n981 vss 0.00413f
C1732 vdd.n982 vss 0.0471f
C1733 vdd.n983 vss 0.0471f
C1734 vdd.n984 vss 0.00324f
C1735 vdd.n985 vss 0.00413f
C1736 vdd.n986 vss 0.00413f
C1737 vdd.n987 vss 0.00679f
C1738 vdd.n988 vss 0.00413f
C1739 vdd.n989 vss 0.0471f
C1740 vdd.n990 vss 0.00324f
C1741 vdd.n992 vss 0.00925f
C1742 vdd.n993 vss 0.0471f
C1743 vdd.n994 vss 0.00425f
C1744 vdd.n995 vss 0.0424f
C1745 vdd.n996 vss 0.0132f
C1746 vdd.n997 vss 0.00324f
C1747 vdd.n998 vss 0.0128f
C1748 vdd.n999 vss 0.02f
C1749 vdd.n1000 vss 0.00425f
C1750 vdd.n1001 vss 0.00413f
C1751 vdd.n1002 vss 0.00251f
C1752 vdd.n1003 vss 0.0471f
C1753 vdd.n1004 vss 0.00251f
C1754 vdd.n1005 vss 0.00517f
C1755 vdd.n1006 vss 0.00679f
C1756 vdd.n1007 vss 0.00324f
C1757 vdd.n1008 vss 0.00324f
C1758 vdd.n1009 vss 0.0132f
C1759 vdd.n1010 vss 0.0424f
C1760 vdd.n1011 vss 0.02f
C1761 vdd.n1012 vss 0.00425f
C1762 vdd.n1013 vss 0.0471f
C1763 vdd.n1015 vss 0.00425f
C1764 vdd.n1016 vss 0.00925f
C1765 vdd.n1017 vss 0.00679f
C1766 vdd.n1018 vss 0.00517f
C1767 vdd.n1019 vss 0.00251f
C1768 vdd.n1020 vss 0.0471f
C1769 vdd.n1021 vss 0.00251f
C1770 vdd.n1022 vss 0.0112f
C1771 vdd.n1023 vss 0.0128f
C1772 vdd.n1024 vss 0.0619f
C1773 vdd.n1025 vss 0.00335f
C1774 vdd.n1026 vss 0.0855f
C1775 vdd.n1027 vss 0.00991f
C1776 vdd.n1028 vss 0.0424f
C1777 vdd.n1029 vss 0.00679f
C1778 vdd.n1030 vss 0.00413f
C1779 vdd.n1031 vss 0.0471f
C1780 vdd.n1032 vss 0.00251f
C1781 vdd.n1033 vss 0.00679f
C1782 vdd.n1034 vss 0.00413f
C1783 vdd.n1035 vss 0.00413f
C1784 vdd.n1036 vss 0.0471f
C1785 vdd.n1037 vss 0.00251f
C1786 vdd.n1038 vss 0.00413f
C1787 vdd.n1039 vss 0.00324f
C1788 vdd.n1040 vss 0.0132f
C1789 vdd.n1041 vss 0.0424f
C1790 vdd.n1042 vss 0.00324f
C1791 vdd.n1043 vss 0.00413f
C1792 vdd.n1044 vss 0.00517f
C1793 vdd.n1045 vss 0.00679f
C1794 vdd.n1046 vss 0.00925f
C1795 vdd.n1047 vss 0.00425f
C1796 vdd.n1048 vss 0.0471f
C1797 vdd.n1050 vss 0.00425f
C1798 vdd.n1051 vss 0.02f
C1799 vdd.n1052 vss 0.0128f
C1800 vdd.n1053 vss 0.0105f
C1801 vdd.n1054 vss 0.00251f
C1802 vdd.n1055 vss 0.0471f
C1803 vdd.n1056 vss 0.00517f
C1804 vdd.n1057 vss 0.00251f
C1805 vdd.n1058 vss 0.0471f
C1806 vdd.n1059 vss 0.0471f
C1807 vdd.n1060 vss 0.00324f
C1808 vdd.n1061 vss 0.00324f
C1809 vdd.n1062 vss 0.00805f
C1810 vdd.n1063 vss 0.0112f
C1811 vdd.n1064 vss 0.0128f
C1812 vdd.n1065 vss 0.00324f
C1813 vdd.n1066 vss 0.00324f
C1814 vdd.n1067 vss 0.00413f
C1815 vdd.n1068 vss 0.00425f
C1816 vdd.n1069 vss 0.0471f
C1817 vdd.n1071 vss 0.00425f
C1818 vdd.n1072 vss 0.00925f
C1819 vdd.n1073 vss 0.0107f
C1820 vdd.n1074 vss 0.0126f
C1821 vdd.n1075 vss 0.0516f
C1822 vdd.n1076 vss 0.00163f
C1823 vdd.n1077 vss 0.00145f
C1824 vdd.n1078 vss 0.0271f
C1825 vdd.n1079 vss 0.00324f
C1826 vdd.n1080 vss 0.0112f
C1827 vdd.n1081 vss 0.0128f
C1828 vdd.n1082 vss 0.00413f
C1829 vdd.n1083 vss 0.00413f
C1830 vdd.n1084 vss 0.0471f
C1831 vdd.n1085 vss 0.0471f
C1832 vdd.n1086 vss 0.00324f
C1833 vdd.n1087 vss 0.00413f
C1834 vdd.n1088 vss 0.00413f
C1835 vdd.n1089 vss 0.00679f
C1836 vdd.n1090 vss 0.00413f
C1837 vdd.n1091 vss 0.0471f
C1838 vdd.n1092 vss 0.00324f
C1839 vdd.n1094 vss 0.00925f
C1840 vdd.n1095 vss 0.0471f
C1841 vdd.n1096 vss 0.00425f
C1842 vdd.n1097 vss 0.0424f
C1843 vdd.n1098 vss 0.0132f
C1844 vdd.n1099 vss 0.00324f
C1845 vdd.n1100 vss 0.0128f
C1846 vdd.n1101 vss 0.02f
C1847 vdd.n1102 vss 0.00425f
C1848 vdd.n1103 vss 0.00413f
C1849 vdd.n1104 vss 0.00251f
C1850 vdd.n1105 vss 0.0471f
C1851 vdd.n1106 vss 0.00251f
C1852 vdd.n1107 vss 0.00517f
C1853 vdd.n1108 vss 0.00679f
C1854 vdd.n1109 vss 0.00324f
C1855 vdd.n1110 vss 0.00324f
C1856 vdd.n1111 vss 0.0132f
C1857 vdd.n1112 vss 0.0424f
C1858 vdd.n1113 vss 0.02f
C1859 vdd.n1114 vss 0.00425f
C1860 vdd.n1115 vss 0.0471f
C1861 vdd.n1117 vss 0.00425f
C1862 vdd.n1118 vss 0.00925f
C1863 vdd.n1119 vss 0.00679f
C1864 vdd.n1120 vss 0.00517f
C1865 vdd.n1121 vss 0.00251f
C1866 vdd.n1122 vss 0.0471f
C1867 vdd.n1123 vss 0.00251f
C1868 vdd.n1124 vss 0.0112f
C1869 vdd.n1125 vss 0.0128f
C1870 vdd.n1126 vss 0.0692f
C1871 vdd.n1127 vss 0.00324f
C1872 vdd.n1128 vss 0.0112f
C1873 vdd.n1129 vss 0.0128f
C1874 vdd.n1130 vss 0.00413f
C1875 vdd.n1131 vss 0.00413f
C1876 vdd.n1132 vss 0.0471f
C1877 vdd.n1133 vss 0.0471f
C1878 vdd.n1134 vss 0.00324f
C1879 vdd.n1135 vss 0.00413f
C1880 vdd.n1136 vss 0.00413f
C1881 vdd.n1137 vss 0.00679f
C1882 vdd.n1138 vss 0.00413f
C1883 vdd.n1139 vss 0.0471f
C1884 vdd.n1140 vss 0.00324f
C1885 vdd.n1141 vss 0.0424f
C1886 vdd.n1142 vss 0.00324f
C1887 vdd.n1143 vss 0.0128f
C1888 vdd.n1144 vss 0.02f
C1889 vdd.n1145 vss 0.0132f
C1890 vdd.n1146 vss 0.00925f
C1891 vdd.n1147 vss 0.00425f
C1892 vdd.n1149 vss 0.0471f
C1893 vdd.n1150 vss 0.00425f
C1894 vdd.n1151 vss 0.00413f
C1895 vdd.n1152 vss 0.00251f
C1896 vdd.n1153 vss 0.0471f
C1897 vdd.n1154 vss 0.00251f
C1898 vdd.n1155 vss 0.00517f
C1899 vdd.n1156 vss 0.00679f
C1900 vdd.n1157 vss 0.00324f
C1901 vdd.n1158 vss 0.00324f
C1902 vdd.n1159 vss 0.0132f
C1903 vdd.n1160 vss 0.0424f
C1904 vdd.n1161 vss 0.02f
C1905 vdd.n1162 vss 0.00425f
C1906 vdd.n1164 vss 0.0471f
C1907 vdd.n1165 vss 0.00425f
C1908 vdd.n1166 vss 0.00925f
C1909 vdd.n1167 vss 0.00679f
C1910 vdd.n1168 vss 0.00517f
C1911 vdd.n1169 vss 0.00251f
C1912 vdd.n1170 vss 0.0471f
C1913 vdd.n1171 vss 0.00251f
C1914 vdd.n1172 vss 0.0112f
C1915 vdd.n1173 vss 0.0128f
C1916 vdd.n1174 vss 0.0666f
C1917 vdd.n1175 vss 0.00324f
C1918 vdd.n1176 vss 0.0112f
C1919 vdd.n1177 vss 0.0128f
C1920 vdd.n1178 vss 0.00413f
C1921 vdd.n1179 vss 0.00413f
C1922 vdd.n1180 vss 0.0471f
C1923 vdd.n1181 vss 0.0471f
C1924 vdd.n1182 vss 0.00324f
C1925 vdd.n1183 vss 0.00413f
C1926 vdd.n1184 vss 0.00413f
C1927 vdd.n1185 vss 0.00679f
C1928 vdd.n1186 vss 0.00413f
C1929 vdd.n1187 vss 0.0471f
C1930 vdd.n1188 vss 0.00324f
C1931 vdd.n1189 vss 0.0424f
C1932 vdd.n1190 vss 0.00324f
C1933 vdd.n1191 vss 0.0128f
C1934 vdd.n1192 vss 0.02f
C1935 vdd.n1193 vss 0.0132f
C1936 vdd.n1194 vss 0.00925f
C1937 vdd.n1195 vss 0.00425f
C1938 vdd.n1197 vss 0.0471f
C1939 vdd.n1198 vss 0.00425f
C1940 vdd.n1199 vss 0.00413f
C1941 vdd.n1200 vss 0.00251f
C1942 vdd.n1201 vss 0.0471f
C1943 vdd.n1202 vss 0.00251f
C1944 vdd.n1203 vss 0.00517f
C1945 vdd.n1204 vss 0.00679f
C1946 vdd.n1205 vss 0.00324f
C1947 vdd.n1206 vss 0.00324f
C1948 vdd.n1207 vss 0.0132f
C1949 vdd.n1208 vss 0.0424f
C1950 vdd.n1209 vss 0.02f
C1951 vdd.n1210 vss 0.00425f
C1952 vdd.n1212 vss 0.0471f
C1953 vdd.n1213 vss 0.00425f
C1954 vdd.n1214 vss 0.00925f
C1955 vdd.n1215 vss 0.00679f
C1956 vdd.n1216 vss 0.00517f
C1957 vdd.n1217 vss 0.00251f
C1958 vdd.n1218 vss 0.0471f
C1959 vdd.n1219 vss 0.00251f
C1960 vdd.n1220 vss 0.0112f
C1961 vdd.n1221 vss 0.0128f
C1962 vdd.n1222 vss 0.0617f
C1963 vdd.n1223 vss 0.00335f
C1964 vdd.n1224 vss 0.0855f
C1965 vdd.n1225 vss 0.0107f
C1966 vdd.n1226 vss 0.0128f
C1967 vdd.n1227 vss 0.0424f
C1968 vdd.n1228 vss 0.00413f
C1969 vdd.n1229 vss 0.0471f
C1970 vdd.n1230 vss 0.00413f
C1971 vdd.n1231 vss 0.00324f
C1972 vdd.n1232 vss 0.00324f
C1973 vdd.n1233 vss 0.00679f
C1974 vdd.n1234 vss 0.00413f
C1975 vdd.n1235 vss 0.0471f
C1976 vdd.n1236 vss 0.00413f
C1977 vdd.n1237 vss 0.0105f
C1978 vdd.n1238 vss 0.0471f
C1979 vdd.n1239 vss 0.00413f
C1980 vdd.n1240 vss 0.00324f
C1981 vdd.n1241 vss 0.00324f
C1982 vdd.n1242 vss 0.0132f
C1983 vdd.n1243 vss 0.0424f
C1984 vdd.n1244 vss 0.0128f
C1985 vdd.n1245 vss 0.02f
C1986 vdd.n1246 vss 0.00425f
C1987 vdd.n1248 vss 0.0471f
C1988 vdd.n1249 vss 0.00425f
C1989 vdd.n1250 vss 0.00925f
C1990 vdd.n1251 vss 0.00679f
C1991 vdd.n1252 vss 0.00517f
C1992 vdd.n1253 vss 0.00251f
C1993 vdd.n1254 vss 0.0471f
C1994 vdd.n1255 vss 0.00251f
C1995 vdd.n1256 vss 0.00413f
C1996 vdd.n1257 vss 0.00324f
C1997 vdd.n1258 vss 0.00324f
C1998 vdd.n1259 vss 0.00805f
C1999 vdd.n1260 vss 0.0112f
C2000 vdd.n1261 vss 0.00251f
C2001 vdd.n1262 vss 0.0471f
C2002 vdd.n1263 vss 0.00251f
C2003 vdd.n1264 vss 0.00517f
C2004 vdd.n1265 vss 0.00679f
C2005 vdd.n1266 vss 0.00925f
C2006 vdd.n1267 vss 0.00425f
C2007 vdd.n1269 vss 0.0471f
C2008 vdd.n1270 vss 0.00425f
C2009 vdd.n1271 vss 0.00991f
C2010 vdd.n1272 vss 0.0126f
C2011 vdd.n1273 vss 0.0516f
C2012 vdd.n1274 vss 0.0011f
C2013 vdd.n1275 vss 0.0271f
C2014 vdd.n1276 vss 0.00324f
C2015 vdd.n1277 vss 0.0112f
C2016 vdd.n1278 vss 0.0128f
C2017 vdd.n1279 vss 0.00413f
C2018 vdd.n1280 vss 0.00413f
C2019 vdd.n1281 vss 0.0471f
C2020 vdd.n1282 vss 0.0471f
C2021 vdd.n1283 vss 0.00324f
C2022 vdd.n1284 vss 0.00413f
C2023 vdd.n1285 vss 0.00413f
C2024 vdd.n1286 vss 0.00679f
C2025 vdd.n1287 vss 0.00413f
C2026 vdd.n1288 vss 0.0471f
C2027 vdd.n1289 vss 0.00324f
C2028 vdd.n1290 vss 0.0424f
C2029 vdd.n1291 vss 0.00324f
C2030 vdd.n1292 vss 0.0128f
C2031 vdd.n1293 vss 0.02f
C2032 vdd.n1294 vss 0.0132f
C2033 vdd.n1295 vss 0.00925f
C2034 vdd.n1296 vss 0.00425f
C2035 vdd.n1298 vss 0.0471f
C2036 vdd.n1299 vss 0.00425f
C2037 vdd.n1300 vss 0.00413f
C2038 vdd.n1301 vss 0.00251f
C2039 vdd.n1302 vss 0.0471f
C2040 vdd.n1303 vss 0.00251f
C2041 vdd.n1304 vss 0.00517f
C2042 vdd.n1305 vss 0.00679f
C2043 vdd.n1306 vss 0.00324f
C2044 vdd.n1307 vss 0.00324f
C2045 vdd.n1308 vss 0.0132f
C2046 vdd.n1309 vss 0.0424f
C2047 vdd.n1310 vss 0.02f
C2048 vdd.n1311 vss 0.00425f
C2049 vdd.n1313 vss 0.0471f
C2050 vdd.n1314 vss 0.00425f
C2051 vdd.n1315 vss 0.00925f
C2052 vdd.n1316 vss 0.00679f
C2053 vdd.n1317 vss 0.00517f
C2054 vdd.n1318 vss 0.00251f
C2055 vdd.n1319 vss 0.0471f
C2056 vdd.n1320 vss 0.00251f
C2057 vdd.n1321 vss 0.0112f
C2058 vdd.n1322 vss 0.0128f
C2059 vdd.n1323 vss 0.0666f
C2060 vdd.n1324 vss 0.00324f
C2061 vdd.n1325 vss 0.0112f
C2062 vdd.n1326 vss 0.0128f
C2063 vdd.n1327 vss 0.00413f
C2064 vdd.n1328 vss 0.00413f
C2065 vdd.n1329 vss 0.0471f
C2066 vdd.n1330 vss 0.0471f
C2067 vdd.n1331 vss 0.00324f
C2068 vdd.n1332 vss 0.00413f
C2069 vdd.n1333 vss 0.00413f
C2070 vdd.n1334 vss 0.00679f
C2071 vdd.n1335 vss 0.00413f
C2072 vdd.n1336 vss 0.0471f
C2073 vdd.n1337 vss 0.00324f
C2074 vdd.n1338 vss 0.0424f
C2075 vdd.n1339 vss 0.00324f
C2076 vdd.n1340 vss 0.0128f
C2077 vdd.n1341 vss 0.02f
C2078 vdd.n1342 vss 0.0132f
C2079 vdd.n1343 vss 0.00925f
C2080 vdd.n1344 vss 0.00425f
C2081 vdd.n1346 vss 0.0471f
C2082 vdd.n1347 vss 0.00425f
C2083 vdd.n1348 vss 0.00413f
C2084 vdd.n1349 vss 0.00251f
C2085 vdd.n1350 vss 0.0471f
C2086 vdd.n1351 vss 0.00251f
C2087 vdd.n1352 vss 0.00517f
C2088 vdd.n1353 vss 0.00679f
C2089 vdd.n1354 vss 0.00324f
C2090 vdd.n1355 vss 0.00324f
C2091 vdd.n1356 vss 0.0132f
C2092 vdd.n1357 vss 0.0424f
C2093 vdd.n1358 vss 0.02f
C2094 vdd.n1359 vss 0.00425f
C2095 vdd.n1361 vss 0.0471f
C2096 vdd.n1362 vss 0.00425f
C2097 vdd.n1363 vss 0.00925f
C2098 vdd.n1364 vss 0.00679f
C2099 vdd.n1365 vss 0.00517f
C2100 vdd.n1366 vss 0.00251f
C2101 vdd.n1367 vss 0.0471f
C2102 vdd.n1368 vss 0.00251f
C2103 vdd.n1369 vss 0.0112f
C2104 vdd.n1370 vss 0.0128f
C2105 vdd.n1371 vss 0.0613f
C2106 vdd.n1372 vss 0.00324f
C2107 vdd.n1373 vss 0.0112f
C2108 vdd.n1374 vss 0.0128f
C2109 vdd.n1375 vss 0.00413f
C2110 vdd.n1376 vss 0.00413f
C2111 vdd.n1377 vss 0.0471f
C2112 vdd.n1378 vss 0.0471f
C2113 vdd.n1379 vss 0.00324f
C2114 vdd.n1380 vss 0.00413f
C2115 vdd.n1381 vss 0.00413f
C2116 vdd.n1382 vss 0.00679f
C2117 vdd.n1383 vss 0.00413f
C2118 vdd.n1384 vss 0.0471f
C2119 vdd.n1385 vss 0.00324f
C2120 vdd.n1386 vss 0.0424f
C2121 vdd.n1387 vss 0.00324f
C2122 vdd.n1388 vss 0.0128f
C2123 vdd.n1389 vss 0.02f
C2124 vdd.n1390 vss 0.0132f
C2125 vdd.n1391 vss 0.00925f
C2126 vdd.n1392 vss 0.00425f
C2127 vdd.n1394 vss 0.0471f
C2128 vdd.n1395 vss 0.00425f
C2129 vdd.n1396 vss 0.00413f
C2130 vdd.n1397 vss 0.00251f
C2131 vdd.n1398 vss 0.0471f
C2132 vdd.n1399 vss 0.00251f
C2133 vdd.n1400 vss 0.00517f
C2134 vdd.n1401 vss 0.00679f
C2135 vdd.n1402 vss 0.00324f
C2136 vdd.n1403 vss 0.00324f
C2137 vdd.n1404 vss 0.0132f
C2138 vdd.n1405 vss 0.0424f
C2139 vdd.n1406 vss 0.02f
C2140 vdd.n1407 vss 0.00425f
C2141 vdd.n1409 vss 0.0471f
C2142 vdd.n1410 vss 0.00425f
C2143 vdd.n1411 vss 0.00925f
C2144 vdd.n1412 vss 0.00679f
C2145 vdd.n1413 vss 0.00517f
C2146 vdd.n1414 vss 0.00251f
C2147 vdd.n1415 vss 0.0471f
C2148 vdd.n1416 vss 0.00251f
C2149 vdd.n1417 vss 0.0112f
C2150 vdd.n1418 vss 0.0128f
C2151 vdd.n1419 vss 0.0666f
C2152 vdd.n1420 vss 0.00324f
C2153 vdd.n1421 vss 0.0112f
C2154 vdd.n1422 vss 0.0128f
C2155 vdd.n1423 vss 0.00413f
C2156 vdd.n1424 vss 0.00413f
C2157 vdd.n1425 vss 0.0471f
C2158 vdd.n1426 vss 0.0471f
C2159 vdd.n1427 vss 0.00324f
C2160 vdd.n1428 vss 0.00413f
C2161 vdd.n1429 vss 0.00413f
C2162 vdd.n1430 vss 0.00679f
C2163 vdd.n1431 vss 0.00413f
C2164 vdd.n1432 vss 0.0471f
C2165 vdd.n1433 vss 0.00324f
C2166 vdd.n1434 vss 0.0424f
C2167 vdd.n1435 vss 0.00324f
C2168 vdd.n1436 vss 0.0128f
C2169 vdd.n1437 vss 0.02f
C2170 vdd.n1438 vss 0.0132f
C2171 vdd.n1439 vss 0.00925f
C2172 vdd.n1440 vss 0.00425f
C2173 vdd.n1442 vss 0.0471f
C2174 vdd.n1443 vss 0.00425f
C2175 vdd.n1444 vss 0.00413f
C2176 vdd.n1445 vss 0.00251f
C2177 vdd.n1446 vss 0.0471f
C2178 vdd.n1447 vss 0.00251f
C2179 vdd.n1448 vss 0.00517f
C2180 vdd.n1449 vss 0.00679f
C2181 vdd.n1450 vss 0.00324f
C2182 vdd.n1451 vss 0.00324f
C2183 vdd.n1452 vss 0.0132f
C2184 vdd.n1453 vss 0.0424f
C2185 vdd.n1454 vss 0.02f
C2186 vdd.n1455 vss 0.00425f
C2187 vdd.n1457 vss 0.0471f
C2188 vdd.n1458 vss 0.00425f
C2189 vdd.n1459 vss 0.00925f
C2190 vdd.n1460 vss 0.00679f
C2191 vdd.n1461 vss 0.00517f
C2192 vdd.n1462 vss 0.00251f
C2193 vdd.n1463 vss 0.0471f
C2194 vdd.n1464 vss 0.00251f
C2195 vdd.n1465 vss 0.0112f
C2196 vdd.n1466 vss 0.0128f
C2197 vdd.n1467 vss 0.0617f
C2198 vdd.n1468 vss 0.00335f
C2199 vdd.n1469 vss 0.0855f
C2200 vdd.n1470 vss 0.0107f
C2201 vdd.n1471 vss 0.0128f
C2202 vdd.n1472 vss 0.0424f
C2203 vdd.n1473 vss 0.00413f
C2204 vdd.n1474 vss 0.0471f
C2205 vdd.n1475 vss 0.00413f
C2206 vdd.n1476 vss 0.00324f
C2207 vdd.n1477 vss 0.00324f
C2208 vdd.n1478 vss 0.00679f
C2209 vdd.n1479 vss 0.00413f
C2210 vdd.n1480 vss 0.0471f
C2211 vdd.n1481 vss 0.00413f
C2212 vdd.n1482 vss 0.0105f
C2213 vdd.n1483 vss 0.0471f
C2214 vdd.n1484 vss 0.00413f
C2215 vdd.n1485 vss 0.00324f
C2216 vdd.n1486 vss 0.00324f
C2217 vdd.n1487 vss 0.0132f
C2218 vdd.n1488 vss 0.0424f
C2219 vdd.n1489 vss 0.0128f
C2220 vdd.n1490 vss 0.02f
C2221 vdd.n1491 vss 0.00425f
C2222 vdd.n1493 vss 0.0471f
C2223 vdd.n1494 vss 0.00425f
C2224 vdd.n1495 vss 0.00925f
C2225 vdd.n1496 vss 0.00679f
C2226 vdd.n1497 vss 0.00517f
C2227 vdd.n1498 vss 0.00251f
C2228 vdd.n1499 vss 0.0471f
C2229 vdd.n1500 vss 0.00251f
C2230 vdd.n1501 vss 0.00413f
C2231 vdd.n1502 vss 0.00324f
C2232 vdd.n1503 vss 0.00324f
C2233 vdd.n1504 vss 0.00805f
C2234 vdd.n1505 vss 0.0112f
C2235 vdd.n1506 vss 0.00251f
C2236 vdd.n1507 vss 0.0471f
C2237 vdd.n1508 vss 0.00251f
C2238 vdd.n1509 vss 0.00517f
C2239 vdd.n1510 vss 0.00679f
C2240 vdd.n1511 vss 0.00925f
C2241 vdd.n1512 vss 0.00425f
C2242 vdd.n1514 vss 0.0471f
C2243 vdd.n1515 vss 0.00425f
C2244 vdd.n1516 vss 0.00991f
C2245 vdd.n1517 vss 0.0126f
C2246 vdd.n1518 vss 0.0516f
C2247 vdd.n1519 vss 0.0011f
C2248 vdd.n1520 vss 0.0271f
C2249 vdd.n1521 vss 0.00324f
C2250 vdd.n1522 vss 0.0112f
C2251 vdd.n1523 vss 0.0128f
C2252 vdd.n1524 vss 0.00413f
C2253 vdd.n1525 vss 0.00413f
C2254 vdd.n1526 vss 0.0471f
C2255 vdd.n1527 vss 0.0471f
C2256 vdd.n1528 vss 0.00324f
C2257 vdd.n1529 vss 0.00413f
C2258 vdd.n1530 vss 0.00413f
C2259 vdd.n1531 vss 0.00679f
C2260 vdd.n1532 vss 0.00413f
C2261 vdd.n1533 vss 0.0471f
C2262 vdd.n1534 vss 0.00324f
C2263 vdd.n1535 vss 0.0424f
C2264 vdd.n1536 vss 0.00324f
C2265 vdd.n1537 vss 0.0128f
C2266 vdd.n1538 vss 0.02f
C2267 vdd.n1539 vss 0.0132f
C2268 vdd.n1540 vss 0.00925f
C2269 vdd.n1541 vss 0.00425f
C2270 vdd.n1543 vss 0.0471f
C2271 vdd.n1544 vss 0.00425f
C2272 vdd.n1545 vss 0.00413f
C2273 vdd.n1546 vss 0.00251f
C2274 vdd.n1547 vss 0.0471f
C2275 vdd.n1548 vss 0.00251f
C2276 vdd.n1549 vss 0.00517f
C2277 vdd.n1550 vss 0.00679f
C2278 vdd.n1551 vss 0.00324f
C2279 vdd.n1552 vss 0.00324f
C2280 vdd.n1553 vss 0.0132f
C2281 vdd.n1554 vss 0.0424f
C2282 vdd.n1555 vss 0.02f
C2283 vdd.n1556 vss 0.00425f
C2284 vdd.n1558 vss 0.0471f
C2285 vdd.n1559 vss 0.00425f
C2286 vdd.n1560 vss 0.00925f
C2287 vdd.n1561 vss 0.00679f
C2288 vdd.n1562 vss 0.00517f
C2289 vdd.n1563 vss 0.00251f
C2290 vdd.n1564 vss 0.0471f
C2291 vdd.n1565 vss 0.00251f
C2292 vdd.n1566 vss 0.0112f
C2293 vdd.n1567 vss 0.0128f
C2294 vdd.n1568 vss 0.0666f
C2295 vdd.n1569 vss 0.00324f
C2296 vdd.n1570 vss 0.0112f
C2297 vdd.n1571 vss 0.0128f
C2298 vdd.n1572 vss 0.00413f
C2299 vdd.n1573 vss 0.00413f
C2300 vdd.n1574 vss 0.0471f
C2301 vdd.n1575 vss 0.0471f
C2302 vdd.n1576 vss 0.00324f
C2303 vdd.n1577 vss 0.00413f
C2304 vdd.n1578 vss 0.00413f
C2305 vdd.n1579 vss 0.00679f
C2306 vdd.n1580 vss 0.00413f
C2307 vdd.n1581 vss 0.0471f
C2308 vdd.n1582 vss 0.00324f
C2309 vdd.n1583 vss 0.0424f
C2310 vdd.n1584 vss 0.00324f
C2311 vdd.n1585 vss 0.0128f
C2312 vdd.n1586 vss 0.02f
C2313 vdd.n1587 vss 0.0132f
C2314 vdd.n1588 vss 0.00925f
C2315 vdd.n1589 vss 0.00425f
C2316 vdd.n1591 vss 0.0471f
C2317 vdd.n1592 vss 0.00425f
C2318 vdd.n1593 vss 0.00413f
C2319 vdd.n1594 vss 0.00251f
C2320 vdd.n1595 vss 0.0471f
C2321 vdd.n1596 vss 0.00251f
C2322 vdd.n1597 vss 0.00517f
C2323 vdd.n1598 vss 0.00679f
C2324 vdd.n1599 vss 0.00324f
C2325 vdd.n1600 vss 0.00324f
C2326 vdd.n1601 vss 0.0132f
C2327 vdd.n1602 vss 0.0424f
C2328 vdd.n1603 vss 0.02f
C2329 vdd.n1604 vss 0.00425f
C2330 vdd.n1606 vss 0.0471f
C2331 vdd.n1607 vss 0.00425f
C2332 vdd.n1608 vss 0.00925f
C2333 vdd.n1609 vss 0.00679f
C2334 vdd.n1610 vss 0.00517f
C2335 vdd.n1611 vss 0.00251f
C2336 vdd.n1612 vss 0.0471f
C2337 vdd.n1613 vss 0.00251f
C2338 vdd.n1614 vss 0.0112f
C2339 vdd.n1615 vss 0.0128f
C2340 vdd.n1616 vss 0.00324f
C2341 vdd.n1617 vss 0.0112f
C2342 vdd.n1618 vss 0.0128f
C2343 vdd.n1619 vss 0.00413f
C2344 vdd.n1620 vss 0.00413f
C2345 vdd.n1621 vss 0.0471f
C2346 vdd.n1622 vss 0.0471f
C2347 vdd.n1623 vss 0.00324f
C2348 vdd.n1624 vss 0.00413f
C2349 vdd.n1625 vss 0.00413f
C2350 vdd.n1626 vss 0.00679f
C2351 vdd.n1627 vss 0.00413f
C2352 vdd.n1628 vss 0.0471f
C2353 vdd.n1629 vss 0.00324f
C2354 vdd.n1630 vss 0.0424f
C2355 vdd.n1631 vss 0.00324f
C2356 vdd.n1632 vss 0.0128f
C2357 vdd.n1633 vss 0.02f
C2358 vdd.n1634 vss 0.0132f
C2359 vdd.n1635 vss 0.00925f
C2360 vdd.n1636 vss 0.00425f
C2361 vdd.n1638 vss 0.0471f
C2362 vdd.n1639 vss 0.00425f
C2363 vdd.n1640 vss 0.00413f
C2364 vdd.n1641 vss 0.00251f
C2365 vdd.n1642 vss 0.0471f
C2366 vdd.n1643 vss 0.00251f
C2367 vdd.n1644 vss 0.00517f
C2368 vdd.n1645 vss 0.00679f
C2369 vdd.n1646 vss 0.00324f
C2370 vdd.n1647 vss 0.00324f
C2371 vdd.n1648 vss 0.0132f
C2372 vdd.n1649 vss 0.0424f
C2373 vdd.n1650 vss 0.02f
C2374 vdd.n1651 vss 0.00425f
C2375 vdd.n1653 vss 0.0471f
C2376 vdd.n1654 vss 0.00425f
C2377 vdd.n1655 vss 0.00925f
C2378 vdd.n1656 vss 0.00679f
C2379 vdd.n1657 vss 0.00517f
C2380 vdd.n1658 vss 0.00251f
C2381 vdd.n1659 vss 0.0471f
C2382 vdd.n1660 vss 0.00251f
C2383 vdd.n1661 vss 0.0112f
C2384 vdd.n1662 vss 0.0128f
C2385 vdd.n1663 vss 0.144f
C2386 vdd.n1664 vss 0.143f
C2387 vdd.n1665 vss 0.0608f
C2388 vdd.n1666 vss 0.00324f
C2389 vdd.n1667 vss 0.0112f
C2390 vdd.n1668 vss 0.0128f
C2391 vdd.n1669 vss 0.00413f
C2392 vdd.n1670 vss 0.00413f
C2393 vdd.n1671 vss 0.0471f
C2394 vdd.n1672 vss 0.0471f
C2395 vdd.n1673 vss 0.00324f
C2396 vdd.n1674 vss 0.00413f
C2397 vdd.n1675 vss 0.00413f
C2398 vdd.n1676 vss 0.00679f
C2399 vdd.n1677 vss 0.00413f
C2400 vdd.n1678 vss 0.0471f
C2401 vdd.n1679 vss 0.00324f
C2402 vdd.n1680 vss 0.0424f
C2403 vdd.n1681 vss 0.00324f
C2404 vdd.n1682 vss 0.0128f
C2405 vdd.n1683 vss 0.02f
C2406 vdd.n1684 vss 0.0132f
C2407 vdd.n1685 vss 0.00925f
C2408 vdd.n1686 vss 0.00425f
C2409 vdd.n1688 vss 0.0471f
C2410 vdd.n1689 vss 0.00425f
C2411 vdd.n1690 vss 0.00413f
C2412 vdd.n1691 vss 0.00251f
C2413 vdd.n1692 vss 0.0471f
C2414 vdd.n1693 vss 0.00251f
C2415 vdd.n1694 vss 0.00517f
C2416 vdd.n1695 vss 0.00679f
C2417 vdd.n1696 vss 0.00324f
C2418 vdd.n1697 vss 0.00324f
C2419 vdd.n1698 vss 0.0132f
C2420 vdd.n1699 vss 0.0424f
C2421 vdd.n1700 vss 0.02f
C2422 vdd.n1701 vss 0.00425f
C2423 vdd.n1703 vss 0.0471f
C2424 vdd.n1704 vss 0.00425f
C2425 vdd.n1705 vss 0.00925f
C2426 vdd.n1706 vss 0.00679f
C2427 vdd.n1707 vss 0.00517f
C2428 vdd.n1708 vss 0.00251f
C2429 vdd.n1709 vss 0.0471f
C2430 vdd.n1710 vss 0.00251f
C2431 vdd.n1711 vss 0.0112f
C2432 vdd.n1712 vss 0.0128f
C2433 vdd.n1713 vss 0.0666f
C2434 vdd.n1714 vss 0.118f
C2435 vdd.n1715 vss 0.121f
C2436 vdd.n1716 vss 0.00324f
C2437 vdd.n1717 vss 0.0112f
C2438 vdd.n1718 vss 0.0128f
C2439 vdd.n1719 vss 0.00413f
C2440 vdd.n1720 vss 0.00413f
C2441 vdd.n1721 vss 0.0471f
C2442 vdd.n1722 vss 0.0471f
C2443 vdd.n1723 vss 0.00324f
C2444 vdd.n1724 vss 0.00413f
C2445 vdd.n1725 vss 0.00413f
C2446 vdd.n1726 vss 0.00679f
C2447 vdd.n1727 vss 0.00413f
C2448 vdd.n1728 vss 0.0471f
C2449 vdd.n1729 vss 0.00324f
C2450 vdd.n1730 vss 0.0424f
C2451 vdd.n1731 vss 0.00324f
C2452 vdd.n1732 vss 0.0128f
C2453 vdd.n1733 vss 0.02f
C2454 vdd.n1734 vss 0.0132f
C2455 vdd.n1735 vss 0.00925f
C2456 vdd.n1736 vss 0.00425f
C2457 vdd.n1738 vss 0.0471f
C2458 vdd.n1739 vss 0.00425f
C2459 vdd.n1740 vss 0.00413f
C2460 vdd.n1741 vss 0.00251f
C2461 vdd.n1742 vss 0.0471f
C2462 vdd.n1743 vss 0.00251f
C2463 vdd.n1744 vss 0.00517f
C2464 vdd.n1745 vss 0.00679f
C2465 vdd.n1746 vss 0.00324f
C2466 vdd.n1747 vss 0.00324f
C2467 vdd.n1748 vss 0.0132f
C2468 vdd.n1749 vss 0.0424f
C2469 vdd.n1750 vss 0.02f
C2470 vdd.n1751 vss 0.00425f
C2471 vdd.n1753 vss 0.0471f
C2472 vdd.n1754 vss 0.00425f
C2473 vdd.n1755 vss 0.00925f
C2474 vdd.n1756 vss 0.00679f
C2475 vdd.n1757 vss 0.00517f
C2476 vdd.n1758 vss 0.00251f
C2477 vdd.n1759 vss 0.0471f
C2478 vdd.n1760 vss 0.00251f
C2479 vdd.n1761 vss 0.0112f
C2480 vdd.n1762 vss 0.0955f
C2481 vdd.n1763 vss 0.0608f
C2482 vdd.n1764 vss 0.00324f
C2483 vdd.n1765 vss 0.0112f
C2484 vdd.n1766 vss 0.0128f
C2485 vdd.n1767 vss 0.00413f
C2486 vdd.n1768 vss 0.00413f
C2487 vdd.n1769 vss 0.0471f
C2488 vdd.n1770 vss 0.0471f
C2489 vdd.n1771 vss 0.00324f
C2490 vdd.n1772 vss 0.00413f
C2491 vdd.n1773 vss 0.00413f
C2492 vdd.n1774 vss 0.00679f
C2493 vdd.n1775 vss 0.00413f
C2494 vdd.n1776 vss 0.0471f
C2495 vdd.n1777 vss 0.00324f
C2496 vdd.n1778 vss 0.0424f
C2497 vdd.n1779 vss 0.00324f
C2498 vdd.n1780 vss 0.0128f
C2499 vdd.n1781 vss 0.02f
C2500 vdd.n1782 vss 0.0132f
C2501 vdd.n1783 vss 0.00925f
C2502 vdd.n1784 vss 0.00425f
C2503 vdd.n1786 vss 0.0471f
C2504 vdd.n1787 vss 0.00425f
C2505 vdd.n1788 vss 0.00413f
C2506 vdd.n1789 vss 0.00251f
C2507 vdd.n1790 vss 0.0471f
C2508 vdd.n1791 vss 0.00251f
C2509 vdd.n1792 vss 0.00517f
C2510 vdd.n1793 vss 0.00679f
C2511 vdd.n1794 vss 0.00324f
C2512 vdd.n1795 vss 0.00324f
C2513 vdd.n1796 vss 0.0132f
C2514 vdd.n1797 vss 0.0424f
C2515 vdd.n1798 vss 0.02f
C2516 vdd.n1799 vss 0.00425f
C2517 vdd.n1801 vss 0.0471f
C2518 vdd.n1802 vss 0.00425f
C2519 vdd.n1803 vss 0.00925f
C2520 vdd.n1804 vss 0.00679f
C2521 vdd.n1805 vss 0.00517f
C2522 vdd.n1806 vss 0.00251f
C2523 vdd.n1807 vss 0.0471f
C2524 vdd.n1808 vss 0.00251f
C2525 vdd.n1809 vss 0.0112f
C2526 vdd.n1810 vss 0.0128f
C2527 vdd.n1811 vss 0.0666f
C2528 vdd.n1812 vss 0.0912f
C2529 vdd.n1813 vss 0.0824f
C2530 vdd.n1814 vss 0.0567f
C2531 vdd.n1815 vss 0.00324f
C2532 vdd.n1816 vss 0.0112f
C2533 vdd.n1817 vss 0.0128f
C2534 vdd.n1818 vss 0.00413f
C2535 vdd.n1819 vss 0.00413f
C2536 vdd.n1820 vss 0.0471f
C2537 vdd.n1821 vss 0.0471f
C2538 vdd.n1822 vss 0.00324f
C2539 vdd.n1823 vss 0.00413f
C2540 vdd.n1824 vss 0.00413f
C2541 vdd.n1825 vss 0.00679f
C2542 vdd.n1826 vss 0.00413f
C2543 vdd.n1827 vss 0.0471f
C2544 vdd.n1828 vss 0.00324f
C2545 vdd.n1829 vss 0.0424f
C2546 vdd.n1830 vss 0.00324f
C2547 vdd.n1831 vss 0.0128f
C2548 vdd.n1832 vss 0.02f
C2549 vdd.n1833 vss 0.0132f
C2550 vdd.n1834 vss 0.00925f
C2551 vdd.n1835 vss 0.00425f
C2552 vdd.n1837 vss 0.0471f
C2553 vdd.n1838 vss 0.00425f
C2554 vdd.n1839 vss 0.00413f
C2555 vdd.n1840 vss 0.00251f
C2556 vdd.n1841 vss 0.0471f
C2557 vdd.n1842 vss 0.00251f
C2558 vdd.n1843 vss 0.00517f
C2559 vdd.n1844 vss 0.00679f
C2560 vdd.n1845 vss 0.00324f
C2561 vdd.n1846 vss 0.00324f
C2562 vdd.n1847 vss 0.0132f
C2563 vdd.n1848 vss 0.0424f
C2564 vdd.n1849 vss 0.02f
C2565 vdd.n1850 vss 0.00425f
C2566 vdd.n1852 vss 0.0471f
C2567 vdd.n1853 vss 0.00425f
C2568 vdd.n1854 vss 0.00925f
C2569 vdd.n1855 vss 0.00679f
C2570 vdd.n1856 vss 0.00517f
C2571 vdd.n1857 vss 0.00251f
C2572 vdd.n1858 vss 0.0471f
C2573 vdd.n1859 vss 0.00251f
C2574 vdd.n1860 vss 0.0112f
C2575 vdd.n1861 vss 0.0128f
C2576 vdd.n1862 vss 0.00324f
C2577 vdd.n1863 vss 0.0112f
C2578 vdd.n1864 vss 0.0128f
C2579 vdd.n1865 vss 0.00413f
C2580 vdd.n1866 vss 0.00413f
C2581 vdd.n1867 vss 0.0471f
C2582 vdd.n1868 vss 0.0471f
C2583 vdd.n1869 vss 0.00324f
C2584 vdd.n1870 vss 0.00413f
C2585 vdd.n1871 vss 0.00413f
C2586 vdd.n1872 vss 0.00679f
C2587 vdd.n1873 vss 0.00413f
C2588 vdd.n1874 vss 0.0471f
C2589 vdd.n1875 vss 0.00324f
C2590 vdd.n1876 vss 0.0424f
C2591 vdd.n1877 vss 0.00324f
C2592 vdd.n1878 vss 0.0128f
C2593 vdd.n1879 vss 0.02f
C2594 vdd.n1880 vss 0.0132f
C2595 vdd.n1881 vss 0.00925f
C2596 vdd.n1882 vss 0.00425f
C2597 vdd.n1884 vss 0.0471f
C2598 vdd.n1885 vss 0.00425f
C2599 vdd.n1886 vss 0.00413f
C2600 vdd.n1887 vss 0.00251f
C2601 vdd.n1888 vss 0.0471f
C2602 vdd.n1889 vss 0.00251f
C2603 vdd.n1890 vss 0.00517f
C2604 vdd.n1891 vss 0.00679f
C2605 vdd.n1892 vss 0.00324f
C2606 vdd.n1893 vss 0.00324f
C2607 vdd.n1894 vss 0.0132f
C2608 vdd.n1895 vss 0.0424f
C2609 vdd.n1896 vss 0.02f
C2610 vdd.n1897 vss 0.00425f
C2611 vdd.n1899 vss 0.0471f
C2612 vdd.n1900 vss 0.00425f
C2613 vdd.n1901 vss 0.00925f
C2614 vdd.n1902 vss 0.00679f
C2615 vdd.n1903 vss 0.00517f
C2616 vdd.n1904 vss 0.00251f
C2617 vdd.n1905 vss 0.0471f
C2618 vdd.n1906 vss 0.00251f
C2619 vdd.n1907 vss 0.0112f
C2620 vdd.n1908 vss 0.0128f
C2621 vdd.n1909 vss 0.0564f
C2622 vdd.n1910 vss 0.00324f
C2623 vdd.n1911 vss 0.0112f
C2624 vdd.n1912 vss 0.0128f
C2625 vdd.n1913 vss 0.00413f
C2626 vdd.n1914 vss 0.00413f
C2627 vdd.n1915 vss 0.0471f
C2628 vdd.n1916 vss 0.0471f
C2629 vdd.n1917 vss 0.00324f
C2630 vdd.n1918 vss 0.00413f
C2631 vdd.n1919 vss 0.00413f
C2632 vdd.n1920 vss 0.00679f
C2633 vdd.n1921 vss 0.00413f
C2634 vdd.n1922 vss 0.0471f
C2635 vdd.n1923 vss 0.00324f
C2636 vdd.n1924 vss 0.0424f
C2637 vdd.n1925 vss 0.00324f
C2638 vdd.n1926 vss 0.0128f
C2639 vdd.n1927 vss 0.02f
C2640 vdd.n1928 vss 0.0132f
C2641 vdd.n1929 vss 0.00925f
C2642 vdd.n1930 vss 0.00425f
C2643 vdd.n1932 vss 0.0471f
C2644 vdd.n1933 vss 0.00425f
C2645 vdd.n1934 vss 0.00413f
C2646 vdd.n1935 vss 0.00251f
C2647 vdd.n1936 vss 0.0471f
C2648 vdd.n1937 vss 0.00251f
C2649 vdd.n1938 vss 0.00517f
C2650 vdd.n1939 vss 0.00679f
C2651 vdd.n1940 vss 0.00324f
C2652 vdd.n1941 vss 0.00324f
C2653 vdd.n1942 vss 0.0132f
C2654 vdd.n1943 vss 0.0424f
C2655 vdd.n1944 vss 0.02f
C2656 vdd.n1945 vss 0.00425f
C2657 vdd.n1947 vss 0.0471f
C2658 vdd.n1948 vss 0.00425f
C2659 vdd.n1949 vss 0.00925f
C2660 vdd.n1950 vss 0.00679f
C2661 vdd.n1951 vss 0.00517f
C2662 vdd.n1952 vss 0.00251f
C2663 vdd.n1953 vss 0.0471f
C2664 vdd.n1954 vss 0.00251f
C2665 vdd.n1955 vss 0.0112f
C2666 vdd.n1956 vss 0.0128f
C2667 vdd.n1957 vss 0.183f
C2668 vdd.n1958 vss 0.256f
C2669 vdd.n1959 vss 0.12f
C2670 vdd.n1960 vss 0.0608f
C2671 vdd.n1961 vss 0.00324f
C2672 vdd.n1962 vss 0.0112f
C2673 vdd.n1963 vss 0.0128f
C2674 vdd.n1964 vss 0.00413f
C2675 vdd.n1965 vss 0.00413f
C2676 vdd.n1966 vss 0.0471f
C2677 vdd.n1967 vss 0.0471f
C2678 vdd.n1968 vss 0.00324f
C2679 vdd.n1969 vss 0.00413f
C2680 vdd.n1970 vss 0.00413f
C2681 vdd.n1971 vss 0.00679f
C2682 vdd.n1972 vss 0.00413f
C2683 vdd.n1973 vss 0.0471f
C2684 vdd.n1974 vss 0.00324f
C2685 vdd.n1975 vss 0.0424f
C2686 vdd.n1976 vss 0.00324f
C2687 vdd.n1977 vss 0.0128f
C2688 vdd.n1978 vss 0.02f
C2689 vdd.n1979 vss 0.0132f
C2690 vdd.n1980 vss 0.00925f
C2691 vdd.n1981 vss 0.00425f
C2692 vdd.n1983 vss 0.0471f
C2693 vdd.n1984 vss 0.00425f
C2694 vdd.n1985 vss 0.00413f
C2695 vdd.n1986 vss 0.00251f
C2696 vdd.n1987 vss 0.0471f
C2697 vdd.n1988 vss 0.00251f
C2698 vdd.n1989 vss 0.00517f
C2699 vdd.n1990 vss 0.00679f
C2700 vdd.n1991 vss 0.00324f
C2701 vdd.n1992 vss 0.00324f
C2702 vdd.n1993 vss 0.0132f
C2703 vdd.n1994 vss 0.0424f
C2704 vdd.n1995 vss 0.02f
C2705 vdd.n1996 vss 0.00425f
C2706 vdd.n1998 vss 0.0471f
C2707 vdd.n1999 vss 0.00425f
C2708 vdd.n2000 vss 0.00925f
C2709 vdd.n2001 vss 0.00679f
C2710 vdd.n2002 vss 0.00517f
C2711 vdd.n2003 vss 0.00251f
C2712 vdd.n2004 vss 0.0471f
C2713 vdd.n2005 vss 0.00251f
C2714 vdd.n2006 vss 0.0112f
C2715 vdd.n2007 vss 0.0128f
C2716 vdd.n2008 vss 0.0666f
C2717 vdd.n2009 vss 0.118f
C2718 vdd.n2010 vss 0.121f
C2719 vdd.n2011 vss 0.00324f
C2720 vdd.n2012 vss 0.0112f
C2721 vdd.n2013 vss 0.0128f
C2722 vdd.n2014 vss 0.00413f
C2723 vdd.n2015 vss 0.00413f
C2724 vdd.n2016 vss 0.0471f
C2725 vdd.n2017 vss 0.0471f
C2726 vdd.n2018 vss 0.00324f
C2727 vdd.n2019 vss 0.00413f
C2728 vdd.n2020 vss 0.00413f
C2729 vdd.n2021 vss 0.00679f
C2730 vdd.n2022 vss 0.00413f
C2731 vdd.n2023 vss 0.0471f
C2732 vdd.n2024 vss 0.00324f
C2733 vdd.n2025 vss 0.0424f
C2734 vdd.n2026 vss 0.00324f
C2735 vdd.n2027 vss 0.0128f
C2736 vdd.n2028 vss 0.02f
C2737 vdd.n2029 vss 0.0132f
C2738 vdd.n2030 vss 0.00925f
C2739 vdd.n2031 vss 0.00425f
C2740 vdd.n2033 vss 0.0471f
C2741 vdd.n2034 vss 0.00425f
C2742 vdd.n2035 vss 0.00413f
C2743 vdd.n2036 vss 0.00251f
C2744 vdd.n2037 vss 0.0471f
C2745 vdd.n2038 vss 0.00251f
C2746 vdd.n2039 vss 0.00517f
C2747 vdd.n2040 vss 0.00679f
C2748 vdd.n2041 vss 0.00324f
C2749 vdd.n2042 vss 0.00324f
C2750 vdd.n2043 vss 0.0132f
C2751 vdd.n2044 vss 0.0424f
C2752 vdd.n2045 vss 0.02f
C2753 vdd.n2046 vss 0.00425f
C2754 vdd.n2048 vss 0.0471f
C2755 vdd.n2049 vss 0.00425f
C2756 vdd.n2050 vss 0.00925f
C2757 vdd.n2051 vss 0.00679f
C2758 vdd.n2052 vss 0.00517f
C2759 vdd.n2053 vss 0.00251f
C2760 vdd.n2054 vss 0.0471f
C2761 vdd.n2055 vss 0.00251f
C2762 vdd.n2056 vss 0.0112f
C2763 vdd.n2057 vss 0.0955f
C2764 vdd.n2058 vss 0.0608f
C2765 vdd.n2059 vss 0.00324f
C2766 vdd.n2060 vss 0.0112f
C2767 vdd.n2061 vss 0.0128f
C2768 vdd.n2062 vss 0.00413f
C2769 vdd.n2063 vss 0.00413f
C2770 vdd.n2064 vss 0.0471f
C2771 vdd.n2065 vss 0.0471f
C2772 vdd.n2066 vss 0.00324f
C2773 vdd.n2067 vss 0.00413f
C2774 vdd.n2068 vss 0.00413f
C2775 vdd.n2069 vss 0.00679f
C2776 vdd.n2070 vss 0.00413f
C2777 vdd.n2071 vss 0.0471f
C2778 vdd.n2072 vss 0.00324f
C2779 vdd.n2073 vss 0.0424f
C2780 vdd.n2074 vss 0.00324f
C2781 vdd.n2075 vss 0.0128f
C2782 vdd.n2076 vss 0.02f
C2783 vdd.n2077 vss 0.0132f
C2784 vdd.n2078 vss 0.00925f
C2785 vdd.n2079 vss 0.00425f
C2786 vdd.n2081 vss 0.0471f
C2787 vdd.n2082 vss 0.00425f
C2788 vdd.n2083 vss 0.00413f
C2789 vdd.n2084 vss 0.00251f
C2790 vdd.n2085 vss 0.0471f
C2791 vdd.n2086 vss 0.00251f
C2792 vdd.n2087 vss 0.00517f
C2793 vdd.n2088 vss 0.00679f
C2794 vdd.n2089 vss 0.00324f
C2795 vdd.n2090 vss 0.00324f
C2796 vdd.n2091 vss 0.0132f
C2797 vdd.n2092 vss 0.0424f
C2798 vdd.n2093 vss 0.02f
C2799 vdd.n2094 vss 0.00425f
C2800 vdd.n2096 vss 0.0471f
C2801 vdd.n2097 vss 0.00425f
C2802 vdd.n2098 vss 0.00925f
C2803 vdd.n2099 vss 0.00679f
C2804 vdd.n2100 vss 0.00517f
C2805 vdd.n2101 vss 0.00251f
C2806 vdd.n2102 vss 0.0471f
C2807 vdd.n2103 vss 0.00251f
C2808 vdd.n2104 vss 0.0112f
C2809 vdd.n2105 vss 0.0128f
C2810 vdd.n2106 vss 0.0666f
C2811 vdd.n2107 vss 0.118f
C2812 vdd.n2108 vss 0.0935f
C2813 vdd.n2109 vss 0.00324f
C2814 vdd.n2110 vss 0.0112f
C2815 vdd.n2111 vss 0.0128f
C2816 vdd.n2112 vss 0.00413f
C2817 vdd.n2113 vss 0.00413f
C2818 vdd.n2114 vss 0.0471f
C2819 vdd.n2115 vss 0.0471f
C2820 vdd.n2116 vss 0.00324f
C2821 vdd.n2117 vss 0.00413f
C2822 vdd.n2118 vss 0.00413f
C2823 vdd.n2119 vss 0.00679f
C2824 vdd.n2120 vss 0.00413f
C2825 vdd.n2121 vss 0.0471f
C2826 vdd.n2122 vss 0.00324f
C2827 vdd.n2123 vss 0.0424f
C2828 vdd.n2124 vss 0.00324f
C2829 vdd.n2125 vss 0.0128f
C2830 vdd.n2126 vss 0.02f
C2831 vdd.n2127 vss 0.0132f
C2832 vdd.n2128 vss 0.00925f
C2833 vdd.n2129 vss 0.00425f
C2834 vdd.n2131 vss 0.0471f
C2835 vdd.n2132 vss 0.00425f
C2836 vdd.n2133 vss 0.00413f
C2837 vdd.n2134 vss 0.00251f
C2838 vdd.n2135 vss 0.0471f
C2839 vdd.n2136 vss 0.00251f
C2840 vdd.n2137 vss 0.00517f
C2841 vdd.n2138 vss 0.00679f
C2842 vdd.n2139 vss 0.00324f
C2843 vdd.n2140 vss 0.00324f
C2844 vdd.n2141 vss 0.0132f
C2845 vdd.n2142 vss 0.0424f
C2846 vdd.n2143 vss 0.02f
C2847 vdd.n2144 vss 0.00425f
C2848 vdd.n2146 vss 0.0471f
C2849 vdd.n2147 vss 0.00425f
C2850 vdd.n2148 vss 0.00925f
C2851 vdd.n2149 vss 0.00679f
C2852 vdd.n2150 vss 0.00517f
C2853 vdd.n2151 vss 0.00251f
C2854 vdd.n2152 vss 0.0471f
C2855 vdd.n2153 vss 0.00251f
C2856 vdd.n2154 vss 0.0112f
C2857 vdd.n2155 vss 0.0128f
C2858 vdd.n2156 vss 0.00324f
C2859 vdd.n2157 vss 0.0112f
C2860 vdd.n2158 vss 0.0128f
C2861 vdd.n2159 vss 0.00413f
C2862 vdd.n2160 vss 0.00413f
C2863 vdd.n2161 vss 0.0471f
C2864 vdd.n2162 vss 0.0471f
C2865 vdd.n2163 vss 0.00324f
C2866 vdd.n2164 vss 0.00413f
C2867 vdd.n2165 vss 0.00413f
C2868 vdd.n2166 vss 0.00679f
C2869 vdd.n2167 vss 0.00413f
C2870 vdd.n2168 vss 0.0471f
C2871 vdd.n2169 vss 0.00324f
C2872 vdd.n2170 vss 0.0424f
C2873 vdd.n2171 vss 0.00324f
C2874 vdd.n2172 vss 0.0128f
C2875 vdd.n2173 vss 0.02f
C2876 vdd.n2174 vss 0.0132f
C2877 vdd.n2175 vss 0.00925f
C2878 vdd.n2176 vss 0.00425f
C2879 vdd.n2178 vss 0.0471f
C2880 vdd.n2179 vss 0.00425f
C2881 vdd.n2180 vss 0.00413f
C2882 vdd.n2181 vss 0.00251f
C2883 vdd.n2182 vss 0.0471f
C2884 vdd.n2183 vss 0.00251f
C2885 vdd.n2184 vss 0.00517f
C2886 vdd.n2185 vss 0.00679f
C2887 vdd.n2186 vss 0.00324f
C2888 vdd.n2187 vss 0.00324f
C2889 vdd.n2188 vss 0.0132f
C2890 vdd.n2189 vss 0.0424f
C2891 vdd.n2190 vss 0.02f
C2892 vdd.n2191 vss 0.00425f
C2893 vdd.n2193 vss 0.0471f
C2894 vdd.n2194 vss 0.00425f
C2895 vdd.n2195 vss 0.00925f
C2896 vdd.n2196 vss 0.00679f
C2897 vdd.n2197 vss 0.00517f
C2898 vdd.n2198 vss 0.00251f
C2899 vdd.n2199 vss 0.0471f
C2900 vdd.n2200 vss 0.00251f
C2901 vdd.n2201 vss 0.0112f
C2902 vdd.n2202 vss 0.0128f
C2903 vdd.n2203 vss 0.144f
C2904 vdd.n2204 vss 0.143f
C2905 vdd.n2205 vss 0.0608f
C2906 vdd.n2206 vss 0.00324f
C2907 vdd.n2207 vss 0.0112f
C2908 vdd.n2208 vss 0.0128f
C2909 vdd.n2209 vss 0.00413f
C2910 vdd.n2210 vss 0.00413f
C2911 vdd.n2211 vss 0.0471f
C2912 vdd.n2212 vss 0.0471f
C2913 vdd.n2213 vss 0.00324f
C2914 vdd.n2214 vss 0.00413f
C2915 vdd.n2215 vss 0.00413f
C2916 vdd.n2216 vss 0.00679f
C2917 vdd.n2217 vss 0.00413f
C2918 vdd.n2218 vss 0.0471f
C2919 vdd.n2219 vss 0.00324f
C2920 vdd.n2220 vss 0.0424f
C2921 vdd.n2221 vss 0.00324f
C2922 vdd.n2222 vss 0.0128f
C2923 vdd.n2223 vss 0.02f
C2924 vdd.n2224 vss 0.0132f
C2925 vdd.n2225 vss 0.00925f
C2926 vdd.n2226 vss 0.00425f
C2927 vdd.n2228 vss 0.0471f
C2928 vdd.n2229 vss 0.00425f
C2929 vdd.n2230 vss 0.00413f
C2930 vdd.n2231 vss 0.00251f
C2931 vdd.n2232 vss 0.0471f
C2932 vdd.n2233 vss 0.00251f
C2933 vdd.n2234 vss 0.00517f
C2934 vdd.n2235 vss 0.00679f
C2935 vdd.n2236 vss 0.00324f
C2936 vdd.n2237 vss 0.00324f
C2937 vdd.n2238 vss 0.0132f
C2938 vdd.n2239 vss 0.0424f
C2939 vdd.n2240 vss 0.02f
C2940 vdd.n2241 vss 0.00425f
C2941 vdd.n2243 vss 0.0471f
C2942 vdd.n2244 vss 0.00425f
C2943 vdd.n2245 vss 0.00925f
C2944 vdd.n2246 vss 0.00679f
C2945 vdd.n2247 vss 0.00517f
C2946 vdd.n2248 vss 0.00251f
C2947 vdd.n2249 vss 0.0471f
C2948 vdd.n2250 vss 0.00251f
C2949 vdd.n2251 vss 0.0112f
C2950 vdd.n2252 vss 0.0128f
C2951 vdd.n2253 vss 0.0666f
C2952 vdd.n2254 vss 0.118f
C2953 vdd.n2255 vss 0.121f
C2954 vdd.n2256 vss 0.00324f
C2955 vdd.n2257 vss 0.0112f
C2956 vdd.n2258 vss 0.0128f
C2957 vdd.n2259 vss 0.00413f
C2958 vdd.n2260 vss 0.00413f
C2959 vdd.n2261 vss 0.0471f
C2960 vdd.n2262 vss 0.0471f
C2961 vdd.n2263 vss 0.00324f
C2962 vdd.n2264 vss 0.00413f
C2963 vdd.n2265 vss 0.00413f
C2964 vdd.n2266 vss 0.00679f
C2965 vdd.n2267 vss 0.00413f
C2966 vdd.n2268 vss 0.0471f
C2967 vdd.n2269 vss 0.00324f
C2968 vdd.n2270 vss 0.0424f
C2969 vdd.n2271 vss 0.00324f
C2970 vdd.n2272 vss 0.0128f
C2971 vdd.n2273 vss 0.02f
C2972 vdd.n2274 vss 0.0132f
C2973 vdd.n2275 vss 0.00925f
C2974 vdd.n2276 vss 0.00425f
C2975 vdd.n2278 vss 0.0471f
C2976 vdd.n2279 vss 0.00425f
C2977 vdd.n2280 vss 0.00413f
C2978 vdd.n2281 vss 0.00251f
C2979 vdd.n2282 vss 0.0471f
C2980 vdd.n2283 vss 0.00251f
C2981 vdd.n2284 vss 0.00517f
C2982 vdd.n2285 vss 0.00679f
C2983 vdd.n2286 vss 0.00324f
C2984 vdd.n2287 vss 0.00324f
C2985 vdd.n2288 vss 0.0132f
C2986 vdd.n2289 vss 0.0424f
C2987 vdd.n2290 vss 0.02f
C2988 vdd.n2291 vss 0.00425f
C2989 vdd.n2293 vss 0.0471f
C2990 vdd.n2294 vss 0.00425f
C2991 vdd.n2295 vss 0.00925f
C2992 vdd.n2296 vss 0.00679f
C2993 vdd.n2297 vss 0.00517f
C2994 vdd.n2298 vss 0.00251f
C2995 vdd.n2299 vss 0.0471f
C2996 vdd.n2300 vss 0.00251f
C2997 vdd.n2301 vss 0.0112f
C2998 vdd.n2302 vss 0.0955f
C2999 vdd.n2303 vss 0.0608f
C3000 vdd.n2304 vss 0.00324f
C3001 vdd.n2305 vss 0.0112f
C3002 vdd.n2306 vss 0.0128f
C3003 vdd.n2307 vss 0.00413f
C3004 vdd.n2308 vss 0.00413f
C3005 vdd.n2309 vss 0.0471f
C3006 vdd.n2310 vss 0.0471f
C3007 vdd.n2311 vss 0.00324f
C3008 vdd.n2312 vss 0.00413f
C3009 vdd.n2313 vss 0.00413f
C3010 vdd.n2314 vss 0.00679f
C3011 vdd.n2315 vss 0.00413f
C3012 vdd.n2316 vss 0.0471f
C3013 vdd.n2317 vss 0.00324f
C3014 vdd.n2318 vss 0.0424f
C3015 vdd.n2319 vss 0.00324f
C3016 vdd.n2320 vss 0.0128f
C3017 vdd.n2321 vss 0.02f
C3018 vdd.n2322 vss 0.0132f
C3019 vdd.n2323 vss 0.00925f
C3020 vdd.n2324 vss 0.00425f
C3021 vdd.n2326 vss 0.0471f
C3022 vdd.n2327 vss 0.00425f
C3023 vdd.n2328 vss 0.00413f
C3024 vdd.n2329 vss 0.00251f
C3025 vdd.n2330 vss 0.0471f
C3026 vdd.n2331 vss 0.00251f
C3027 vdd.n2332 vss 0.00517f
C3028 vdd.n2333 vss 0.00679f
C3029 vdd.n2334 vss 0.00324f
C3030 vdd.n2335 vss 0.00324f
C3031 vdd.n2336 vss 0.0132f
C3032 vdd.n2337 vss 0.0424f
C3033 vdd.n2338 vss 0.02f
C3034 vdd.n2339 vss 0.00425f
C3035 vdd.n2341 vss 0.0471f
C3036 vdd.n2342 vss 0.00425f
C3037 vdd.n2343 vss 0.00925f
C3038 vdd.n2344 vss 0.00679f
C3039 vdd.n2345 vss 0.00517f
C3040 vdd.n2346 vss 0.00251f
C3041 vdd.n2347 vss 0.0471f
C3042 vdd.n2348 vss 0.00251f
C3043 vdd.n2349 vss 0.0112f
C3044 vdd.n2350 vss 0.0128f
C3045 vdd.n2351 vss 0.0666f
C3046 vdd.n2352 vss 0.0912f
C3047 vdd.n2353 vss 0.0824f
C3048 vdd.n2354 vss 0.0567f
C3049 vdd.n2355 vss 0.00324f
C3050 vdd.n2356 vss 0.0112f
C3051 vdd.n2357 vss 0.0128f
C3052 vdd.n2358 vss 0.00413f
C3053 vdd.n2359 vss 0.00413f
C3054 vdd.n2360 vss 0.0471f
C3055 vdd.n2361 vss 0.0471f
C3056 vdd.n2362 vss 0.00324f
C3057 vdd.n2363 vss 0.00413f
C3058 vdd.n2364 vss 0.00413f
C3059 vdd.n2365 vss 0.00679f
C3060 vdd.n2366 vss 0.00413f
C3061 vdd.n2367 vss 0.0471f
C3062 vdd.n2368 vss 0.00324f
C3063 vdd.n2369 vss 0.0424f
C3064 vdd.n2370 vss 0.00324f
C3065 vdd.n2371 vss 0.0128f
C3066 vdd.n2372 vss 0.02f
C3067 vdd.n2373 vss 0.0132f
C3068 vdd.n2374 vss 0.00925f
C3069 vdd.n2375 vss 0.00425f
C3070 vdd.n2377 vss 0.0471f
C3071 vdd.n2378 vss 0.00425f
C3072 vdd.n2379 vss 0.00413f
C3073 vdd.n2380 vss 0.00251f
C3074 vdd.n2381 vss 0.0471f
C3075 vdd.n2382 vss 0.00251f
C3076 vdd.n2383 vss 0.00517f
C3077 vdd.n2384 vss 0.00679f
C3078 vdd.n2385 vss 0.00324f
C3079 vdd.n2386 vss 0.00324f
C3080 vdd.n2387 vss 0.0132f
C3081 vdd.n2388 vss 0.0424f
C3082 vdd.n2389 vss 0.02f
C3083 vdd.n2390 vss 0.00425f
C3084 vdd.n2392 vss 0.0471f
C3085 vdd.n2393 vss 0.00425f
C3086 vdd.n2394 vss 0.00925f
C3087 vdd.n2395 vss 0.00679f
C3088 vdd.n2396 vss 0.00517f
C3089 vdd.n2397 vss 0.00251f
C3090 vdd.n2398 vss 0.0471f
C3091 vdd.n2399 vss 0.00251f
C3092 vdd.n2400 vss 0.0112f
C3093 vdd.n2401 vss 0.0128f
C3094 vdd.n2402 vss 0.00324f
C3095 vdd.n2403 vss 0.0112f
C3096 vdd.n2404 vss 0.0128f
C3097 vdd.n2405 vss 0.00413f
C3098 vdd.n2406 vss 0.00413f
C3099 vdd.n2407 vss 0.0471f
C3100 vdd.n2408 vss 0.0471f
C3101 vdd.n2409 vss 0.00324f
C3102 vdd.n2410 vss 0.00413f
C3103 vdd.n2411 vss 0.00413f
C3104 vdd.n2412 vss 0.00679f
C3105 vdd.n2413 vss 0.00413f
C3106 vdd.n2414 vss 0.0471f
C3107 vdd.n2415 vss 0.00324f
C3108 vdd.n2416 vss 0.0424f
C3109 vdd.n2417 vss 0.00324f
C3110 vdd.n2418 vss 0.0128f
C3111 vdd.n2419 vss 0.02f
C3112 vdd.n2420 vss 0.0132f
C3113 vdd.n2421 vss 0.00925f
C3114 vdd.n2422 vss 0.00425f
C3115 vdd.n2424 vss 0.0471f
C3116 vdd.n2425 vss 0.00425f
C3117 vdd.n2426 vss 0.00413f
C3118 vdd.n2427 vss 0.00251f
C3119 vdd.n2428 vss 0.0471f
C3120 vdd.n2429 vss 0.00251f
C3121 vdd.n2430 vss 0.00517f
C3122 vdd.n2431 vss 0.00679f
C3123 vdd.n2432 vss 0.00324f
C3124 vdd.n2433 vss 0.00324f
C3125 vdd.n2434 vss 0.0132f
C3126 vdd.n2435 vss 0.0424f
C3127 vdd.n2436 vss 0.02f
C3128 vdd.n2437 vss 0.00425f
C3129 vdd.n2439 vss 0.0471f
C3130 vdd.n2440 vss 0.00425f
C3131 vdd.n2441 vss 0.00925f
C3132 vdd.n2442 vss 0.00679f
C3133 vdd.n2443 vss 0.00517f
C3134 vdd.n2444 vss 0.00251f
C3135 vdd.n2445 vss 0.0471f
C3136 vdd.n2446 vss 0.00251f
C3137 vdd.n2447 vss 0.0112f
C3138 vdd.n2448 vss 0.0128f
C3139 vdd.n2449 vss 0.144f
C3140 vdd.n2450 vss 0.143f
C3141 vdd.n2451 vss 0.0608f
C3142 vdd.n2452 vss 0.00324f
C3143 vdd.n2453 vss 0.0112f
C3144 vdd.n2454 vss 0.0128f
C3145 vdd.n2455 vss 0.00413f
C3146 vdd.n2456 vss 0.00413f
C3147 vdd.n2457 vss 0.0471f
C3148 vdd.n2458 vss 0.0471f
C3149 vdd.n2459 vss 0.00324f
C3150 vdd.n2460 vss 0.00413f
C3151 vdd.n2461 vss 0.00413f
C3152 vdd.n2462 vss 0.00679f
C3153 vdd.n2463 vss 0.00413f
C3154 vdd.n2464 vss 0.0471f
C3155 vdd.n2465 vss 0.00324f
C3156 vdd.n2466 vss 0.0424f
C3157 vdd.n2467 vss 0.00324f
C3158 vdd.n2468 vss 0.0128f
C3159 vdd.n2469 vss 0.02f
C3160 vdd.n2470 vss 0.0132f
C3161 vdd.n2471 vss 0.00925f
C3162 vdd.n2472 vss 0.00425f
C3163 vdd.n2474 vss 0.0471f
C3164 vdd.n2475 vss 0.00425f
C3165 vdd.n2476 vss 0.00413f
C3166 vdd.n2477 vss 0.00251f
C3167 vdd.n2478 vss 0.0471f
C3168 vdd.n2479 vss 0.00251f
C3169 vdd.n2480 vss 0.00517f
C3170 vdd.n2481 vss 0.00679f
C3171 vdd.n2482 vss 0.00324f
C3172 vdd.n2483 vss 0.00324f
C3173 vdd.n2484 vss 0.0132f
C3174 vdd.n2485 vss 0.0424f
C3175 vdd.n2486 vss 0.02f
C3176 vdd.n2487 vss 0.00425f
C3177 vdd.n2489 vss 0.0471f
C3178 vdd.n2490 vss 0.00425f
C3179 vdd.n2491 vss 0.00925f
C3180 vdd.n2492 vss 0.00679f
C3181 vdd.n2493 vss 0.00517f
C3182 vdd.n2494 vss 0.00251f
C3183 vdd.n2495 vss 0.0471f
C3184 vdd.n2496 vss 0.00251f
C3185 vdd.n2497 vss 0.0112f
C3186 vdd.n2498 vss 0.0128f
C3187 vdd.n2499 vss 0.0666f
C3188 vdd.n2500 vss 0.118f
C3189 vdd.n2501 vss 0.121f
C3190 vdd.n2502 vss 0.00324f
C3191 vdd.n2503 vss 0.0112f
C3192 vdd.n2504 vss 0.0128f
C3193 vdd.n2505 vss 0.00413f
C3194 vdd.n2506 vss 0.00413f
C3195 vdd.n2507 vss 0.0471f
C3196 vdd.n2508 vss 0.0471f
C3197 vdd.n2509 vss 0.00324f
C3198 vdd.n2510 vss 0.00413f
C3199 vdd.n2511 vss 0.00413f
C3200 vdd.n2512 vss 0.00679f
C3201 vdd.n2513 vss 0.00413f
C3202 vdd.n2514 vss 0.0471f
C3203 vdd.n2515 vss 0.00324f
C3204 vdd.n2516 vss 0.0424f
C3205 vdd.n2517 vss 0.00324f
C3206 vdd.n2518 vss 0.0128f
C3207 vdd.n2519 vss 0.02f
C3208 vdd.n2520 vss 0.0132f
C3209 vdd.n2521 vss 0.00925f
C3210 vdd.n2522 vss 0.00425f
C3211 vdd.n2524 vss 0.0471f
C3212 vdd.n2525 vss 0.00425f
C3213 vdd.n2526 vss 0.00413f
C3214 vdd.n2527 vss 0.00251f
C3215 vdd.n2528 vss 0.0471f
C3216 vdd.n2529 vss 0.00251f
C3217 vdd.n2530 vss 0.00517f
C3218 vdd.n2531 vss 0.00679f
C3219 vdd.n2532 vss 0.00324f
C3220 vdd.n2533 vss 0.00324f
C3221 vdd.n2534 vss 0.0132f
C3222 vdd.n2535 vss 0.0424f
C3223 vdd.n2536 vss 0.02f
C3224 vdd.n2537 vss 0.00425f
C3225 vdd.n2539 vss 0.0471f
C3226 vdd.n2540 vss 0.00425f
C3227 vdd.n2541 vss 0.00925f
C3228 vdd.n2542 vss 0.00679f
C3229 vdd.n2543 vss 0.00517f
C3230 vdd.n2544 vss 0.00251f
C3231 vdd.n2545 vss 0.0471f
C3232 vdd.n2546 vss 0.00251f
C3233 vdd.n2547 vss 0.0112f
C3234 vdd.n2548 vss 0.0955f
C3235 vdd.n2549 vss 0.0608f
C3236 vdd.n2550 vss 0.00324f
C3237 vdd.n2551 vss 0.0112f
C3238 vdd.n2552 vss 0.0128f
C3239 vdd.n2553 vss 0.00413f
C3240 vdd.n2554 vss 0.00413f
C3241 vdd.n2555 vss 0.0471f
C3242 vdd.n2556 vss 0.0471f
C3243 vdd.n2557 vss 0.00324f
C3244 vdd.n2558 vss 0.00413f
C3245 vdd.n2559 vss 0.00413f
C3246 vdd.n2560 vss 0.00679f
C3247 vdd.n2561 vss 0.00413f
C3248 vdd.n2562 vss 0.0471f
C3249 vdd.n2563 vss 0.00324f
C3250 vdd.n2564 vss 0.0424f
C3251 vdd.n2565 vss 0.00324f
C3252 vdd.n2566 vss 0.0128f
C3253 vdd.n2567 vss 0.02f
C3254 vdd.n2568 vss 0.0132f
C3255 vdd.n2569 vss 0.00925f
C3256 vdd.n2570 vss 0.00425f
C3257 vdd.n2572 vss 0.0471f
C3258 vdd.n2573 vss 0.00425f
C3259 vdd.n2574 vss 0.00413f
C3260 vdd.n2575 vss 0.00251f
C3261 vdd.n2576 vss 0.0471f
C3262 vdd.n2577 vss 0.00251f
C3263 vdd.n2578 vss 0.00517f
C3264 vdd.n2579 vss 0.00679f
C3265 vdd.n2580 vss 0.00324f
C3266 vdd.n2581 vss 0.00324f
C3267 vdd.n2582 vss 0.0132f
C3268 vdd.n2583 vss 0.0424f
C3269 vdd.n2584 vss 0.02f
C3270 vdd.n2585 vss 0.00425f
C3271 vdd.n2587 vss 0.0471f
C3272 vdd.n2588 vss 0.00425f
C3273 vdd.n2589 vss 0.00925f
C3274 vdd.n2590 vss 0.00679f
C3275 vdd.n2591 vss 0.00517f
C3276 vdd.n2592 vss 0.00251f
C3277 vdd.n2593 vss 0.0471f
C3278 vdd.n2594 vss 0.00251f
C3279 vdd.n2595 vss 0.0112f
C3280 vdd.n2596 vss 0.0128f
C3281 vdd.n2597 vss 0.0666f
C3282 vdd.n2598 vss 0.299f
C3283 vdd.n2599 vss 0.00324f
C3284 vdd.n2600 vss 0.0112f
C3285 vdd.n2601 vss 0.0128f
C3286 vdd.n2602 vss 0.00413f
C3287 vdd.n2603 vss 0.00413f
C3288 vdd.n2604 vss 0.0471f
C3289 vdd.n2605 vss 0.0471f
C3290 vdd.n2606 vss 0.00324f
C3291 vdd.n2607 vss 0.00413f
C3292 vdd.n2608 vss 0.00413f
C3293 vdd.n2609 vss 0.00679f
C3294 vdd.n2610 vss 0.00413f
C3295 vdd.n2611 vss 0.0471f
C3296 vdd.n2612 vss 0.00324f
C3297 vdd.n2614 vss 0.00925f
C3298 vdd.n2615 vss 0.0471f
C3299 vdd.n2616 vss 0.00425f
C3300 vdd.n2617 vss 0.0424f
C3301 vdd.n2618 vss 0.0132f
C3302 vdd.n2619 vss 0.00324f
C3303 vdd.n2620 vss 0.0128f
C3304 vdd.n2621 vss 0.02f
C3305 vdd.n2622 vss 0.00425f
C3306 vdd.n2623 vss 0.00413f
C3307 vdd.n2624 vss 0.00251f
C3308 vdd.n2625 vss 0.0471f
C3309 vdd.n2626 vss 0.00251f
C3310 vdd.n2627 vss 0.00517f
C3311 vdd.n2628 vss 0.00679f
C3312 vdd.n2629 vss 0.00324f
C3313 vdd.n2630 vss 0.00324f
C3314 vdd.n2631 vss 0.0132f
C3315 vdd.n2632 vss 0.0424f
C3316 vdd.n2633 vss 0.02f
C3317 vdd.n2634 vss 0.00425f
C3318 vdd.n2635 vss 0.0471f
C3319 vdd.n2637 vss 0.00425f
C3320 vdd.n2638 vss 0.00925f
C3321 vdd.n2639 vss 0.00679f
C3322 vdd.n2640 vss 0.00517f
C3323 vdd.n2641 vss 0.00251f
C3324 vdd.n2642 vss 0.0471f
C3325 vdd.n2643 vss 0.00251f
C3326 vdd.n2644 vss 0.0112f
C3327 vdd.n2645 vss 0.0128f
C3328 vdd.n2646 vss 0.0619f
C3329 vdd.n2647 vss 0.262f
C3330 vdd.n2648 vss 0.00324f
C3331 vdd.n2649 vss 0.0112f
C3332 vdd.n2650 vss 0.0128f
C3333 vdd.n2651 vss 0.00413f
C3334 vdd.n2652 vss 0.00413f
C3335 vdd.n2653 vss 0.0471f
C3336 vdd.n2654 vss 0.0471f
C3337 vdd.n2655 vss 0.00324f
C3338 vdd.n2656 vss 0.00413f
C3339 vdd.n2657 vss 0.00413f
C3340 vdd.n2658 vss 0.00679f
C3341 vdd.n2659 vss 0.00413f
C3342 vdd.n2660 vss 0.0471f
C3343 vdd.n2661 vss 0.00324f
C3344 vdd.n2663 vss 0.00925f
C3345 vdd.n2664 vss 0.0471f
C3346 vdd.n2665 vss 0.00425f
C3347 vdd.n2666 vss 0.0424f
C3348 vdd.n2667 vss 0.0132f
C3349 vdd.n2668 vss 0.00324f
C3350 vdd.n2669 vss 0.0128f
C3351 vdd.n2670 vss 0.02f
C3352 vdd.n2671 vss 0.00425f
C3353 vdd.n2672 vss 0.00413f
C3354 vdd.n2673 vss 0.00251f
C3355 vdd.n2674 vss 0.0471f
C3356 vdd.n2675 vss 0.00251f
C3357 vdd.n2676 vss 0.00517f
C3358 vdd.n2677 vss 0.00679f
C3359 vdd.n2678 vss 0.00324f
C3360 vdd.n2679 vss 0.00324f
C3361 vdd.n2680 vss 0.0132f
C3362 vdd.n2681 vss 0.0424f
C3363 vdd.n2682 vss 0.02f
C3364 vdd.n2683 vss 0.00425f
C3365 vdd.n2684 vss 0.0471f
C3366 vdd.n2686 vss 0.00425f
C3367 vdd.n2687 vss 0.00925f
C3368 vdd.n2688 vss 0.00679f
C3369 vdd.n2689 vss 0.00517f
C3370 vdd.n2690 vss 0.00251f
C3371 vdd.n2691 vss 0.0471f
C3372 vdd.n2692 vss 0.00251f
C3373 vdd.n2693 vss 0.0112f
C3374 vdd.n2694 vss 0.0128f
C3375 vdd.n2695 vss 0.146f
C3376 vdd.n2696 vss 0.00324f
C3377 vdd.n2697 vss 0.0112f
C3378 vdd.n2698 vss 0.0128f
C3379 vdd.n2699 vss 0.00413f
C3380 vdd.n2700 vss 0.00413f
C3381 vdd.n2701 vss 0.0471f
C3382 vdd.n2702 vss 0.0471f
C3383 vdd.n2703 vss 0.00324f
C3384 vdd.n2704 vss 0.00413f
C3385 vdd.n2705 vss 0.00413f
C3386 vdd.n2706 vss 0.00679f
C3387 vdd.n2707 vss 0.00413f
C3388 vdd.n2708 vss 0.0471f
C3389 vdd.n2709 vss 0.00324f
C3390 vdd.n2711 vss 0.00925f
C3391 vdd.n2712 vss 0.0471f
C3392 vdd.n2713 vss 0.00425f
C3393 vdd.n2714 vss 0.0424f
C3394 vdd.n2715 vss 0.0132f
C3395 vdd.n2716 vss 0.00324f
C3396 vdd.n2717 vss 0.0128f
C3397 vdd.n2718 vss 0.02f
C3398 vdd.n2719 vss 0.00425f
C3399 vdd.n2720 vss 0.00413f
C3400 vdd.n2721 vss 0.00251f
C3401 vdd.n2722 vss 0.0471f
C3402 vdd.n2723 vss 0.00251f
C3403 vdd.n2724 vss 0.00517f
C3404 vdd.n2725 vss 0.00679f
C3405 vdd.n2726 vss 0.00324f
C3406 vdd.n2727 vss 0.00324f
C3407 vdd.n2728 vss 0.0132f
C3408 vdd.n2729 vss 0.0424f
C3409 vdd.n2730 vss 0.02f
C3410 vdd.n2731 vss 0.00425f
C3411 vdd.n2732 vss 0.0471f
C3412 vdd.n2734 vss 0.00425f
C3413 vdd.n2735 vss 0.00925f
C3414 vdd.n2736 vss 0.00679f
C3415 vdd.n2737 vss 0.00517f
C3416 vdd.n2738 vss 0.00251f
C3417 vdd.n2739 vss 0.0471f
C3418 vdd.n2740 vss 0.00251f
C3419 vdd.n2741 vss 0.0112f
C3420 vdd.n2742 vss 0.0128f
C3421 vdd.n2743 vss 0.146f
C3422 vdd.n2744 vss 0.0596f
C3423 vdd.n2745 vss 0.00324f
C3424 vdd.n2746 vss 0.0112f
C3425 vdd.n2747 vss 0.0128f
C3426 vdd.n2748 vss 0.00413f
C3427 vdd.n2749 vss 0.00413f
C3428 vdd.n2750 vss 0.0471f
C3429 vdd.n2751 vss 0.0471f
C3430 vdd.n2752 vss 0.00324f
C3431 vdd.n2753 vss 0.00413f
C3432 vdd.n2754 vss 0.00413f
C3433 vdd.n2755 vss 0.00679f
C3434 vdd.n2756 vss 0.00413f
C3435 vdd.n2757 vss 0.0471f
C3436 vdd.n2758 vss 0.00324f
C3437 vdd.n2760 vss 0.00925f
C3438 vdd.n2761 vss 0.0471f
C3439 vdd.n2762 vss 0.00425f
C3440 vdd.n2763 vss 0.0424f
C3441 vdd.n2764 vss 0.0132f
C3442 vdd.n2765 vss 0.00324f
C3443 vdd.n2766 vss 0.0128f
C3444 vdd.n2767 vss 0.02f
C3445 vdd.n2768 vss 0.00425f
C3446 vdd.n2769 vss 0.00413f
C3447 vdd.n2770 vss 0.00251f
C3448 vdd.n2771 vss 0.0471f
C3449 vdd.n2772 vss 0.00251f
C3450 vdd.n2773 vss 0.00517f
C3451 vdd.n2774 vss 0.00679f
C3452 vdd.n2775 vss 0.00324f
C3453 vdd.n2776 vss 0.00324f
C3454 vdd.n2777 vss 0.0132f
C3455 vdd.n2778 vss 0.0424f
C3456 vdd.n2779 vss 0.02f
C3457 vdd.n2780 vss 0.00425f
C3458 vdd.n2781 vss 0.0471f
C3459 vdd.n2783 vss 0.00425f
C3460 vdd.n2784 vss 0.00925f
C3461 vdd.n2785 vss 0.00679f
C3462 vdd.n2786 vss 0.00517f
C3463 vdd.n2787 vss 0.00251f
C3464 vdd.n2788 vss 0.0471f
C3465 vdd.n2789 vss 0.00251f
C3466 vdd.n2790 vss 0.0112f
C3467 vdd.n2791 vss 0.0128f
C3468 vdd.n2792 vss 0.0692f
C3469 vdd.n2793 vss 0.118f
C3470 vdd.n2794 vss 0.121f
C3471 vdd.n2795 vss 0.00324f
C3472 vdd.n2796 vss 0.0112f
C3473 vdd.n2797 vss 0.0128f
C3474 vdd.n2798 vss 0.00413f
C3475 vdd.n2799 vss 0.00413f
C3476 vdd.n2800 vss 0.0471f
C3477 vdd.n2801 vss 0.0471f
C3478 vdd.n2802 vss 0.00324f
C3479 vdd.n2803 vss 0.00413f
C3480 vdd.n2804 vss 0.00413f
C3481 vdd.n2805 vss 0.00679f
C3482 vdd.n2806 vss 0.00413f
C3483 vdd.n2807 vss 0.0471f
C3484 vdd.n2808 vss 0.00324f
C3485 vdd.n2810 vss 0.00925f
C3486 vdd.n2811 vss 0.0471f
C3487 vdd.n2812 vss 0.00425f
C3488 vdd.n2813 vss 0.0424f
C3489 vdd.n2814 vss 0.0132f
C3490 vdd.n2815 vss 0.00324f
C3491 vdd.n2816 vss 0.0128f
C3492 vdd.n2817 vss 0.02f
C3493 vdd.n2818 vss 0.00425f
C3494 vdd.n2819 vss 0.00413f
C3495 vdd.n2820 vss 0.00251f
C3496 vdd.n2821 vss 0.0471f
C3497 vdd.n2822 vss 0.00251f
C3498 vdd.n2823 vss 0.00517f
C3499 vdd.n2824 vss 0.00679f
C3500 vdd.n2825 vss 0.00324f
C3501 vdd.n2826 vss 0.00324f
C3502 vdd.n2827 vss 0.0132f
C3503 vdd.n2828 vss 0.0424f
C3504 vdd.n2829 vss 0.02f
C3505 vdd.n2830 vss 0.00425f
C3506 vdd.n2831 vss 0.0471f
C3507 vdd.n2833 vss 0.00425f
C3508 vdd.n2834 vss 0.00925f
C3509 vdd.n2835 vss 0.00679f
C3510 vdd.n2836 vss 0.00517f
C3511 vdd.n2837 vss 0.00251f
C3512 vdd.n2838 vss 0.0471f
C3513 vdd.n2839 vss 0.00251f
C3514 vdd.n2840 vss 0.0112f
C3515 vdd.n2841 vss 0.098f
C3516 vdd.n2842 vss 0.0596f
C3517 vdd.n2843 vss 0.00324f
C3518 vdd.n2844 vss 0.0112f
C3519 vdd.n2845 vss 0.0128f
C3520 vdd.n2846 vss 0.00413f
C3521 vdd.n2847 vss 0.00413f
C3522 vdd.n2848 vss 0.0471f
C3523 vdd.n2849 vss 0.0471f
C3524 vdd.n2850 vss 0.00324f
C3525 vdd.n2851 vss 0.00413f
C3526 vdd.n2852 vss 0.00413f
C3527 vdd.n2853 vss 0.00679f
C3528 vdd.n2854 vss 0.00413f
C3529 vdd.n2855 vss 0.0471f
C3530 vdd.n2856 vss 0.00324f
C3531 vdd.n2858 vss 0.00925f
C3532 vdd.n2859 vss 0.0471f
C3533 vdd.n2860 vss 0.00425f
C3534 vdd.n2861 vss 0.0424f
C3535 vdd.n2862 vss 0.0132f
C3536 vdd.n2863 vss 0.00324f
C3537 vdd.n2864 vss 0.0128f
C3538 vdd.n2865 vss 0.02f
C3539 vdd.n2866 vss 0.00425f
C3540 vdd.n2867 vss 0.00413f
C3541 vdd.n2868 vss 0.00251f
C3542 vdd.n2869 vss 0.0471f
C3543 vdd.n2870 vss 0.00251f
C3544 vdd.n2871 vss 0.00517f
C3545 vdd.n2872 vss 0.00679f
C3546 vdd.n2873 vss 0.00324f
C3547 vdd.n2874 vss 0.00324f
C3548 vdd.n2875 vss 0.0132f
C3549 vdd.n2876 vss 0.0424f
C3550 vdd.n2877 vss 0.02f
C3551 vdd.n2878 vss 0.00425f
C3552 vdd.n2879 vss 0.0471f
C3553 vdd.n2881 vss 0.00425f
C3554 vdd.n2882 vss 0.00925f
C3555 vdd.n2883 vss 0.00679f
C3556 vdd.n2884 vss 0.00517f
C3557 vdd.n2885 vss 0.00251f
C3558 vdd.n2886 vss 0.0471f
C3559 vdd.n2887 vss 0.00251f
C3560 vdd.n2888 vss 0.0112f
C3561 vdd.n2889 vss 0.0128f
C3562 vdd.n2890 vss 0.0692f
C3563 vdd.n2891 vss 0.0912f
C3564 vdd.n2892 vss 0.0824f
C3565 vdd.n2893 vss 0.059f
C3566 vdd.n2894 vss 0.00324f
C3567 vdd.n2895 vss 0.0112f
C3568 vdd.n2896 vss 0.0128f
C3569 vdd.n2897 vss 0.00413f
C3570 vdd.n2898 vss 0.00413f
C3571 vdd.n2899 vss 0.0471f
C3572 vdd.n2900 vss 0.0471f
C3573 vdd.n2901 vss 0.00324f
C3574 vdd.n2902 vss 0.00413f
C3575 vdd.n2903 vss 0.00413f
C3576 vdd.n2904 vss 0.00679f
C3577 vdd.n2905 vss 0.00413f
C3578 vdd.n2906 vss 0.0471f
C3579 vdd.n2907 vss 0.00324f
C3580 vdd.n2909 vss 0.00925f
C3581 vdd.n2910 vss 0.0471f
C3582 vdd.n2911 vss 0.00425f
C3583 vdd.n2912 vss 0.0424f
C3584 vdd.n2913 vss 0.0132f
C3585 vdd.n2914 vss 0.00324f
C3586 vdd.n2915 vss 0.0128f
C3587 vdd.n2916 vss 0.02f
C3588 vdd.n2917 vss 0.00425f
C3589 vdd.n2918 vss 0.00413f
C3590 vdd.n2919 vss 0.00251f
C3591 vdd.n2920 vss 0.0471f
C3592 vdd.n2921 vss 0.00251f
C3593 vdd.n2922 vss 0.00517f
C3594 vdd.n2923 vss 0.00679f
C3595 vdd.n2924 vss 0.00324f
C3596 vdd.n2925 vss 0.00324f
C3597 vdd.n2926 vss 0.0132f
C3598 vdd.n2927 vss 0.0424f
C3599 vdd.n2928 vss 0.02f
C3600 vdd.n2929 vss 0.00425f
C3601 vdd.n2930 vss 0.0471f
C3602 vdd.n2932 vss 0.00425f
C3603 vdd.n2933 vss 0.00925f
C3604 vdd.n2934 vss 0.00679f
C3605 vdd.n2935 vss 0.00517f
C3606 vdd.n2936 vss 0.00251f
C3607 vdd.n2937 vss 0.0471f
C3608 vdd.n2938 vss 0.00251f
C3609 vdd.n2939 vss 0.0112f
C3610 vdd.n2940 vss 0.0128f
C3611 vdd.n2941 vss 0.185f
C3612 vdd.n2942 vss 0.00324f
C3613 vdd.n2943 vss 0.0112f
C3614 vdd.n2944 vss 0.0128f
C3615 vdd.n2945 vss 0.00413f
C3616 vdd.n2946 vss 0.00413f
C3617 vdd.n2947 vss 0.0471f
C3618 vdd.n2948 vss 0.0471f
C3619 vdd.n2949 vss 0.00324f
C3620 vdd.n2950 vss 0.00413f
C3621 vdd.n2951 vss 0.00413f
C3622 vdd.n2952 vss 0.00679f
C3623 vdd.n2953 vss 0.00413f
C3624 vdd.n2954 vss 0.0471f
C3625 vdd.n2955 vss 0.00324f
C3626 vdd.n2957 vss 0.00925f
C3627 vdd.n2958 vss 0.0471f
C3628 vdd.n2959 vss 0.00425f
C3629 vdd.n2960 vss 0.0424f
C3630 vdd.n2961 vss 0.0132f
C3631 vdd.n2962 vss 0.00324f
C3632 vdd.n2963 vss 0.0128f
C3633 vdd.n2964 vss 0.02f
C3634 vdd.n2965 vss 0.00425f
C3635 vdd.n2966 vss 0.00413f
C3636 vdd.n2967 vss 0.00251f
C3637 vdd.n2968 vss 0.0471f
C3638 vdd.n2969 vss 0.00251f
C3639 vdd.n2970 vss 0.00517f
C3640 vdd.n2971 vss 0.00679f
C3641 vdd.n2972 vss 0.00324f
C3642 vdd.n2973 vss 0.00324f
C3643 vdd.n2974 vss 0.0132f
C3644 vdd.n2975 vss 0.0424f
C3645 vdd.n2976 vss 0.02f
C3646 vdd.n2977 vss 0.00425f
C3647 vdd.n2978 vss 0.0471f
C3648 vdd.n2980 vss 0.00425f
C3649 vdd.n2981 vss 0.00925f
C3650 vdd.n2982 vss 0.00679f
C3651 vdd.n2983 vss 0.00517f
C3652 vdd.n2984 vss 0.00251f
C3653 vdd.n2985 vss 0.0471f
C3654 vdd.n2986 vss 0.00251f
C3655 vdd.n2987 vss 0.0112f
C3656 vdd.n2988 vss 0.0128f
C3657 vdd.n2989 vss 0.059f
C3658 vdd.n2990 vss 0.256f
C3659 vdd.n2991 vss 0.00324f
C3660 vdd.n2992 vss 0.0112f
C3661 vdd.n2993 vss 0.0128f
C3662 vdd.n2994 vss 0.00413f
C3663 vdd.n2995 vss 0.00413f
C3664 vdd.n2996 vss 0.0471f
C3665 vdd.n2997 vss 0.0471f
C3666 vdd.n2998 vss 0.00324f
C3667 vdd.n2999 vss 0.00413f
C3668 vdd.n3000 vss 0.00413f
C3669 vdd.n3001 vss 0.00679f
C3670 vdd.n3002 vss 0.00413f
C3671 vdd.n3003 vss 0.0471f
C3672 vdd.n3004 vss 0.00324f
C3673 vdd.n3006 vss 0.00925f
C3674 vdd.n3007 vss 0.0471f
C3675 vdd.n3008 vss 0.00425f
C3676 vdd.n3009 vss 0.0424f
C3677 vdd.n3010 vss 0.0132f
C3678 vdd.n3011 vss 0.00324f
C3679 vdd.n3012 vss 0.0128f
C3680 vdd.n3013 vss 0.02f
C3681 vdd.n3014 vss 0.00425f
C3682 vdd.n3015 vss 0.00413f
C3683 vdd.n3016 vss 0.00251f
C3684 vdd.n3017 vss 0.0471f
C3685 vdd.n3018 vss 0.00251f
C3686 vdd.n3019 vss 0.00517f
C3687 vdd.n3020 vss 0.00679f
C3688 vdd.n3021 vss 0.00324f
C3689 vdd.n3022 vss 0.00324f
C3690 vdd.n3023 vss 0.0132f
C3691 vdd.n3024 vss 0.0424f
C3692 vdd.n3025 vss 0.02f
C3693 vdd.n3026 vss 0.00425f
C3694 vdd.n3027 vss 0.0471f
C3695 vdd.n3029 vss 0.00425f
C3696 vdd.n3030 vss 0.00925f
C3697 vdd.n3031 vss 0.00679f
C3698 vdd.n3032 vss 0.00517f
C3699 vdd.n3033 vss 0.00251f
C3700 vdd.n3034 vss 0.0471f
C3701 vdd.n3035 vss 0.00251f
C3702 vdd.n3036 vss 0.0112f
C3703 vdd.n3037 vss 0.0128f
C3704 vdd.n3038 vss 0.123f
C3705 vdd.n3039 vss 0.0596f
C3706 vdd.n3040 vss 0.00324f
C3707 vdd.n3041 vss 0.0112f
C3708 vdd.n3042 vss 0.0128f
C3709 vdd.n3043 vss 0.00413f
C3710 vdd.n3044 vss 0.00413f
C3711 vdd.n3045 vss 0.0471f
C3712 vdd.n3046 vss 0.0471f
C3713 vdd.n3047 vss 0.00324f
C3714 vdd.n3048 vss 0.00413f
C3715 vdd.n3049 vss 0.00413f
C3716 vdd.n3050 vss 0.00679f
C3717 vdd.n3051 vss 0.00413f
C3718 vdd.n3052 vss 0.0471f
C3719 vdd.n3053 vss 0.00324f
C3720 vdd.n3055 vss 0.00925f
C3721 vdd.n3056 vss 0.0471f
C3722 vdd.n3057 vss 0.00425f
C3723 vdd.n3058 vss 0.0424f
C3724 vdd.n3059 vss 0.0132f
C3725 vdd.n3060 vss 0.00324f
C3726 vdd.n3061 vss 0.0128f
C3727 vdd.n3062 vss 0.02f
C3728 vdd.n3063 vss 0.00425f
C3729 vdd.n3064 vss 0.00413f
C3730 vdd.n3065 vss 0.00251f
C3731 vdd.n3066 vss 0.0471f
C3732 vdd.n3067 vss 0.00251f
C3733 vdd.n3068 vss 0.00517f
C3734 vdd.n3069 vss 0.00679f
C3735 vdd.n3070 vss 0.00324f
C3736 vdd.n3071 vss 0.00324f
C3737 vdd.n3072 vss 0.0132f
C3738 vdd.n3073 vss 0.0424f
C3739 vdd.n3074 vss 0.02f
C3740 vdd.n3075 vss 0.00425f
C3741 vdd.n3076 vss 0.0471f
C3742 vdd.n3078 vss 0.00425f
C3743 vdd.n3079 vss 0.00925f
C3744 vdd.n3080 vss 0.00679f
C3745 vdd.n3081 vss 0.00517f
C3746 vdd.n3082 vss 0.00251f
C3747 vdd.n3083 vss 0.0471f
C3748 vdd.n3084 vss 0.00251f
C3749 vdd.n3085 vss 0.0112f
C3750 vdd.n3086 vss 0.0128f
C3751 vdd.n3087 vss 0.0692f
C3752 vdd.n3088 vss 0.118f
C3753 vdd.n3089 vss 0.121f
C3754 vdd.n3090 vss 0.00324f
C3755 vdd.n3091 vss 0.0112f
C3756 vdd.n3092 vss 0.0128f
C3757 vdd.n3093 vss 0.00413f
C3758 vdd.n3094 vss 0.00413f
C3759 vdd.n3095 vss 0.0471f
C3760 vdd.n3096 vss 0.0471f
C3761 vdd.n3097 vss 0.00324f
C3762 vdd.n3098 vss 0.00413f
C3763 vdd.n3099 vss 0.00413f
C3764 vdd.n3100 vss 0.00679f
C3765 vdd.n3101 vss 0.00413f
C3766 vdd.n3102 vss 0.0471f
C3767 vdd.n3103 vss 0.00324f
C3768 vdd.n3105 vss 0.00925f
C3769 vdd.n3106 vss 0.0471f
C3770 vdd.n3107 vss 0.00425f
C3771 vdd.n3108 vss 0.0424f
C3772 vdd.n3109 vss 0.0132f
C3773 vdd.n3110 vss 0.00324f
C3774 vdd.n3111 vss 0.0128f
C3775 vdd.n3112 vss 0.02f
C3776 vdd.n3113 vss 0.00425f
C3777 vdd.n3114 vss 0.00413f
C3778 vdd.n3115 vss 0.00251f
C3779 vdd.n3116 vss 0.0471f
C3780 vdd.n3117 vss 0.00251f
C3781 vdd.n3118 vss 0.00517f
C3782 vdd.n3119 vss 0.00679f
C3783 vdd.n3120 vss 0.00324f
C3784 vdd.n3121 vss 0.00324f
C3785 vdd.n3122 vss 0.0132f
C3786 vdd.n3123 vss 0.0424f
C3787 vdd.n3124 vss 0.02f
C3788 vdd.n3125 vss 0.00425f
C3789 vdd.n3126 vss 0.0471f
C3790 vdd.n3128 vss 0.00425f
C3791 vdd.n3129 vss 0.00925f
C3792 vdd.n3130 vss 0.00679f
C3793 vdd.n3131 vss 0.00517f
C3794 vdd.n3132 vss 0.00251f
C3795 vdd.n3133 vss 0.0471f
C3796 vdd.n3134 vss 0.00251f
C3797 vdd.n3135 vss 0.0112f
C3798 vdd.n3136 vss 0.098f
C3799 vdd.n3137 vss 0.0596f
C3800 vdd.n3138 vss 0.00324f
C3801 vdd.n3139 vss 0.0112f
C3802 vdd.n3140 vss 0.0128f
C3803 vdd.n3141 vss 0.00413f
C3804 vdd.n3142 vss 0.00413f
C3805 vdd.n3143 vss 0.0471f
C3806 vdd.n3144 vss 0.0471f
C3807 vdd.n3145 vss 0.00324f
C3808 vdd.n3146 vss 0.00413f
C3809 vdd.n3147 vss 0.00413f
C3810 vdd.n3148 vss 0.00679f
C3811 vdd.n3149 vss 0.00413f
C3812 vdd.n3150 vss 0.0471f
C3813 vdd.n3151 vss 0.00324f
C3814 vdd.n3153 vss 0.00925f
C3815 vdd.n3154 vss 0.0471f
C3816 vdd.n3155 vss 0.00425f
C3817 vdd.n3156 vss 0.0424f
C3818 vdd.n3157 vss 0.0132f
C3819 vdd.n3158 vss 0.00324f
C3820 vdd.n3159 vss 0.0128f
C3821 vdd.n3160 vss 0.02f
C3822 vdd.n3161 vss 0.00425f
C3823 vdd.n3162 vss 0.00413f
C3824 vdd.n3163 vss 0.00251f
C3825 vdd.n3164 vss 0.0471f
C3826 vdd.n3165 vss 0.00251f
C3827 vdd.n3166 vss 0.00517f
C3828 vdd.n3167 vss 0.00679f
C3829 vdd.n3168 vss 0.00324f
C3830 vdd.n3169 vss 0.00324f
C3831 vdd.n3170 vss 0.0132f
C3832 vdd.n3171 vss 0.0424f
C3833 vdd.n3172 vss 0.02f
C3834 vdd.n3173 vss 0.00425f
C3835 vdd.n3174 vss 0.0471f
C3836 vdd.n3176 vss 0.00425f
C3837 vdd.n3177 vss 0.00925f
C3838 vdd.n3178 vss 0.00679f
C3839 vdd.n3179 vss 0.00517f
C3840 vdd.n3180 vss 0.00251f
C3841 vdd.n3181 vss 0.0471f
C3842 vdd.n3182 vss 0.00251f
C3843 vdd.n3183 vss 0.0112f
C3844 vdd.n3184 vss 0.0128f
C3845 vdd.n3185 vss 0.0692f
C3846 vdd.n3186 vss 0.118f
C3847 vdd.n3187 vss 0.0951f
C3848 vdd.n3188 vss 0.00324f
C3849 vdd.n3189 vss 0.0112f
C3850 vdd.n3190 vss 0.0128f
C3851 vdd.n3191 vss 0.00413f
C3852 vdd.n3192 vss 0.00413f
C3853 vdd.n3193 vss 0.0471f
C3854 vdd.n3194 vss 0.0471f
C3855 vdd.n3195 vss 0.00324f
C3856 vdd.n3196 vss 0.00413f
C3857 vdd.n3197 vss 0.00413f
C3858 vdd.n3198 vss 0.00679f
C3859 vdd.n3199 vss 0.00413f
C3860 vdd.n3200 vss 0.0471f
C3861 vdd.n3201 vss 0.00324f
C3862 vdd.n3203 vss 0.00925f
C3863 vdd.n3204 vss 0.0471f
C3864 vdd.n3205 vss 0.00425f
C3865 vdd.n3206 vss 0.0424f
C3866 vdd.n3207 vss 0.0132f
C3867 vdd.n3208 vss 0.00324f
C3868 vdd.n3209 vss 0.0128f
C3869 vdd.n3210 vss 0.02f
C3870 vdd.n3211 vss 0.00425f
C3871 vdd.n3212 vss 0.00413f
C3872 vdd.n3213 vss 0.00251f
C3873 vdd.n3214 vss 0.0471f
C3874 vdd.n3215 vss 0.00251f
C3875 vdd.n3216 vss 0.00517f
C3876 vdd.n3217 vss 0.00679f
C3877 vdd.n3218 vss 0.00324f
C3878 vdd.n3219 vss 0.00324f
C3879 vdd.n3220 vss 0.0132f
C3880 vdd.n3221 vss 0.0424f
C3881 vdd.n3222 vss 0.02f
C3882 vdd.n3223 vss 0.00425f
C3883 vdd.n3224 vss 0.0471f
C3884 vdd.n3226 vss 0.00425f
C3885 vdd.n3227 vss 0.00925f
C3886 vdd.n3228 vss 0.00679f
C3887 vdd.n3229 vss 0.00517f
C3888 vdd.n3230 vss 0.00251f
C3889 vdd.n3231 vss 0.0471f
C3890 vdd.n3232 vss 0.00251f
C3891 vdd.n3233 vss 0.0112f
C3892 vdd.n3234 vss 0.0128f
C3893 vdd.n3235 vss 0.146f
C3894 vdd.n3236 vss 0.00324f
C3895 vdd.n3237 vss 0.0112f
C3896 vdd.n3238 vss 0.0128f
C3897 vdd.n3239 vss 0.00413f
C3898 vdd.n3240 vss 0.00413f
C3899 vdd.n3241 vss 0.0471f
C3900 vdd.n3242 vss 0.0471f
C3901 vdd.n3243 vss 0.00324f
C3902 vdd.n3244 vss 0.00413f
C3903 vdd.n3245 vss 0.00413f
C3904 vdd.n3246 vss 0.00679f
C3905 vdd.n3247 vss 0.00413f
C3906 vdd.n3248 vss 0.0471f
C3907 vdd.n3249 vss 0.00324f
C3908 vdd.n3251 vss 0.00925f
C3909 vdd.n3252 vss 0.0471f
C3910 vdd.n3253 vss 0.00425f
C3911 vdd.n3254 vss 0.0424f
C3912 vdd.n3255 vss 0.0132f
C3913 vdd.n3256 vss 0.00324f
C3914 vdd.n3257 vss 0.0128f
C3915 vdd.n3258 vss 0.02f
C3916 vdd.n3259 vss 0.00425f
C3917 vdd.n3260 vss 0.00413f
C3918 vdd.n3261 vss 0.00251f
C3919 vdd.n3262 vss 0.0471f
C3920 vdd.n3263 vss 0.00251f
C3921 vdd.n3264 vss 0.00517f
C3922 vdd.n3265 vss 0.00679f
C3923 vdd.n3266 vss 0.00324f
C3924 vdd.n3267 vss 0.00324f
C3925 vdd.n3268 vss 0.0132f
C3926 vdd.n3269 vss 0.0424f
C3927 vdd.n3270 vss 0.02f
C3928 vdd.n3271 vss 0.00425f
C3929 vdd.n3272 vss 0.0471f
C3930 vdd.n3274 vss 0.00425f
C3931 vdd.n3275 vss 0.00925f
C3932 vdd.n3276 vss 0.00679f
C3933 vdd.n3277 vss 0.00517f
C3934 vdd.n3278 vss 0.00251f
C3935 vdd.n3279 vss 0.0471f
C3936 vdd.n3280 vss 0.00251f
C3937 vdd.n3281 vss 0.0112f
C3938 vdd.n3282 vss 0.0128f
C3939 vdd.n3283 vss 0.146f
C3940 vdd.n3284 vss 0.0596f
C3941 vdd.n3285 vss 0.00324f
C3942 vdd.n3286 vss 0.0112f
C3943 vdd.n3287 vss 0.0128f
C3944 vdd.n3288 vss 0.00413f
C3945 vdd.n3289 vss 0.00413f
C3946 vdd.n3290 vss 0.0471f
C3947 vdd.n3291 vss 0.0471f
C3948 vdd.n3292 vss 0.00324f
C3949 vdd.n3293 vss 0.00413f
C3950 vdd.n3294 vss 0.00413f
C3951 vdd.n3295 vss 0.00679f
C3952 vdd.n3296 vss 0.00413f
C3953 vdd.n3297 vss 0.0471f
C3954 vdd.n3298 vss 0.00324f
C3955 vdd.n3300 vss 0.00925f
C3956 vdd.n3301 vss 0.0471f
C3957 vdd.n3302 vss 0.00425f
C3958 vdd.n3303 vss 0.0424f
C3959 vdd.n3304 vss 0.0132f
C3960 vdd.n3305 vss 0.00324f
C3961 vdd.n3306 vss 0.0128f
C3962 vdd.n3307 vss 0.02f
C3963 vdd.n3308 vss 0.00425f
C3964 vdd.n3309 vss 0.00413f
C3965 vdd.n3310 vss 0.00251f
C3966 vdd.n3311 vss 0.0471f
C3967 vdd.n3312 vss 0.00251f
C3968 vdd.n3313 vss 0.00517f
C3969 vdd.n3314 vss 0.00679f
C3970 vdd.n3315 vss 0.00324f
C3971 vdd.n3316 vss 0.00324f
C3972 vdd.n3317 vss 0.0132f
C3973 vdd.n3318 vss 0.0424f
C3974 vdd.n3319 vss 0.02f
C3975 vdd.n3320 vss 0.00425f
C3976 vdd.n3321 vss 0.0471f
C3977 vdd.n3323 vss 0.00425f
C3978 vdd.n3324 vss 0.00925f
C3979 vdd.n3325 vss 0.00679f
C3980 vdd.n3326 vss 0.00517f
C3981 vdd.n3327 vss 0.00251f
C3982 vdd.n3328 vss 0.0471f
C3983 vdd.n3329 vss 0.00251f
C3984 vdd.n3330 vss 0.0112f
C3985 vdd.n3331 vss 0.0128f
C3986 vdd.n3332 vss 0.0692f
C3987 vdd.n3333 vss 0.118f
C3988 vdd.n3334 vss 0.121f
C3989 vdd.n3335 vss 0.00324f
C3990 vdd.n3336 vss 0.0112f
C3991 vdd.n3337 vss 0.0128f
C3992 vdd.n3338 vss 0.00413f
C3993 vdd.n3339 vss 0.00413f
C3994 vdd.n3340 vss 0.0471f
C3995 vdd.n3341 vss 0.0471f
C3996 vdd.n3342 vss 0.00324f
C3997 vdd.n3343 vss 0.00413f
C3998 vdd.n3344 vss 0.00413f
C3999 vdd.n3345 vss 0.00679f
C4000 vdd.n3346 vss 0.00413f
C4001 vdd.n3347 vss 0.0471f
C4002 vdd.n3348 vss 0.00324f
C4003 vdd.n3350 vss 0.00925f
C4004 vdd.n3351 vss 0.0471f
C4005 vdd.n3352 vss 0.00425f
C4006 vdd.n3353 vss 0.0424f
C4007 vdd.n3354 vss 0.0132f
C4008 vdd.n3355 vss 0.00324f
C4009 vdd.n3356 vss 0.0128f
C4010 vdd.n3357 vss 0.02f
C4011 vdd.n3358 vss 0.00425f
C4012 vdd.n3359 vss 0.00413f
C4013 vdd.n3360 vss 0.00251f
C4014 vdd.n3361 vss 0.0471f
C4015 vdd.n3362 vss 0.00251f
C4016 vdd.n3363 vss 0.00517f
C4017 vdd.n3364 vss 0.00679f
C4018 vdd.n3365 vss 0.00324f
C4019 vdd.n3366 vss 0.00324f
C4020 vdd.n3367 vss 0.0132f
C4021 vdd.n3368 vss 0.0424f
C4022 vdd.n3369 vss 0.02f
C4023 vdd.n3370 vss 0.00425f
C4024 vdd.n3371 vss 0.0471f
C4025 vdd.n3373 vss 0.00425f
C4026 vdd.n3374 vss 0.00925f
C4027 vdd.n3375 vss 0.00679f
C4028 vdd.n3376 vss 0.00517f
C4029 vdd.n3377 vss 0.00251f
C4030 vdd.n3378 vss 0.0471f
C4031 vdd.n3379 vss 0.00251f
C4032 vdd.n3380 vss 0.0112f
C4033 vdd.n3381 vss 0.098f
C4034 vdd.n3382 vss 0.0596f
C4035 vdd.n3383 vss 0.00324f
C4036 vdd.n3384 vss 0.0112f
C4037 vdd.n3385 vss 0.0128f
C4038 vdd.n3386 vss 0.00413f
C4039 vdd.n3387 vss 0.00413f
C4040 vdd.n3388 vss 0.0471f
C4041 vdd.n3389 vss 0.0471f
C4042 vdd.n3390 vss 0.00324f
C4043 vdd.n3391 vss 0.00413f
C4044 vdd.n3392 vss 0.00413f
C4045 vdd.n3393 vss 0.00679f
C4046 vdd.n3394 vss 0.00413f
C4047 vdd.n3395 vss 0.0471f
C4048 vdd.n3396 vss 0.00324f
C4049 vdd.n3398 vss 0.00925f
C4050 vdd.n3399 vss 0.0471f
C4051 vdd.n3400 vss 0.00425f
C4052 vdd.n3401 vss 0.0424f
C4053 vdd.n3402 vss 0.0132f
C4054 vdd.n3403 vss 0.00324f
C4055 vdd.n3404 vss 0.0128f
C4056 vdd.n3405 vss 0.02f
C4057 vdd.n3406 vss 0.00425f
C4058 vdd.n3407 vss 0.00413f
C4059 vdd.n3408 vss 0.00251f
C4060 vdd.n3409 vss 0.0471f
C4061 vdd.n3410 vss 0.00251f
C4062 vdd.n3411 vss 0.00517f
C4063 vdd.n3412 vss 0.00679f
C4064 vdd.n3413 vss 0.00324f
C4065 vdd.n3414 vss 0.00324f
C4066 vdd.n3415 vss 0.0132f
C4067 vdd.n3416 vss 0.0424f
C4068 vdd.n3417 vss 0.02f
C4069 vdd.n3418 vss 0.00425f
C4070 vdd.n3419 vss 0.0471f
C4071 vdd.n3421 vss 0.00425f
C4072 vdd.n3422 vss 0.00925f
C4073 vdd.n3423 vss 0.00679f
C4074 vdd.n3424 vss 0.00517f
C4075 vdd.n3425 vss 0.00251f
C4076 vdd.n3426 vss 0.0471f
C4077 vdd.n3427 vss 0.00251f
C4078 vdd.n3428 vss 0.0112f
C4079 vdd.n3429 vss 0.0128f
C4080 vdd.n3430 vss 0.0692f
C4081 vdd.n3431 vss 0.0912f
C4082 vdd.n3432 vss 0.0824f
C4083 vdd.n3433 vss 0.059f
C4084 vdd.n3434 vss 0.00324f
C4085 vdd.n3435 vss 0.0112f
C4086 vdd.n3436 vss 0.0128f
C4087 vdd.n3437 vss 0.00413f
C4088 vdd.n3438 vss 0.00413f
C4089 vdd.n3439 vss 0.0471f
C4090 vdd.n3440 vss 0.0471f
C4091 vdd.n3441 vss 0.00324f
C4092 vdd.n3442 vss 0.00413f
C4093 vdd.n3443 vss 0.00413f
C4094 vdd.n3444 vss 0.00679f
C4095 vdd.n3445 vss 0.00413f
C4096 vdd.n3446 vss 0.0471f
C4097 vdd.n3447 vss 0.00324f
C4098 vdd.n3449 vss 0.00925f
C4099 vdd.n3450 vss 0.0471f
C4100 vdd.n3451 vss 0.00425f
C4101 vdd.n3452 vss 0.0424f
C4102 vdd.n3453 vss 0.0132f
C4103 vdd.n3454 vss 0.00324f
C4104 vdd.n3455 vss 0.0128f
C4105 vdd.n3456 vss 0.02f
C4106 vdd.n3457 vss 0.00425f
C4107 vdd.n3458 vss 0.00413f
C4108 vdd.n3459 vss 0.00251f
C4109 vdd.n3460 vss 0.0471f
C4110 vdd.n3461 vss 0.00251f
C4111 vdd.n3462 vss 0.00517f
C4112 vdd.n3463 vss 0.00679f
C4113 vdd.n3464 vss 0.00324f
C4114 vdd.n3465 vss 0.00324f
C4115 vdd.n3466 vss 0.0132f
C4116 vdd.n3467 vss 0.0424f
C4117 vdd.n3468 vss 0.02f
C4118 vdd.n3469 vss 0.00425f
C4119 vdd.n3470 vss 0.0471f
C4120 vdd.n3472 vss 0.00425f
C4121 vdd.n3473 vss 0.00925f
C4122 vdd.n3474 vss 0.00679f
C4123 vdd.n3475 vss 0.00517f
C4124 vdd.n3476 vss 0.00251f
C4125 vdd.n3477 vss 0.0471f
C4126 vdd.n3478 vss 0.00251f
C4127 vdd.n3479 vss 0.0112f
C4128 vdd.n3480 vss 0.0128f
C4129 vdd.n3481 vss 0.146f
C4130 vdd.n3482 vss 0.00324f
C4131 vdd.n3483 vss 0.0112f
C4132 vdd.n3484 vss 0.0128f
C4133 vdd.n3485 vss 0.00413f
C4134 vdd.n3486 vss 0.00413f
C4135 vdd.n3487 vss 0.0471f
C4136 vdd.n3488 vss 0.0471f
C4137 vdd.n3489 vss 0.00324f
C4138 vdd.n3490 vss 0.00413f
C4139 vdd.n3491 vss 0.00413f
C4140 vdd.n3492 vss 0.00679f
C4141 vdd.n3493 vss 0.00413f
C4142 vdd.n3494 vss 0.0471f
C4143 vdd.n3495 vss 0.00324f
C4144 vdd.n3497 vss 0.00925f
C4145 vdd.n3498 vss 0.0471f
C4146 vdd.n3499 vss 0.00425f
C4147 vdd.n3500 vss 0.0424f
C4148 vdd.n3501 vss 0.0132f
C4149 vdd.n3502 vss 0.00324f
C4150 vdd.n3503 vss 0.0128f
C4151 vdd.n3504 vss 0.02f
C4152 vdd.n3505 vss 0.00425f
C4153 vdd.n3506 vss 0.00413f
C4154 vdd.n3507 vss 0.00251f
C4155 vdd.n3508 vss 0.0471f
C4156 vdd.n3509 vss 0.00251f
C4157 vdd.n3510 vss 0.00517f
C4158 vdd.n3511 vss 0.00679f
C4159 vdd.n3512 vss 0.00324f
C4160 vdd.n3513 vss 0.00324f
C4161 vdd.n3514 vss 0.0132f
C4162 vdd.n3515 vss 0.0424f
C4163 vdd.n3516 vss 0.02f
C4164 vdd.n3517 vss 0.00425f
C4165 vdd.n3518 vss 0.0471f
C4166 vdd.n3520 vss 0.00425f
C4167 vdd.n3521 vss 0.00925f
C4168 vdd.n3522 vss 0.00679f
C4169 vdd.n3523 vss 0.00517f
C4170 vdd.n3524 vss 0.00251f
C4171 vdd.n3525 vss 0.0471f
C4172 vdd.n3526 vss 0.00251f
C4173 vdd.n3527 vss 0.0112f
C4174 vdd.n3528 vss 0.0128f
C4175 vdd.n3529 vss 0.146f
C4176 vdd.n3530 vss 0.0596f
C4177 vdd.n3531 vss 0.00324f
C4178 vdd.n3532 vss 0.0112f
C4179 vdd.n3533 vss 0.0128f
C4180 vdd.n3534 vss 0.00413f
C4181 vdd.n3535 vss 0.00413f
C4182 vdd.n3536 vss 0.0471f
C4183 vdd.n3537 vss 0.0471f
C4184 vdd.n3538 vss 0.00324f
C4185 vdd.n3539 vss 0.00413f
C4186 vdd.n3540 vss 0.00413f
C4187 vdd.n3541 vss 0.00679f
C4188 vdd.n3542 vss 0.00413f
C4189 vdd.n3543 vss 0.0471f
C4190 vdd.n3544 vss 0.00324f
C4191 vdd.n3546 vss 0.00925f
C4192 vdd.n3547 vss 0.0471f
C4193 vdd.n3548 vss 0.00425f
C4194 vdd.n3549 vss 0.0424f
C4195 vdd.n3550 vss 0.0132f
C4196 vdd.n3551 vss 0.00324f
C4197 vdd.n3552 vss 0.0128f
C4198 vdd.n3553 vss 0.02f
C4199 vdd.n3554 vss 0.00425f
C4200 vdd.n3555 vss 0.00413f
C4201 vdd.n3556 vss 0.00251f
C4202 vdd.n3557 vss 0.0471f
C4203 vdd.n3558 vss 0.00251f
C4204 vdd.n3559 vss 0.00517f
C4205 vdd.n3560 vss 0.00679f
C4206 vdd.n3561 vss 0.00324f
C4207 vdd.n3562 vss 0.00324f
C4208 vdd.n3563 vss 0.0132f
C4209 vdd.n3564 vss 0.0424f
C4210 vdd.n3565 vss 0.02f
C4211 vdd.n3566 vss 0.00425f
C4212 vdd.n3567 vss 0.0471f
C4213 vdd.n3569 vss 0.00425f
C4214 vdd.n3570 vss 0.00925f
C4215 vdd.n3571 vss 0.00679f
C4216 vdd.n3572 vss 0.00517f
C4217 vdd.n3573 vss 0.00251f
C4218 vdd.n3574 vss 0.0471f
C4219 vdd.n3575 vss 0.00251f
C4220 vdd.n3576 vss 0.0112f
C4221 vdd.n3577 vss 0.0128f
C4222 vdd.n3578 vss 0.0692f
C4223 vdd.n3579 vss 0.118f
C4224 vdd.n3580 vss 0.121f
C4225 vdd.n3581 vss 0.00324f
C4226 vdd.n3582 vss 0.0112f
C4227 vdd.n3583 vss 0.0128f
C4228 vdd.n3584 vss 0.00413f
C4229 vdd.n3585 vss 0.00413f
C4230 vdd.n3586 vss 0.0471f
C4231 vdd.n3587 vss 0.0471f
C4232 vdd.n3588 vss 0.00324f
C4233 vdd.n3589 vss 0.00413f
C4234 vdd.n3590 vss 0.00413f
C4235 vdd.n3591 vss 0.00679f
C4236 vdd.n3592 vss 0.00413f
C4237 vdd.n3593 vss 0.0471f
C4238 vdd.n3594 vss 0.00324f
C4239 vdd.n3596 vss 0.00925f
C4240 vdd.n3597 vss 0.0471f
C4241 vdd.n3598 vss 0.00425f
C4242 vdd.n3599 vss 0.0424f
C4243 vdd.n3600 vss 0.0132f
C4244 vdd.n3601 vss 0.00324f
C4245 vdd.n3602 vss 0.0128f
C4246 vdd.n3603 vss 0.02f
C4247 vdd.n3604 vss 0.00425f
C4248 vdd.n3605 vss 0.00413f
C4249 vdd.n3606 vss 0.00251f
C4250 vdd.n3607 vss 0.0471f
C4251 vdd.n3608 vss 0.00251f
C4252 vdd.n3609 vss 0.00517f
C4253 vdd.n3610 vss 0.00679f
C4254 vdd.n3611 vss 0.00324f
C4255 vdd.n3612 vss 0.00324f
C4256 vdd.n3613 vss 0.0132f
C4257 vdd.n3614 vss 0.0424f
C4258 vdd.n3615 vss 0.02f
C4259 vdd.n3616 vss 0.00425f
C4260 vdd.n3617 vss 0.0471f
C4261 vdd.n3619 vss 0.00425f
C4262 vdd.n3620 vss 0.00925f
C4263 vdd.n3621 vss 0.00679f
C4264 vdd.n3622 vss 0.00517f
C4265 vdd.n3623 vss 0.00251f
C4266 vdd.n3624 vss 0.0471f
C4267 vdd.n3625 vss 0.00251f
C4268 vdd.n3626 vss 0.0112f
C4269 vdd.n3627 vss 0.098f
C4270 vdd.n3628 vss 0.0596f
C4271 vdd.n3629 vss 0.00324f
C4272 vdd.n3630 vss 0.0112f
C4273 vdd.n3631 vss 0.0128f
C4274 vdd.n3632 vss 0.00413f
C4275 vdd.n3633 vss 0.00413f
C4276 vdd.n3634 vss 0.0471f
C4277 vdd.n3635 vss 0.0471f
C4278 vdd.n3636 vss 0.00324f
C4279 vdd.n3637 vss 0.00413f
C4280 vdd.n3638 vss 0.00413f
C4281 vdd.n3639 vss 0.00679f
C4282 vdd.n3640 vss 0.00413f
C4283 vdd.n3641 vss 0.0471f
C4284 vdd.n3642 vss 0.00324f
C4285 vdd.n3644 vss 0.00925f
C4286 vdd.n3645 vss 0.0471f
C4287 vdd.n3646 vss 0.00425f
C4288 vdd.n3647 vss 0.0424f
C4289 vdd.n3648 vss 0.0132f
C4290 vdd.n3649 vss 0.00324f
C4291 vdd.n3650 vss 0.0128f
C4292 vdd.n3651 vss 0.02f
C4293 vdd.n3652 vss 0.00425f
C4294 vdd.n3653 vss 0.00413f
C4295 vdd.n3654 vss 0.00251f
C4296 vdd.n3655 vss 0.0471f
C4297 vdd.n3656 vss 0.00251f
C4298 vdd.n3657 vss 0.00517f
C4299 vdd.n3658 vss 0.00679f
C4300 vdd.n3659 vss 0.00324f
C4301 vdd.n3660 vss 0.00324f
C4302 vdd.n3661 vss 0.0132f
C4303 vdd.n3662 vss 0.0424f
C4304 vdd.n3663 vss 0.02f
C4305 vdd.n3664 vss 0.00425f
C4306 vdd.n3665 vss 0.0471f
C4307 vdd.n3667 vss 0.00425f
C4308 vdd.n3668 vss 0.00925f
C4309 vdd.n3669 vss 0.00679f
C4310 vdd.n3670 vss 0.00517f
C4311 vdd.n3671 vss 0.00251f
C4312 vdd.n3672 vss 0.0471f
C4313 vdd.n3673 vss 0.00251f
C4314 vdd.n3674 vss 0.0112f
C4315 vdd.n3675 vss 0.0128f
C4316 vdd.n3676 vss 0.0692f
C4317 vdd.n3677 vss 0.121f
C4318 vdd.n3678 vss 0.291f
C4319 vdd.n3679 vss 0.227f
C4320 vdd.n3680 vss 0.00324f
C4321 vdd.n3681 vss 0.0112f
C4322 vdd.n3682 vss 0.0128f
C4323 vdd.n3683 vss 0.00413f
C4324 vdd.n3684 vss 0.00413f
C4325 vdd.n3685 vss 0.0471f
C4326 vdd.n3686 vss 0.0471f
C4327 vdd.n3687 vss 0.00324f
C4328 vdd.n3688 vss 0.00413f
C4329 vdd.n3689 vss 0.00413f
C4330 vdd.n3690 vss 0.00679f
C4331 vdd.n3691 vss 0.00413f
C4332 vdd.n3692 vss 0.0471f
C4333 vdd.n3693 vss 0.00324f
C4334 vdd.n3695 vss 0.00925f
C4335 vdd.n3696 vss 0.0471f
C4336 vdd.n3697 vss 0.00425f
C4337 vdd.n3698 vss 0.0424f
C4338 vdd.n3699 vss 0.0132f
C4339 vdd.n3700 vss 0.00324f
C4340 vdd.n3701 vss 0.0128f
C4341 vdd.n3702 vss 0.02f
C4342 vdd.n3703 vss 0.00425f
C4343 vdd.n3704 vss 0.00413f
C4344 vdd.n3705 vss 0.00251f
C4345 vdd.n3706 vss 0.0471f
C4346 vdd.n3707 vss 0.00251f
C4347 vdd.n3708 vss 0.00517f
C4348 vdd.n3709 vss 0.00679f
C4349 vdd.n3710 vss 0.00324f
C4350 vdd.n3711 vss 0.00324f
C4351 vdd.n3712 vss 0.0132f
C4352 vdd.n3713 vss 0.0424f
C4353 vdd.n3714 vss 0.02f
C4354 vdd.n3715 vss 0.00425f
C4355 vdd.n3716 vss 0.0471f
C4356 vdd.n3718 vss 0.00425f
C4357 vdd.n3719 vss 0.00925f
C4358 vdd.n3720 vss 0.00679f
C4359 vdd.n3721 vss 0.00517f
C4360 vdd.n3722 vss 0.00251f
C4361 vdd.n3723 vss 0.0471f
C4362 vdd.n3724 vss 0.00251f
C4363 vdd.n3725 vss 0.0112f
C4364 vdd.n3726 vss 0.0128f
C4365 vdd.n3727 vss 0.18f
C4366 vdd.n3728 vss 0.00324f
C4367 vdd.n3729 vss 0.0112f
C4368 vdd.n3730 vss 0.0128f
C4369 vdd.n3731 vss 0.00413f
C4370 vdd.n3732 vss 0.00413f
C4371 vdd.n3733 vss 0.0471f
C4372 vdd.n3734 vss 0.0471f
C4373 vdd.n3735 vss 0.00324f
C4374 vdd.n3736 vss 0.00413f
C4375 vdd.n3737 vss 0.00413f
C4376 vdd.n3738 vss 0.00679f
C4377 vdd.n3739 vss 0.00413f
C4378 vdd.n3740 vss 0.0471f
C4379 vdd.n3741 vss 0.00324f
C4380 vdd.n3743 vss 0.00925f
C4381 vdd.n3744 vss 0.0471f
C4382 vdd.n3745 vss 0.00425f
C4383 vdd.n3746 vss 0.0424f
C4384 vdd.n3747 vss 0.0132f
C4385 vdd.n3748 vss 0.00324f
C4386 vdd.n3749 vss 0.0128f
C4387 vdd.n3750 vss 0.02f
C4388 vdd.n3751 vss 0.00425f
C4389 vdd.n3752 vss 0.00413f
C4390 vdd.n3753 vss 0.00251f
C4391 vdd.n3754 vss 0.0471f
C4392 vdd.n3755 vss 0.00251f
C4393 vdd.n3756 vss 0.00517f
C4394 vdd.n3757 vss 0.00679f
C4395 vdd.n3758 vss 0.00324f
C4396 vdd.n3759 vss 0.00324f
C4397 vdd.n3760 vss 0.0132f
C4398 vdd.n3761 vss 0.0424f
C4399 vdd.n3762 vss 0.02f
C4400 vdd.n3763 vss 0.00425f
C4401 vdd.n3764 vss 0.0471f
C4402 vdd.n3766 vss 0.00425f
C4403 vdd.n3767 vss 0.00925f
C4404 vdd.n3768 vss 0.00679f
C4405 vdd.n3769 vss 0.00517f
C4406 vdd.n3770 vss 0.00251f
C4407 vdd.n3771 vss 0.0471f
C4408 vdd.n3772 vss 0.00251f
C4409 vdd.n3773 vss 0.0112f
C4410 vdd.n3774 vss 0.0128f
C4411 vdd.n3775 vss 0.248f
C4412 vdd.n3776 vss 0.00324f
C4413 vdd.n3777 vss 0.0112f
C4414 vdd.n3778 vss 0.0128f
C4415 vdd.n3779 vss 0.00413f
C4416 vdd.n3780 vss 0.00413f
C4417 vdd.n3781 vss 0.0471f
C4418 vdd.n3782 vss 0.0471f
C4419 vdd.n3783 vss 0.00324f
C4420 vdd.n3784 vss 0.00413f
C4421 vdd.n3785 vss 0.00413f
C4422 vdd.n3786 vss 0.00679f
C4423 vdd.n3787 vss 0.00413f
C4424 vdd.n3788 vss 0.0471f
C4425 vdd.n3789 vss 0.00324f
C4426 vdd.n3790 vss 0.0424f
C4427 vdd.n3791 vss 0.00324f
C4428 vdd.n3792 vss 0.0128f
C4429 vdd.n3793 vss 0.02f
C4430 vdd.n3794 vss 0.0132f
C4431 vdd.n3795 vss 0.00925f
C4432 vdd.n3796 vss 0.00425f
C4433 vdd.n3798 vss 0.0471f
C4434 vdd.n3799 vss 0.00425f
C4435 vdd.n3800 vss 0.00413f
C4436 vdd.n3801 vss 0.00251f
C4437 vdd.n3802 vss 0.0471f
C4438 vdd.n3803 vss 0.00251f
C4439 vdd.n3804 vss 0.00517f
C4440 vdd.n3805 vss 0.00679f
C4441 vdd.n3806 vss 0.00324f
C4442 vdd.n3807 vss 0.00324f
C4443 vdd.n3808 vss 0.0132f
C4444 vdd.n3809 vss 0.0424f
C4445 vdd.n3810 vss 0.02f
C4446 vdd.n3811 vss 0.00425f
C4447 vdd.n3813 vss 0.0471f
C4448 vdd.n3814 vss 0.00425f
C4449 vdd.n3815 vss 0.00925f
C4450 vdd.n3816 vss 0.00679f
C4451 vdd.n3817 vss 0.00517f
C4452 vdd.n3818 vss 0.00251f
C4453 vdd.n3819 vss 0.0471f
C4454 vdd.n3820 vss 0.00251f
C4455 vdd.n3821 vss 0.0112f
C4456 vdd.n3822 vss 0.0128f
C4457 vdd.n3823 vss 0.0599f
C4458 vdd.n3824 vss 0.202f
C4459 vdd.n3825 vss 0.00324f
C4460 vdd.n3826 vss 0.0112f
C4461 vdd.n3827 vss 0.0128f
C4462 vdd.n3828 vss 0.00413f
C4463 vdd.n3829 vss 0.00413f
C4464 vdd.n3830 vss 0.0471f
C4465 vdd.n3831 vss 0.0471f
C4466 vdd.n3832 vss 0.00324f
C4467 vdd.n3833 vss 0.00413f
C4468 vdd.n3834 vss 0.00413f
C4469 vdd.n3835 vss 0.00679f
C4470 vdd.n3836 vss 0.00413f
C4471 vdd.n3837 vss 0.0471f
C4472 vdd.n3838 vss 0.00324f
C4473 vdd.n3840 vss 0.00925f
C4474 vdd.n3841 vss 0.0471f
C4475 vdd.n3842 vss 0.00425f
C4476 vdd.n3843 vss 0.0424f
C4477 vdd.n3844 vss 0.0132f
C4478 vdd.n3845 vss 0.00324f
C4479 vdd.n3846 vss 0.0128f
C4480 vdd.n3847 vss 0.02f
C4481 vdd.n3848 vss 0.00425f
C4482 vdd.n3849 vss 0.00413f
C4483 vdd.n3850 vss 0.00251f
C4484 vdd.n3851 vss 0.0471f
C4485 vdd.n3852 vss 0.00251f
C4486 vdd.n3853 vss 0.00517f
C4487 vdd.n3854 vss 0.00679f
C4488 vdd.n3855 vss 0.00324f
C4489 vdd.n3856 vss 0.00324f
C4490 vdd.n3857 vss 0.0132f
C4491 vdd.n3858 vss 0.0424f
C4492 vdd.n3859 vss 0.02f
C4493 vdd.n3860 vss 0.00425f
C4494 vdd.n3861 vss 0.0471f
C4495 vdd.n3863 vss 0.00425f
C4496 vdd.n3864 vss 0.00925f
C4497 vdd.n3865 vss 0.00679f
C4498 vdd.n3866 vss 0.00517f
C4499 vdd.n3867 vss 0.00251f
C4500 vdd.n3868 vss 0.0471f
C4501 vdd.n3869 vss 0.00251f
C4502 vdd.n3870 vss 0.0112f
C4503 vdd.n3871 vss 0.0128f
C4504 vdd.n3872 vss 0.0692f
C4505 vdd.n3873 vss 0.00324f
C4506 vdd.n3874 vss 0.0112f
C4507 vdd.n3875 vss 0.0128f
C4508 vdd.n3876 vss 0.00413f
C4509 vdd.n3877 vss 0.00413f
C4510 vdd.n3878 vss 0.0471f
C4511 vdd.n3879 vss 0.0471f
C4512 vdd.n3880 vss 0.00324f
C4513 vdd.n3881 vss 0.00413f
C4514 vdd.n3882 vss 0.00413f
C4515 vdd.n3883 vss 0.00679f
C4516 vdd.n3884 vss 0.00413f
C4517 vdd.n3885 vss 0.0471f
C4518 vdd.n3886 vss 0.00324f
C4519 vdd.n3888 vss 0.00925f
C4520 vdd.n3889 vss 0.0471f
C4521 vdd.n3890 vss 0.00425f
C4522 vdd.n3891 vss 0.0424f
C4523 vdd.n3892 vss 0.0132f
C4524 vdd.n3893 vss 0.00324f
C4525 vdd.n3894 vss 0.0128f
C4526 vdd.n3895 vss 0.02f
C4527 vdd.n3896 vss 0.00425f
C4528 vdd.n3897 vss 0.00413f
C4529 vdd.n3898 vss 0.00251f
C4530 vdd.n3899 vss 0.0471f
C4531 vdd.n3900 vss 0.00251f
C4532 vdd.n3901 vss 0.00517f
C4533 vdd.n3902 vss 0.00679f
C4534 vdd.n3903 vss 0.00324f
C4535 vdd.n3904 vss 0.00324f
C4536 vdd.n3905 vss 0.0132f
C4537 vdd.n3906 vss 0.0424f
C4538 vdd.n3907 vss 0.02f
C4539 vdd.n3908 vss 0.00425f
C4540 vdd.n3909 vss 0.0471f
C4541 vdd.n3911 vss 0.00425f
C4542 vdd.n3912 vss 0.00925f
C4543 vdd.n3913 vss 0.00679f
C4544 vdd.n3914 vss 0.00517f
C4545 vdd.n3915 vss 0.00251f
C4546 vdd.n3916 vss 0.0471f
C4547 vdd.n3917 vss 0.00251f
C4548 vdd.n3918 vss 0.0112f
C4549 vdd.n3919 vss 0.0128f
C4550 vdd.n3920 vss 0.0619f
C4551 vdd.n3921 vss 0.00335f
C4552 vdd.n3922 vss 0.0855f
C4553 vdd.n3923 vss 0.00991f
C4554 vdd.n3924 vss 0.0424f
C4555 vdd.n3925 vss 0.00679f
C4556 vdd.n3926 vss 0.00413f
C4557 vdd.n3927 vss 0.0471f
C4558 vdd.n3928 vss 0.00251f
C4559 vdd.n3929 vss 0.00679f
C4560 vdd.n3930 vss 0.00413f
C4561 vdd.n3931 vss 0.00413f
C4562 vdd.n3932 vss 0.0471f
C4563 vdd.n3933 vss 0.00251f
C4564 vdd.n3934 vss 0.00413f
C4565 vdd.n3935 vss 0.00324f
C4566 vdd.n3936 vss 0.0132f
C4567 vdd.n3937 vss 0.0424f
C4568 vdd.n3938 vss 0.00324f
C4569 vdd.n3939 vss 0.00413f
C4570 vdd.n3940 vss 0.00517f
C4571 vdd.n3941 vss 0.00679f
C4572 vdd.n3942 vss 0.00925f
C4573 vdd.n3943 vss 0.00425f
C4574 vdd.n3944 vss 0.0471f
C4575 vdd.n3946 vss 0.00425f
C4576 vdd.n3947 vss 0.02f
C4577 vdd.n3948 vss 0.0128f
C4578 vdd.n3949 vss 0.0105f
C4579 vdd.n3950 vss 0.00251f
C4580 vdd.n3951 vss 0.0471f
C4581 vdd.n3952 vss 0.00517f
C4582 vdd.n3953 vss 0.00251f
C4583 vdd.n3954 vss 0.0471f
C4584 vdd.n3955 vss 0.0471f
C4585 vdd.n3956 vss 0.00324f
C4586 vdd.n3957 vss 0.00324f
C4587 vdd.n3958 vss 0.00805f
C4588 vdd.n3959 vss 0.0112f
C4589 vdd.n3960 vss 0.0128f
C4590 vdd.n3961 vss 0.00324f
C4591 vdd.n3962 vss 0.00324f
C4592 vdd.n3963 vss 0.00413f
C4593 vdd.n3964 vss 0.00425f
C4594 vdd.n3965 vss 0.0471f
C4595 vdd.n3967 vss 0.00425f
C4596 vdd.n3968 vss 0.00925f
C4597 vdd.n3969 vss 0.0107f
C4598 vdd.n3970 vss 0.0126f
C4599 vdd.n3971 vss 0.0516f
C4600 vdd.n3972 vss 0.00163f
C4601 vdd.n3973 vss 0.00145f
C4602 vdd.n3974 vss 0.0271f
C4603 vdd.n3975 vss 0.00324f
C4604 vdd.n3976 vss 0.0112f
C4605 vdd.n3977 vss 0.0128f
C4606 vdd.n3978 vss 0.00413f
C4607 vdd.n3979 vss 0.00413f
C4608 vdd.n3980 vss 0.0471f
C4609 vdd.n3981 vss 0.0471f
C4610 vdd.n3982 vss 0.00324f
C4611 vdd.n3983 vss 0.00413f
C4612 vdd.n3984 vss 0.00413f
C4613 vdd.n3985 vss 0.00679f
C4614 vdd.n3986 vss 0.00413f
C4615 vdd.n3987 vss 0.0471f
C4616 vdd.n3988 vss 0.00324f
C4617 vdd.n3990 vss 0.00925f
C4618 vdd.n3991 vss 0.0471f
C4619 vdd.n3992 vss 0.00425f
C4620 vdd.n3993 vss 0.0424f
C4621 vdd.n3994 vss 0.0132f
C4622 vdd.n3995 vss 0.00324f
C4623 vdd.n3996 vss 0.0128f
C4624 vdd.n3997 vss 0.02f
C4625 vdd.n3998 vss 0.00425f
C4626 vdd.n3999 vss 0.00413f
C4627 vdd.n4000 vss 0.00251f
C4628 vdd.n4001 vss 0.0471f
C4629 vdd.n4002 vss 0.00251f
C4630 vdd.n4003 vss 0.00517f
C4631 vdd.n4004 vss 0.00679f
C4632 vdd.n4005 vss 0.00324f
C4633 vdd.n4006 vss 0.00324f
C4634 vdd.n4007 vss 0.0132f
C4635 vdd.n4008 vss 0.0424f
C4636 vdd.n4009 vss 0.02f
C4637 vdd.n4010 vss 0.00425f
C4638 vdd.n4011 vss 0.0471f
C4639 vdd.n4013 vss 0.00425f
C4640 vdd.n4014 vss 0.00925f
C4641 vdd.n4015 vss 0.00679f
C4642 vdd.n4016 vss 0.00517f
C4643 vdd.n4017 vss 0.00251f
C4644 vdd.n4018 vss 0.0471f
C4645 vdd.n4019 vss 0.00251f
C4646 vdd.n4020 vss 0.0112f
C4647 vdd.n4021 vss 0.0128f
C4648 vdd.n4022 vss 0.0692f
C4649 vdd.n4023 vss 0.00324f
C4650 vdd.n4024 vss 0.0112f
C4651 vdd.n4025 vss 0.0128f
C4652 vdd.n4026 vss 0.00413f
C4653 vdd.n4027 vss 0.00413f
C4654 vdd.n4028 vss 0.0471f
C4655 vdd.n4029 vss 0.0471f
C4656 vdd.n4030 vss 0.00324f
C4657 vdd.n4031 vss 0.00413f
C4658 vdd.n4032 vss 0.00413f
C4659 vdd.n4033 vss 0.00679f
C4660 vdd.n4034 vss 0.00413f
C4661 vdd.n4035 vss 0.0471f
C4662 vdd.n4036 vss 0.00324f
C4663 vdd.n4038 vss 0.00925f
C4664 vdd.n4039 vss 0.0471f
C4665 vdd.n4040 vss 0.00425f
C4666 vdd.n4041 vss 0.0424f
C4667 vdd.n4042 vss 0.0132f
C4668 vdd.n4043 vss 0.00324f
C4669 vdd.n4044 vss 0.0128f
C4670 vdd.n4045 vss 0.02f
C4671 vdd.n4046 vss 0.00425f
C4672 vdd.n4047 vss 0.00413f
C4673 vdd.n4048 vss 0.00251f
C4674 vdd.n4049 vss 0.0471f
C4675 vdd.n4050 vss 0.00251f
C4676 vdd.n4051 vss 0.00517f
C4677 vdd.n4052 vss 0.00679f
C4678 vdd.n4053 vss 0.00324f
C4679 vdd.n4054 vss 0.00324f
C4680 vdd.n4055 vss 0.0132f
C4681 vdd.n4056 vss 0.0424f
C4682 vdd.n4057 vss 0.02f
C4683 vdd.n4058 vss 0.00425f
C4684 vdd.n4059 vss 0.0471f
C4685 vdd.n4061 vss 0.00425f
C4686 vdd.n4062 vss 0.00925f
C4687 vdd.n4063 vss 0.00679f
C4688 vdd.n4064 vss 0.00517f
C4689 vdd.n4065 vss 0.00251f
C4690 vdd.n4066 vss 0.0471f
C4691 vdd.n4067 vss 0.00251f
C4692 vdd.n4068 vss 0.0112f
C4693 vdd.n4069 vss 0.0128f
C4694 vdd.n4070 vss 0.0619f
C4695 vdd.n4071 vss 0.00324f
C4696 vdd.n4072 vss 0.0112f
C4697 vdd.n4073 vss 0.0128f
C4698 vdd.n4074 vss 0.00413f
C4699 vdd.n4075 vss 0.00413f
C4700 vdd.n4076 vss 0.0471f
C4701 vdd.n4077 vss 0.0471f
C4702 vdd.n4078 vss 0.00324f
C4703 vdd.n4079 vss 0.00413f
C4704 vdd.n4080 vss 0.00413f
C4705 vdd.n4081 vss 0.00679f
C4706 vdd.n4082 vss 0.00413f
C4707 vdd.n4083 vss 0.0471f
C4708 vdd.n4084 vss 0.00324f
C4709 vdd.n4086 vss 0.00925f
C4710 vdd.n4087 vss 0.0471f
C4711 vdd.n4088 vss 0.00425f
C4712 vdd.n4089 vss 0.0424f
C4713 vdd.n4090 vss 0.0132f
C4714 vdd.n4091 vss 0.00324f
C4715 vdd.n4092 vss 0.0128f
C4716 vdd.n4093 vss 0.02f
C4717 vdd.n4094 vss 0.00425f
C4718 vdd.n4095 vss 0.00413f
C4719 vdd.n4096 vss 0.00251f
C4720 vdd.n4097 vss 0.0471f
C4721 vdd.n4098 vss 0.00251f
C4722 vdd.n4099 vss 0.00517f
C4723 vdd.n4100 vss 0.00679f
C4724 vdd.n4101 vss 0.00324f
C4725 vdd.n4102 vss 0.00324f
C4726 vdd.n4103 vss 0.0132f
C4727 vdd.n4104 vss 0.0424f
C4728 vdd.n4105 vss 0.02f
C4729 vdd.n4106 vss 0.00425f
C4730 vdd.n4107 vss 0.0471f
C4731 vdd.n4109 vss 0.00425f
C4732 vdd.n4110 vss 0.00925f
C4733 vdd.n4111 vss 0.00679f
C4734 vdd.n4112 vss 0.00517f
C4735 vdd.n4113 vss 0.00251f
C4736 vdd.n4114 vss 0.0471f
C4737 vdd.n4115 vss 0.00251f
C4738 vdd.n4116 vss 0.0112f
C4739 vdd.n4117 vss 0.0128f
C4740 vdd.n4118 vss 0.0692f
C4741 vdd.n4119 vss 0.00324f
C4742 vdd.n4120 vss 0.0112f
C4743 vdd.n4121 vss 0.0128f
C4744 vdd.n4122 vss 0.00413f
C4745 vdd.n4123 vss 0.00413f
C4746 vdd.n4124 vss 0.0471f
C4747 vdd.n4125 vss 0.0471f
C4748 vdd.n4126 vss 0.00324f
C4749 vdd.n4127 vss 0.00413f
C4750 vdd.n4128 vss 0.00413f
C4751 vdd.n4129 vss 0.00679f
C4752 vdd.n4130 vss 0.00413f
C4753 vdd.n4131 vss 0.0471f
C4754 vdd.n4132 vss 0.00324f
C4755 vdd.n4134 vss 0.00925f
C4756 vdd.n4135 vss 0.0471f
C4757 vdd.n4136 vss 0.00425f
C4758 vdd.n4137 vss 0.0424f
C4759 vdd.n4138 vss 0.0132f
C4760 vdd.n4139 vss 0.00324f
C4761 vdd.n4140 vss 0.0128f
C4762 vdd.n4141 vss 0.02f
C4763 vdd.n4142 vss 0.00425f
C4764 vdd.n4143 vss 0.00413f
C4765 vdd.n4144 vss 0.00251f
C4766 vdd.n4145 vss 0.0471f
C4767 vdd.n4146 vss 0.00251f
C4768 vdd.n4147 vss 0.00517f
C4769 vdd.n4148 vss 0.00679f
C4770 vdd.n4149 vss 0.00324f
C4771 vdd.n4150 vss 0.00324f
C4772 vdd.n4151 vss 0.0132f
C4773 vdd.n4152 vss 0.0424f
C4774 vdd.n4153 vss 0.02f
C4775 vdd.n4154 vss 0.00425f
C4776 vdd.n4155 vss 0.0471f
C4777 vdd.n4157 vss 0.00425f
C4778 vdd.n4158 vss 0.00925f
C4779 vdd.n4159 vss 0.00679f
C4780 vdd.n4160 vss 0.00517f
C4781 vdd.n4161 vss 0.00251f
C4782 vdd.n4162 vss 0.0471f
C4783 vdd.n4163 vss 0.00251f
C4784 vdd.n4164 vss 0.0112f
C4785 vdd.n4165 vss 0.0128f
C4786 vdd.n4166 vss 0.0619f
C4787 vdd.n4167 vss 0.00335f
C4788 vdd.n4168 vss 0.0855f
C4789 vdd.n4169 vss 0.00991f
C4790 vdd.n4170 vss 0.0424f
C4791 vdd.n4171 vss 0.00679f
C4792 vdd.n4172 vss 0.00413f
C4793 vdd.n4173 vss 0.0471f
C4794 vdd.n4174 vss 0.00251f
C4795 vdd.n4175 vss 0.00679f
C4796 vdd.n4176 vss 0.00413f
C4797 vdd.n4177 vss 0.00413f
C4798 vdd.n4178 vss 0.0471f
C4799 vdd.n4179 vss 0.00251f
C4800 vdd.n4180 vss 0.00413f
C4801 vdd.n4181 vss 0.00324f
C4802 vdd.n4182 vss 0.0132f
C4803 vdd.n4183 vss 0.0424f
C4804 vdd.n4184 vss 0.00324f
C4805 vdd.n4185 vss 0.00413f
C4806 vdd.n4186 vss 0.00517f
C4807 vdd.n4187 vss 0.00679f
C4808 vdd.n4188 vss 0.00925f
C4809 vdd.n4189 vss 0.00425f
C4810 vdd.n4190 vss 0.0471f
C4811 vdd.n4192 vss 0.00425f
C4812 vdd.n4193 vss 0.02f
C4813 vdd.n4194 vss 0.0128f
C4814 vdd.n4195 vss 0.0105f
C4815 vdd.n4196 vss 0.00251f
C4816 vdd.n4197 vss 0.0471f
C4817 vdd.n4198 vss 0.00517f
C4818 vdd.n4199 vss 0.00251f
C4819 vdd.n4200 vss 0.0471f
C4820 vdd.n4201 vss 0.0471f
C4821 vdd.n4202 vss 0.00324f
C4822 vdd.n4203 vss 0.00324f
C4823 vdd.n4204 vss 0.00805f
C4824 vdd.n4205 vss 0.0112f
C4825 vdd.n4206 vss 0.0128f
C4826 vdd.n4207 vss 0.00324f
C4827 vdd.n4208 vss 0.00324f
C4828 vdd.n4209 vss 0.00413f
C4829 vdd.n4210 vss 0.00425f
C4830 vdd.n4211 vss 0.0471f
C4831 vdd.n4213 vss 0.00425f
C4832 vdd.n4214 vss 0.00925f
C4833 vdd.n4215 vss 0.0107f
C4834 vdd.n4216 vss 0.0126f
C4835 vdd.n4217 vss 0.0516f
C4836 vdd.n4218 vss 0.00163f
C4837 vdd.n4219 vss 0.00145f
C4838 vdd.n4220 vss 0.0271f
C4839 vdd.n4221 vss 0.00324f
C4840 vdd.n4222 vss 0.0112f
C4841 vdd.n4223 vss 0.0128f
C4842 vdd.n4224 vss 0.00413f
C4843 vdd.n4225 vss 0.00413f
C4844 vdd.n4226 vss 0.0471f
C4845 vdd.n4227 vss 0.0471f
C4846 vdd.n4228 vss 0.00324f
C4847 vdd.n4229 vss 0.00413f
C4848 vdd.n4230 vss 0.00413f
C4849 vdd.n4231 vss 0.00679f
C4850 vdd.n4232 vss 0.00413f
C4851 vdd.n4233 vss 0.0471f
C4852 vdd.n4234 vss 0.00324f
C4853 vdd.n4236 vss 0.00925f
C4854 vdd.n4237 vss 0.0471f
C4855 vdd.n4238 vss 0.00425f
C4856 vdd.n4239 vss 0.0424f
C4857 vdd.n4240 vss 0.0132f
C4858 vdd.n4241 vss 0.00324f
C4859 vdd.n4242 vss 0.0128f
C4860 vdd.n4243 vss 0.02f
C4861 vdd.n4244 vss 0.00425f
C4862 vdd.n4245 vss 0.00413f
C4863 vdd.n4246 vss 0.00251f
C4864 vdd.n4247 vss 0.0471f
C4865 vdd.n4248 vss 0.00251f
C4866 vdd.n4249 vss 0.00517f
C4867 vdd.n4250 vss 0.00679f
C4868 vdd.n4251 vss 0.00324f
C4869 vdd.n4252 vss 0.00324f
C4870 vdd.n4253 vss 0.0132f
C4871 vdd.n4254 vss 0.0424f
C4872 vdd.n4255 vss 0.02f
C4873 vdd.n4256 vss 0.00425f
C4874 vdd.n4257 vss 0.0471f
C4875 vdd.n4259 vss 0.00425f
C4876 vdd.n4260 vss 0.00925f
C4877 vdd.n4261 vss 0.00679f
C4878 vdd.n4262 vss 0.00517f
C4879 vdd.n4263 vss 0.00251f
C4880 vdd.n4264 vss 0.0471f
C4881 vdd.n4265 vss 0.00251f
C4882 vdd.n4266 vss 0.0112f
C4883 vdd.n4267 vss 0.0128f
C4884 vdd.n4268 vss 0.0692f
C4885 vdd.n4269 vss 0.00324f
C4886 vdd.n4270 vss 0.0112f
C4887 vdd.n4271 vss 0.0128f
C4888 vdd.n4272 vss 0.00413f
C4889 vdd.n4273 vss 0.00413f
C4890 vdd.n4274 vss 0.0471f
C4891 vdd.n4275 vss 0.0471f
C4892 vdd.n4276 vss 0.00324f
C4893 vdd.n4277 vss 0.00413f
C4894 vdd.n4278 vss 0.00413f
C4895 vdd.n4279 vss 0.00679f
C4896 vdd.n4280 vss 0.00413f
C4897 vdd.n4281 vss 0.0471f
C4898 vdd.n4282 vss 0.00324f
C4899 vdd.n4283 vss 0.0424f
C4900 vdd.n4284 vss 0.00324f
C4901 vdd.n4285 vss 0.0128f
C4902 vdd.n4286 vss 0.02f
C4903 vdd.n4287 vss 0.0132f
C4904 vdd.n4288 vss 0.00925f
C4905 vdd.n4289 vss 0.00425f
C4906 vdd.n4291 vss 0.0471f
C4907 vdd.n4292 vss 0.00425f
C4908 vdd.n4293 vss 0.00413f
C4909 vdd.n4294 vss 0.00251f
C4910 vdd.n4295 vss 0.0471f
C4911 vdd.n4296 vss 0.00251f
C4912 vdd.n4297 vss 0.00517f
C4913 vdd.n4298 vss 0.00679f
C4914 vdd.n4299 vss 0.00324f
C4915 vdd.n4300 vss 0.00324f
C4916 vdd.n4301 vss 0.0132f
C4917 vdd.n4302 vss 0.0424f
C4918 vdd.n4303 vss 0.02f
C4919 vdd.n4304 vss 0.00425f
C4920 vdd.n4306 vss 0.0471f
C4921 vdd.n4307 vss 0.00425f
C4922 vdd.n4308 vss 0.00925f
C4923 vdd.n4309 vss 0.00679f
C4924 vdd.n4310 vss 0.00517f
C4925 vdd.n4311 vss 0.00251f
C4926 vdd.n4312 vss 0.0471f
C4927 vdd.n4313 vss 0.00251f
C4928 vdd.n4314 vss 0.0112f
C4929 vdd.n4315 vss 0.0128f
C4930 vdd.n4316 vss 0.0666f
C4931 vdd.n4317 vss 0.00324f
C4932 vdd.n4318 vss 0.0112f
C4933 vdd.n4319 vss 0.0128f
C4934 vdd.n4320 vss 0.00413f
C4935 vdd.n4321 vss 0.00413f
C4936 vdd.n4322 vss 0.0471f
C4937 vdd.n4323 vss 0.0471f
C4938 vdd.n4324 vss 0.00324f
C4939 vdd.n4325 vss 0.00413f
C4940 vdd.n4326 vss 0.00413f
C4941 vdd.n4327 vss 0.00679f
C4942 vdd.n4328 vss 0.00413f
C4943 vdd.n4329 vss 0.0471f
C4944 vdd.n4330 vss 0.00324f
C4945 vdd.n4331 vss 0.0424f
C4946 vdd.n4332 vss 0.00324f
C4947 vdd.n4333 vss 0.0128f
C4948 vdd.n4334 vss 0.02f
C4949 vdd.n4335 vss 0.0132f
C4950 vdd.n4336 vss 0.00925f
C4951 vdd.n4337 vss 0.00425f
C4952 vdd.n4339 vss 0.0471f
C4953 vdd.n4340 vss 0.00425f
C4954 vdd.n4341 vss 0.00413f
C4955 vdd.n4342 vss 0.00251f
C4956 vdd.n4343 vss 0.0471f
C4957 vdd.n4344 vss 0.00251f
C4958 vdd.n4345 vss 0.00517f
C4959 vdd.n4346 vss 0.00679f
C4960 vdd.n4347 vss 0.00324f
C4961 vdd.n4348 vss 0.00324f
C4962 vdd.n4349 vss 0.0132f
C4963 vdd.n4350 vss 0.0424f
C4964 vdd.n4351 vss 0.02f
C4965 vdd.n4352 vss 0.00425f
C4966 vdd.n4354 vss 0.0471f
C4967 vdd.n4355 vss 0.00425f
C4968 vdd.n4356 vss 0.00925f
C4969 vdd.n4357 vss 0.00679f
C4970 vdd.n4358 vss 0.00517f
C4971 vdd.n4359 vss 0.00251f
C4972 vdd.n4360 vss 0.0471f
C4973 vdd.n4361 vss 0.00251f
C4974 vdd.n4362 vss 0.0112f
C4975 vdd.n4363 vss 0.0128f
C4976 vdd.n4364 vss 0.0617f
C4977 vdd.n4365 vss 0.00335f
C4978 vdd.n4366 vss 0.0855f
C4979 vdd.n4367 vss 0.0107f
C4980 vdd.n4368 vss 0.0128f
C4981 vdd.n4369 vss 0.0424f
C4982 vdd.n4370 vss 0.00413f
C4983 vdd.n4371 vss 0.0471f
C4984 vdd.n4372 vss 0.00413f
C4985 vdd.n4373 vss 0.00324f
C4986 vdd.n4374 vss 0.00324f
C4987 vdd.n4375 vss 0.00679f
C4988 vdd.n4376 vss 0.00413f
C4989 vdd.n4377 vss 0.0471f
C4990 vdd.n4378 vss 0.00413f
C4991 vdd.n4379 vss 0.0105f
C4992 vdd.n4380 vss 0.0471f
C4993 vdd.n4381 vss 0.00413f
C4994 vdd.n4382 vss 0.00324f
C4995 vdd.n4383 vss 0.00324f
C4996 vdd.n4384 vss 0.0132f
C4997 vdd.n4385 vss 0.0424f
C4998 vdd.n4386 vss 0.0128f
C4999 vdd.n4387 vss 0.02f
C5000 vdd.n4388 vss 0.00425f
C5001 vdd.n4390 vss 0.0471f
C5002 vdd.n4391 vss 0.00425f
C5003 vdd.n4392 vss 0.00925f
C5004 vdd.n4393 vss 0.00679f
C5005 vdd.n4394 vss 0.00517f
C5006 vdd.n4395 vss 0.00251f
C5007 vdd.n4396 vss 0.0471f
C5008 vdd.n4397 vss 0.00251f
C5009 vdd.n4398 vss 0.00413f
C5010 vdd.n4399 vss 0.00324f
C5011 vdd.n4400 vss 0.00324f
C5012 vdd.n4401 vss 0.00805f
C5013 vdd.n4402 vss 0.0112f
C5014 vdd.n4403 vss 0.00251f
C5015 vdd.n4404 vss 0.0471f
C5016 vdd.n4405 vss 0.00251f
C5017 vdd.n4406 vss 0.00517f
C5018 vdd.n4407 vss 0.00679f
C5019 vdd.n4408 vss 0.00925f
C5020 vdd.n4409 vss 0.00425f
C5021 vdd.n4411 vss 0.0471f
C5022 vdd.n4412 vss 0.00425f
C5023 vdd.n4413 vss 0.00991f
C5024 vdd.n4414 vss 0.0126f
C5025 vdd.n4415 vss 0.0516f
C5026 vdd.n4416 vss 0.0011f
C5027 vdd.n4417 vss 0.0271f
C5028 vdd.n4418 vss 0.00324f
C5029 vdd.n4419 vss 0.0112f
C5030 vdd.n4420 vss 0.0128f
C5031 vdd.n4421 vss 0.00413f
C5032 vdd.n4422 vss 0.00413f
C5033 vdd.n4423 vss 0.0471f
C5034 vdd.n4424 vss 0.0471f
C5035 vdd.n4425 vss 0.00324f
C5036 vdd.n4426 vss 0.00413f
C5037 vdd.n4427 vss 0.00413f
C5038 vdd.n4428 vss 0.00679f
C5039 vdd.n4429 vss 0.00413f
C5040 vdd.n4430 vss 0.0471f
C5041 vdd.n4431 vss 0.00324f
C5042 vdd.n4432 vss 0.0424f
C5043 vdd.n4433 vss 0.00324f
C5044 vdd.n4434 vss 0.0128f
C5045 vdd.n4435 vss 0.02f
C5046 vdd.n4436 vss 0.0132f
C5047 vdd.n4437 vss 0.00925f
C5048 vdd.n4438 vss 0.00425f
C5049 vdd.n4440 vss 0.0471f
C5050 vdd.n4441 vss 0.00425f
C5051 vdd.n4442 vss 0.00413f
C5052 vdd.n4443 vss 0.00251f
C5053 vdd.n4444 vss 0.0471f
C5054 vdd.n4445 vss 0.00251f
C5055 vdd.n4446 vss 0.00517f
C5056 vdd.n4447 vss 0.00679f
C5057 vdd.n4448 vss 0.00324f
C5058 vdd.n4449 vss 0.00324f
C5059 vdd.n4450 vss 0.0132f
C5060 vdd.n4451 vss 0.0424f
C5061 vdd.n4452 vss 0.02f
C5062 vdd.n4453 vss 0.00425f
C5063 vdd.n4455 vss 0.0471f
C5064 vdd.n4456 vss 0.00425f
C5065 vdd.n4457 vss 0.00925f
C5066 vdd.n4458 vss 0.00679f
C5067 vdd.n4459 vss 0.00517f
C5068 vdd.n4460 vss 0.00251f
C5069 vdd.n4461 vss 0.0471f
C5070 vdd.n4462 vss 0.00251f
C5071 vdd.n4463 vss 0.0112f
C5072 vdd.n4464 vss 0.0128f
C5073 vdd.n4465 vss 0.0666f
C5074 vdd.n4466 vss 0.00324f
C5075 vdd.n4467 vss 0.0112f
C5076 vdd.n4468 vss 0.0128f
C5077 vdd.n4469 vss 0.00413f
C5078 vdd.n4470 vss 0.00413f
C5079 vdd.n4471 vss 0.0471f
C5080 vdd.n4472 vss 0.0471f
C5081 vdd.n4473 vss 0.00324f
C5082 vdd.n4474 vss 0.00413f
C5083 vdd.n4475 vss 0.00413f
C5084 vdd.n4476 vss 0.00679f
C5085 vdd.n4477 vss 0.00413f
C5086 vdd.n4478 vss 0.0471f
C5087 vdd.n4479 vss 0.00324f
C5088 vdd.n4480 vss 0.0424f
C5089 vdd.n4481 vss 0.00324f
C5090 vdd.n4482 vss 0.0128f
C5091 vdd.n4483 vss 0.02f
C5092 vdd.n4484 vss 0.0132f
C5093 vdd.n4485 vss 0.00925f
C5094 vdd.n4486 vss 0.00425f
C5095 vdd.n4488 vss 0.0471f
C5096 vdd.n4489 vss 0.00425f
C5097 vdd.n4490 vss 0.00413f
C5098 vdd.n4491 vss 0.00251f
C5099 vdd.n4492 vss 0.0471f
C5100 vdd.n4493 vss 0.00251f
C5101 vdd.n4494 vss 0.00517f
C5102 vdd.n4495 vss 0.00679f
C5103 vdd.n4496 vss 0.00324f
C5104 vdd.n4497 vss 0.00324f
C5105 vdd.n4498 vss 0.0132f
C5106 vdd.n4499 vss 0.0424f
C5107 vdd.n4500 vss 0.02f
C5108 vdd.n4501 vss 0.00425f
C5109 vdd.n4503 vss 0.0471f
C5110 vdd.n4504 vss 0.00425f
C5111 vdd.n4505 vss 0.00925f
C5112 vdd.n4506 vss 0.00679f
C5113 vdd.n4507 vss 0.00517f
C5114 vdd.n4508 vss 0.00251f
C5115 vdd.n4509 vss 0.0471f
C5116 vdd.n4510 vss 0.00251f
C5117 vdd.n4511 vss 0.0112f
C5118 vdd.n4512 vss 0.0128f
C5119 vdd.n4513 vss 0.0613f
C5120 vdd.n4514 vss 0.00324f
C5121 vdd.n4515 vss 0.0112f
C5122 vdd.n4516 vss 0.0128f
C5123 vdd.n4517 vss 0.00413f
C5124 vdd.n4518 vss 0.00413f
C5125 vdd.n4519 vss 0.0471f
C5126 vdd.n4520 vss 0.0471f
C5127 vdd.n4521 vss 0.00324f
C5128 vdd.n4522 vss 0.00413f
C5129 vdd.n4523 vss 0.00413f
C5130 vdd.n4524 vss 0.00679f
C5131 vdd.n4525 vss 0.00413f
C5132 vdd.n4526 vss 0.0471f
C5133 vdd.n4527 vss 0.00324f
C5134 vdd.n4528 vss 0.0424f
C5135 vdd.n4529 vss 0.00324f
C5136 vdd.n4530 vss 0.0128f
C5137 vdd.n4531 vss 0.02f
C5138 vdd.n4532 vss 0.0132f
C5139 vdd.n4533 vss 0.00925f
C5140 vdd.n4534 vss 0.00425f
C5141 vdd.n4536 vss 0.0471f
C5142 vdd.n4537 vss 0.00425f
C5143 vdd.n4538 vss 0.00413f
C5144 vdd.n4539 vss 0.00251f
C5145 vdd.n4540 vss 0.0471f
C5146 vdd.n4541 vss 0.00251f
C5147 vdd.n4542 vss 0.00517f
C5148 vdd.n4543 vss 0.00679f
C5149 vdd.n4544 vss 0.00324f
C5150 vdd.n4545 vss 0.00324f
C5151 vdd.n4546 vss 0.0132f
C5152 vdd.n4547 vss 0.0424f
C5153 vdd.n4548 vss 0.02f
C5154 vdd.n4549 vss 0.00425f
C5155 vdd.n4551 vss 0.0471f
C5156 vdd.n4552 vss 0.00425f
C5157 vdd.n4553 vss 0.00925f
C5158 vdd.n4554 vss 0.00679f
C5159 vdd.n4555 vss 0.00517f
C5160 vdd.n4556 vss 0.00251f
C5161 vdd.n4557 vss 0.0471f
C5162 vdd.n4558 vss 0.00251f
C5163 vdd.n4559 vss 0.0112f
C5164 vdd.n4560 vss 0.0128f
C5165 vdd.n4561 vss 0.0666f
C5166 vdd.n4562 vss 0.00324f
C5167 vdd.n4563 vss 0.0112f
C5168 vdd.n4564 vss 0.0128f
C5169 vdd.n4565 vss 0.00413f
C5170 vdd.n4566 vss 0.00413f
C5171 vdd.n4567 vss 0.0471f
C5172 vdd.n4568 vss 0.0471f
C5173 vdd.n4569 vss 0.00324f
C5174 vdd.n4570 vss 0.00413f
C5175 vdd.n4571 vss 0.00413f
C5176 vdd.n4572 vss 0.00679f
C5177 vdd.n4573 vss 0.00413f
C5178 vdd.n4574 vss 0.0471f
C5179 vdd.n4575 vss 0.00324f
C5180 vdd.n4576 vss 0.0424f
C5181 vdd.n4577 vss 0.00324f
C5182 vdd.n4578 vss 0.0128f
C5183 vdd.n4579 vss 0.02f
C5184 vdd.n4580 vss 0.0132f
C5185 vdd.n4581 vss 0.00925f
C5186 vdd.n4582 vss 0.00425f
C5187 vdd.n4584 vss 0.0471f
C5188 vdd.n4585 vss 0.00425f
C5189 vdd.n4586 vss 0.00413f
C5190 vdd.n4587 vss 0.00251f
C5191 vdd.n4588 vss 0.0471f
C5192 vdd.n4589 vss 0.00251f
C5193 vdd.n4590 vss 0.00517f
C5194 vdd.n4591 vss 0.00679f
C5195 vdd.n4592 vss 0.00324f
C5196 vdd.n4593 vss 0.00324f
C5197 vdd.n4594 vss 0.0132f
C5198 vdd.n4595 vss 0.0424f
C5199 vdd.n4596 vss 0.02f
C5200 vdd.n4597 vss 0.00425f
C5201 vdd.n4599 vss 0.0471f
C5202 vdd.n4600 vss 0.00425f
C5203 vdd.n4601 vss 0.00925f
C5204 vdd.n4602 vss 0.00679f
C5205 vdd.n4603 vss 0.00517f
C5206 vdd.n4604 vss 0.00251f
C5207 vdd.n4605 vss 0.0471f
C5208 vdd.n4606 vss 0.00251f
C5209 vdd.n4607 vss 0.0112f
C5210 vdd.n4608 vss 0.0128f
C5211 vdd.n4609 vss 0.0617f
C5212 vdd.n4610 vss 0.00335f
C5213 vdd.n4611 vss 0.0855f
C5214 vdd.n4612 vss 0.0107f
C5215 vdd.n4613 vss 0.0128f
C5216 vdd.n4614 vss 0.0424f
C5217 vdd.n4615 vss 0.00413f
C5218 vdd.n4616 vss 0.0471f
C5219 vdd.n4617 vss 0.00413f
C5220 vdd.n4618 vss 0.00324f
C5221 vdd.n4619 vss 0.00324f
C5222 vdd.n4620 vss 0.00679f
C5223 vdd.n4621 vss 0.00413f
C5224 vdd.n4622 vss 0.0471f
C5225 vdd.n4623 vss 0.00413f
C5226 vdd.n4624 vss 0.0105f
C5227 vdd.n4625 vss 0.0471f
C5228 vdd.n4626 vss 0.00413f
C5229 vdd.n4627 vss 0.00324f
C5230 vdd.n4628 vss 0.00324f
C5231 vdd.n4629 vss 0.0132f
C5232 vdd.n4630 vss 0.0424f
C5233 vdd.n4631 vss 0.0128f
C5234 vdd.n4632 vss 0.02f
C5235 vdd.n4633 vss 0.00425f
C5236 vdd.n4635 vss 0.0471f
C5237 vdd.n4636 vss 0.00425f
C5238 vdd.n4637 vss 0.00925f
C5239 vdd.n4638 vss 0.00679f
C5240 vdd.n4639 vss 0.00517f
C5241 vdd.n4640 vss 0.00251f
C5242 vdd.n4641 vss 0.0471f
C5243 vdd.n4642 vss 0.00251f
C5244 vdd.n4643 vss 0.00413f
C5245 vdd.n4644 vss 0.00324f
C5246 vdd.n4645 vss 0.00324f
C5247 vdd.n4646 vss 0.00805f
C5248 vdd.n4647 vss 0.0112f
C5249 vdd.n4648 vss 0.00251f
C5250 vdd.n4649 vss 0.0471f
C5251 vdd.n4650 vss 0.00251f
C5252 vdd.n4651 vss 0.00517f
C5253 vdd.n4652 vss 0.00679f
C5254 vdd.n4653 vss 0.00925f
C5255 vdd.n4654 vss 0.00425f
C5256 vdd.n4656 vss 0.0471f
C5257 vdd.n4657 vss 0.00425f
C5258 vdd.n4658 vss 0.00991f
C5259 vdd.n4659 vss 0.0126f
C5260 vdd.n4660 vss 0.0516f
C5261 vdd.n4661 vss 0.0011f
C5262 vdd.n4662 vss 0.0271f
C5263 vdd.n4663 vss 0.00324f
C5264 vdd.n4664 vss 0.0112f
C5265 vdd.n4665 vss 0.0128f
C5266 vdd.n4666 vss 0.00413f
C5267 vdd.n4667 vss 0.00413f
C5268 vdd.n4668 vss 0.0471f
C5269 vdd.n4669 vss 0.0471f
C5270 vdd.n4670 vss 0.00324f
C5271 vdd.n4671 vss 0.00413f
C5272 vdd.n4672 vss 0.00413f
C5273 vdd.n4673 vss 0.00679f
C5274 vdd.n4674 vss 0.00413f
C5275 vdd.n4675 vss 0.0471f
C5276 vdd.n4676 vss 0.00324f
C5277 vdd.n4677 vss 0.0424f
C5278 vdd.n4678 vss 0.00324f
C5279 vdd.n4679 vss 0.0128f
C5280 vdd.n4680 vss 0.02f
C5281 vdd.n4681 vss 0.0132f
C5282 vdd.n4682 vss 0.00925f
C5283 vdd.n4683 vss 0.00425f
C5284 vdd.n4685 vss 0.0471f
C5285 vdd.n4686 vss 0.00425f
C5286 vdd.n4687 vss 0.00413f
C5287 vdd.n4688 vss 0.00251f
C5288 vdd.n4689 vss 0.0471f
C5289 vdd.n4690 vss 0.00251f
C5290 vdd.n4691 vss 0.00517f
C5291 vdd.n4692 vss 0.00679f
C5292 vdd.n4693 vss 0.00324f
C5293 vdd.n4694 vss 0.00324f
C5294 vdd.n4695 vss 0.0132f
C5295 vdd.n4696 vss 0.0424f
C5296 vdd.n4697 vss 0.02f
C5297 vdd.n4698 vss 0.00425f
C5298 vdd.n4700 vss 0.0471f
C5299 vdd.n4701 vss 0.00425f
C5300 vdd.n4702 vss 0.00925f
C5301 vdd.n4703 vss 0.00679f
C5302 vdd.n4704 vss 0.00517f
C5303 vdd.n4705 vss 0.00251f
C5304 vdd.n4706 vss 0.0471f
C5305 vdd.n4707 vss 0.00251f
C5306 vdd.n4708 vss 0.0112f
C5307 vdd.n4709 vss 0.0128f
C5308 vdd.n4710 vss 0.0666f
C5309 vdd.n4711 vss 0.00324f
C5310 vdd.n4712 vss 0.0112f
C5311 vdd.n4713 vss 0.0128f
C5312 vdd.n4714 vss 0.00413f
C5313 vdd.n4715 vss 0.00413f
C5314 vdd.n4716 vss 0.0471f
C5315 vdd.n4717 vss 0.0471f
C5316 vdd.n4718 vss 0.00324f
C5317 vdd.n4719 vss 0.00413f
C5318 vdd.n4720 vss 0.00413f
C5319 vdd.n4721 vss 0.00679f
C5320 vdd.n4722 vss 0.00413f
C5321 vdd.n4723 vss 0.0471f
C5322 vdd.n4724 vss 0.00324f
C5323 vdd.n4725 vss 0.0424f
C5324 vdd.n4726 vss 0.00324f
C5325 vdd.n4727 vss 0.0128f
C5326 vdd.n4728 vss 0.02f
C5327 vdd.n4729 vss 0.0132f
C5328 vdd.n4730 vss 0.00925f
C5329 vdd.n4731 vss 0.00425f
C5330 vdd.n4733 vss 0.0471f
C5331 vdd.n4734 vss 0.00425f
C5332 vdd.n4735 vss 0.00413f
C5333 vdd.n4736 vss 0.00251f
C5334 vdd.n4737 vss 0.0471f
C5335 vdd.n4738 vss 0.00251f
C5336 vdd.n4739 vss 0.00517f
C5337 vdd.n4740 vss 0.00679f
C5338 vdd.n4741 vss 0.00324f
C5339 vdd.n4742 vss 0.00324f
C5340 vdd.n4743 vss 0.0132f
C5341 vdd.n4744 vss 0.0424f
C5342 vdd.n4745 vss 0.02f
C5343 vdd.n4746 vss 0.00425f
C5344 vdd.n4748 vss 0.0471f
C5345 vdd.n4749 vss 0.00425f
C5346 vdd.n4750 vss 0.00925f
C5347 vdd.n4751 vss 0.00679f
C5348 vdd.n4752 vss 0.00517f
C5349 vdd.n4753 vss 0.00251f
C5350 vdd.n4754 vss 0.0471f
C5351 vdd.n4755 vss 0.00251f
C5352 vdd.n4756 vss 0.0112f
C5353 vdd.n4757 vss 0.0128f
C5354 vdd.n4758 vss 0.00324f
C5355 vdd.n4759 vss 0.0112f
C5356 vdd.n4760 vss 0.0128f
C5357 vdd.n4761 vss 0.00413f
C5358 vdd.n4762 vss 0.00413f
C5359 vdd.n4763 vss 0.0471f
C5360 vdd.n4764 vss 0.0471f
C5361 vdd.n4765 vss 0.00324f
C5362 vdd.n4766 vss 0.00413f
C5363 vdd.n4767 vss 0.00413f
C5364 vdd.n4768 vss 0.00679f
C5365 vdd.n4769 vss 0.00413f
C5366 vdd.n4770 vss 0.0471f
C5367 vdd.n4771 vss 0.00324f
C5368 vdd.n4772 vss 0.0424f
C5369 vdd.n4773 vss 0.00324f
C5370 vdd.n4774 vss 0.0128f
C5371 vdd.n4775 vss 0.02f
C5372 vdd.n4776 vss 0.0132f
C5373 vdd.n4777 vss 0.00925f
C5374 vdd.n4778 vss 0.00425f
C5375 vdd.n4780 vss 0.0471f
C5376 vdd.n4781 vss 0.00425f
C5377 vdd.n4782 vss 0.00413f
C5378 vdd.n4783 vss 0.00251f
C5379 vdd.n4784 vss 0.0471f
C5380 vdd.n4785 vss 0.00251f
C5381 vdd.n4786 vss 0.00517f
C5382 vdd.n4787 vss 0.00679f
C5383 vdd.n4788 vss 0.00324f
C5384 vdd.n4789 vss 0.00324f
C5385 vdd.n4790 vss 0.0132f
C5386 vdd.n4791 vss 0.0424f
C5387 vdd.n4792 vss 0.02f
C5388 vdd.n4793 vss 0.00425f
C5389 vdd.n4795 vss 0.0471f
C5390 vdd.n4796 vss 0.00425f
C5391 vdd.n4797 vss 0.00925f
C5392 vdd.n4798 vss 0.00679f
C5393 vdd.n4799 vss 0.00517f
C5394 vdd.n4800 vss 0.00251f
C5395 vdd.n4801 vss 0.0471f
C5396 vdd.n4802 vss 0.00251f
C5397 vdd.n4803 vss 0.0112f
C5398 vdd.n4804 vss 0.0128f
C5399 vdd.n4805 vss 0.144f
C5400 vdd.n4806 vss 0.143f
C5401 vdd.n4807 vss 0.0608f
C5402 vdd.n4808 vss 0.00324f
C5403 vdd.n4809 vss 0.0112f
C5404 vdd.n4810 vss 0.0128f
C5405 vdd.n4811 vss 0.00413f
C5406 vdd.n4812 vss 0.00413f
C5407 vdd.n4813 vss 0.0471f
C5408 vdd.n4814 vss 0.0471f
C5409 vdd.n4815 vss 0.00324f
C5410 vdd.n4816 vss 0.00413f
C5411 vdd.n4817 vss 0.00413f
C5412 vdd.n4818 vss 0.00679f
C5413 vdd.n4819 vss 0.00413f
C5414 vdd.n4820 vss 0.0471f
C5415 vdd.n4821 vss 0.00324f
C5416 vdd.n4822 vss 0.0424f
C5417 vdd.n4823 vss 0.00324f
C5418 vdd.n4824 vss 0.0128f
C5419 vdd.n4825 vss 0.02f
C5420 vdd.n4826 vss 0.0132f
C5421 vdd.n4827 vss 0.00925f
C5422 vdd.n4828 vss 0.00425f
C5423 vdd.n4830 vss 0.0471f
C5424 vdd.n4831 vss 0.00425f
C5425 vdd.n4832 vss 0.00413f
C5426 vdd.n4833 vss 0.00251f
C5427 vdd.n4834 vss 0.0471f
C5428 vdd.n4835 vss 0.00251f
C5429 vdd.n4836 vss 0.00517f
C5430 vdd.n4837 vss 0.00679f
C5431 vdd.n4838 vss 0.00324f
C5432 vdd.n4839 vss 0.00324f
C5433 vdd.n4840 vss 0.0132f
C5434 vdd.n4841 vss 0.0424f
C5435 vdd.n4842 vss 0.02f
C5436 vdd.n4843 vss 0.00425f
C5437 vdd.n4845 vss 0.0471f
C5438 vdd.n4846 vss 0.00425f
C5439 vdd.n4847 vss 0.00925f
C5440 vdd.n4848 vss 0.00679f
C5441 vdd.n4849 vss 0.00517f
C5442 vdd.n4850 vss 0.00251f
C5443 vdd.n4851 vss 0.0471f
C5444 vdd.n4852 vss 0.00251f
C5445 vdd.n4853 vss 0.0112f
C5446 vdd.n4854 vss 0.0128f
C5447 vdd.n4855 vss 0.0666f
C5448 vdd.n4856 vss 0.118f
C5449 vdd.n4857 vss 0.121f
C5450 vdd.n4858 vss 0.00324f
C5451 vdd.n4859 vss 0.0112f
C5452 vdd.n4860 vss 0.0128f
C5453 vdd.n4861 vss 0.00413f
C5454 vdd.n4862 vss 0.00413f
C5455 vdd.n4863 vss 0.0471f
C5456 vdd.n4864 vss 0.0471f
C5457 vdd.n4865 vss 0.00324f
C5458 vdd.n4866 vss 0.00413f
C5459 vdd.n4867 vss 0.00413f
C5460 vdd.n4868 vss 0.00679f
C5461 vdd.n4869 vss 0.00413f
C5462 vdd.n4870 vss 0.0471f
C5463 vdd.n4871 vss 0.00324f
C5464 vdd.n4872 vss 0.0424f
C5465 vdd.n4873 vss 0.00324f
C5466 vdd.n4874 vss 0.0128f
C5467 vdd.n4875 vss 0.02f
C5468 vdd.n4876 vss 0.0132f
C5469 vdd.n4877 vss 0.00925f
C5470 vdd.n4878 vss 0.00425f
C5471 vdd.n4880 vss 0.0471f
C5472 vdd.n4881 vss 0.00425f
C5473 vdd.n4882 vss 0.00413f
C5474 vdd.n4883 vss 0.00251f
C5475 vdd.n4884 vss 0.0471f
C5476 vdd.n4885 vss 0.00251f
C5477 vdd.n4886 vss 0.00517f
C5478 vdd.n4887 vss 0.00679f
C5479 vdd.n4888 vss 0.00324f
C5480 vdd.n4889 vss 0.00324f
C5481 vdd.n4890 vss 0.0132f
C5482 vdd.n4891 vss 0.0424f
C5483 vdd.n4892 vss 0.02f
C5484 vdd.n4893 vss 0.00425f
C5485 vdd.n4895 vss 0.0471f
C5486 vdd.n4896 vss 0.00425f
C5487 vdd.n4897 vss 0.00925f
C5488 vdd.n4898 vss 0.00679f
C5489 vdd.n4899 vss 0.00517f
C5490 vdd.n4900 vss 0.00251f
C5491 vdd.n4901 vss 0.0471f
C5492 vdd.n4902 vss 0.00251f
C5493 vdd.n4903 vss 0.0112f
C5494 vdd.n4904 vss 0.0955f
C5495 vdd.n4905 vss 0.0608f
C5496 vdd.n4906 vss 0.00324f
C5497 vdd.n4907 vss 0.0112f
C5498 vdd.n4908 vss 0.0128f
C5499 vdd.n4909 vss 0.00413f
C5500 vdd.n4910 vss 0.00413f
C5501 vdd.n4911 vss 0.0471f
C5502 vdd.n4912 vss 0.0471f
C5503 vdd.n4913 vss 0.00324f
C5504 vdd.n4914 vss 0.00413f
C5505 vdd.n4915 vss 0.00413f
C5506 vdd.n4916 vss 0.00679f
C5507 vdd.n4917 vss 0.00413f
C5508 vdd.n4918 vss 0.0471f
C5509 vdd.n4919 vss 0.00324f
C5510 vdd.n4920 vss 0.0424f
C5511 vdd.n4921 vss 0.00324f
C5512 vdd.n4922 vss 0.0128f
C5513 vdd.n4923 vss 0.02f
C5514 vdd.n4924 vss 0.0132f
C5515 vdd.n4925 vss 0.00925f
C5516 vdd.n4926 vss 0.00425f
C5517 vdd.n4928 vss 0.0471f
C5518 vdd.n4929 vss 0.00425f
C5519 vdd.n4930 vss 0.00413f
C5520 vdd.n4931 vss 0.00251f
C5521 vdd.n4932 vss 0.0471f
C5522 vdd.n4933 vss 0.00251f
C5523 vdd.n4934 vss 0.00517f
C5524 vdd.n4935 vss 0.00679f
C5525 vdd.n4936 vss 0.00324f
C5526 vdd.n4937 vss 0.00324f
C5527 vdd.n4938 vss 0.0132f
C5528 vdd.n4939 vss 0.0424f
C5529 vdd.n4940 vss 0.02f
C5530 vdd.n4941 vss 0.00425f
C5531 vdd.n4943 vss 0.0471f
C5532 vdd.n4944 vss 0.00425f
C5533 vdd.n4945 vss 0.00925f
C5534 vdd.n4946 vss 0.00679f
C5535 vdd.n4947 vss 0.00517f
C5536 vdd.n4948 vss 0.00251f
C5537 vdd.n4949 vss 0.0471f
C5538 vdd.n4950 vss 0.00251f
C5539 vdd.n4951 vss 0.0112f
C5540 vdd.n4952 vss 0.0128f
C5541 vdd.n4953 vss 0.0666f
C5542 vdd.n4954 vss 0.0912f
C5543 vdd.n4955 vss 0.0824f
C5544 vdd.n4956 vss 0.0567f
C5545 vdd.n4957 vss 0.00324f
C5546 vdd.n4958 vss 0.0112f
C5547 vdd.n4959 vss 0.0128f
C5548 vdd.n4960 vss 0.00413f
C5549 vdd.n4961 vss 0.00413f
C5550 vdd.n4962 vss 0.0471f
C5551 vdd.n4963 vss 0.0471f
C5552 vdd.n4964 vss 0.00324f
C5553 vdd.n4965 vss 0.00413f
C5554 vdd.n4966 vss 0.00413f
C5555 vdd.n4967 vss 0.00679f
C5556 vdd.n4968 vss 0.00413f
C5557 vdd.n4969 vss 0.0471f
C5558 vdd.n4970 vss 0.00324f
C5559 vdd.n4971 vss 0.0424f
C5560 vdd.n4972 vss 0.00324f
C5561 vdd.n4973 vss 0.0128f
C5562 vdd.n4974 vss 0.02f
C5563 vdd.n4975 vss 0.0132f
C5564 vdd.n4976 vss 0.00925f
C5565 vdd.n4977 vss 0.00425f
C5566 vdd.n4979 vss 0.0471f
C5567 vdd.n4980 vss 0.00425f
C5568 vdd.n4981 vss 0.00413f
C5569 vdd.n4982 vss 0.00251f
C5570 vdd.n4983 vss 0.0471f
C5571 vdd.n4984 vss 0.00251f
C5572 vdd.n4985 vss 0.00517f
C5573 vdd.n4986 vss 0.00679f
C5574 vdd.n4987 vss 0.00324f
C5575 vdd.n4988 vss 0.00324f
C5576 vdd.n4989 vss 0.0132f
C5577 vdd.n4990 vss 0.0424f
C5578 vdd.n4991 vss 0.02f
C5579 vdd.n4992 vss 0.00425f
C5580 vdd.n4994 vss 0.0471f
C5581 vdd.n4995 vss 0.00425f
C5582 vdd.n4996 vss 0.00925f
C5583 vdd.n4997 vss 0.00679f
C5584 vdd.n4998 vss 0.00517f
C5585 vdd.n4999 vss 0.00251f
C5586 vdd.n5000 vss 0.0471f
C5587 vdd.n5001 vss 0.00251f
C5588 vdd.n5002 vss 0.0112f
C5589 vdd.n5003 vss 0.0128f
C5590 vdd.n5004 vss 0.00324f
C5591 vdd.n5005 vss 0.0112f
C5592 vdd.n5006 vss 0.0128f
C5593 vdd.n5007 vss 0.00413f
C5594 vdd.n5008 vss 0.00413f
C5595 vdd.n5009 vss 0.0471f
C5596 vdd.n5010 vss 0.0471f
C5597 vdd.n5011 vss 0.00324f
C5598 vdd.n5012 vss 0.00413f
C5599 vdd.n5013 vss 0.00413f
C5600 vdd.n5014 vss 0.00679f
C5601 vdd.n5015 vss 0.00413f
C5602 vdd.n5016 vss 0.0471f
C5603 vdd.n5017 vss 0.00324f
C5604 vdd.n5018 vss 0.0424f
C5605 vdd.n5019 vss 0.00324f
C5606 vdd.n5020 vss 0.0128f
C5607 vdd.n5021 vss 0.02f
C5608 vdd.n5022 vss 0.0132f
C5609 vdd.n5023 vss 0.00925f
C5610 vdd.n5024 vss 0.00425f
C5611 vdd.n5026 vss 0.0471f
C5612 vdd.n5027 vss 0.00425f
C5613 vdd.n5028 vss 0.00413f
C5614 vdd.n5029 vss 0.00251f
C5615 vdd.n5030 vss 0.0471f
C5616 vdd.n5031 vss 0.00251f
C5617 vdd.n5032 vss 0.00517f
C5618 vdd.n5033 vss 0.00679f
C5619 vdd.n5034 vss 0.00324f
C5620 vdd.n5035 vss 0.00324f
C5621 vdd.n5036 vss 0.0132f
C5622 vdd.n5037 vss 0.0424f
C5623 vdd.n5038 vss 0.02f
C5624 vdd.n5039 vss 0.00425f
C5625 vdd.n5041 vss 0.0471f
C5626 vdd.n5042 vss 0.00425f
C5627 vdd.n5043 vss 0.00925f
C5628 vdd.n5044 vss 0.00679f
C5629 vdd.n5045 vss 0.00517f
C5630 vdd.n5046 vss 0.00251f
C5631 vdd.n5047 vss 0.0471f
C5632 vdd.n5048 vss 0.00251f
C5633 vdd.n5049 vss 0.0112f
C5634 vdd.n5050 vss 0.0128f
C5635 vdd.n5051 vss 0.0564f
C5636 vdd.n5052 vss 0.00324f
C5637 vdd.n5053 vss 0.0112f
C5638 vdd.n5054 vss 0.0128f
C5639 vdd.n5055 vss 0.00413f
C5640 vdd.n5056 vss 0.00413f
C5641 vdd.n5057 vss 0.0471f
C5642 vdd.n5058 vss 0.0471f
C5643 vdd.n5059 vss 0.00324f
C5644 vdd.n5060 vss 0.00413f
C5645 vdd.n5061 vss 0.00413f
C5646 vdd.n5062 vss 0.00679f
C5647 vdd.n5063 vss 0.00413f
C5648 vdd.n5064 vss 0.0471f
C5649 vdd.n5065 vss 0.00324f
C5650 vdd.n5066 vss 0.0424f
C5651 vdd.n5067 vss 0.00324f
C5652 vdd.n5068 vss 0.0128f
C5653 vdd.n5069 vss 0.02f
C5654 vdd.n5070 vss 0.0132f
C5655 vdd.n5071 vss 0.00925f
C5656 vdd.n5072 vss 0.00425f
C5657 vdd.n5074 vss 0.0471f
C5658 vdd.n5075 vss 0.00425f
C5659 vdd.n5076 vss 0.00413f
C5660 vdd.n5077 vss 0.00251f
C5661 vdd.n5078 vss 0.0471f
C5662 vdd.n5079 vss 0.00251f
C5663 vdd.n5080 vss 0.00517f
C5664 vdd.n5081 vss 0.00679f
C5665 vdd.n5082 vss 0.00324f
C5666 vdd.n5083 vss 0.00324f
C5667 vdd.n5084 vss 0.0132f
C5668 vdd.n5085 vss 0.0424f
C5669 vdd.n5086 vss 0.02f
C5670 vdd.n5087 vss 0.00425f
C5671 vdd.n5089 vss 0.0471f
C5672 vdd.n5090 vss 0.00425f
C5673 vdd.n5091 vss 0.00925f
C5674 vdd.n5092 vss 0.00679f
C5675 vdd.n5093 vss 0.00517f
C5676 vdd.n5094 vss 0.00251f
C5677 vdd.n5095 vss 0.0471f
C5678 vdd.n5096 vss 0.00251f
C5679 vdd.n5097 vss 0.0112f
C5680 vdd.n5098 vss 0.0128f
C5681 vdd.n5099 vss 0.183f
C5682 vdd.n5100 vss 0.256f
C5683 vdd.n5101 vss 0.12f
C5684 vdd.n5102 vss 0.0608f
C5685 vdd.n5103 vss 0.00324f
C5686 vdd.n5104 vss 0.0112f
C5687 vdd.n5105 vss 0.0128f
C5688 vdd.n5106 vss 0.00413f
C5689 vdd.n5107 vss 0.00413f
C5690 vdd.n5108 vss 0.0471f
C5691 vdd.n5109 vss 0.0471f
C5692 vdd.n5110 vss 0.00324f
C5693 vdd.n5111 vss 0.00413f
C5694 vdd.n5112 vss 0.00413f
C5695 vdd.n5113 vss 0.00679f
C5696 vdd.n5114 vss 0.00413f
C5697 vdd.n5115 vss 0.0471f
C5698 vdd.n5116 vss 0.00324f
C5699 vdd.n5117 vss 0.0424f
C5700 vdd.n5118 vss 0.00324f
C5701 vdd.n5119 vss 0.0128f
C5702 vdd.n5120 vss 0.02f
C5703 vdd.n5121 vss 0.0132f
C5704 vdd.n5122 vss 0.00925f
C5705 vdd.n5123 vss 0.00425f
C5706 vdd.n5125 vss 0.0471f
C5707 vdd.n5126 vss 0.00425f
C5708 vdd.n5127 vss 0.00413f
C5709 vdd.n5128 vss 0.00251f
C5710 vdd.n5129 vss 0.0471f
C5711 vdd.n5130 vss 0.00251f
C5712 vdd.n5131 vss 0.00517f
C5713 vdd.n5132 vss 0.00679f
C5714 vdd.n5133 vss 0.00324f
C5715 vdd.n5134 vss 0.00324f
C5716 vdd.n5135 vss 0.0132f
C5717 vdd.n5136 vss 0.0424f
C5718 vdd.n5137 vss 0.02f
C5719 vdd.n5138 vss 0.00425f
C5720 vdd.n5140 vss 0.0471f
C5721 vdd.n5141 vss 0.00425f
C5722 vdd.n5142 vss 0.00925f
C5723 vdd.n5143 vss 0.00679f
C5724 vdd.n5144 vss 0.00517f
C5725 vdd.n5145 vss 0.00251f
C5726 vdd.n5146 vss 0.0471f
C5727 vdd.n5147 vss 0.00251f
C5728 vdd.n5148 vss 0.0112f
C5729 vdd.n5149 vss 0.0128f
C5730 vdd.n5150 vss 0.0666f
C5731 vdd.n5151 vss 0.118f
C5732 vdd.n5152 vss 0.121f
C5733 vdd.n5153 vss 0.00324f
C5734 vdd.n5154 vss 0.0112f
C5735 vdd.n5155 vss 0.0128f
C5736 vdd.n5156 vss 0.00413f
C5737 vdd.n5157 vss 0.00413f
C5738 vdd.n5158 vss 0.0471f
C5739 vdd.n5159 vss 0.0471f
C5740 vdd.n5160 vss 0.00324f
C5741 vdd.n5161 vss 0.00413f
C5742 vdd.n5162 vss 0.00413f
C5743 vdd.n5163 vss 0.00679f
C5744 vdd.n5164 vss 0.00413f
C5745 vdd.n5165 vss 0.0471f
C5746 vdd.n5166 vss 0.00324f
C5747 vdd.n5167 vss 0.0424f
C5748 vdd.n5168 vss 0.00324f
C5749 vdd.n5169 vss 0.0128f
C5750 vdd.n5170 vss 0.02f
C5751 vdd.n5171 vss 0.0132f
C5752 vdd.n5172 vss 0.00925f
C5753 vdd.n5173 vss 0.00425f
C5754 vdd.n5175 vss 0.0471f
C5755 vdd.n5176 vss 0.00425f
C5756 vdd.n5177 vss 0.00413f
C5757 vdd.n5178 vss 0.00251f
C5758 vdd.n5179 vss 0.0471f
C5759 vdd.n5180 vss 0.00251f
C5760 vdd.n5181 vss 0.00517f
C5761 vdd.n5182 vss 0.00679f
C5762 vdd.n5183 vss 0.00324f
C5763 vdd.n5184 vss 0.00324f
C5764 vdd.n5185 vss 0.0132f
C5765 vdd.n5186 vss 0.0424f
C5766 vdd.n5187 vss 0.02f
C5767 vdd.n5188 vss 0.00425f
C5768 vdd.n5190 vss 0.0471f
C5769 vdd.n5191 vss 0.00425f
C5770 vdd.n5192 vss 0.00925f
C5771 vdd.n5193 vss 0.00679f
C5772 vdd.n5194 vss 0.00517f
C5773 vdd.n5195 vss 0.00251f
C5774 vdd.n5196 vss 0.0471f
C5775 vdd.n5197 vss 0.00251f
C5776 vdd.n5198 vss 0.0112f
C5777 vdd.n5199 vss 0.0955f
C5778 vdd.n5200 vss 0.0608f
C5779 vdd.n5201 vss 0.00324f
C5780 vdd.n5202 vss 0.0112f
C5781 vdd.n5203 vss 0.0128f
C5782 vdd.n5204 vss 0.00413f
C5783 vdd.n5205 vss 0.00413f
C5784 vdd.n5206 vss 0.0471f
C5785 vdd.n5207 vss 0.0471f
C5786 vdd.n5208 vss 0.00324f
C5787 vdd.n5209 vss 0.00413f
C5788 vdd.n5210 vss 0.00413f
C5789 vdd.n5211 vss 0.00679f
C5790 vdd.n5212 vss 0.00413f
C5791 vdd.n5213 vss 0.0471f
C5792 vdd.n5214 vss 0.00324f
C5793 vdd.n5215 vss 0.0424f
C5794 vdd.n5216 vss 0.00324f
C5795 vdd.n5217 vss 0.0128f
C5796 vdd.n5218 vss 0.02f
C5797 vdd.n5219 vss 0.0132f
C5798 vdd.n5220 vss 0.00925f
C5799 vdd.n5221 vss 0.00425f
C5800 vdd.n5223 vss 0.0471f
C5801 vdd.n5224 vss 0.00425f
C5802 vdd.n5225 vss 0.00413f
C5803 vdd.n5226 vss 0.00251f
C5804 vdd.n5227 vss 0.0471f
C5805 vdd.n5228 vss 0.00251f
C5806 vdd.n5229 vss 0.00517f
C5807 vdd.n5230 vss 0.00679f
C5808 vdd.n5231 vss 0.00324f
C5809 vdd.n5232 vss 0.00324f
C5810 vdd.n5233 vss 0.0132f
C5811 vdd.n5234 vss 0.0424f
C5812 vdd.n5235 vss 0.02f
C5813 vdd.n5236 vss 0.00425f
C5814 vdd.n5238 vss 0.0471f
C5815 vdd.n5239 vss 0.00425f
C5816 vdd.n5240 vss 0.00925f
C5817 vdd.n5241 vss 0.00679f
C5818 vdd.n5242 vss 0.00517f
C5819 vdd.n5243 vss 0.00251f
C5820 vdd.n5244 vss 0.0471f
C5821 vdd.n5245 vss 0.00251f
C5822 vdd.n5246 vss 0.0112f
C5823 vdd.n5247 vss 0.0128f
C5824 vdd.n5248 vss 0.0666f
C5825 vdd.n5249 vss 0.118f
C5826 vdd.n5250 vss 0.0935f
C5827 vdd.n5251 vss 0.00324f
C5828 vdd.n5252 vss 0.0112f
C5829 vdd.n5253 vss 0.0128f
C5830 vdd.n5254 vss 0.00413f
C5831 vdd.n5255 vss 0.00413f
C5832 vdd.n5256 vss 0.0471f
C5833 vdd.n5257 vss 0.0471f
C5834 vdd.n5258 vss 0.00324f
C5835 vdd.n5259 vss 0.00413f
C5836 vdd.n5260 vss 0.00413f
C5837 vdd.n5261 vss 0.00679f
C5838 vdd.n5262 vss 0.00413f
C5839 vdd.n5263 vss 0.0471f
C5840 vdd.n5264 vss 0.00324f
C5841 vdd.n5265 vss 0.0424f
C5842 vdd.n5266 vss 0.00324f
C5843 vdd.n5267 vss 0.0128f
C5844 vdd.n5268 vss 0.02f
C5845 vdd.n5269 vss 0.0132f
C5846 vdd.n5270 vss 0.00925f
C5847 vdd.n5271 vss 0.00425f
C5848 vdd.n5273 vss 0.0471f
C5849 vdd.n5274 vss 0.00425f
C5850 vdd.n5275 vss 0.00413f
C5851 vdd.n5276 vss 0.00251f
C5852 vdd.n5277 vss 0.0471f
C5853 vdd.n5278 vss 0.00251f
C5854 vdd.n5279 vss 0.00517f
C5855 vdd.n5280 vss 0.00679f
C5856 vdd.n5281 vss 0.00324f
C5857 vdd.n5282 vss 0.00324f
C5858 vdd.n5283 vss 0.0132f
C5859 vdd.n5284 vss 0.0424f
C5860 vdd.n5285 vss 0.02f
C5861 vdd.n5286 vss 0.00425f
C5862 vdd.n5288 vss 0.0471f
C5863 vdd.n5289 vss 0.00425f
C5864 vdd.n5290 vss 0.00925f
C5865 vdd.n5291 vss 0.00679f
C5866 vdd.n5292 vss 0.00517f
C5867 vdd.n5293 vss 0.00251f
C5868 vdd.n5294 vss 0.0471f
C5869 vdd.n5295 vss 0.00251f
C5870 vdd.n5296 vss 0.0112f
C5871 vdd.n5297 vss 0.0128f
C5872 vdd.n5298 vss 0.00324f
C5873 vdd.n5299 vss 0.0112f
C5874 vdd.n5300 vss 0.0128f
C5875 vdd.n5301 vss 0.00413f
C5876 vdd.n5302 vss 0.00413f
C5877 vdd.n5303 vss 0.0471f
C5878 vdd.n5304 vss 0.0471f
C5879 vdd.n5305 vss 0.00324f
C5880 vdd.n5306 vss 0.00413f
C5881 vdd.n5307 vss 0.00413f
C5882 vdd.n5308 vss 0.00679f
C5883 vdd.n5309 vss 0.00413f
C5884 vdd.n5310 vss 0.0471f
C5885 vdd.n5311 vss 0.00324f
C5886 vdd.n5312 vss 0.0424f
C5887 vdd.n5313 vss 0.00324f
C5888 vdd.n5314 vss 0.0128f
C5889 vdd.n5315 vss 0.02f
C5890 vdd.n5316 vss 0.0132f
C5891 vdd.n5317 vss 0.00925f
C5892 vdd.n5318 vss 0.00425f
C5893 vdd.n5320 vss 0.0471f
C5894 vdd.n5321 vss 0.00425f
C5895 vdd.n5322 vss 0.00413f
C5896 vdd.n5323 vss 0.00251f
C5897 vdd.n5324 vss 0.0471f
C5898 vdd.n5325 vss 0.00251f
C5899 vdd.n5326 vss 0.00517f
C5900 vdd.n5327 vss 0.00679f
C5901 vdd.n5328 vss 0.00324f
C5902 vdd.n5329 vss 0.00324f
C5903 vdd.n5330 vss 0.0132f
C5904 vdd.n5331 vss 0.0424f
C5905 vdd.n5332 vss 0.02f
C5906 vdd.n5333 vss 0.00425f
C5907 vdd.n5335 vss 0.0471f
C5908 vdd.n5336 vss 0.00425f
C5909 vdd.n5337 vss 0.00925f
C5910 vdd.n5338 vss 0.00679f
C5911 vdd.n5339 vss 0.00517f
C5912 vdd.n5340 vss 0.00251f
C5913 vdd.n5341 vss 0.0471f
C5914 vdd.n5342 vss 0.00251f
C5915 vdd.n5343 vss 0.0112f
C5916 vdd.n5344 vss 0.0128f
C5917 vdd.n5345 vss 0.144f
C5918 vdd.n5346 vss 0.143f
C5919 vdd.n5347 vss 0.0608f
C5920 vdd.n5348 vss 0.00324f
C5921 vdd.n5349 vss 0.0112f
C5922 vdd.n5350 vss 0.0128f
C5923 vdd.n5351 vss 0.00413f
C5924 vdd.n5352 vss 0.00413f
C5925 vdd.n5353 vss 0.0471f
C5926 vdd.n5354 vss 0.0471f
C5927 vdd.n5355 vss 0.00324f
C5928 vdd.n5356 vss 0.00413f
C5929 vdd.n5357 vss 0.00413f
C5930 vdd.n5358 vss 0.00679f
C5931 vdd.n5359 vss 0.00413f
C5932 vdd.n5360 vss 0.0471f
C5933 vdd.n5361 vss 0.00324f
C5934 vdd.n5362 vss 0.0424f
C5935 vdd.n5363 vss 0.00324f
C5936 vdd.n5364 vss 0.0128f
C5937 vdd.n5365 vss 0.02f
C5938 vdd.n5366 vss 0.0132f
C5939 vdd.n5367 vss 0.00925f
C5940 vdd.n5368 vss 0.00425f
C5941 vdd.n5370 vss 0.0471f
C5942 vdd.n5371 vss 0.00425f
C5943 vdd.n5372 vss 0.00413f
C5944 vdd.n5373 vss 0.00251f
C5945 vdd.n5374 vss 0.0471f
C5946 vdd.n5375 vss 0.00251f
C5947 vdd.n5376 vss 0.00517f
C5948 vdd.n5377 vss 0.00679f
C5949 vdd.n5378 vss 0.00324f
C5950 vdd.n5379 vss 0.00324f
C5951 vdd.n5380 vss 0.0132f
C5952 vdd.n5381 vss 0.0424f
C5953 vdd.n5382 vss 0.02f
C5954 vdd.n5383 vss 0.00425f
C5955 vdd.n5385 vss 0.0471f
C5956 vdd.n5386 vss 0.00425f
C5957 vdd.n5387 vss 0.00925f
C5958 vdd.n5388 vss 0.00679f
C5959 vdd.n5389 vss 0.00517f
C5960 vdd.n5390 vss 0.00251f
C5961 vdd.n5391 vss 0.0471f
C5962 vdd.n5392 vss 0.00251f
C5963 vdd.n5393 vss 0.0112f
C5964 vdd.n5394 vss 0.0128f
C5965 vdd.n5395 vss 0.0666f
C5966 vdd.n5396 vss 0.118f
C5967 vdd.n5397 vss 0.121f
C5968 vdd.n5398 vss 0.00324f
C5969 vdd.n5399 vss 0.0112f
C5970 vdd.n5400 vss 0.0128f
C5971 vdd.n5401 vss 0.00413f
C5972 vdd.n5402 vss 0.00413f
C5973 vdd.n5403 vss 0.0471f
C5974 vdd.n5404 vss 0.0471f
C5975 vdd.n5405 vss 0.00324f
C5976 vdd.n5406 vss 0.00413f
C5977 vdd.n5407 vss 0.00413f
C5978 vdd.n5408 vss 0.00679f
C5979 vdd.n5409 vss 0.00413f
C5980 vdd.n5410 vss 0.0471f
C5981 vdd.n5411 vss 0.00324f
C5982 vdd.n5412 vss 0.0424f
C5983 vdd.n5413 vss 0.00324f
C5984 vdd.n5414 vss 0.0128f
C5985 vdd.n5415 vss 0.02f
C5986 vdd.n5416 vss 0.0132f
C5987 vdd.n5417 vss 0.00925f
C5988 vdd.n5418 vss 0.00425f
C5989 vdd.n5420 vss 0.0471f
C5990 vdd.n5421 vss 0.00425f
C5991 vdd.n5422 vss 0.00413f
C5992 vdd.n5423 vss 0.00251f
C5993 vdd.n5424 vss 0.0471f
C5994 vdd.n5425 vss 0.00251f
C5995 vdd.n5426 vss 0.00517f
C5996 vdd.n5427 vss 0.00679f
C5997 vdd.n5428 vss 0.00324f
C5998 vdd.n5429 vss 0.00324f
C5999 vdd.n5430 vss 0.0132f
C6000 vdd.n5431 vss 0.0424f
C6001 vdd.n5432 vss 0.02f
C6002 vdd.n5433 vss 0.00425f
C6003 vdd.n5435 vss 0.0471f
C6004 vdd.n5436 vss 0.00425f
C6005 vdd.n5437 vss 0.00925f
C6006 vdd.n5438 vss 0.00679f
C6007 vdd.n5439 vss 0.00517f
C6008 vdd.n5440 vss 0.00251f
C6009 vdd.n5441 vss 0.0471f
C6010 vdd.n5442 vss 0.00251f
C6011 vdd.n5443 vss 0.0112f
C6012 vdd.n5444 vss 0.0955f
C6013 vdd.n5445 vss 0.0608f
C6014 vdd.n5446 vss 0.00324f
C6015 vdd.n5447 vss 0.0112f
C6016 vdd.n5448 vss 0.0128f
C6017 vdd.n5449 vss 0.00413f
C6018 vdd.n5450 vss 0.00413f
C6019 vdd.n5451 vss 0.0471f
C6020 vdd.n5452 vss 0.0471f
C6021 vdd.n5453 vss 0.00324f
C6022 vdd.n5454 vss 0.00413f
C6023 vdd.n5455 vss 0.00413f
C6024 vdd.n5456 vss 0.00679f
C6025 vdd.n5457 vss 0.00413f
C6026 vdd.n5458 vss 0.0471f
C6027 vdd.n5459 vss 0.00324f
C6028 vdd.n5460 vss 0.0424f
C6029 vdd.n5461 vss 0.00324f
C6030 vdd.n5462 vss 0.0128f
C6031 vdd.n5463 vss 0.02f
C6032 vdd.n5464 vss 0.0132f
C6033 vdd.n5465 vss 0.00925f
C6034 vdd.n5466 vss 0.00425f
C6035 vdd.n5468 vss 0.0471f
C6036 vdd.n5469 vss 0.00425f
C6037 vdd.n5470 vss 0.00413f
C6038 vdd.n5471 vss 0.00251f
C6039 vdd.n5472 vss 0.0471f
C6040 vdd.n5473 vss 0.00251f
C6041 vdd.n5474 vss 0.00517f
C6042 vdd.n5475 vss 0.00679f
C6043 vdd.n5476 vss 0.00324f
C6044 vdd.n5477 vss 0.00324f
C6045 vdd.n5478 vss 0.0132f
C6046 vdd.n5479 vss 0.0424f
C6047 vdd.n5480 vss 0.02f
C6048 vdd.n5481 vss 0.00425f
C6049 vdd.n5483 vss 0.0471f
C6050 vdd.n5484 vss 0.00425f
C6051 vdd.n5485 vss 0.00925f
C6052 vdd.n5486 vss 0.00679f
C6053 vdd.n5487 vss 0.00517f
C6054 vdd.n5488 vss 0.00251f
C6055 vdd.n5489 vss 0.0471f
C6056 vdd.n5490 vss 0.00251f
C6057 vdd.n5491 vss 0.0112f
C6058 vdd.n5492 vss 0.0128f
C6059 vdd.n5493 vss 0.0666f
C6060 vdd.n5494 vss 0.0912f
C6061 vdd.n5495 vss 0.0824f
C6062 vdd.n5496 vss 0.0567f
C6063 vdd.n5497 vss 0.00324f
C6064 vdd.n5498 vss 0.0112f
C6065 vdd.n5499 vss 0.0128f
C6066 vdd.n5500 vss 0.00413f
C6067 vdd.n5501 vss 0.00413f
C6068 vdd.n5502 vss 0.0471f
C6069 vdd.n5503 vss 0.0471f
C6070 vdd.n5504 vss 0.00324f
C6071 vdd.n5505 vss 0.00413f
C6072 vdd.n5506 vss 0.00413f
C6073 vdd.n5507 vss 0.00679f
C6074 vdd.n5508 vss 0.00413f
C6075 vdd.n5509 vss 0.0471f
C6076 vdd.n5510 vss 0.00324f
C6077 vdd.n5511 vss 0.0424f
C6078 vdd.n5512 vss 0.00324f
C6079 vdd.n5513 vss 0.0128f
C6080 vdd.n5514 vss 0.02f
C6081 vdd.n5515 vss 0.0132f
C6082 vdd.n5516 vss 0.00925f
C6083 vdd.n5517 vss 0.00425f
C6084 vdd.n5519 vss 0.0471f
C6085 vdd.n5520 vss 0.00425f
C6086 vdd.n5521 vss 0.00413f
C6087 vdd.n5522 vss 0.00251f
C6088 vdd.n5523 vss 0.0471f
C6089 vdd.n5524 vss 0.00251f
C6090 vdd.n5525 vss 0.00517f
C6091 vdd.n5526 vss 0.00679f
C6092 vdd.n5527 vss 0.00324f
C6093 vdd.n5528 vss 0.00324f
C6094 vdd.n5529 vss 0.0132f
C6095 vdd.n5530 vss 0.0424f
C6096 vdd.n5531 vss 0.02f
C6097 vdd.n5532 vss 0.00425f
C6098 vdd.n5534 vss 0.0471f
C6099 vdd.n5535 vss 0.00425f
C6100 vdd.n5536 vss 0.00925f
C6101 vdd.n5537 vss 0.00679f
C6102 vdd.n5538 vss 0.00517f
C6103 vdd.n5539 vss 0.00251f
C6104 vdd.n5540 vss 0.0471f
C6105 vdd.n5541 vss 0.00251f
C6106 vdd.n5542 vss 0.0112f
C6107 vdd.n5543 vss 0.0128f
C6108 vdd.n5544 vss 0.00324f
C6109 vdd.n5545 vss 0.0112f
C6110 vdd.n5546 vss 0.0128f
C6111 vdd.n5547 vss 0.00413f
C6112 vdd.n5548 vss 0.00413f
C6113 vdd.n5549 vss 0.0471f
C6114 vdd.n5550 vss 0.0471f
C6115 vdd.n5551 vss 0.00324f
C6116 vdd.n5552 vss 0.00413f
C6117 vdd.n5553 vss 0.00413f
C6118 vdd.n5554 vss 0.00679f
C6119 vdd.n5555 vss 0.00413f
C6120 vdd.n5556 vss 0.0471f
C6121 vdd.n5557 vss 0.00324f
C6122 vdd.n5558 vss 0.0424f
C6123 vdd.n5559 vss 0.00324f
C6124 vdd.n5560 vss 0.0128f
C6125 vdd.n5561 vss 0.02f
C6126 vdd.n5562 vss 0.0132f
C6127 vdd.n5563 vss 0.00925f
C6128 vdd.n5564 vss 0.00425f
C6129 vdd.n5566 vss 0.0471f
C6130 vdd.n5567 vss 0.00425f
C6131 vdd.n5568 vss 0.00413f
C6132 vdd.n5569 vss 0.00251f
C6133 vdd.n5570 vss 0.0471f
C6134 vdd.n5571 vss 0.00251f
C6135 vdd.n5572 vss 0.00517f
C6136 vdd.n5573 vss 0.00679f
C6137 vdd.n5574 vss 0.00324f
C6138 vdd.n5575 vss 0.00324f
C6139 vdd.n5576 vss 0.0132f
C6140 vdd.n5577 vss 0.0424f
C6141 vdd.n5578 vss 0.02f
C6142 vdd.n5579 vss 0.00425f
C6143 vdd.n5581 vss 0.0471f
C6144 vdd.n5582 vss 0.00425f
C6145 vdd.n5583 vss 0.00925f
C6146 vdd.n5584 vss 0.00679f
C6147 vdd.n5585 vss 0.00517f
C6148 vdd.n5586 vss 0.00251f
C6149 vdd.n5587 vss 0.0471f
C6150 vdd.n5588 vss 0.00251f
C6151 vdd.n5589 vss 0.0112f
C6152 vdd.n5590 vss 0.0128f
C6153 vdd.n5591 vss 0.144f
C6154 vdd.n5592 vss 0.143f
C6155 vdd.n5593 vss 0.0608f
C6156 vdd.n5594 vss 0.00324f
C6157 vdd.n5595 vss 0.0112f
C6158 vdd.n5596 vss 0.0128f
C6159 vdd.n5597 vss 0.00413f
C6160 vdd.n5598 vss 0.00413f
C6161 vdd.n5599 vss 0.0471f
C6162 vdd.n5600 vss 0.0471f
C6163 vdd.n5601 vss 0.00324f
C6164 vdd.n5602 vss 0.00413f
C6165 vdd.n5603 vss 0.00413f
C6166 vdd.n5604 vss 0.00679f
C6167 vdd.n5605 vss 0.00413f
C6168 vdd.n5606 vss 0.0471f
C6169 vdd.n5607 vss 0.00324f
C6170 vdd.n5608 vss 0.0424f
C6171 vdd.n5609 vss 0.00324f
C6172 vdd.n5610 vss 0.0128f
C6173 vdd.n5611 vss 0.02f
C6174 vdd.n5612 vss 0.0132f
C6175 vdd.n5613 vss 0.00925f
C6176 vdd.n5614 vss 0.00425f
C6177 vdd.n5616 vss 0.0471f
C6178 vdd.n5617 vss 0.00425f
C6179 vdd.n5618 vss 0.00413f
C6180 vdd.n5619 vss 0.00251f
C6181 vdd.n5620 vss 0.0471f
C6182 vdd.n5621 vss 0.00251f
C6183 vdd.n5622 vss 0.00517f
C6184 vdd.n5623 vss 0.00679f
C6185 vdd.n5624 vss 0.00324f
C6186 vdd.n5625 vss 0.00324f
C6187 vdd.n5626 vss 0.0132f
C6188 vdd.n5627 vss 0.0424f
C6189 vdd.n5628 vss 0.02f
C6190 vdd.n5629 vss 0.00425f
C6191 vdd.n5631 vss 0.0471f
C6192 vdd.n5632 vss 0.00425f
C6193 vdd.n5633 vss 0.00925f
C6194 vdd.n5634 vss 0.00679f
C6195 vdd.n5635 vss 0.00517f
C6196 vdd.n5636 vss 0.00251f
C6197 vdd.n5637 vss 0.0471f
C6198 vdd.n5638 vss 0.00251f
C6199 vdd.n5639 vss 0.0112f
C6200 vdd.n5640 vss 0.0128f
C6201 vdd.n5641 vss 0.0666f
C6202 vdd.n5642 vss 0.118f
C6203 vdd.n5643 vss 0.121f
C6204 vdd.n5644 vss 0.00324f
C6205 vdd.n5645 vss 0.0112f
C6206 vdd.n5646 vss 0.0128f
C6207 vdd.n5647 vss 0.00413f
C6208 vdd.n5648 vss 0.00413f
C6209 vdd.n5649 vss 0.0471f
C6210 vdd.n5650 vss 0.0471f
C6211 vdd.n5651 vss 0.00324f
C6212 vdd.n5652 vss 0.00413f
C6213 vdd.n5653 vss 0.00413f
C6214 vdd.n5654 vss 0.00679f
C6215 vdd.n5655 vss 0.00413f
C6216 vdd.n5656 vss 0.0471f
C6217 vdd.n5657 vss 0.00324f
C6218 vdd.n5658 vss 0.0424f
C6219 vdd.n5659 vss 0.00324f
C6220 vdd.n5660 vss 0.0128f
C6221 vdd.n5661 vss 0.02f
C6222 vdd.n5662 vss 0.0132f
C6223 vdd.n5663 vss 0.00925f
C6224 vdd.n5664 vss 0.00425f
C6225 vdd.n5666 vss 0.0471f
C6226 vdd.n5667 vss 0.00425f
C6227 vdd.n5668 vss 0.00413f
C6228 vdd.n5669 vss 0.00251f
C6229 vdd.n5670 vss 0.0471f
C6230 vdd.n5671 vss 0.00251f
C6231 vdd.n5672 vss 0.00517f
C6232 vdd.n5673 vss 0.00679f
C6233 vdd.n5674 vss 0.00324f
C6234 vdd.n5675 vss 0.00324f
C6235 vdd.n5676 vss 0.0132f
C6236 vdd.n5677 vss 0.0424f
C6237 vdd.n5678 vss 0.02f
C6238 vdd.n5679 vss 0.00425f
C6239 vdd.n5681 vss 0.0471f
C6240 vdd.n5682 vss 0.00425f
C6241 vdd.n5683 vss 0.00925f
C6242 vdd.n5684 vss 0.00679f
C6243 vdd.n5685 vss 0.00517f
C6244 vdd.n5686 vss 0.00251f
C6245 vdd.n5687 vss 0.0471f
C6246 vdd.n5688 vss 0.00251f
C6247 vdd.n5689 vss 0.0112f
C6248 vdd.n5690 vss 0.0955f
C6249 vdd.n5691 vss 0.0608f
C6250 vdd.n5692 vss 0.00324f
C6251 vdd.n5693 vss 0.0112f
C6252 vdd.n5694 vss 0.0128f
C6253 vdd.n5695 vss 0.00413f
C6254 vdd.n5696 vss 0.00413f
C6255 vdd.n5697 vss 0.0471f
C6256 vdd.n5698 vss 0.0471f
C6257 vdd.n5699 vss 0.00324f
C6258 vdd.n5700 vss 0.00413f
C6259 vdd.n5701 vss 0.00413f
C6260 vdd.n5702 vss 0.00679f
C6261 vdd.n5703 vss 0.00413f
C6262 vdd.n5704 vss 0.0471f
C6263 vdd.n5705 vss 0.00324f
C6264 vdd.n5706 vss 0.0424f
C6265 vdd.n5707 vss 0.00324f
C6266 vdd.n5708 vss 0.0128f
C6267 vdd.n5709 vss 0.02f
C6268 vdd.n5710 vss 0.0132f
C6269 vdd.n5711 vss 0.00925f
C6270 vdd.n5712 vss 0.00425f
C6271 vdd.n5714 vss 0.0471f
C6272 vdd.n5715 vss 0.00425f
C6273 vdd.n5716 vss 0.00413f
C6274 vdd.n5717 vss 0.00251f
C6275 vdd.n5718 vss 0.0471f
C6276 vdd.n5719 vss 0.00251f
C6277 vdd.n5720 vss 0.00517f
C6278 vdd.n5721 vss 0.00679f
C6279 vdd.n5722 vss 0.00324f
C6280 vdd.n5723 vss 0.00324f
C6281 vdd.n5724 vss 0.0132f
C6282 vdd.n5725 vss 0.0424f
C6283 vdd.n5726 vss 0.02f
C6284 vdd.n5727 vss 0.00425f
C6285 vdd.n5729 vss 0.0471f
C6286 vdd.n5730 vss 0.00425f
C6287 vdd.n5731 vss 0.00925f
C6288 vdd.n5732 vss 0.00679f
C6289 vdd.n5733 vss 0.00517f
C6290 vdd.n5734 vss 0.00251f
C6291 vdd.n5735 vss 0.0471f
C6292 vdd.n5736 vss 0.00251f
C6293 vdd.n5737 vss 0.0112f
C6294 vdd.n5738 vss 0.0128f
C6295 vdd.n5739 vss 0.0666f
C6296 vdd.n5740 vss 0.299f
C6297 vdd.n5741 vss 0.00324f
C6298 vdd.n5742 vss 0.0112f
C6299 vdd.n5743 vss 0.0128f
C6300 vdd.n5744 vss 0.00413f
C6301 vdd.n5745 vss 0.00413f
C6302 vdd.n5746 vss 0.0471f
C6303 vdd.n5747 vss 0.0471f
C6304 vdd.n5748 vss 0.00324f
C6305 vdd.n5749 vss 0.00413f
C6306 vdd.n5750 vss 0.00413f
C6307 vdd.n5751 vss 0.00679f
C6308 vdd.n5752 vss 0.00413f
C6309 vdd.n5753 vss 0.0471f
C6310 vdd.n5754 vss 0.00324f
C6311 vdd.n5756 vss 0.00925f
C6312 vdd.n5757 vss 0.0471f
C6313 vdd.n5758 vss 0.00425f
C6314 vdd.n5759 vss 0.0424f
C6315 vdd.n5760 vss 0.0132f
C6316 vdd.n5761 vss 0.00324f
C6317 vdd.n5762 vss 0.0128f
C6318 vdd.n5763 vss 0.02f
C6319 vdd.n5764 vss 0.00425f
C6320 vdd.n5765 vss 0.00413f
C6321 vdd.n5766 vss 0.00251f
C6322 vdd.n5767 vss 0.0471f
C6323 vdd.n5768 vss 0.00251f
C6324 vdd.n5769 vss 0.00517f
C6325 vdd.n5770 vss 0.00679f
C6326 vdd.n5771 vss 0.00324f
C6327 vdd.n5772 vss 0.00324f
C6328 vdd.n5773 vss 0.0132f
C6329 vdd.n5774 vss 0.0424f
C6330 vdd.n5775 vss 0.02f
C6331 vdd.n5776 vss 0.00425f
C6332 vdd.n5777 vss 0.0471f
C6333 vdd.n5779 vss 0.00425f
C6334 vdd.n5780 vss 0.00925f
C6335 vdd.n5781 vss 0.00679f
C6336 vdd.n5782 vss 0.00517f
C6337 vdd.n5783 vss 0.00251f
C6338 vdd.n5784 vss 0.0471f
C6339 vdd.n5785 vss 0.00251f
C6340 vdd.n5786 vss 0.0112f
C6341 vdd.n5787 vss 0.0128f
C6342 vdd.n5788 vss 0.0619f
C6343 vdd.n5789 vss 0.262f
C6344 vdd.n5790 vss 0.00324f
C6345 vdd.n5791 vss 0.0112f
C6346 vdd.n5792 vss 0.0128f
C6347 vdd.n5793 vss 0.00413f
C6348 vdd.n5794 vss 0.00413f
C6349 vdd.n5795 vss 0.0471f
C6350 vdd.n5796 vss 0.0471f
C6351 vdd.n5797 vss 0.00324f
C6352 vdd.n5798 vss 0.00413f
C6353 vdd.n5799 vss 0.00413f
C6354 vdd.n5800 vss 0.00679f
C6355 vdd.n5801 vss 0.00413f
C6356 vdd.n5802 vss 0.0471f
C6357 vdd.n5803 vss 0.00324f
C6358 vdd.n5805 vss 0.00925f
C6359 vdd.n5806 vss 0.0471f
C6360 vdd.n5807 vss 0.00425f
C6361 vdd.n5808 vss 0.0424f
C6362 vdd.n5809 vss 0.0132f
C6363 vdd.n5810 vss 0.00324f
C6364 vdd.n5811 vss 0.0128f
C6365 vdd.n5812 vss 0.02f
C6366 vdd.n5813 vss 0.00425f
C6367 vdd.n5814 vss 0.00413f
C6368 vdd.n5815 vss 0.00251f
C6369 vdd.n5816 vss 0.0471f
C6370 vdd.n5817 vss 0.00251f
C6371 vdd.n5818 vss 0.00517f
C6372 vdd.n5819 vss 0.00679f
C6373 vdd.n5820 vss 0.00324f
C6374 vdd.n5821 vss 0.00324f
C6375 vdd.n5822 vss 0.0132f
C6376 vdd.n5823 vss 0.0424f
C6377 vdd.n5824 vss 0.02f
C6378 vdd.n5825 vss 0.00425f
C6379 vdd.n5826 vss 0.0471f
C6380 vdd.n5828 vss 0.00425f
C6381 vdd.n5829 vss 0.00925f
C6382 vdd.n5830 vss 0.00679f
C6383 vdd.n5831 vss 0.00517f
C6384 vdd.n5832 vss 0.00251f
C6385 vdd.n5833 vss 0.0471f
C6386 vdd.n5834 vss 0.00251f
C6387 vdd.n5835 vss 0.0112f
C6388 vdd.n5836 vss 0.0128f
C6389 vdd.n5837 vss 0.146f
C6390 vdd.n5838 vss 0.00324f
C6391 vdd.n5839 vss 0.0112f
C6392 vdd.n5840 vss 0.0128f
C6393 vdd.n5841 vss 0.00413f
C6394 vdd.n5842 vss 0.00413f
C6395 vdd.n5843 vss 0.0471f
C6396 vdd.n5844 vss 0.0471f
C6397 vdd.n5845 vss 0.00324f
C6398 vdd.n5846 vss 0.00413f
C6399 vdd.n5847 vss 0.00413f
C6400 vdd.n5848 vss 0.00679f
C6401 vdd.n5849 vss 0.00413f
C6402 vdd.n5850 vss 0.0471f
C6403 vdd.n5851 vss 0.00324f
C6404 vdd.n5853 vss 0.00925f
C6405 vdd.n5854 vss 0.0471f
C6406 vdd.n5855 vss 0.00425f
C6407 vdd.n5856 vss 0.0424f
C6408 vdd.n5857 vss 0.0132f
C6409 vdd.n5858 vss 0.00324f
C6410 vdd.n5859 vss 0.0128f
C6411 vdd.n5860 vss 0.02f
C6412 vdd.n5861 vss 0.00425f
C6413 vdd.n5862 vss 0.00413f
C6414 vdd.n5863 vss 0.00251f
C6415 vdd.n5864 vss 0.0471f
C6416 vdd.n5865 vss 0.00251f
C6417 vdd.n5866 vss 0.00517f
C6418 vdd.n5867 vss 0.00679f
C6419 vdd.n5868 vss 0.00324f
C6420 vdd.n5869 vss 0.00324f
C6421 vdd.n5870 vss 0.0132f
C6422 vdd.n5871 vss 0.0424f
C6423 vdd.n5872 vss 0.02f
C6424 vdd.n5873 vss 0.00425f
C6425 vdd.n5874 vss 0.0471f
C6426 vdd.n5876 vss 0.00425f
C6427 vdd.n5877 vss 0.00925f
C6428 vdd.n5878 vss 0.00679f
C6429 vdd.n5879 vss 0.00517f
C6430 vdd.n5880 vss 0.00251f
C6431 vdd.n5881 vss 0.0471f
C6432 vdd.n5882 vss 0.00251f
C6433 vdd.n5883 vss 0.0112f
C6434 vdd.n5884 vss 0.0128f
C6435 vdd.n5885 vss 0.146f
C6436 vdd.n5886 vss 0.0596f
C6437 vdd.n5887 vss 0.00324f
C6438 vdd.n5888 vss 0.0112f
C6439 vdd.n5889 vss 0.0128f
C6440 vdd.n5890 vss 0.00413f
C6441 vdd.n5891 vss 0.00413f
C6442 vdd.n5892 vss 0.0471f
C6443 vdd.n5893 vss 0.0471f
C6444 vdd.n5894 vss 0.00324f
C6445 vdd.n5895 vss 0.00413f
C6446 vdd.n5896 vss 0.00413f
C6447 vdd.n5897 vss 0.00679f
C6448 vdd.n5898 vss 0.00413f
C6449 vdd.n5899 vss 0.0471f
C6450 vdd.n5900 vss 0.00324f
C6451 vdd.n5902 vss 0.00925f
C6452 vdd.n5903 vss 0.0471f
C6453 vdd.n5904 vss 0.00425f
C6454 vdd.n5905 vss 0.0424f
C6455 vdd.n5906 vss 0.0132f
C6456 vdd.n5907 vss 0.00324f
C6457 vdd.n5908 vss 0.0128f
C6458 vdd.n5909 vss 0.02f
C6459 vdd.n5910 vss 0.00425f
C6460 vdd.n5911 vss 0.00413f
C6461 vdd.n5912 vss 0.00251f
C6462 vdd.n5913 vss 0.0471f
C6463 vdd.n5914 vss 0.00251f
C6464 vdd.n5915 vss 0.00517f
C6465 vdd.n5916 vss 0.00679f
C6466 vdd.n5917 vss 0.00324f
C6467 vdd.n5918 vss 0.00324f
C6468 vdd.n5919 vss 0.0132f
C6469 vdd.n5920 vss 0.0424f
C6470 vdd.n5921 vss 0.02f
C6471 vdd.n5922 vss 0.00425f
C6472 vdd.n5923 vss 0.0471f
C6473 vdd.n5925 vss 0.00425f
C6474 vdd.n5926 vss 0.00925f
C6475 vdd.n5927 vss 0.00679f
C6476 vdd.n5928 vss 0.00517f
C6477 vdd.n5929 vss 0.00251f
C6478 vdd.n5930 vss 0.0471f
C6479 vdd.n5931 vss 0.00251f
C6480 vdd.n5932 vss 0.0112f
C6481 vdd.n5933 vss 0.0128f
C6482 vdd.n5934 vss 0.0692f
C6483 vdd.n5935 vss 0.118f
C6484 vdd.n5936 vss 0.121f
C6485 vdd.n5937 vss 0.00324f
C6486 vdd.n5938 vss 0.0112f
C6487 vdd.n5939 vss 0.0128f
C6488 vdd.n5940 vss 0.00413f
C6489 vdd.n5941 vss 0.00413f
C6490 vdd.n5942 vss 0.0471f
C6491 vdd.n5943 vss 0.0471f
C6492 vdd.n5944 vss 0.00324f
C6493 vdd.n5945 vss 0.00413f
C6494 vdd.n5946 vss 0.00413f
C6495 vdd.n5947 vss 0.00679f
C6496 vdd.n5948 vss 0.00413f
C6497 vdd.n5949 vss 0.0471f
C6498 vdd.n5950 vss 0.00324f
C6499 vdd.n5952 vss 0.00925f
C6500 vdd.n5953 vss 0.0471f
C6501 vdd.n5954 vss 0.00425f
C6502 vdd.n5955 vss 0.0424f
C6503 vdd.n5956 vss 0.0132f
C6504 vdd.n5957 vss 0.00324f
C6505 vdd.n5958 vss 0.0128f
C6506 vdd.n5959 vss 0.02f
C6507 vdd.n5960 vss 0.00425f
C6508 vdd.n5961 vss 0.00413f
C6509 vdd.n5962 vss 0.00251f
C6510 vdd.n5963 vss 0.0471f
C6511 vdd.n5964 vss 0.00251f
C6512 vdd.n5965 vss 0.00517f
C6513 vdd.n5966 vss 0.00679f
C6514 vdd.n5967 vss 0.00324f
C6515 vdd.n5968 vss 0.00324f
C6516 vdd.n5969 vss 0.0132f
C6517 vdd.n5970 vss 0.0424f
C6518 vdd.n5971 vss 0.02f
C6519 vdd.n5972 vss 0.00425f
C6520 vdd.n5973 vss 0.0471f
C6521 vdd.n5975 vss 0.00425f
C6522 vdd.n5976 vss 0.00925f
C6523 vdd.n5977 vss 0.00679f
C6524 vdd.n5978 vss 0.00517f
C6525 vdd.n5979 vss 0.00251f
C6526 vdd.n5980 vss 0.0471f
C6527 vdd.n5981 vss 0.00251f
C6528 vdd.n5982 vss 0.0112f
C6529 vdd.n5983 vss 0.098f
C6530 vdd.n5984 vss 0.0596f
C6531 vdd.n5985 vss 0.00324f
C6532 vdd.n5986 vss 0.0112f
C6533 vdd.n5987 vss 0.0128f
C6534 vdd.n5988 vss 0.00413f
C6535 vdd.n5989 vss 0.00413f
C6536 vdd.n5990 vss 0.0471f
C6537 vdd.n5991 vss 0.0471f
C6538 vdd.n5992 vss 0.00324f
C6539 vdd.n5993 vss 0.00413f
C6540 vdd.n5994 vss 0.00413f
C6541 vdd.n5995 vss 0.00679f
C6542 vdd.n5996 vss 0.00413f
C6543 vdd.n5997 vss 0.0471f
C6544 vdd.n5998 vss 0.00324f
C6545 vdd.n6000 vss 0.00925f
C6546 vdd.n6001 vss 0.0471f
C6547 vdd.n6002 vss 0.00425f
C6548 vdd.n6003 vss 0.0424f
C6549 vdd.n6004 vss 0.0132f
C6550 vdd.n6005 vss 0.00324f
C6551 vdd.n6006 vss 0.0128f
C6552 vdd.n6007 vss 0.02f
C6553 vdd.n6008 vss 0.00425f
C6554 vdd.n6009 vss 0.00413f
C6555 vdd.n6010 vss 0.00251f
C6556 vdd.n6011 vss 0.0471f
C6557 vdd.n6012 vss 0.00251f
C6558 vdd.n6013 vss 0.00517f
C6559 vdd.n6014 vss 0.00679f
C6560 vdd.n6015 vss 0.00324f
C6561 vdd.n6016 vss 0.00324f
C6562 vdd.n6017 vss 0.0132f
C6563 vdd.n6018 vss 0.0424f
C6564 vdd.n6019 vss 0.02f
C6565 vdd.n6020 vss 0.00425f
C6566 vdd.n6021 vss 0.0471f
C6567 vdd.n6023 vss 0.00425f
C6568 vdd.n6024 vss 0.00925f
C6569 vdd.n6025 vss 0.00679f
C6570 vdd.n6026 vss 0.00517f
C6571 vdd.n6027 vss 0.00251f
C6572 vdd.n6028 vss 0.0471f
C6573 vdd.n6029 vss 0.00251f
C6574 vdd.n6030 vss 0.0112f
C6575 vdd.n6031 vss 0.0128f
C6576 vdd.n6032 vss 0.0692f
C6577 vdd.n6033 vss 0.0912f
C6578 vdd.n6034 vss 0.0824f
C6579 vdd.n6035 vss 0.059f
C6580 vdd.n6036 vss 0.00324f
C6581 vdd.n6037 vss 0.0112f
C6582 vdd.n6038 vss 0.0128f
C6583 vdd.n6039 vss 0.00413f
C6584 vdd.n6040 vss 0.00413f
C6585 vdd.n6041 vss 0.0471f
C6586 vdd.n6042 vss 0.0471f
C6587 vdd.n6043 vss 0.00324f
C6588 vdd.n6044 vss 0.00413f
C6589 vdd.n6045 vss 0.00413f
C6590 vdd.n6046 vss 0.00679f
C6591 vdd.n6047 vss 0.00413f
C6592 vdd.n6048 vss 0.0471f
C6593 vdd.n6049 vss 0.00324f
C6594 vdd.n6051 vss 0.00925f
C6595 vdd.n6052 vss 0.0471f
C6596 vdd.n6053 vss 0.00425f
C6597 vdd.n6054 vss 0.0424f
C6598 vdd.n6055 vss 0.0132f
C6599 vdd.n6056 vss 0.00324f
C6600 vdd.n6057 vss 0.0128f
C6601 vdd.n6058 vss 0.02f
C6602 vdd.n6059 vss 0.00425f
C6603 vdd.n6060 vss 0.00413f
C6604 vdd.n6061 vss 0.00251f
C6605 vdd.n6062 vss 0.0471f
C6606 vdd.n6063 vss 0.00251f
C6607 vdd.n6064 vss 0.00517f
C6608 vdd.n6065 vss 0.00679f
C6609 vdd.n6066 vss 0.00324f
C6610 vdd.n6067 vss 0.00324f
C6611 vdd.n6068 vss 0.0132f
C6612 vdd.n6069 vss 0.0424f
C6613 vdd.n6070 vss 0.02f
C6614 vdd.n6071 vss 0.00425f
C6615 vdd.n6072 vss 0.0471f
C6616 vdd.n6074 vss 0.00425f
C6617 vdd.n6075 vss 0.00925f
C6618 vdd.n6076 vss 0.00679f
C6619 vdd.n6077 vss 0.00517f
C6620 vdd.n6078 vss 0.00251f
C6621 vdd.n6079 vss 0.0471f
C6622 vdd.n6080 vss 0.00251f
C6623 vdd.n6081 vss 0.0112f
C6624 vdd.n6082 vss 0.0128f
C6625 vdd.n6083 vss 0.185f
C6626 vdd.n6084 vss 0.00324f
C6627 vdd.n6085 vss 0.0112f
C6628 vdd.n6086 vss 0.0128f
C6629 vdd.n6087 vss 0.00413f
C6630 vdd.n6088 vss 0.00413f
C6631 vdd.n6089 vss 0.0471f
C6632 vdd.n6090 vss 0.0471f
C6633 vdd.n6091 vss 0.00324f
C6634 vdd.n6092 vss 0.00413f
C6635 vdd.n6093 vss 0.00413f
C6636 vdd.n6094 vss 0.00679f
C6637 vdd.n6095 vss 0.00413f
C6638 vdd.n6096 vss 0.0471f
C6639 vdd.n6097 vss 0.00324f
C6640 vdd.n6099 vss 0.00925f
C6641 vdd.n6100 vss 0.0471f
C6642 vdd.n6101 vss 0.00425f
C6643 vdd.n6102 vss 0.0424f
C6644 vdd.n6103 vss 0.0132f
C6645 vdd.n6104 vss 0.00324f
C6646 vdd.n6105 vss 0.0128f
C6647 vdd.n6106 vss 0.02f
C6648 vdd.n6107 vss 0.00425f
C6649 vdd.n6108 vss 0.00413f
C6650 vdd.n6109 vss 0.00251f
C6651 vdd.n6110 vss 0.0471f
C6652 vdd.n6111 vss 0.00251f
C6653 vdd.n6112 vss 0.00517f
C6654 vdd.n6113 vss 0.00679f
C6655 vdd.n6114 vss 0.00324f
C6656 vdd.n6115 vss 0.00324f
C6657 vdd.n6116 vss 0.0132f
C6658 vdd.n6117 vss 0.0424f
C6659 vdd.n6118 vss 0.02f
C6660 vdd.n6119 vss 0.00425f
C6661 vdd.n6120 vss 0.0471f
C6662 vdd.n6122 vss 0.00425f
C6663 vdd.n6123 vss 0.00925f
C6664 vdd.n6124 vss 0.00679f
C6665 vdd.n6125 vss 0.00517f
C6666 vdd.n6126 vss 0.00251f
C6667 vdd.n6127 vss 0.0471f
C6668 vdd.n6128 vss 0.00251f
C6669 vdd.n6129 vss 0.0112f
C6670 vdd.n6130 vss 0.0128f
C6671 vdd.n6131 vss 0.059f
C6672 vdd.n6132 vss 0.256f
C6673 vdd.n6133 vss 0.00324f
C6674 vdd.n6134 vss 0.0112f
C6675 vdd.n6135 vss 0.0128f
C6676 vdd.n6136 vss 0.00413f
C6677 vdd.n6137 vss 0.00413f
C6678 vdd.n6138 vss 0.0471f
C6679 vdd.n6139 vss 0.0471f
C6680 vdd.n6140 vss 0.00324f
C6681 vdd.n6141 vss 0.00413f
C6682 vdd.n6142 vss 0.00413f
C6683 vdd.n6143 vss 0.00679f
C6684 vdd.n6144 vss 0.00413f
C6685 vdd.n6145 vss 0.0471f
C6686 vdd.n6146 vss 0.00324f
C6687 vdd.n6148 vss 0.00925f
C6688 vdd.n6149 vss 0.0471f
C6689 vdd.n6150 vss 0.00425f
C6690 vdd.n6151 vss 0.0424f
C6691 vdd.n6152 vss 0.0132f
C6692 vdd.n6153 vss 0.00324f
C6693 vdd.n6154 vss 0.0128f
C6694 vdd.n6155 vss 0.02f
C6695 vdd.n6156 vss 0.00425f
C6696 vdd.n6157 vss 0.00413f
C6697 vdd.n6158 vss 0.00251f
C6698 vdd.n6159 vss 0.0471f
C6699 vdd.n6160 vss 0.00251f
C6700 vdd.n6161 vss 0.00517f
C6701 vdd.n6162 vss 0.00679f
C6702 vdd.n6163 vss 0.00324f
C6703 vdd.n6164 vss 0.00324f
C6704 vdd.n6165 vss 0.0132f
C6705 vdd.n6166 vss 0.0424f
C6706 vdd.n6167 vss 0.02f
C6707 vdd.n6168 vss 0.00425f
C6708 vdd.n6169 vss 0.0471f
C6709 vdd.n6171 vss 0.00425f
C6710 vdd.n6172 vss 0.00925f
C6711 vdd.n6173 vss 0.00679f
C6712 vdd.n6174 vss 0.00517f
C6713 vdd.n6175 vss 0.00251f
C6714 vdd.n6176 vss 0.0471f
C6715 vdd.n6177 vss 0.00251f
C6716 vdd.n6178 vss 0.0112f
C6717 vdd.n6179 vss 0.0128f
C6718 vdd.n6180 vss 0.123f
C6719 vdd.n6181 vss 0.0596f
C6720 vdd.n6182 vss 0.00324f
C6721 vdd.n6183 vss 0.0112f
C6722 vdd.n6184 vss 0.0128f
C6723 vdd.n6185 vss 0.00413f
C6724 vdd.n6186 vss 0.00413f
C6725 vdd.n6187 vss 0.0471f
C6726 vdd.n6188 vss 0.0471f
C6727 vdd.n6189 vss 0.00324f
C6728 vdd.n6190 vss 0.00413f
C6729 vdd.n6191 vss 0.00413f
C6730 vdd.n6192 vss 0.00679f
C6731 vdd.n6193 vss 0.00413f
C6732 vdd.n6194 vss 0.0471f
C6733 vdd.n6195 vss 0.00324f
C6734 vdd.n6197 vss 0.00925f
C6735 vdd.n6198 vss 0.0471f
C6736 vdd.n6199 vss 0.00425f
C6737 vdd.n6200 vss 0.0424f
C6738 vdd.n6201 vss 0.0132f
C6739 vdd.n6202 vss 0.00324f
C6740 vdd.n6203 vss 0.0128f
C6741 vdd.n6204 vss 0.02f
C6742 vdd.n6205 vss 0.00425f
C6743 vdd.n6206 vss 0.00413f
C6744 vdd.n6207 vss 0.00251f
C6745 vdd.n6208 vss 0.0471f
C6746 vdd.n6209 vss 0.00251f
C6747 vdd.n6210 vss 0.00517f
C6748 vdd.n6211 vss 0.00679f
C6749 vdd.n6212 vss 0.00324f
C6750 vdd.n6213 vss 0.00324f
C6751 vdd.n6214 vss 0.0132f
C6752 vdd.n6215 vss 0.0424f
C6753 vdd.n6216 vss 0.02f
C6754 vdd.n6217 vss 0.00425f
C6755 vdd.n6218 vss 0.0471f
C6756 vdd.n6220 vss 0.00425f
C6757 vdd.n6221 vss 0.00925f
C6758 vdd.n6222 vss 0.00679f
C6759 vdd.n6223 vss 0.00517f
C6760 vdd.n6224 vss 0.00251f
C6761 vdd.n6225 vss 0.0471f
C6762 vdd.n6226 vss 0.00251f
C6763 vdd.n6227 vss 0.0112f
C6764 vdd.n6228 vss 0.0128f
C6765 vdd.n6229 vss 0.0692f
C6766 vdd.n6230 vss 0.118f
C6767 vdd.n6231 vss 0.121f
C6768 vdd.n6232 vss 0.00324f
C6769 vdd.n6233 vss 0.0112f
C6770 vdd.n6234 vss 0.0128f
C6771 vdd.n6235 vss 0.00413f
C6772 vdd.n6236 vss 0.00413f
C6773 vdd.n6237 vss 0.0471f
C6774 vdd.n6238 vss 0.0471f
C6775 vdd.n6239 vss 0.00324f
C6776 vdd.n6240 vss 0.00413f
C6777 vdd.n6241 vss 0.00413f
C6778 vdd.n6242 vss 0.00679f
C6779 vdd.n6243 vss 0.00413f
C6780 vdd.n6244 vss 0.0471f
C6781 vdd.n6245 vss 0.00324f
C6782 vdd.n6247 vss 0.00925f
C6783 vdd.n6248 vss 0.0471f
C6784 vdd.n6249 vss 0.00425f
C6785 vdd.n6250 vss 0.0424f
C6786 vdd.n6251 vss 0.0132f
C6787 vdd.n6252 vss 0.00324f
C6788 vdd.n6253 vss 0.0128f
C6789 vdd.n6254 vss 0.02f
C6790 vdd.n6255 vss 0.00425f
C6791 vdd.n6256 vss 0.00413f
C6792 vdd.n6257 vss 0.00251f
C6793 vdd.n6258 vss 0.0471f
C6794 vdd.n6259 vss 0.00251f
C6795 vdd.n6260 vss 0.00517f
C6796 vdd.n6261 vss 0.00679f
C6797 vdd.n6262 vss 0.00324f
C6798 vdd.n6263 vss 0.00324f
C6799 vdd.n6264 vss 0.0132f
C6800 vdd.n6265 vss 0.0424f
C6801 vdd.n6266 vss 0.02f
C6802 vdd.n6267 vss 0.00425f
C6803 vdd.n6268 vss 0.0471f
C6804 vdd.n6270 vss 0.00425f
C6805 vdd.n6271 vss 0.00925f
C6806 vdd.n6272 vss 0.00679f
C6807 vdd.n6273 vss 0.00517f
C6808 vdd.n6274 vss 0.00251f
C6809 vdd.n6275 vss 0.0471f
C6810 vdd.n6276 vss 0.00251f
C6811 vdd.n6277 vss 0.0112f
C6812 vdd.n6278 vss 0.098f
C6813 vdd.n6279 vss 0.0596f
C6814 vdd.n6280 vss 0.00324f
C6815 vdd.n6281 vss 0.0112f
C6816 vdd.n6282 vss 0.0128f
C6817 vdd.n6283 vss 0.00413f
C6818 vdd.n6284 vss 0.00413f
C6819 vdd.n6285 vss 0.0471f
C6820 vdd.n6286 vss 0.0471f
C6821 vdd.n6287 vss 0.00324f
C6822 vdd.n6288 vss 0.00413f
C6823 vdd.n6289 vss 0.00413f
C6824 vdd.n6290 vss 0.00679f
C6825 vdd.n6291 vss 0.00413f
C6826 vdd.n6292 vss 0.0471f
C6827 vdd.n6293 vss 0.00324f
C6828 vdd.n6295 vss 0.00925f
C6829 vdd.n6296 vss 0.0471f
C6830 vdd.n6297 vss 0.00425f
C6831 vdd.n6298 vss 0.0424f
C6832 vdd.n6299 vss 0.0132f
C6833 vdd.n6300 vss 0.00324f
C6834 vdd.n6301 vss 0.0128f
C6835 vdd.n6302 vss 0.02f
C6836 vdd.n6303 vss 0.00425f
C6837 vdd.n6304 vss 0.00413f
C6838 vdd.n6305 vss 0.00251f
C6839 vdd.n6306 vss 0.0471f
C6840 vdd.n6307 vss 0.00251f
C6841 vdd.n6308 vss 0.00517f
C6842 vdd.n6309 vss 0.00679f
C6843 vdd.n6310 vss 0.00324f
C6844 vdd.n6311 vss 0.00324f
C6845 vdd.n6312 vss 0.0132f
C6846 vdd.n6313 vss 0.0424f
C6847 vdd.n6314 vss 0.02f
C6848 vdd.n6315 vss 0.00425f
C6849 vdd.n6316 vss 0.0471f
C6850 vdd.n6318 vss 0.00425f
C6851 vdd.n6319 vss 0.00925f
C6852 vdd.n6320 vss 0.00679f
C6853 vdd.n6321 vss 0.00517f
C6854 vdd.n6322 vss 0.00251f
C6855 vdd.n6323 vss 0.0471f
C6856 vdd.n6324 vss 0.00251f
C6857 vdd.n6325 vss 0.0112f
C6858 vdd.n6326 vss 0.0128f
C6859 vdd.n6327 vss 0.0692f
C6860 vdd.n6328 vss 0.118f
C6861 vdd.n6329 vss 0.0951f
C6862 vdd.n6330 vss 0.00324f
C6863 vdd.n6331 vss 0.0112f
C6864 vdd.n6332 vss 0.0128f
C6865 vdd.n6333 vss 0.00413f
C6866 vdd.n6334 vss 0.00413f
C6867 vdd.n6335 vss 0.0471f
C6868 vdd.n6336 vss 0.0471f
C6869 vdd.n6337 vss 0.00324f
C6870 vdd.n6338 vss 0.00413f
C6871 vdd.n6339 vss 0.00413f
C6872 vdd.n6340 vss 0.00679f
C6873 vdd.n6341 vss 0.00413f
C6874 vdd.n6342 vss 0.0471f
C6875 vdd.n6343 vss 0.00324f
C6876 vdd.n6345 vss 0.00925f
C6877 vdd.n6346 vss 0.0471f
C6878 vdd.n6347 vss 0.00425f
C6879 vdd.n6348 vss 0.0424f
C6880 vdd.n6349 vss 0.0132f
C6881 vdd.n6350 vss 0.00324f
C6882 vdd.n6351 vss 0.0128f
C6883 vdd.n6352 vss 0.02f
C6884 vdd.n6353 vss 0.00425f
C6885 vdd.n6354 vss 0.00413f
C6886 vdd.n6355 vss 0.00251f
C6887 vdd.n6356 vss 0.0471f
C6888 vdd.n6357 vss 0.00251f
C6889 vdd.n6358 vss 0.00517f
C6890 vdd.n6359 vss 0.00679f
C6891 vdd.n6360 vss 0.00324f
C6892 vdd.n6361 vss 0.00324f
C6893 vdd.n6362 vss 0.0132f
C6894 vdd.n6363 vss 0.0424f
C6895 vdd.n6364 vss 0.02f
C6896 vdd.n6365 vss 0.00425f
C6897 vdd.n6366 vss 0.0471f
C6898 vdd.n6368 vss 0.00425f
C6899 vdd.n6369 vss 0.00925f
C6900 vdd.n6370 vss 0.00679f
C6901 vdd.n6371 vss 0.00517f
C6902 vdd.n6372 vss 0.00251f
C6903 vdd.n6373 vss 0.0471f
C6904 vdd.n6374 vss 0.00251f
C6905 vdd.n6375 vss 0.0112f
C6906 vdd.n6376 vss 0.0128f
C6907 vdd.n6377 vss 0.146f
C6908 vdd.n6378 vss 0.00324f
C6909 vdd.n6379 vss 0.0112f
C6910 vdd.n6380 vss 0.0128f
C6911 vdd.n6381 vss 0.00413f
C6912 vdd.n6382 vss 0.00413f
C6913 vdd.n6383 vss 0.0471f
C6914 vdd.n6384 vss 0.0471f
C6915 vdd.n6385 vss 0.00324f
C6916 vdd.n6386 vss 0.00413f
C6917 vdd.n6387 vss 0.00413f
C6918 vdd.n6388 vss 0.00679f
C6919 vdd.n6389 vss 0.00413f
C6920 vdd.n6390 vss 0.0471f
C6921 vdd.n6391 vss 0.00324f
C6922 vdd.n6393 vss 0.00925f
C6923 vdd.n6394 vss 0.0471f
C6924 vdd.n6395 vss 0.00425f
C6925 vdd.n6396 vss 0.0424f
C6926 vdd.n6397 vss 0.0132f
C6927 vdd.n6398 vss 0.00324f
C6928 vdd.n6399 vss 0.0128f
C6929 vdd.n6400 vss 0.02f
C6930 vdd.n6401 vss 0.00425f
C6931 vdd.n6402 vss 0.00413f
C6932 vdd.n6403 vss 0.00251f
C6933 vdd.n6404 vss 0.0471f
C6934 vdd.n6405 vss 0.00251f
C6935 vdd.n6406 vss 0.00517f
C6936 vdd.n6407 vss 0.00679f
C6937 vdd.n6408 vss 0.00324f
C6938 vdd.n6409 vss 0.00324f
C6939 vdd.n6410 vss 0.0132f
C6940 vdd.n6411 vss 0.0424f
C6941 vdd.n6412 vss 0.02f
C6942 vdd.n6413 vss 0.00425f
C6943 vdd.n6414 vss 0.0471f
C6944 vdd.n6416 vss 0.00425f
C6945 vdd.n6417 vss 0.00925f
C6946 vdd.n6418 vss 0.00679f
C6947 vdd.n6419 vss 0.00517f
C6948 vdd.n6420 vss 0.00251f
C6949 vdd.n6421 vss 0.0471f
C6950 vdd.n6422 vss 0.00251f
C6951 vdd.n6423 vss 0.0112f
C6952 vdd.n6424 vss 0.0128f
C6953 vdd.n6425 vss 0.146f
C6954 vdd.n6426 vss 0.0596f
C6955 vdd.n6427 vss 0.00324f
C6956 vdd.n6428 vss 0.0112f
C6957 vdd.n6429 vss 0.0128f
C6958 vdd.n6430 vss 0.00413f
C6959 vdd.n6431 vss 0.00413f
C6960 vdd.n6432 vss 0.0471f
C6961 vdd.n6433 vss 0.0471f
C6962 vdd.n6434 vss 0.00324f
C6963 vdd.n6435 vss 0.00413f
C6964 vdd.n6436 vss 0.00413f
C6965 vdd.n6437 vss 0.00679f
C6966 vdd.n6438 vss 0.00413f
C6967 vdd.n6439 vss 0.0471f
C6968 vdd.n6440 vss 0.00324f
C6969 vdd.n6442 vss 0.00925f
C6970 vdd.n6443 vss 0.0471f
C6971 vdd.n6444 vss 0.00425f
C6972 vdd.n6445 vss 0.0424f
C6973 vdd.n6446 vss 0.0132f
C6974 vdd.n6447 vss 0.00324f
C6975 vdd.n6448 vss 0.0128f
C6976 vdd.n6449 vss 0.02f
C6977 vdd.n6450 vss 0.00425f
C6978 vdd.n6451 vss 0.00413f
C6979 vdd.n6452 vss 0.00251f
C6980 vdd.n6453 vss 0.0471f
C6981 vdd.n6454 vss 0.00251f
C6982 vdd.n6455 vss 0.00517f
C6983 vdd.n6456 vss 0.00679f
C6984 vdd.n6457 vss 0.00324f
C6985 vdd.n6458 vss 0.00324f
C6986 vdd.n6459 vss 0.0132f
C6987 vdd.n6460 vss 0.0424f
C6988 vdd.n6461 vss 0.02f
C6989 vdd.n6462 vss 0.00425f
C6990 vdd.n6463 vss 0.0471f
C6991 vdd.n6465 vss 0.00425f
C6992 vdd.n6466 vss 0.00925f
C6993 vdd.n6467 vss 0.00679f
C6994 vdd.n6468 vss 0.00517f
C6995 vdd.n6469 vss 0.00251f
C6996 vdd.n6470 vss 0.0471f
C6997 vdd.n6471 vss 0.00251f
C6998 vdd.n6472 vss 0.0112f
C6999 vdd.n6473 vss 0.0128f
C7000 vdd.n6474 vss 0.0692f
C7001 vdd.n6475 vss 0.118f
C7002 vdd.n6476 vss 0.121f
C7003 vdd.n6477 vss 0.00324f
C7004 vdd.n6478 vss 0.0112f
C7005 vdd.n6479 vss 0.0128f
C7006 vdd.n6480 vss 0.00413f
C7007 vdd.n6481 vss 0.00413f
C7008 vdd.n6482 vss 0.0471f
C7009 vdd.n6483 vss 0.0471f
C7010 vdd.n6484 vss 0.00324f
C7011 vdd.n6485 vss 0.00413f
C7012 vdd.n6486 vss 0.00413f
C7013 vdd.n6487 vss 0.00679f
C7014 vdd.n6488 vss 0.00413f
C7015 vdd.n6489 vss 0.0471f
C7016 vdd.n6490 vss 0.00324f
C7017 vdd.n6492 vss 0.00925f
C7018 vdd.n6493 vss 0.0471f
C7019 vdd.n6494 vss 0.00425f
C7020 vdd.n6495 vss 0.0424f
C7021 vdd.n6496 vss 0.0132f
C7022 vdd.n6497 vss 0.00324f
C7023 vdd.n6498 vss 0.0128f
C7024 vdd.n6499 vss 0.02f
C7025 vdd.n6500 vss 0.00425f
C7026 vdd.n6501 vss 0.00413f
C7027 vdd.n6502 vss 0.00251f
C7028 vdd.n6503 vss 0.0471f
C7029 vdd.n6504 vss 0.00251f
C7030 vdd.n6505 vss 0.00517f
C7031 vdd.n6506 vss 0.00679f
C7032 vdd.n6507 vss 0.00324f
C7033 vdd.n6508 vss 0.00324f
C7034 vdd.n6509 vss 0.0132f
C7035 vdd.n6510 vss 0.0424f
C7036 vdd.n6511 vss 0.02f
C7037 vdd.n6512 vss 0.00425f
C7038 vdd.n6513 vss 0.0471f
C7039 vdd.n6515 vss 0.00425f
C7040 vdd.n6516 vss 0.00925f
C7041 vdd.n6517 vss 0.00679f
C7042 vdd.n6518 vss 0.00517f
C7043 vdd.n6519 vss 0.00251f
C7044 vdd.n6520 vss 0.0471f
C7045 vdd.n6521 vss 0.00251f
C7046 vdd.n6522 vss 0.0112f
C7047 vdd.n6523 vss 0.098f
C7048 vdd.n6524 vss 0.0596f
C7049 vdd.n6525 vss 0.00324f
C7050 vdd.n6526 vss 0.0112f
C7051 vdd.n6527 vss 0.0128f
C7052 vdd.n6528 vss 0.00413f
C7053 vdd.n6529 vss 0.00413f
C7054 vdd.n6530 vss 0.0471f
C7055 vdd.n6531 vss 0.0471f
C7056 vdd.n6532 vss 0.00324f
C7057 vdd.n6533 vss 0.00413f
C7058 vdd.n6534 vss 0.00413f
C7059 vdd.n6535 vss 0.00679f
C7060 vdd.n6536 vss 0.00413f
C7061 vdd.n6537 vss 0.0471f
C7062 vdd.n6538 vss 0.00324f
C7063 vdd.n6540 vss 0.00925f
C7064 vdd.n6541 vss 0.0471f
C7065 vdd.n6542 vss 0.00425f
C7066 vdd.n6543 vss 0.0424f
C7067 vdd.n6544 vss 0.0132f
C7068 vdd.n6545 vss 0.00324f
C7069 vdd.n6546 vss 0.0128f
C7070 vdd.n6547 vss 0.02f
C7071 vdd.n6548 vss 0.00425f
C7072 vdd.n6549 vss 0.00413f
C7073 vdd.n6550 vss 0.00251f
C7074 vdd.n6551 vss 0.0471f
C7075 vdd.n6552 vss 0.00251f
C7076 vdd.n6553 vss 0.00517f
C7077 vdd.n6554 vss 0.00679f
C7078 vdd.n6555 vss 0.00324f
C7079 vdd.n6556 vss 0.00324f
C7080 vdd.n6557 vss 0.0132f
C7081 vdd.n6558 vss 0.0424f
C7082 vdd.n6559 vss 0.02f
C7083 vdd.n6560 vss 0.00425f
C7084 vdd.n6561 vss 0.0471f
C7085 vdd.n6563 vss 0.00425f
C7086 vdd.n6564 vss 0.00925f
C7087 vdd.n6565 vss 0.00679f
C7088 vdd.n6566 vss 0.00517f
C7089 vdd.n6567 vss 0.00251f
C7090 vdd.n6568 vss 0.0471f
C7091 vdd.n6569 vss 0.00251f
C7092 vdd.n6570 vss 0.0112f
C7093 vdd.n6571 vss 0.0128f
C7094 vdd.n6572 vss 0.0692f
C7095 vdd.n6573 vss 0.0912f
C7096 vdd.n6574 vss 0.0824f
C7097 vdd.n6575 vss 0.059f
C7098 vdd.n6576 vss 0.00324f
C7099 vdd.n6577 vss 0.0112f
C7100 vdd.n6578 vss 0.0128f
C7101 vdd.n6579 vss 0.00413f
C7102 vdd.n6580 vss 0.00413f
C7103 vdd.n6581 vss 0.0471f
C7104 vdd.n6582 vss 0.0471f
C7105 vdd.n6583 vss 0.00324f
C7106 vdd.n6584 vss 0.00413f
C7107 vdd.n6585 vss 0.00413f
C7108 vdd.n6586 vss 0.00679f
C7109 vdd.n6587 vss 0.00413f
C7110 vdd.n6588 vss 0.0471f
C7111 vdd.n6589 vss 0.00324f
C7112 vdd.n6591 vss 0.00925f
C7113 vdd.n6592 vss 0.0471f
C7114 vdd.n6593 vss 0.00425f
C7115 vdd.n6594 vss 0.0424f
C7116 vdd.n6595 vss 0.0132f
C7117 vdd.n6596 vss 0.00324f
C7118 vdd.n6597 vss 0.0128f
C7119 vdd.n6598 vss 0.02f
C7120 vdd.n6599 vss 0.00425f
C7121 vdd.n6600 vss 0.00413f
C7122 vdd.n6601 vss 0.00251f
C7123 vdd.n6602 vss 0.0471f
C7124 vdd.n6603 vss 0.00251f
C7125 vdd.n6604 vss 0.00517f
C7126 vdd.n6605 vss 0.00679f
C7127 vdd.n6606 vss 0.00324f
C7128 vdd.n6607 vss 0.00324f
C7129 vdd.n6608 vss 0.0132f
C7130 vdd.n6609 vss 0.0424f
C7131 vdd.n6610 vss 0.02f
C7132 vdd.n6611 vss 0.00425f
C7133 vdd.n6612 vss 0.0471f
C7134 vdd.n6614 vss 0.00425f
C7135 vdd.n6615 vss 0.00925f
C7136 vdd.n6616 vss 0.00679f
C7137 vdd.n6617 vss 0.00517f
C7138 vdd.n6618 vss 0.00251f
C7139 vdd.n6619 vss 0.0471f
C7140 vdd.n6620 vss 0.00251f
C7141 vdd.n6621 vss 0.0112f
C7142 vdd.n6622 vss 0.0128f
C7143 vdd.n6623 vss 0.146f
C7144 vdd.n6624 vss 0.00324f
C7145 vdd.n6625 vss 0.0112f
C7146 vdd.n6626 vss 0.0128f
C7147 vdd.n6627 vss 0.00413f
C7148 vdd.n6628 vss 0.00413f
C7149 vdd.n6629 vss 0.0471f
C7150 vdd.n6630 vss 0.0471f
C7151 vdd.n6631 vss 0.00324f
C7152 vdd.n6632 vss 0.00413f
C7153 vdd.n6633 vss 0.00413f
C7154 vdd.n6634 vss 0.00679f
C7155 vdd.n6635 vss 0.00413f
C7156 vdd.n6636 vss 0.0471f
C7157 vdd.n6637 vss 0.00324f
C7158 vdd.n6639 vss 0.00925f
C7159 vdd.n6640 vss 0.0471f
C7160 vdd.n6641 vss 0.00425f
C7161 vdd.n6642 vss 0.0424f
C7162 vdd.n6643 vss 0.0132f
C7163 vdd.n6644 vss 0.00324f
C7164 vdd.n6645 vss 0.0128f
C7165 vdd.n6646 vss 0.02f
C7166 vdd.n6647 vss 0.00425f
C7167 vdd.n6648 vss 0.00413f
C7168 vdd.n6649 vss 0.00251f
C7169 vdd.n6650 vss 0.0471f
C7170 vdd.n6651 vss 0.00251f
C7171 vdd.n6652 vss 0.00517f
C7172 vdd.n6653 vss 0.00679f
C7173 vdd.n6654 vss 0.00324f
C7174 vdd.n6655 vss 0.00324f
C7175 vdd.n6656 vss 0.0132f
C7176 vdd.n6657 vss 0.0424f
C7177 vdd.n6658 vss 0.02f
C7178 vdd.n6659 vss 0.00425f
C7179 vdd.n6660 vss 0.0471f
C7180 vdd.n6662 vss 0.00425f
C7181 vdd.n6663 vss 0.00925f
C7182 vdd.n6664 vss 0.00679f
C7183 vdd.n6665 vss 0.00517f
C7184 vdd.n6666 vss 0.00251f
C7185 vdd.n6667 vss 0.0471f
C7186 vdd.n6668 vss 0.00251f
C7187 vdd.n6669 vss 0.0112f
C7188 vdd.n6670 vss 0.0128f
C7189 vdd.n6671 vss 0.146f
C7190 vdd.n6672 vss 0.0596f
C7191 vdd.n6673 vss 0.00324f
C7192 vdd.n6674 vss 0.0112f
C7193 vdd.n6675 vss 0.0128f
C7194 vdd.n6676 vss 0.00413f
C7195 vdd.n6677 vss 0.00413f
C7196 vdd.n6678 vss 0.0471f
C7197 vdd.n6679 vss 0.0471f
C7198 vdd.n6680 vss 0.00324f
C7199 vdd.n6681 vss 0.00413f
C7200 vdd.n6682 vss 0.00413f
C7201 vdd.n6683 vss 0.00679f
C7202 vdd.n6684 vss 0.00413f
C7203 vdd.n6685 vss 0.0471f
C7204 vdd.n6686 vss 0.00324f
C7205 vdd.n6688 vss 0.00925f
C7206 vdd.n6689 vss 0.0471f
C7207 vdd.n6690 vss 0.00425f
C7208 vdd.n6691 vss 0.0424f
C7209 vdd.n6692 vss 0.0132f
C7210 vdd.n6693 vss 0.00324f
C7211 vdd.n6694 vss 0.0128f
C7212 vdd.n6695 vss 0.02f
C7213 vdd.n6696 vss 0.00425f
C7214 vdd.n6697 vss 0.00413f
C7215 vdd.n6698 vss 0.00251f
C7216 vdd.n6699 vss 0.0471f
C7217 vdd.n6700 vss 0.00251f
C7218 vdd.n6701 vss 0.00517f
C7219 vdd.n6702 vss 0.00679f
C7220 vdd.n6703 vss 0.00324f
C7221 vdd.n6704 vss 0.00324f
C7222 vdd.n6705 vss 0.0132f
C7223 vdd.n6706 vss 0.0424f
C7224 vdd.n6707 vss 0.02f
C7225 vdd.n6708 vss 0.00425f
C7226 vdd.n6709 vss 0.0471f
C7227 vdd.n6711 vss 0.00425f
C7228 vdd.n6712 vss 0.00925f
C7229 vdd.n6713 vss 0.00679f
C7230 vdd.n6714 vss 0.00517f
C7231 vdd.n6715 vss 0.00251f
C7232 vdd.n6716 vss 0.0471f
C7233 vdd.n6717 vss 0.00251f
C7234 vdd.n6718 vss 0.0112f
C7235 vdd.n6719 vss 0.0128f
C7236 vdd.n6720 vss 0.0692f
C7237 vdd.n6721 vss 0.118f
C7238 vdd.n6722 vss 0.121f
C7239 vdd.n6723 vss 0.00324f
C7240 vdd.n6724 vss 0.0112f
C7241 vdd.n6725 vss 0.0128f
C7242 vdd.n6726 vss 0.00413f
C7243 vdd.n6727 vss 0.00413f
C7244 vdd.n6728 vss 0.0471f
C7245 vdd.n6729 vss 0.0471f
C7246 vdd.n6730 vss 0.00324f
C7247 vdd.n6731 vss 0.00413f
C7248 vdd.n6732 vss 0.00413f
C7249 vdd.n6733 vss 0.00679f
C7250 vdd.n6734 vss 0.00413f
C7251 vdd.n6735 vss 0.0471f
C7252 vdd.n6736 vss 0.00324f
C7253 vdd.n6738 vss 0.00925f
C7254 vdd.n6739 vss 0.0471f
C7255 vdd.n6740 vss 0.00425f
C7256 vdd.n6741 vss 0.0424f
C7257 vdd.n6742 vss 0.0132f
C7258 vdd.n6743 vss 0.00324f
C7259 vdd.n6744 vss 0.0128f
C7260 vdd.n6745 vss 0.02f
C7261 vdd.n6746 vss 0.00425f
C7262 vdd.n6747 vss 0.00413f
C7263 vdd.n6748 vss 0.00251f
C7264 vdd.n6749 vss 0.0471f
C7265 vdd.n6750 vss 0.00251f
C7266 vdd.n6751 vss 0.00517f
C7267 vdd.n6752 vss 0.00679f
C7268 vdd.n6753 vss 0.00324f
C7269 vdd.n6754 vss 0.00324f
C7270 vdd.n6755 vss 0.0132f
C7271 vdd.n6756 vss 0.0424f
C7272 vdd.n6757 vss 0.02f
C7273 vdd.n6758 vss 0.00425f
C7274 vdd.n6759 vss 0.0471f
C7275 vdd.n6761 vss 0.00425f
C7276 vdd.n6762 vss 0.00925f
C7277 vdd.n6763 vss 0.00679f
C7278 vdd.n6764 vss 0.00517f
C7279 vdd.n6765 vss 0.00251f
C7280 vdd.n6766 vss 0.0471f
C7281 vdd.n6767 vss 0.00251f
C7282 vdd.n6768 vss 0.0112f
C7283 vdd.n6769 vss 0.098f
C7284 vdd.n6770 vss 0.0596f
C7285 vdd.n6771 vss 0.00324f
C7286 vdd.n6772 vss 0.0112f
C7287 vdd.n6773 vss 0.0128f
C7288 vdd.n6774 vss 0.00413f
C7289 vdd.n6775 vss 0.00413f
C7290 vdd.n6776 vss 0.0471f
C7291 vdd.n6777 vss 0.0471f
C7292 vdd.n6778 vss 0.00324f
C7293 vdd.n6779 vss 0.00413f
C7294 vdd.n6780 vss 0.00413f
C7295 vdd.n6781 vss 0.00679f
C7296 vdd.n6782 vss 0.00413f
C7297 vdd.n6783 vss 0.0471f
C7298 vdd.n6784 vss 0.00324f
C7299 vdd.n6786 vss 0.00925f
C7300 vdd.n6787 vss 0.0471f
C7301 vdd.n6788 vss 0.00425f
C7302 vdd.n6789 vss 0.0424f
C7303 vdd.n6790 vss 0.0132f
C7304 vdd.n6791 vss 0.00324f
C7305 vdd.n6792 vss 0.0128f
C7306 vdd.n6793 vss 0.02f
C7307 vdd.n6794 vss 0.00425f
C7308 vdd.n6795 vss 0.00413f
C7309 vdd.n6796 vss 0.00251f
C7310 vdd.n6797 vss 0.0471f
C7311 vdd.n6798 vss 0.00251f
C7312 vdd.n6799 vss 0.00517f
C7313 vdd.n6800 vss 0.00679f
C7314 vdd.n6801 vss 0.00324f
C7315 vdd.n6802 vss 0.00324f
C7316 vdd.n6803 vss 0.0132f
C7317 vdd.n6804 vss 0.0424f
C7318 vdd.n6805 vss 0.02f
C7319 vdd.n6806 vss 0.00425f
C7320 vdd.n6807 vss 0.0471f
C7321 vdd.n6809 vss 0.00425f
C7322 vdd.n6810 vss 0.00925f
C7323 vdd.n6811 vss 0.00679f
C7324 vdd.n6812 vss 0.00517f
C7325 vdd.n6813 vss 0.00251f
C7326 vdd.n6814 vss 0.0471f
C7327 vdd.n6815 vss 0.00251f
C7328 vdd.n6816 vss 0.0112f
C7329 vdd.n6817 vss 0.0128f
C7330 vdd.n6818 vss 0.0692f
C7331 vdd.n6819 vss 0.121f
C7332 vdd.n6820 vss 0.291f
C7333 vdd.n6821 vss 0.234f
C7334 vdd.n6822 vss 0.00324f
C7335 vdd.n6823 vss 0.0112f
C7336 vdd.n6824 vss 0.0128f
C7337 vdd.n6825 vss 0.00413f
C7338 vdd.n6826 vss 0.00413f
C7339 vdd.n6827 vss 0.0471f
C7340 vdd.n6828 vss 0.0471f
C7341 vdd.n6829 vss 0.00324f
C7342 vdd.n6830 vss 0.00413f
C7343 vdd.n6831 vss 0.00413f
C7344 vdd.n6832 vss 0.00679f
C7345 vdd.n6833 vss 0.00413f
C7346 vdd.n6834 vss 0.0471f
C7347 vdd.n6835 vss 0.00324f
C7348 vdd.n6837 vss 0.00925f
C7349 vdd.n6838 vss 0.0471f
C7350 vdd.n6839 vss 0.00425f
C7351 vdd.n6840 vss 0.0424f
C7352 vdd.n6841 vss 0.0132f
C7353 vdd.n6842 vss 0.00324f
C7354 vdd.n6843 vss 0.0128f
C7355 vdd.n6844 vss 0.02f
C7356 vdd.n6845 vss 0.00425f
C7357 vdd.n6846 vss 0.00413f
C7358 vdd.n6847 vss 0.00251f
C7359 vdd.n6848 vss 0.0471f
C7360 vdd.n6849 vss 0.00251f
C7361 vdd.n6850 vss 0.00517f
C7362 vdd.n6851 vss 0.00679f
C7363 vdd.n6852 vss 0.00324f
C7364 vdd.n6853 vss 0.00324f
C7365 vdd.n6854 vss 0.0132f
C7366 vdd.n6855 vss 0.0424f
C7367 vdd.n6856 vss 0.02f
C7368 vdd.n6857 vss 0.00425f
C7369 vdd.n6858 vss 0.0471f
C7370 vdd.n6860 vss 0.00425f
C7371 vdd.n6861 vss 0.00925f
C7372 vdd.n6862 vss 0.00679f
C7373 vdd.n6863 vss 0.00517f
C7374 vdd.n6864 vss 0.00251f
C7375 vdd.n6865 vss 0.0471f
C7376 vdd.n6866 vss 0.00251f
C7377 vdd.n6867 vss 0.0112f
C7378 vdd.n6868 vss 0.0128f
C7379 vdd.n6869 vss 0.187f
C7380 vdd.n6870 vss 0.00324f
C7381 vdd.n6871 vss 0.0112f
C7382 vdd.n6872 vss 0.0128f
C7383 vdd.n6873 vss 0.00413f
C7384 vdd.n6874 vss 0.00413f
C7385 vdd.n6875 vss 0.0471f
C7386 vdd.n6876 vss 0.0471f
C7387 vdd.n6877 vss 0.00324f
C7388 vdd.n6878 vss 0.00413f
C7389 vdd.n6879 vss 0.00413f
C7390 vdd.n6880 vss 0.00679f
C7391 vdd.n6881 vss 0.00413f
C7392 vdd.n6882 vss 0.0471f
C7393 vdd.n6883 vss 0.00324f
C7394 vdd.n6885 vss 0.00925f
C7395 vdd.n6886 vss 0.0471f
C7396 vdd.n6887 vss 0.00425f
C7397 vdd.n6888 vss 0.0424f
C7398 vdd.n6889 vss 0.0132f
C7399 vdd.n6890 vss 0.00324f
C7400 vdd.n6891 vss 0.0128f
C7401 vdd.n6892 vss 0.02f
C7402 vdd.n6893 vss 0.00425f
C7403 vdd.n6894 vss 0.00413f
C7404 vdd.n6895 vss 0.00251f
C7405 vdd.n6896 vss 0.0471f
C7406 vdd.n6897 vss 0.00251f
C7407 vdd.n6898 vss 0.00517f
C7408 vdd.n6899 vss 0.00679f
C7409 vdd.n6900 vss 0.00324f
C7410 vdd.n6901 vss 0.00324f
C7411 vdd.n6902 vss 0.0132f
C7412 vdd.n6903 vss 0.0424f
C7413 vdd.n6904 vss 0.02f
C7414 vdd.n6905 vss 0.00425f
C7415 vdd.n6906 vss 0.0471f
C7416 vdd.n6908 vss 0.00425f
C7417 vdd.n6909 vss 0.00925f
C7418 vdd.n6910 vss 0.00679f
C7419 vdd.n6911 vss 0.00517f
C7420 vdd.n6912 vss 0.00251f
C7421 vdd.n6913 vss 0.0471f
C7422 vdd.n6914 vss 0.00251f
C7423 vdd.n6915 vss 0.0112f
C7424 vdd.n6916 vss 0.0128f
C7425 vdd.n6917 vss 0.241f
C7426 vdd.n6918 vss 0.00324f
C7427 vdd.n6919 vss 0.0112f
C7428 vdd.n6920 vss 0.0128f
C7429 vdd.n6921 vss 0.00413f
C7430 vdd.n6922 vss 0.00413f
C7431 vdd.n6923 vss 0.0471f
C7432 vdd.n6924 vss 0.0471f
C7433 vdd.n6925 vss 0.00324f
C7434 vdd.n6926 vss 0.00413f
C7435 vdd.n6927 vss 0.00413f
C7436 vdd.n6928 vss 0.00679f
C7437 vdd.n6929 vss 0.00413f
C7438 vdd.n6930 vss 0.0471f
C7439 vdd.n6931 vss 0.00324f
C7440 vdd.n6932 vss 0.0424f
C7441 vdd.n6933 vss 0.00324f
C7442 vdd.n6934 vss 0.0128f
C7443 vdd.n6935 vss 0.02f
C7444 vdd.n6936 vss 0.0132f
C7445 vdd.n6937 vss 0.00925f
C7446 vdd.n6938 vss 0.00425f
C7447 vdd.n6940 vss 0.0471f
C7448 vdd.n6941 vss 0.00425f
C7449 vdd.n6942 vss 0.00413f
C7450 vdd.n6943 vss 0.00251f
C7451 vdd.n6944 vss 0.0471f
C7452 vdd.n6945 vss 0.00251f
C7453 vdd.n6946 vss 0.00517f
C7454 vdd.n6947 vss 0.00679f
C7455 vdd.n6948 vss 0.00324f
C7456 vdd.n6949 vss 0.00324f
C7457 vdd.n6950 vss 0.0132f
C7458 vdd.n6951 vss 0.0424f
C7459 vdd.n6952 vss 0.02f
C7460 vdd.n6953 vss 0.00425f
C7461 vdd.n6955 vss 0.0471f
C7462 vdd.n6956 vss 0.00425f
C7463 vdd.n6957 vss 0.00925f
C7464 vdd.n6958 vss 0.00679f
C7465 vdd.n6959 vss 0.00517f
C7466 vdd.n6960 vss 0.00251f
C7467 vdd.n6961 vss 0.0471f
C7468 vdd.n6962 vss 0.00251f
C7469 vdd.n6963 vss 0.0112f
C7470 vdd.n6964 vss 0.0128f
C7471 vdd.n6965 vss 0.0599f
C7472 vdd.n6966 vss 0.202f
C7473 vdd.n6967 vss 0.00324f
C7474 vdd.n6968 vss 0.0112f
C7475 vdd.n6969 vss 0.0128f
C7476 vdd.n6970 vss 0.00413f
C7477 vdd.n6971 vss 0.00413f
C7478 vdd.n6972 vss 0.0471f
C7479 vdd.n6973 vss 0.0471f
C7480 vdd.n6974 vss 0.00324f
C7481 vdd.n6975 vss 0.00413f
C7482 vdd.n6976 vss 0.00413f
C7483 vdd.n6977 vss 0.00679f
C7484 vdd.n6978 vss 0.00413f
C7485 vdd.n6979 vss 0.0471f
C7486 vdd.n6980 vss 0.00324f
C7487 vdd.n6982 vss 0.00925f
C7488 vdd.n6983 vss 0.0471f
C7489 vdd.n6984 vss 0.00425f
C7490 vdd.n6985 vss 0.0424f
C7491 vdd.n6986 vss 0.0132f
C7492 vdd.n6987 vss 0.00324f
C7493 vdd.n6988 vss 0.0128f
C7494 vdd.n6989 vss 0.02f
C7495 vdd.n6990 vss 0.00425f
C7496 vdd.n6991 vss 0.00413f
C7497 vdd.n6992 vss 0.00251f
C7498 vdd.n6993 vss 0.0471f
C7499 vdd.n6994 vss 0.00251f
C7500 vdd.n6995 vss 0.00517f
C7501 vdd.n6996 vss 0.00679f
C7502 vdd.n6997 vss 0.00324f
C7503 vdd.n6998 vss 0.00324f
C7504 vdd.n6999 vss 0.0132f
C7505 vdd.n7000 vss 0.0424f
C7506 vdd.n7001 vss 0.02f
C7507 vdd.n7002 vss 0.00425f
C7508 vdd.n7003 vss 0.0471f
C7509 vdd.n7005 vss 0.00425f
C7510 vdd.n7006 vss 0.00925f
C7511 vdd.n7007 vss 0.00679f
C7512 vdd.n7008 vss 0.00517f
C7513 vdd.n7009 vss 0.00251f
C7514 vdd.n7010 vss 0.0471f
C7515 vdd.n7011 vss 0.00251f
C7516 vdd.n7012 vss 0.0112f
C7517 vdd.n7013 vss 0.0128f
C7518 vdd.n7014 vss 0.0692f
C7519 vdd.n7015 vss 0.00324f
C7520 vdd.n7016 vss 0.0112f
C7521 vdd.n7017 vss 0.0128f
C7522 vdd.n7018 vss 0.00413f
C7523 vdd.n7019 vss 0.00413f
C7524 vdd.n7020 vss 0.0471f
C7525 vdd.n7021 vss 0.0471f
C7526 vdd.n7022 vss 0.00324f
C7527 vdd.n7023 vss 0.00413f
C7528 vdd.n7024 vss 0.00413f
C7529 vdd.n7025 vss 0.00679f
C7530 vdd.n7026 vss 0.00413f
C7531 vdd.n7027 vss 0.0471f
C7532 vdd.n7028 vss 0.00324f
C7533 vdd.n7030 vss 0.00925f
C7534 vdd.n7031 vss 0.0471f
C7535 vdd.n7032 vss 0.00425f
C7536 vdd.n7033 vss 0.0424f
C7537 vdd.n7034 vss 0.0132f
C7538 vdd.n7035 vss 0.00324f
C7539 vdd.n7036 vss 0.0128f
C7540 vdd.n7037 vss 0.02f
C7541 vdd.n7038 vss 0.00425f
C7542 vdd.n7039 vss 0.00413f
C7543 vdd.n7040 vss 0.00251f
C7544 vdd.n7041 vss 0.0471f
C7545 vdd.n7042 vss 0.00251f
C7546 vdd.n7043 vss 0.00517f
C7547 vdd.n7044 vss 0.00679f
C7548 vdd.n7045 vss 0.00324f
C7549 vdd.n7046 vss 0.00324f
C7550 vdd.n7047 vss 0.0132f
C7551 vdd.n7048 vss 0.0424f
C7552 vdd.n7049 vss 0.02f
C7553 vdd.n7050 vss 0.00425f
C7554 vdd.n7051 vss 0.0471f
C7555 vdd.n7053 vss 0.00425f
C7556 vdd.n7054 vss 0.00925f
C7557 vdd.n7055 vss 0.00679f
C7558 vdd.n7056 vss 0.00517f
C7559 vdd.n7057 vss 0.00251f
C7560 vdd.n7058 vss 0.0471f
C7561 vdd.n7059 vss 0.00251f
C7562 vdd.n7060 vss 0.0112f
C7563 vdd.n7061 vss 0.0128f
C7564 vdd.n7062 vss 0.0619f
C7565 vdd.n7063 vss 0.00335f
C7566 vdd.n7064 vss 0.0855f
C7567 vdd.n7065 vss 0.00991f
C7568 vdd.n7066 vss 0.0424f
C7569 vdd.n7067 vss 0.00679f
C7570 vdd.n7068 vss 0.00413f
C7571 vdd.n7069 vss 0.0471f
C7572 vdd.n7070 vss 0.00251f
C7573 vdd.n7071 vss 0.00679f
C7574 vdd.n7072 vss 0.00413f
C7575 vdd.n7073 vss 0.00413f
C7576 vdd.n7074 vss 0.0471f
C7577 vdd.n7075 vss 0.00251f
C7578 vdd.n7076 vss 0.00413f
C7579 vdd.n7077 vss 0.00324f
C7580 vdd.n7078 vss 0.0132f
C7581 vdd.n7079 vss 0.0424f
C7582 vdd.n7080 vss 0.00324f
C7583 vdd.n7081 vss 0.00413f
C7584 vdd.n7082 vss 0.00517f
C7585 vdd.n7083 vss 0.00679f
C7586 vdd.n7084 vss 0.00925f
C7587 vdd.n7085 vss 0.00425f
C7588 vdd.n7086 vss 0.0471f
C7589 vdd.n7088 vss 0.00425f
C7590 vdd.n7089 vss 0.02f
C7591 vdd.n7090 vss 0.0128f
C7592 vdd.n7091 vss 0.0105f
C7593 vdd.n7092 vss 0.00251f
C7594 vdd.n7093 vss 0.0471f
C7595 vdd.n7094 vss 0.00517f
C7596 vdd.n7095 vss 0.00251f
C7597 vdd.n7096 vss 0.0471f
C7598 vdd.n7097 vss 0.0471f
C7599 vdd.n7098 vss 0.00324f
C7600 vdd.n7099 vss 0.00324f
C7601 vdd.n7100 vss 0.00805f
C7602 vdd.n7101 vss 0.0112f
C7603 vdd.n7102 vss 0.0128f
C7604 vdd.n7103 vss 0.00324f
C7605 vdd.n7104 vss 0.00324f
C7606 vdd.n7105 vss 0.00413f
C7607 vdd.n7106 vss 0.00425f
C7608 vdd.n7107 vss 0.0471f
C7609 vdd.n7109 vss 0.00425f
C7610 vdd.n7110 vss 0.00925f
C7611 vdd.n7111 vss 0.0107f
C7612 vdd.n7112 vss 0.0126f
C7613 vdd.n7113 vss 0.0516f
C7614 vdd.n7114 vss 0.00163f
C7615 vdd.n7115 vss 0.00145f
C7616 vdd.n7116 vss 0.0271f
C7617 vdd.n7117 vss 0.00324f
C7618 vdd.n7118 vss 0.0112f
C7619 vdd.n7119 vss 0.0128f
C7620 vdd.n7120 vss 0.00413f
C7621 vdd.n7121 vss 0.00413f
C7622 vdd.n7122 vss 0.0471f
C7623 vdd.n7123 vss 0.0471f
C7624 vdd.n7124 vss 0.00324f
C7625 vdd.n7125 vss 0.00413f
C7626 vdd.n7126 vss 0.00413f
C7627 vdd.n7127 vss 0.00679f
C7628 vdd.n7128 vss 0.00413f
C7629 vdd.n7129 vss 0.0471f
C7630 vdd.n7130 vss 0.00324f
C7631 vdd.n7132 vss 0.00925f
C7632 vdd.n7133 vss 0.0471f
C7633 vdd.n7134 vss 0.00425f
C7634 vdd.n7135 vss 0.0424f
C7635 vdd.n7136 vss 0.0132f
C7636 vdd.n7137 vss 0.00324f
C7637 vdd.n7138 vss 0.0128f
C7638 vdd.n7139 vss 0.02f
C7639 vdd.n7140 vss 0.00425f
C7640 vdd.n7141 vss 0.00413f
C7641 vdd.n7142 vss 0.00251f
C7642 vdd.n7143 vss 0.0471f
C7643 vdd.n7144 vss 0.00251f
C7644 vdd.n7145 vss 0.00517f
C7645 vdd.n7146 vss 0.00679f
C7646 vdd.n7147 vss 0.00324f
C7647 vdd.n7148 vss 0.00324f
C7648 vdd.n7149 vss 0.0132f
C7649 vdd.n7150 vss 0.0424f
C7650 vdd.n7151 vss 0.02f
C7651 vdd.n7152 vss 0.00425f
C7652 vdd.n7153 vss 0.0471f
C7653 vdd.n7155 vss 0.00425f
C7654 vdd.n7156 vss 0.00925f
C7655 vdd.n7157 vss 0.00679f
C7656 vdd.n7158 vss 0.00517f
C7657 vdd.n7159 vss 0.00251f
C7658 vdd.n7160 vss 0.0471f
C7659 vdd.n7161 vss 0.00251f
C7660 vdd.n7162 vss 0.0112f
C7661 vdd.n7163 vss 0.0128f
C7662 vdd.n7164 vss 0.0692f
C7663 vdd.n7165 vss 0.00324f
C7664 vdd.n7166 vss 0.0112f
C7665 vdd.n7167 vss 0.0128f
C7666 vdd.n7168 vss 0.00413f
C7667 vdd.n7169 vss 0.00413f
C7668 vdd.n7170 vss 0.0471f
C7669 vdd.n7171 vss 0.0471f
C7670 vdd.n7172 vss 0.00324f
C7671 vdd.n7173 vss 0.00413f
C7672 vdd.n7174 vss 0.00413f
C7673 vdd.n7175 vss 0.00679f
C7674 vdd.n7176 vss 0.00413f
C7675 vdd.n7177 vss 0.0471f
C7676 vdd.n7178 vss 0.00324f
C7677 vdd.n7180 vss 0.00925f
C7678 vdd.n7181 vss 0.0471f
C7679 vdd.n7182 vss 0.00425f
C7680 vdd.n7183 vss 0.0424f
C7681 vdd.n7184 vss 0.0132f
C7682 vdd.n7185 vss 0.00324f
C7683 vdd.n7186 vss 0.0128f
C7684 vdd.n7187 vss 0.02f
C7685 vdd.n7188 vss 0.00425f
C7686 vdd.n7189 vss 0.00413f
C7687 vdd.n7190 vss 0.00251f
C7688 vdd.n7191 vss 0.0471f
C7689 vdd.n7192 vss 0.00251f
C7690 vdd.n7193 vss 0.00517f
C7691 vdd.n7194 vss 0.00679f
C7692 vdd.n7195 vss 0.00324f
C7693 vdd.n7196 vss 0.00324f
C7694 vdd.n7197 vss 0.0132f
C7695 vdd.n7198 vss 0.0424f
C7696 vdd.n7199 vss 0.02f
C7697 vdd.n7200 vss 0.00425f
C7698 vdd.n7201 vss 0.0471f
C7699 vdd.n7203 vss 0.00425f
C7700 vdd.n7204 vss 0.00925f
C7701 vdd.n7205 vss 0.00679f
C7702 vdd.n7206 vss 0.00517f
C7703 vdd.n7207 vss 0.00251f
C7704 vdd.n7208 vss 0.0471f
C7705 vdd.n7209 vss 0.00251f
C7706 vdd.n7210 vss 0.0112f
C7707 vdd.n7211 vss 0.0128f
C7708 vdd.n7212 vss 0.0619f
C7709 vdd.n7213 vss 0.00324f
C7710 vdd.n7214 vss 0.0112f
C7711 vdd.n7215 vss 0.0128f
C7712 vdd.n7216 vss 0.00413f
C7713 vdd.n7217 vss 0.00413f
C7714 vdd.n7218 vss 0.0471f
C7715 vdd.n7219 vss 0.0471f
C7716 vdd.n7220 vss 0.00324f
C7717 vdd.n7221 vss 0.00413f
C7718 vdd.n7222 vss 0.00413f
C7719 vdd.n7223 vss 0.00679f
C7720 vdd.n7224 vss 0.00413f
C7721 vdd.n7225 vss 0.0471f
C7722 vdd.n7226 vss 0.00324f
C7723 vdd.n7228 vss 0.00925f
C7724 vdd.n7229 vss 0.0471f
C7725 vdd.n7230 vss 0.00425f
C7726 vdd.n7231 vss 0.0424f
C7727 vdd.n7232 vss 0.0132f
C7728 vdd.n7233 vss 0.00324f
C7729 vdd.n7234 vss 0.0128f
C7730 vdd.n7235 vss 0.02f
C7731 vdd.n7236 vss 0.00425f
C7732 vdd.n7237 vss 0.00413f
C7733 vdd.n7238 vss 0.00251f
C7734 vdd.n7239 vss 0.0471f
C7735 vdd.n7240 vss 0.00251f
C7736 vdd.n7241 vss 0.00517f
C7737 vdd.n7242 vss 0.00679f
C7738 vdd.n7243 vss 0.00324f
C7739 vdd.n7244 vss 0.00324f
C7740 vdd.n7245 vss 0.0132f
C7741 vdd.n7246 vss 0.0424f
C7742 vdd.n7247 vss 0.02f
C7743 vdd.n7248 vss 0.00425f
C7744 vdd.n7249 vss 0.0471f
C7745 vdd.n7251 vss 0.00425f
C7746 vdd.n7252 vss 0.00925f
C7747 vdd.n7253 vss 0.00679f
C7748 vdd.n7254 vss 0.00517f
C7749 vdd.n7255 vss 0.00251f
C7750 vdd.n7256 vss 0.0471f
C7751 vdd.n7257 vss 0.00251f
C7752 vdd.n7258 vss 0.0112f
C7753 vdd.n7259 vss 0.0128f
C7754 vdd.n7260 vss 0.0692f
C7755 vdd.n7261 vss 0.00324f
C7756 vdd.n7262 vss 0.0112f
C7757 vdd.n7263 vss 0.0128f
C7758 vdd.n7264 vss 0.00413f
C7759 vdd.n7265 vss 0.00413f
C7760 vdd.n7266 vss 0.0471f
C7761 vdd.n7267 vss 0.0471f
C7762 vdd.n7268 vss 0.00324f
C7763 vdd.n7269 vss 0.00413f
C7764 vdd.n7270 vss 0.00413f
C7765 vdd.n7271 vss 0.00679f
C7766 vdd.n7272 vss 0.00413f
C7767 vdd.n7273 vss 0.0471f
C7768 vdd.n7274 vss 0.00324f
C7769 vdd.n7276 vss 0.00925f
C7770 vdd.n7277 vss 0.0471f
C7771 vdd.n7278 vss 0.00425f
C7772 vdd.n7279 vss 0.0424f
C7773 vdd.n7280 vss 0.0132f
C7774 vdd.n7281 vss 0.00324f
C7775 vdd.n7282 vss 0.0128f
C7776 vdd.n7283 vss 0.02f
C7777 vdd.n7284 vss 0.00425f
C7778 vdd.n7285 vss 0.00413f
C7779 vdd.n7286 vss 0.00251f
C7780 vdd.n7287 vss 0.0471f
C7781 vdd.n7288 vss 0.00251f
C7782 vdd.n7289 vss 0.00517f
C7783 vdd.n7290 vss 0.00679f
C7784 vdd.n7291 vss 0.00324f
C7785 vdd.n7292 vss 0.00324f
C7786 vdd.n7293 vss 0.0132f
C7787 vdd.n7294 vss 0.0424f
C7788 vdd.n7295 vss 0.02f
C7789 vdd.n7296 vss 0.00425f
C7790 vdd.n7297 vss 0.0471f
C7791 vdd.n7299 vss 0.00425f
C7792 vdd.n7300 vss 0.00925f
C7793 vdd.n7301 vss 0.00679f
C7794 vdd.n7302 vss 0.00517f
C7795 vdd.n7303 vss 0.00251f
C7796 vdd.n7304 vss 0.0471f
C7797 vdd.n7305 vss 0.00251f
C7798 vdd.n7306 vss 0.0112f
C7799 vdd.n7307 vss 0.0128f
C7800 vdd.n7308 vss 0.0619f
C7801 vdd.n7309 vss 0.00335f
C7802 vdd.n7310 vss 0.0855f
C7803 vdd.n7311 vss 0.00991f
C7804 vdd.n7312 vss 0.0424f
C7805 vdd.n7313 vss 0.00679f
C7806 vdd.n7314 vss 0.00413f
C7807 vdd.n7315 vss 0.0471f
C7808 vdd.n7316 vss 0.00251f
C7809 vdd.n7317 vss 0.00679f
C7810 vdd.n7318 vss 0.00413f
C7811 vdd.n7319 vss 0.00413f
C7812 vdd.n7320 vss 0.0471f
C7813 vdd.n7321 vss 0.00251f
C7814 vdd.n7322 vss 0.00413f
C7815 vdd.n7323 vss 0.00324f
C7816 vdd.n7324 vss 0.0132f
C7817 vdd.n7325 vss 0.0424f
C7818 vdd.n7326 vss 0.00324f
C7819 vdd.n7327 vss 0.00413f
C7820 vdd.n7328 vss 0.00517f
C7821 vdd.n7329 vss 0.00679f
C7822 vdd.n7330 vss 0.00925f
C7823 vdd.n7331 vss 0.00425f
C7824 vdd.n7332 vss 0.0471f
C7825 vdd.n7334 vss 0.00425f
C7826 vdd.n7335 vss 0.02f
C7827 vdd.n7336 vss 0.0128f
C7828 vdd.n7337 vss 0.0105f
C7829 vdd.n7338 vss 0.00251f
C7830 vdd.n7339 vss 0.0471f
C7831 vdd.n7340 vss 0.00517f
C7832 vdd.n7341 vss 0.00251f
C7833 vdd.n7342 vss 0.0471f
C7834 vdd.n7343 vss 0.0471f
C7835 vdd.n7344 vss 0.00324f
C7836 vdd.n7345 vss 0.00324f
C7837 vdd.n7346 vss 0.00805f
C7838 vdd.n7347 vss 0.0112f
C7839 vdd.n7348 vss 0.0128f
C7840 vdd.n7349 vss 0.00324f
C7841 vdd.n7350 vss 0.00324f
C7842 vdd.n7351 vss 0.00413f
C7843 vdd.n7352 vss 0.00425f
C7844 vdd.n7353 vss 0.0471f
C7845 vdd.n7355 vss 0.00425f
C7846 vdd.n7356 vss 0.00925f
C7847 vdd.n7357 vss 0.0107f
C7848 vdd.n7358 vss 0.0126f
C7849 vdd.n7359 vss 0.0516f
C7850 vdd.n7360 vss 0.00163f
C7851 vdd.n7361 vss 0.00145f
C7852 vdd.n7362 vss 0.0271f
C7853 vdd.n7363 vss 0.00324f
C7854 vdd.n7364 vss 0.0112f
C7855 vdd.n7365 vss 0.0128f
C7856 vdd.n7366 vss 0.00413f
C7857 vdd.n7367 vss 0.00413f
C7858 vdd.n7368 vss 0.0471f
C7859 vdd.n7369 vss 0.0471f
C7860 vdd.n7370 vss 0.00324f
C7861 vdd.n7371 vss 0.00413f
C7862 vdd.n7372 vss 0.00413f
C7863 vdd.n7373 vss 0.00679f
C7864 vdd.n7374 vss 0.00413f
C7865 vdd.n7375 vss 0.0471f
C7866 vdd.n7376 vss 0.00324f
C7867 vdd.n7378 vss 0.00925f
C7868 vdd.n7379 vss 0.0471f
C7869 vdd.n7380 vss 0.00425f
C7870 vdd.n7381 vss 0.0424f
C7871 vdd.n7382 vss 0.0132f
C7872 vdd.n7383 vss 0.00324f
C7873 vdd.n7384 vss 0.0128f
C7874 vdd.n7385 vss 0.02f
C7875 vdd.n7386 vss 0.00425f
C7876 vdd.n7387 vss 0.00413f
C7877 vdd.n7388 vss 0.00251f
C7878 vdd.n7389 vss 0.0471f
C7879 vdd.n7390 vss 0.00251f
C7880 vdd.n7391 vss 0.00517f
C7881 vdd.n7392 vss 0.00679f
C7882 vdd.n7393 vss 0.00324f
C7883 vdd.n7394 vss 0.00324f
C7884 vdd.n7395 vss 0.0132f
C7885 vdd.n7396 vss 0.0424f
C7886 vdd.n7397 vss 0.02f
C7887 vdd.n7398 vss 0.00425f
C7888 vdd.n7399 vss 0.0471f
C7889 vdd.n7401 vss 0.00425f
C7890 vdd.n7402 vss 0.00925f
C7891 vdd.n7403 vss 0.00679f
C7892 vdd.n7404 vss 0.00517f
C7893 vdd.n7405 vss 0.00251f
C7894 vdd.n7406 vss 0.0471f
C7895 vdd.n7407 vss 0.00251f
C7896 vdd.n7408 vss 0.0112f
C7897 vdd.n7409 vss 0.0128f
C7898 vdd.n7410 vss 0.0692f
C7899 vdd.n7411 vss 0.00324f
C7900 vdd.n7412 vss 0.0112f
C7901 vdd.n7413 vss 0.0128f
C7902 vdd.n7414 vss 0.00413f
C7903 vdd.n7415 vss 0.00413f
C7904 vdd.n7416 vss 0.0471f
C7905 vdd.n7417 vss 0.0471f
C7906 vdd.n7418 vss 0.00324f
C7907 vdd.n7419 vss 0.00413f
C7908 vdd.n7420 vss 0.00413f
C7909 vdd.n7421 vss 0.00679f
C7910 vdd.n7422 vss 0.00413f
C7911 vdd.n7423 vss 0.0471f
C7912 vdd.n7424 vss 0.00324f
C7913 vdd.n7425 vss 0.0424f
C7914 vdd.n7426 vss 0.00324f
C7915 vdd.n7427 vss 0.0128f
C7916 vdd.n7428 vss 0.02f
C7917 vdd.n7429 vss 0.0132f
C7918 vdd.n7430 vss 0.00925f
C7919 vdd.n7431 vss 0.00425f
C7920 vdd.n7433 vss 0.0471f
C7921 vdd.n7434 vss 0.00425f
C7922 vdd.n7435 vss 0.00413f
C7923 vdd.n7436 vss 0.00251f
C7924 vdd.n7437 vss 0.0471f
C7925 vdd.n7438 vss 0.00251f
C7926 vdd.n7439 vss 0.00517f
C7927 vdd.n7440 vss 0.00679f
C7928 vdd.n7441 vss 0.00324f
C7929 vdd.n7442 vss 0.00324f
C7930 vdd.n7443 vss 0.0132f
C7931 vdd.n7444 vss 0.0424f
C7932 vdd.n7445 vss 0.02f
C7933 vdd.n7446 vss 0.00425f
C7934 vdd.n7448 vss 0.0471f
C7935 vdd.n7449 vss 0.00425f
C7936 vdd.n7450 vss 0.00925f
C7937 vdd.n7451 vss 0.00679f
C7938 vdd.n7452 vss 0.00517f
C7939 vdd.n7453 vss 0.00251f
C7940 vdd.n7454 vss 0.0471f
C7941 vdd.n7455 vss 0.00251f
C7942 vdd.n7456 vss 0.0112f
C7943 vdd.n7457 vss 0.0128f
C7944 vdd.n7458 vss 0.0666f
C7945 vdd.n7459 vss 0.00324f
C7946 vdd.n7460 vss 0.0112f
C7947 vdd.n7461 vss 0.0128f
C7948 vdd.n7462 vss 0.00413f
C7949 vdd.n7463 vss 0.00413f
C7950 vdd.n7464 vss 0.0471f
C7951 vdd.n7465 vss 0.0471f
C7952 vdd.n7466 vss 0.00324f
C7953 vdd.n7467 vss 0.00413f
C7954 vdd.n7468 vss 0.00413f
C7955 vdd.n7469 vss 0.00679f
C7956 vdd.n7470 vss 0.00413f
C7957 vdd.n7471 vss 0.0471f
C7958 vdd.n7472 vss 0.00324f
C7959 vdd.n7473 vss 0.0424f
C7960 vdd.n7474 vss 0.00324f
C7961 vdd.n7475 vss 0.0128f
C7962 vdd.n7476 vss 0.02f
C7963 vdd.n7477 vss 0.0132f
C7964 vdd.n7478 vss 0.00925f
C7965 vdd.n7479 vss 0.00425f
C7966 vdd.n7481 vss 0.0471f
C7967 vdd.n7482 vss 0.00425f
C7968 vdd.n7483 vss 0.00413f
C7969 vdd.n7484 vss 0.00251f
C7970 vdd.n7485 vss 0.0471f
C7971 vdd.n7486 vss 0.00251f
C7972 vdd.n7487 vss 0.00517f
C7973 vdd.n7488 vss 0.00679f
C7974 vdd.n7489 vss 0.00324f
C7975 vdd.n7490 vss 0.00324f
C7976 vdd.n7491 vss 0.0132f
C7977 vdd.n7492 vss 0.0424f
C7978 vdd.n7493 vss 0.02f
C7979 vdd.n7494 vss 0.00425f
C7980 vdd.n7496 vss 0.0471f
C7981 vdd.n7497 vss 0.00425f
C7982 vdd.n7498 vss 0.00925f
C7983 vdd.n7499 vss 0.00679f
C7984 vdd.n7500 vss 0.00517f
C7985 vdd.n7501 vss 0.00251f
C7986 vdd.n7502 vss 0.0471f
C7987 vdd.n7503 vss 0.00251f
C7988 vdd.n7504 vss 0.0112f
C7989 vdd.n7505 vss 0.0128f
C7990 vdd.n7506 vss 0.0617f
C7991 vdd.n7507 vss 0.00335f
C7992 vdd.n7508 vss 0.0855f
C7993 vdd.n7509 vss 0.0107f
C7994 vdd.n7510 vss 0.0128f
C7995 vdd.n7511 vss 0.0424f
C7996 vdd.n7512 vss 0.00413f
C7997 vdd.n7513 vss 0.0471f
C7998 vdd.n7514 vss 0.00413f
C7999 vdd.n7515 vss 0.00324f
C8000 vdd.n7516 vss 0.00324f
C8001 vdd.n7517 vss 0.00679f
C8002 vdd.n7518 vss 0.00413f
C8003 vdd.n7519 vss 0.0471f
C8004 vdd.n7520 vss 0.00413f
C8005 vdd.n7521 vss 0.0105f
C8006 vdd.n7522 vss 0.0471f
C8007 vdd.n7523 vss 0.00413f
C8008 vdd.n7524 vss 0.00324f
C8009 vdd.n7525 vss 0.00324f
C8010 vdd.n7526 vss 0.0132f
C8011 vdd.n7527 vss 0.0424f
C8012 vdd.n7528 vss 0.0128f
C8013 vdd.n7529 vss 0.02f
C8014 vdd.n7530 vss 0.00425f
C8015 vdd.n7532 vss 0.0471f
C8016 vdd.n7533 vss 0.00425f
C8017 vdd.n7534 vss 0.00925f
C8018 vdd.n7535 vss 0.00679f
C8019 vdd.n7536 vss 0.00517f
C8020 vdd.n7537 vss 0.00251f
C8021 vdd.n7538 vss 0.0471f
C8022 vdd.n7539 vss 0.00251f
C8023 vdd.n7540 vss 0.00413f
C8024 vdd.n7541 vss 0.00324f
C8025 vdd.n7542 vss 0.00324f
C8026 vdd.n7543 vss 0.00805f
C8027 vdd.n7544 vss 0.0112f
C8028 vdd.n7545 vss 0.00251f
C8029 vdd.n7546 vss 0.0471f
C8030 vdd.n7547 vss 0.00251f
C8031 vdd.n7548 vss 0.00517f
C8032 vdd.n7549 vss 0.00679f
C8033 vdd.n7550 vss 0.00925f
C8034 vdd.n7551 vss 0.00425f
C8035 vdd.n7553 vss 0.0471f
C8036 vdd.n7554 vss 0.00425f
C8037 vdd.n7555 vss 0.00991f
C8038 vdd.n7556 vss 0.0126f
C8039 vdd.n7557 vss 0.0516f
C8040 vdd.n7558 vss 0.0011f
C8041 vdd.n7559 vss 0.0271f
C8042 vdd.n7560 vss 0.00324f
C8043 vdd.n7561 vss 0.0112f
C8044 vdd.n7562 vss 0.0128f
C8045 vdd.n7563 vss 0.00413f
C8046 vdd.n7564 vss 0.00413f
C8047 vdd.n7565 vss 0.0471f
C8048 vdd.n7566 vss 0.0471f
C8049 vdd.n7567 vss 0.00324f
C8050 vdd.n7568 vss 0.00413f
C8051 vdd.n7569 vss 0.00413f
C8052 vdd.n7570 vss 0.00679f
C8053 vdd.n7571 vss 0.00413f
C8054 vdd.n7572 vss 0.0471f
C8055 vdd.n7573 vss 0.00324f
C8056 vdd.n7574 vss 0.0424f
C8057 vdd.n7575 vss 0.00324f
C8058 vdd.n7576 vss 0.0128f
C8059 vdd.n7577 vss 0.02f
C8060 vdd.n7578 vss 0.0132f
C8061 vdd.n7579 vss 0.00925f
C8062 vdd.n7580 vss 0.00425f
C8063 vdd.n7582 vss 0.0471f
C8064 vdd.n7583 vss 0.00425f
C8065 vdd.n7584 vss 0.00413f
C8066 vdd.n7585 vss 0.00251f
C8067 vdd.n7586 vss 0.0471f
C8068 vdd.n7587 vss 0.00251f
C8069 vdd.n7588 vss 0.00517f
C8070 vdd.n7589 vss 0.00679f
C8071 vdd.n7590 vss 0.00324f
C8072 vdd.n7591 vss 0.00324f
C8073 vdd.n7592 vss 0.0132f
C8074 vdd.n7593 vss 0.0424f
C8075 vdd.n7594 vss 0.02f
C8076 vdd.n7595 vss 0.00425f
C8077 vdd.n7597 vss 0.0471f
C8078 vdd.n7598 vss 0.00425f
C8079 vdd.n7599 vss 0.00925f
C8080 vdd.n7600 vss 0.00679f
C8081 vdd.n7601 vss 0.00517f
C8082 vdd.n7602 vss 0.00251f
C8083 vdd.n7603 vss 0.0471f
C8084 vdd.n7604 vss 0.00251f
C8085 vdd.n7605 vss 0.0112f
C8086 vdd.n7606 vss 0.0128f
C8087 vdd.n7607 vss 0.0666f
C8088 vdd.n7608 vss 0.00324f
C8089 vdd.n7609 vss 0.0112f
C8090 vdd.n7610 vss 0.0128f
C8091 vdd.n7611 vss 0.00413f
C8092 vdd.n7612 vss 0.00413f
C8093 vdd.n7613 vss 0.0471f
C8094 vdd.n7614 vss 0.0471f
C8095 vdd.n7615 vss 0.00324f
C8096 vdd.n7616 vss 0.00413f
C8097 vdd.n7617 vss 0.00413f
C8098 vdd.n7618 vss 0.00679f
C8099 vdd.n7619 vss 0.00413f
C8100 vdd.n7620 vss 0.0471f
C8101 vdd.n7621 vss 0.00324f
C8102 vdd.n7622 vss 0.0424f
C8103 vdd.n7623 vss 0.00324f
C8104 vdd.n7624 vss 0.0128f
C8105 vdd.n7625 vss 0.02f
C8106 vdd.n7626 vss 0.0132f
C8107 vdd.n7627 vss 0.00925f
C8108 vdd.n7628 vss 0.00425f
C8109 vdd.n7630 vss 0.0471f
C8110 vdd.n7631 vss 0.00425f
C8111 vdd.n7632 vss 0.00413f
C8112 vdd.n7633 vss 0.00251f
C8113 vdd.n7634 vss 0.0471f
C8114 vdd.n7635 vss 0.00251f
C8115 vdd.n7636 vss 0.00517f
C8116 vdd.n7637 vss 0.00679f
C8117 vdd.n7638 vss 0.00324f
C8118 vdd.n7639 vss 0.00324f
C8119 vdd.n7640 vss 0.0132f
C8120 vdd.n7641 vss 0.0424f
C8121 vdd.n7642 vss 0.02f
C8122 vdd.n7643 vss 0.00425f
C8123 vdd.n7645 vss 0.0471f
C8124 vdd.n7646 vss 0.00425f
C8125 vdd.n7647 vss 0.00925f
C8126 vdd.n7648 vss 0.00679f
C8127 vdd.n7649 vss 0.00517f
C8128 vdd.n7650 vss 0.00251f
C8129 vdd.n7651 vss 0.0471f
C8130 vdd.n7652 vss 0.00251f
C8131 vdd.n7653 vss 0.0112f
C8132 vdd.n7654 vss 0.0128f
C8133 vdd.n7655 vss 0.0613f
C8134 vdd.n7656 vss 0.00324f
C8135 vdd.n7657 vss 0.0112f
C8136 vdd.n7658 vss 0.0128f
C8137 vdd.n7659 vss 0.00413f
C8138 vdd.n7660 vss 0.00413f
C8139 vdd.n7661 vss 0.0471f
C8140 vdd.n7662 vss 0.0471f
C8141 vdd.n7663 vss 0.00324f
C8142 vdd.n7664 vss 0.00413f
C8143 vdd.n7665 vss 0.00413f
C8144 vdd.n7666 vss 0.00679f
C8145 vdd.n7667 vss 0.00413f
C8146 vdd.n7668 vss 0.0471f
C8147 vdd.n7669 vss 0.00324f
C8148 vdd.n7670 vss 0.0424f
C8149 vdd.n7671 vss 0.00324f
C8150 vdd.n7672 vss 0.0128f
C8151 vdd.n7673 vss 0.02f
C8152 vdd.n7674 vss 0.0132f
C8153 vdd.n7675 vss 0.00925f
C8154 vdd.n7676 vss 0.00425f
C8155 vdd.n7678 vss 0.0471f
C8156 vdd.n7679 vss 0.00425f
C8157 vdd.n7680 vss 0.00413f
C8158 vdd.n7681 vss 0.00251f
C8159 vdd.n7682 vss 0.0471f
C8160 vdd.n7683 vss 0.00251f
C8161 vdd.n7684 vss 0.00517f
C8162 vdd.n7685 vss 0.00679f
C8163 vdd.n7686 vss 0.00324f
C8164 vdd.n7687 vss 0.00324f
C8165 vdd.n7688 vss 0.0132f
C8166 vdd.n7689 vss 0.0424f
C8167 vdd.n7690 vss 0.02f
C8168 vdd.n7691 vss 0.00425f
C8169 vdd.n7693 vss 0.0471f
C8170 vdd.n7694 vss 0.00425f
C8171 vdd.n7695 vss 0.00925f
C8172 vdd.n7696 vss 0.00679f
C8173 vdd.n7697 vss 0.00517f
C8174 vdd.n7698 vss 0.00251f
C8175 vdd.n7699 vss 0.0471f
C8176 vdd.n7700 vss 0.00251f
C8177 vdd.n7701 vss 0.0112f
C8178 vdd.n7702 vss 0.0128f
C8179 vdd.n7703 vss 0.0666f
C8180 vdd.n7704 vss 0.00324f
C8181 vdd.n7705 vss 0.0112f
C8182 vdd.n7706 vss 0.0128f
C8183 vdd.n7707 vss 0.00413f
C8184 vdd.n7708 vss 0.00413f
C8185 vdd.n7709 vss 0.0471f
C8186 vdd.n7710 vss 0.0471f
C8187 vdd.n7711 vss 0.00324f
C8188 vdd.n7712 vss 0.00413f
C8189 vdd.n7713 vss 0.00413f
C8190 vdd.n7714 vss 0.00679f
C8191 vdd.n7715 vss 0.00413f
C8192 vdd.n7716 vss 0.0471f
C8193 vdd.n7717 vss 0.00324f
C8194 vdd.n7718 vss 0.0424f
C8195 vdd.n7719 vss 0.00324f
C8196 vdd.n7720 vss 0.0128f
C8197 vdd.n7721 vss 0.02f
C8198 vdd.n7722 vss 0.0132f
C8199 vdd.n7723 vss 0.00925f
C8200 vdd.n7724 vss 0.00425f
C8201 vdd.n7726 vss 0.0471f
C8202 vdd.n7727 vss 0.00425f
C8203 vdd.n7728 vss 0.00413f
C8204 vdd.n7729 vss 0.00251f
C8205 vdd.n7730 vss 0.0471f
C8206 vdd.n7731 vss 0.00251f
C8207 vdd.n7732 vss 0.00517f
C8208 vdd.n7733 vss 0.00679f
C8209 vdd.n7734 vss 0.00324f
C8210 vdd.n7735 vss 0.00324f
C8211 vdd.n7736 vss 0.0132f
C8212 vdd.n7737 vss 0.0424f
C8213 vdd.n7738 vss 0.02f
C8214 vdd.n7739 vss 0.00425f
C8215 vdd.n7741 vss 0.0471f
C8216 vdd.n7742 vss 0.00425f
C8217 vdd.n7743 vss 0.00925f
C8218 vdd.n7744 vss 0.00679f
C8219 vdd.n7745 vss 0.00517f
C8220 vdd.n7746 vss 0.00251f
C8221 vdd.n7747 vss 0.0471f
C8222 vdd.n7748 vss 0.00251f
C8223 vdd.n7749 vss 0.0112f
C8224 vdd.n7750 vss 0.0128f
C8225 vdd.n7751 vss 0.0617f
C8226 vdd.n7752 vss 0.00335f
C8227 vdd.n7753 vss 0.0855f
C8228 vdd.n7754 vss 0.0107f
C8229 vdd.n7755 vss 0.0128f
C8230 vdd.n7756 vss 0.0424f
C8231 vdd.n7757 vss 0.00413f
C8232 vdd.n7758 vss 0.0471f
C8233 vdd.n7759 vss 0.00413f
C8234 vdd.n7760 vss 0.00324f
C8235 vdd.n7761 vss 0.00324f
C8236 vdd.n7762 vss 0.00679f
C8237 vdd.n7763 vss 0.00413f
C8238 vdd.n7764 vss 0.0471f
C8239 vdd.n7765 vss 0.00413f
C8240 vdd.n7766 vss 0.0105f
C8241 vdd.n7767 vss 0.0471f
C8242 vdd.n7768 vss 0.00413f
C8243 vdd.n7769 vss 0.00324f
C8244 vdd.n7770 vss 0.00324f
C8245 vdd.n7771 vss 0.0132f
C8246 vdd.n7772 vss 0.0424f
C8247 vdd.n7773 vss 0.0128f
C8248 vdd.n7774 vss 0.02f
C8249 vdd.n7775 vss 0.00425f
C8250 vdd.n7777 vss 0.0471f
C8251 vdd.n7778 vss 0.00425f
C8252 vdd.n7779 vss 0.00925f
C8253 vdd.n7780 vss 0.00679f
C8254 vdd.n7781 vss 0.00517f
C8255 vdd.n7782 vss 0.00251f
C8256 vdd.n7783 vss 0.0471f
C8257 vdd.n7784 vss 0.00251f
C8258 vdd.n7785 vss 0.00413f
C8259 vdd.n7786 vss 0.00324f
C8260 vdd.n7787 vss 0.00324f
C8261 vdd.n7788 vss 0.00805f
C8262 vdd.n7789 vss 0.0112f
C8263 vdd.n7790 vss 0.00251f
C8264 vdd.n7791 vss 0.0471f
C8265 vdd.n7792 vss 0.00251f
C8266 vdd.n7793 vss 0.00517f
C8267 vdd.n7794 vss 0.00679f
C8268 vdd.n7795 vss 0.00925f
C8269 vdd.n7796 vss 0.00425f
C8270 vdd.n7798 vss 0.0471f
C8271 vdd.n7799 vss 0.00425f
C8272 vdd.n7800 vss 0.00991f
C8273 vdd.n7801 vss 0.0126f
C8274 vdd.n7802 vss 0.0516f
C8275 vdd.n7803 vss 0.0011f
C8276 vdd.n7804 vss 0.0271f
C8277 vdd.n7805 vss 0.00324f
C8278 vdd.n7806 vss 0.0112f
C8279 vdd.n7807 vss 0.0128f
C8280 vdd.n7808 vss 0.00413f
C8281 vdd.n7809 vss 0.00413f
C8282 vdd.n7810 vss 0.0471f
C8283 vdd.n7811 vss 0.0471f
C8284 vdd.n7812 vss 0.00324f
C8285 vdd.n7813 vss 0.00413f
C8286 vdd.n7814 vss 0.00413f
C8287 vdd.n7815 vss 0.00679f
C8288 vdd.n7816 vss 0.00413f
C8289 vdd.n7817 vss 0.0471f
C8290 vdd.n7818 vss 0.00324f
C8291 vdd.n7819 vss 0.0424f
C8292 vdd.n7820 vss 0.00324f
C8293 vdd.n7821 vss 0.0128f
C8294 vdd.n7822 vss 0.02f
C8295 vdd.n7823 vss 0.0132f
C8296 vdd.n7824 vss 0.00925f
C8297 vdd.n7825 vss 0.00425f
C8298 vdd.n7827 vss 0.0471f
C8299 vdd.n7828 vss 0.00425f
C8300 vdd.n7829 vss 0.00413f
C8301 vdd.n7830 vss 0.00251f
C8302 vdd.n7831 vss 0.0471f
C8303 vdd.n7832 vss 0.00251f
C8304 vdd.n7833 vss 0.00517f
C8305 vdd.n7834 vss 0.00679f
C8306 vdd.n7835 vss 0.00324f
C8307 vdd.n7836 vss 0.00324f
C8308 vdd.n7837 vss 0.0132f
C8309 vdd.n7838 vss 0.0424f
C8310 vdd.n7839 vss 0.02f
C8311 vdd.n7840 vss 0.00425f
C8312 vdd.n7842 vss 0.0471f
C8313 vdd.n7843 vss 0.00425f
C8314 vdd.n7844 vss 0.00925f
C8315 vdd.n7845 vss 0.00679f
C8316 vdd.n7846 vss 0.00517f
C8317 vdd.n7847 vss 0.00251f
C8318 vdd.n7848 vss 0.0471f
C8319 vdd.n7849 vss 0.00251f
C8320 vdd.n7850 vss 0.0112f
C8321 vdd.n7851 vss 0.0128f
C8322 vdd.n7852 vss 0.0666f
C8323 vdd.n7853 vss 0.00324f
C8324 vdd.n7854 vss 0.0112f
C8325 vdd.n7855 vss 0.0128f
C8326 vdd.n7856 vss 0.00413f
C8327 vdd.n7857 vss 0.00413f
C8328 vdd.n7858 vss 0.0471f
C8329 vdd.n7859 vss 0.0471f
C8330 vdd.n7860 vss 0.00324f
C8331 vdd.n7861 vss 0.00413f
C8332 vdd.n7862 vss 0.00413f
C8333 vdd.n7863 vss 0.00679f
C8334 vdd.n7864 vss 0.00413f
C8335 vdd.n7865 vss 0.0471f
C8336 vdd.n7866 vss 0.00324f
C8337 vdd.n7867 vss 0.0424f
C8338 vdd.n7868 vss 0.00324f
C8339 vdd.n7869 vss 0.0128f
C8340 vdd.n7870 vss 0.02f
C8341 vdd.n7871 vss 0.0132f
C8342 vdd.n7872 vss 0.00925f
C8343 vdd.n7873 vss 0.00425f
C8344 vdd.n7875 vss 0.0471f
C8345 vdd.n7876 vss 0.00425f
C8346 vdd.n7877 vss 0.00413f
C8347 vdd.n7878 vss 0.00251f
C8348 vdd.n7879 vss 0.0471f
C8349 vdd.n7880 vss 0.00251f
C8350 vdd.n7881 vss 0.00517f
C8351 vdd.n7882 vss 0.00679f
C8352 vdd.n7883 vss 0.00324f
C8353 vdd.n7884 vss 0.00324f
C8354 vdd.n7885 vss 0.0132f
C8355 vdd.n7886 vss 0.0424f
C8356 vdd.n7887 vss 0.02f
C8357 vdd.n7888 vss 0.00425f
C8358 vdd.n7890 vss 0.0471f
C8359 vdd.n7891 vss 0.00425f
C8360 vdd.n7892 vss 0.00925f
C8361 vdd.n7893 vss 0.00679f
C8362 vdd.n7894 vss 0.00517f
C8363 vdd.n7895 vss 0.00251f
C8364 vdd.n7896 vss 0.0471f
C8365 vdd.n7897 vss 0.00251f
C8366 vdd.n7898 vss 0.0112f
C8367 vdd.n7899 vss 0.0128f
C8368 vdd.n7900 vss 0.00324f
C8369 vdd.n7901 vss 0.0112f
C8370 vdd.n7902 vss 0.0128f
C8371 vdd.n7903 vss 0.00413f
C8372 vdd.n7904 vss 0.00413f
C8373 vdd.n7905 vss 0.0471f
C8374 vdd.n7906 vss 0.0471f
C8375 vdd.n7907 vss 0.00324f
C8376 vdd.n7908 vss 0.00413f
C8377 vdd.n7909 vss 0.00413f
C8378 vdd.n7910 vss 0.00679f
C8379 vdd.n7911 vss 0.00413f
C8380 vdd.n7912 vss 0.0471f
C8381 vdd.n7913 vss 0.00324f
C8382 vdd.n7914 vss 0.0424f
C8383 vdd.n7915 vss 0.00324f
C8384 vdd.n7916 vss 0.0128f
C8385 vdd.n7917 vss 0.02f
C8386 vdd.n7918 vss 0.0132f
C8387 vdd.n7919 vss 0.00925f
C8388 vdd.n7920 vss 0.00425f
C8389 vdd.n7922 vss 0.0471f
C8390 vdd.n7923 vss 0.00425f
C8391 vdd.n7924 vss 0.00413f
C8392 vdd.n7925 vss 0.00251f
C8393 vdd.n7926 vss 0.0471f
C8394 vdd.n7927 vss 0.00251f
C8395 vdd.n7928 vss 0.00517f
C8396 vdd.n7929 vss 0.00679f
C8397 vdd.n7930 vss 0.00324f
C8398 vdd.n7931 vss 0.00324f
C8399 vdd.n7932 vss 0.0132f
C8400 vdd.n7933 vss 0.0424f
C8401 vdd.n7934 vss 0.02f
C8402 vdd.n7935 vss 0.00425f
C8403 vdd.n7937 vss 0.0471f
C8404 vdd.n7938 vss 0.00425f
C8405 vdd.n7939 vss 0.00925f
C8406 vdd.n7940 vss 0.00679f
C8407 vdd.n7941 vss 0.00517f
C8408 vdd.n7942 vss 0.00251f
C8409 vdd.n7943 vss 0.0471f
C8410 vdd.n7944 vss 0.00251f
C8411 vdd.n7945 vss 0.0112f
C8412 vdd.n7946 vss 0.0128f
C8413 vdd.n7947 vss 0.144f
C8414 vdd.n7948 vss 0.143f
C8415 vdd.n7949 vss 0.0608f
C8416 vdd.n7950 vss 0.00324f
C8417 vdd.n7951 vss 0.0112f
C8418 vdd.n7952 vss 0.0128f
C8419 vdd.n7953 vss 0.00413f
C8420 vdd.n7954 vss 0.00413f
C8421 vdd.n7955 vss 0.0471f
C8422 vdd.n7956 vss 0.0471f
C8423 vdd.n7957 vss 0.00324f
C8424 vdd.n7958 vss 0.00413f
C8425 vdd.n7959 vss 0.00413f
C8426 vdd.n7960 vss 0.00679f
C8427 vdd.n7961 vss 0.00413f
C8428 vdd.n7962 vss 0.0471f
C8429 vdd.n7963 vss 0.00324f
C8430 vdd.n7964 vss 0.0424f
C8431 vdd.n7965 vss 0.00324f
C8432 vdd.n7966 vss 0.0128f
C8433 vdd.n7967 vss 0.02f
C8434 vdd.n7968 vss 0.0132f
C8435 vdd.n7969 vss 0.00925f
C8436 vdd.n7970 vss 0.00425f
C8437 vdd.n7972 vss 0.0471f
C8438 vdd.n7973 vss 0.00425f
C8439 vdd.n7974 vss 0.00413f
C8440 vdd.n7975 vss 0.00251f
C8441 vdd.n7976 vss 0.0471f
C8442 vdd.n7977 vss 0.00251f
C8443 vdd.n7978 vss 0.00517f
C8444 vdd.n7979 vss 0.00679f
C8445 vdd.n7980 vss 0.00324f
C8446 vdd.n7981 vss 0.00324f
C8447 vdd.n7982 vss 0.0132f
C8448 vdd.n7983 vss 0.0424f
C8449 vdd.n7984 vss 0.02f
C8450 vdd.n7985 vss 0.00425f
C8451 vdd.n7987 vss 0.0471f
C8452 vdd.n7988 vss 0.00425f
C8453 vdd.n7989 vss 0.00925f
C8454 vdd.n7990 vss 0.00679f
C8455 vdd.n7991 vss 0.00517f
C8456 vdd.n7992 vss 0.00251f
C8457 vdd.n7993 vss 0.0471f
C8458 vdd.n7994 vss 0.00251f
C8459 vdd.n7995 vss 0.0112f
C8460 vdd.n7996 vss 0.0128f
C8461 vdd.n7997 vss 0.0666f
C8462 vdd.n7998 vss 0.118f
C8463 vdd.n7999 vss 0.121f
C8464 vdd.n8000 vss 0.00324f
C8465 vdd.n8001 vss 0.0112f
C8466 vdd.n8002 vss 0.0128f
C8467 vdd.n8003 vss 0.00413f
C8468 vdd.n8004 vss 0.00413f
C8469 vdd.n8005 vss 0.0471f
C8470 vdd.n8006 vss 0.0471f
C8471 vdd.n8007 vss 0.00324f
C8472 vdd.n8008 vss 0.00413f
C8473 vdd.n8009 vss 0.00413f
C8474 vdd.n8010 vss 0.00679f
C8475 vdd.n8011 vss 0.00413f
C8476 vdd.n8012 vss 0.0471f
C8477 vdd.n8013 vss 0.00324f
C8478 vdd.n8014 vss 0.0424f
C8479 vdd.n8015 vss 0.00324f
C8480 vdd.n8016 vss 0.0128f
C8481 vdd.n8017 vss 0.02f
C8482 vdd.n8018 vss 0.0132f
C8483 vdd.n8019 vss 0.00925f
C8484 vdd.n8020 vss 0.00425f
C8485 vdd.n8022 vss 0.0471f
C8486 vdd.n8023 vss 0.00425f
C8487 vdd.n8024 vss 0.00413f
C8488 vdd.n8025 vss 0.00251f
C8489 vdd.n8026 vss 0.0471f
C8490 vdd.n8027 vss 0.00251f
C8491 vdd.n8028 vss 0.00517f
C8492 vdd.n8029 vss 0.00679f
C8493 vdd.n8030 vss 0.00324f
C8494 vdd.n8031 vss 0.00324f
C8495 vdd.n8032 vss 0.0132f
C8496 vdd.n8033 vss 0.0424f
C8497 vdd.n8034 vss 0.02f
C8498 vdd.n8035 vss 0.00425f
C8499 vdd.n8037 vss 0.0471f
C8500 vdd.n8038 vss 0.00425f
C8501 vdd.n8039 vss 0.00925f
C8502 vdd.n8040 vss 0.00679f
C8503 vdd.n8041 vss 0.00517f
C8504 vdd.n8042 vss 0.00251f
C8505 vdd.n8043 vss 0.0471f
C8506 vdd.n8044 vss 0.00251f
C8507 vdd.n8045 vss 0.0112f
C8508 vdd.n8046 vss 0.0955f
C8509 vdd.n8047 vss 0.0608f
C8510 vdd.n8048 vss 0.00324f
C8511 vdd.n8049 vss 0.0112f
C8512 vdd.n8050 vss 0.0128f
C8513 vdd.n8051 vss 0.00413f
C8514 vdd.n8052 vss 0.00413f
C8515 vdd.n8053 vss 0.0471f
C8516 vdd.n8054 vss 0.0471f
C8517 vdd.n8055 vss 0.00324f
C8518 vdd.n8056 vss 0.00413f
C8519 vdd.n8057 vss 0.00413f
C8520 vdd.n8058 vss 0.00679f
C8521 vdd.n8059 vss 0.00413f
C8522 vdd.n8060 vss 0.0471f
C8523 vdd.n8061 vss 0.00324f
C8524 vdd.n8062 vss 0.0424f
C8525 vdd.n8063 vss 0.00324f
C8526 vdd.n8064 vss 0.0128f
C8527 vdd.n8065 vss 0.02f
C8528 vdd.n8066 vss 0.0132f
C8529 vdd.n8067 vss 0.00925f
C8530 vdd.n8068 vss 0.00425f
C8531 vdd.n8070 vss 0.0471f
C8532 vdd.n8071 vss 0.00425f
C8533 vdd.n8072 vss 0.00413f
C8534 vdd.n8073 vss 0.00251f
C8535 vdd.n8074 vss 0.0471f
C8536 vdd.n8075 vss 0.00251f
C8537 vdd.n8076 vss 0.00517f
C8538 vdd.n8077 vss 0.00679f
C8539 vdd.n8078 vss 0.00324f
C8540 vdd.n8079 vss 0.00324f
C8541 vdd.n8080 vss 0.0132f
C8542 vdd.n8081 vss 0.0424f
C8543 vdd.n8082 vss 0.02f
C8544 vdd.n8083 vss 0.00425f
C8545 vdd.n8085 vss 0.0471f
C8546 vdd.n8086 vss 0.00425f
C8547 vdd.n8087 vss 0.00925f
C8548 vdd.n8088 vss 0.00679f
C8549 vdd.n8089 vss 0.00517f
C8550 vdd.n8090 vss 0.00251f
C8551 vdd.n8091 vss 0.0471f
C8552 vdd.n8092 vss 0.00251f
C8553 vdd.n8093 vss 0.0112f
C8554 vdd.n8094 vss 0.0128f
C8555 vdd.n8095 vss 0.0666f
C8556 vdd.n8096 vss 0.0912f
C8557 vdd.n8097 vss 0.0824f
C8558 vdd.n8098 vss 0.0567f
C8559 vdd.n8099 vss 0.00324f
C8560 vdd.n8100 vss 0.0112f
C8561 vdd.n8101 vss 0.0128f
C8562 vdd.n8102 vss 0.00413f
C8563 vdd.n8103 vss 0.00413f
C8564 vdd.n8104 vss 0.0471f
C8565 vdd.n8105 vss 0.0471f
C8566 vdd.n8106 vss 0.00324f
C8567 vdd.n8107 vss 0.00413f
C8568 vdd.n8108 vss 0.00413f
C8569 vdd.n8109 vss 0.00679f
C8570 vdd.n8110 vss 0.00413f
C8571 vdd.n8111 vss 0.0471f
C8572 vdd.n8112 vss 0.00324f
C8573 vdd.n8113 vss 0.0424f
C8574 vdd.n8114 vss 0.00324f
C8575 vdd.n8115 vss 0.0128f
C8576 vdd.n8116 vss 0.02f
C8577 vdd.n8117 vss 0.0132f
C8578 vdd.n8118 vss 0.00925f
C8579 vdd.n8119 vss 0.00425f
C8580 vdd.n8121 vss 0.0471f
C8581 vdd.n8122 vss 0.00425f
C8582 vdd.n8123 vss 0.00413f
C8583 vdd.n8124 vss 0.00251f
C8584 vdd.n8125 vss 0.0471f
C8585 vdd.n8126 vss 0.00251f
C8586 vdd.n8127 vss 0.00517f
C8587 vdd.n8128 vss 0.00679f
C8588 vdd.n8129 vss 0.00324f
C8589 vdd.n8130 vss 0.00324f
C8590 vdd.n8131 vss 0.0132f
C8591 vdd.n8132 vss 0.0424f
C8592 vdd.n8133 vss 0.02f
C8593 vdd.n8134 vss 0.00425f
C8594 vdd.n8136 vss 0.0471f
C8595 vdd.n8137 vss 0.00425f
C8596 vdd.n8138 vss 0.00925f
C8597 vdd.n8139 vss 0.00679f
C8598 vdd.n8140 vss 0.00517f
C8599 vdd.n8141 vss 0.00251f
C8600 vdd.n8142 vss 0.0471f
C8601 vdd.n8143 vss 0.00251f
C8602 vdd.n8144 vss 0.0112f
C8603 vdd.n8145 vss 0.0128f
C8604 vdd.n8146 vss 0.00324f
C8605 vdd.n8147 vss 0.0112f
C8606 vdd.n8148 vss 0.0128f
C8607 vdd.n8149 vss 0.00413f
C8608 vdd.n8150 vss 0.00413f
C8609 vdd.n8151 vss 0.0471f
C8610 vdd.n8152 vss 0.0471f
C8611 vdd.n8153 vss 0.00324f
C8612 vdd.n8154 vss 0.00413f
C8613 vdd.n8155 vss 0.00413f
C8614 vdd.n8156 vss 0.00679f
C8615 vdd.n8157 vss 0.00413f
C8616 vdd.n8158 vss 0.0471f
C8617 vdd.n8159 vss 0.00324f
C8618 vdd.n8160 vss 0.0424f
C8619 vdd.n8161 vss 0.00324f
C8620 vdd.n8162 vss 0.0128f
C8621 vdd.n8163 vss 0.02f
C8622 vdd.n8164 vss 0.0132f
C8623 vdd.n8165 vss 0.00925f
C8624 vdd.n8166 vss 0.00425f
C8625 vdd.n8168 vss 0.0471f
C8626 vdd.n8169 vss 0.00425f
C8627 vdd.n8170 vss 0.00413f
C8628 vdd.n8171 vss 0.00251f
C8629 vdd.n8172 vss 0.0471f
C8630 vdd.n8173 vss 0.00251f
C8631 vdd.n8174 vss 0.00517f
C8632 vdd.n8175 vss 0.00679f
C8633 vdd.n8176 vss 0.00324f
C8634 vdd.n8177 vss 0.00324f
C8635 vdd.n8178 vss 0.0132f
C8636 vdd.n8179 vss 0.0424f
C8637 vdd.n8180 vss 0.02f
C8638 vdd.n8181 vss 0.00425f
C8639 vdd.n8183 vss 0.0471f
C8640 vdd.n8184 vss 0.00425f
C8641 vdd.n8185 vss 0.00925f
C8642 vdd.n8186 vss 0.00679f
C8643 vdd.n8187 vss 0.00517f
C8644 vdd.n8188 vss 0.00251f
C8645 vdd.n8189 vss 0.0471f
C8646 vdd.n8190 vss 0.00251f
C8647 vdd.n8191 vss 0.0112f
C8648 vdd.n8192 vss 0.0128f
C8649 vdd.n8193 vss 0.0564f
C8650 vdd.n8194 vss 0.00324f
C8651 vdd.n8195 vss 0.0112f
C8652 vdd.n8196 vss 0.0128f
C8653 vdd.n8197 vss 0.00413f
C8654 vdd.n8198 vss 0.00413f
C8655 vdd.n8199 vss 0.0471f
C8656 vdd.n8200 vss 0.0471f
C8657 vdd.n8201 vss 0.00324f
C8658 vdd.n8202 vss 0.00413f
C8659 vdd.n8203 vss 0.00413f
C8660 vdd.n8204 vss 0.00679f
C8661 vdd.n8205 vss 0.00413f
C8662 vdd.n8206 vss 0.0471f
C8663 vdd.n8207 vss 0.00324f
C8664 vdd.n8208 vss 0.0424f
C8665 vdd.n8209 vss 0.00324f
C8666 vdd.n8210 vss 0.0128f
C8667 vdd.n8211 vss 0.02f
C8668 vdd.n8212 vss 0.0132f
C8669 vdd.n8213 vss 0.00925f
C8670 vdd.n8214 vss 0.00425f
C8671 vdd.n8216 vss 0.0471f
C8672 vdd.n8217 vss 0.00425f
C8673 vdd.n8218 vss 0.00413f
C8674 vdd.n8219 vss 0.00251f
C8675 vdd.n8220 vss 0.0471f
C8676 vdd.n8221 vss 0.00251f
C8677 vdd.n8222 vss 0.00517f
C8678 vdd.n8223 vss 0.00679f
C8679 vdd.n8224 vss 0.00324f
C8680 vdd.n8225 vss 0.00324f
C8681 vdd.n8226 vss 0.0132f
C8682 vdd.n8227 vss 0.0424f
C8683 vdd.n8228 vss 0.02f
C8684 vdd.n8229 vss 0.00425f
C8685 vdd.n8231 vss 0.0471f
C8686 vdd.n8232 vss 0.00425f
C8687 vdd.n8233 vss 0.00925f
C8688 vdd.n8234 vss 0.00679f
C8689 vdd.n8235 vss 0.00517f
C8690 vdd.n8236 vss 0.00251f
C8691 vdd.n8237 vss 0.0471f
C8692 vdd.n8238 vss 0.00251f
C8693 vdd.n8239 vss 0.0112f
C8694 vdd.n8240 vss 0.0128f
C8695 vdd.n8241 vss 0.183f
C8696 vdd.n8242 vss 0.256f
C8697 vdd.n8243 vss 0.12f
C8698 vdd.n8244 vss 0.0608f
C8699 vdd.n8245 vss 0.00324f
C8700 vdd.n8246 vss 0.0112f
C8701 vdd.n8247 vss 0.0128f
C8702 vdd.n8248 vss 0.00413f
C8703 vdd.n8249 vss 0.00413f
C8704 vdd.n8250 vss 0.0471f
C8705 vdd.n8251 vss 0.0471f
C8706 vdd.n8252 vss 0.00324f
C8707 vdd.n8253 vss 0.00413f
C8708 vdd.n8254 vss 0.00413f
C8709 vdd.n8255 vss 0.00679f
C8710 vdd.n8256 vss 0.00413f
C8711 vdd.n8257 vss 0.0471f
C8712 vdd.n8258 vss 0.00324f
C8713 vdd.n8259 vss 0.0424f
C8714 vdd.n8260 vss 0.00324f
C8715 vdd.n8261 vss 0.0128f
C8716 vdd.n8262 vss 0.02f
C8717 vdd.n8263 vss 0.0132f
C8718 vdd.n8264 vss 0.00925f
C8719 vdd.n8265 vss 0.00425f
C8720 vdd.n8267 vss 0.0471f
C8721 vdd.n8268 vss 0.00425f
C8722 vdd.n8269 vss 0.00413f
C8723 vdd.n8270 vss 0.00251f
C8724 vdd.n8271 vss 0.0471f
C8725 vdd.n8272 vss 0.00251f
C8726 vdd.n8273 vss 0.00517f
C8727 vdd.n8274 vss 0.00679f
C8728 vdd.n8275 vss 0.00324f
C8729 vdd.n8276 vss 0.00324f
C8730 vdd.n8277 vss 0.0132f
C8731 vdd.n8278 vss 0.0424f
C8732 vdd.n8279 vss 0.02f
C8733 vdd.n8280 vss 0.00425f
C8734 vdd.n8282 vss 0.0471f
C8735 vdd.n8283 vss 0.00425f
C8736 vdd.n8284 vss 0.00925f
C8737 vdd.n8285 vss 0.00679f
C8738 vdd.n8286 vss 0.00517f
C8739 vdd.n8287 vss 0.00251f
C8740 vdd.n8288 vss 0.0471f
C8741 vdd.n8289 vss 0.00251f
C8742 vdd.n8290 vss 0.0112f
C8743 vdd.n8291 vss 0.0128f
C8744 vdd.n8292 vss 0.0666f
C8745 vdd.n8293 vss 0.118f
C8746 vdd.n8294 vss 0.121f
C8747 vdd.n8295 vss 0.00324f
C8748 vdd.n8296 vss 0.0112f
C8749 vdd.n8297 vss 0.0128f
C8750 vdd.n8298 vss 0.00413f
C8751 vdd.n8299 vss 0.00413f
C8752 vdd.n8300 vss 0.0471f
C8753 vdd.n8301 vss 0.0471f
C8754 vdd.n8302 vss 0.00324f
C8755 vdd.n8303 vss 0.00413f
C8756 vdd.n8304 vss 0.00413f
C8757 vdd.n8305 vss 0.00679f
C8758 vdd.n8306 vss 0.00413f
C8759 vdd.n8307 vss 0.0471f
C8760 vdd.n8308 vss 0.00324f
C8761 vdd.n8309 vss 0.0424f
C8762 vdd.n8310 vss 0.00324f
C8763 vdd.n8311 vss 0.0128f
C8764 vdd.n8312 vss 0.02f
C8765 vdd.n8313 vss 0.0132f
C8766 vdd.n8314 vss 0.00925f
C8767 vdd.n8315 vss 0.00425f
C8768 vdd.n8317 vss 0.0471f
C8769 vdd.n8318 vss 0.00425f
C8770 vdd.n8319 vss 0.00413f
C8771 vdd.n8320 vss 0.00251f
C8772 vdd.n8321 vss 0.0471f
C8773 vdd.n8322 vss 0.00251f
C8774 vdd.n8323 vss 0.00517f
C8775 vdd.n8324 vss 0.00679f
C8776 vdd.n8325 vss 0.00324f
C8777 vdd.n8326 vss 0.00324f
C8778 vdd.n8327 vss 0.0132f
C8779 vdd.n8328 vss 0.0424f
C8780 vdd.n8329 vss 0.02f
C8781 vdd.n8330 vss 0.00425f
C8782 vdd.n8332 vss 0.0471f
C8783 vdd.n8333 vss 0.00425f
C8784 vdd.n8334 vss 0.00925f
C8785 vdd.n8335 vss 0.00679f
C8786 vdd.n8336 vss 0.00517f
C8787 vdd.n8337 vss 0.00251f
C8788 vdd.n8338 vss 0.0471f
C8789 vdd.n8339 vss 0.00251f
C8790 vdd.n8340 vss 0.0112f
C8791 vdd.n8341 vss 0.0955f
C8792 vdd.n8342 vss 0.0608f
C8793 vdd.n8343 vss 0.00324f
C8794 vdd.n8344 vss 0.0112f
C8795 vdd.n8345 vss 0.0128f
C8796 vdd.n8346 vss 0.00413f
C8797 vdd.n8347 vss 0.00413f
C8798 vdd.n8348 vss 0.0471f
C8799 vdd.n8349 vss 0.0471f
C8800 vdd.n8350 vss 0.00324f
C8801 vdd.n8351 vss 0.00413f
C8802 vdd.n8352 vss 0.00413f
C8803 vdd.n8353 vss 0.00679f
C8804 vdd.n8354 vss 0.00413f
C8805 vdd.n8355 vss 0.0471f
C8806 vdd.n8356 vss 0.00324f
C8807 vdd.n8357 vss 0.0424f
C8808 vdd.n8358 vss 0.00324f
C8809 vdd.n8359 vss 0.0128f
C8810 vdd.n8360 vss 0.02f
C8811 vdd.n8361 vss 0.0132f
C8812 vdd.n8362 vss 0.00925f
C8813 vdd.n8363 vss 0.00425f
C8814 vdd.n8365 vss 0.0471f
C8815 vdd.n8366 vss 0.00425f
C8816 vdd.n8367 vss 0.00413f
C8817 vdd.n8368 vss 0.00251f
C8818 vdd.n8369 vss 0.0471f
C8819 vdd.n8370 vss 0.00251f
C8820 vdd.n8371 vss 0.00517f
C8821 vdd.n8372 vss 0.00679f
C8822 vdd.n8373 vss 0.00324f
C8823 vdd.n8374 vss 0.00324f
C8824 vdd.n8375 vss 0.0132f
C8825 vdd.n8376 vss 0.0424f
C8826 vdd.n8377 vss 0.02f
C8827 vdd.n8378 vss 0.00425f
C8828 vdd.n8380 vss 0.0471f
C8829 vdd.n8381 vss 0.00425f
C8830 vdd.n8382 vss 0.00925f
C8831 vdd.n8383 vss 0.00679f
C8832 vdd.n8384 vss 0.00517f
C8833 vdd.n8385 vss 0.00251f
C8834 vdd.n8386 vss 0.0471f
C8835 vdd.n8387 vss 0.00251f
C8836 vdd.n8388 vss 0.0112f
C8837 vdd.n8389 vss 0.0128f
C8838 vdd.n8390 vss 0.0666f
C8839 vdd.n8391 vss 0.118f
C8840 vdd.n8392 vss 0.0935f
C8841 vdd.n8393 vss 0.00324f
C8842 vdd.n8394 vss 0.0112f
C8843 vdd.n8395 vss 0.0128f
C8844 vdd.n8396 vss 0.00413f
C8845 vdd.n8397 vss 0.00413f
C8846 vdd.n8398 vss 0.0471f
C8847 vdd.n8399 vss 0.0471f
C8848 vdd.n8400 vss 0.00324f
C8849 vdd.n8401 vss 0.00413f
C8850 vdd.n8402 vss 0.00413f
C8851 vdd.n8403 vss 0.00679f
C8852 vdd.n8404 vss 0.00413f
C8853 vdd.n8405 vss 0.0471f
C8854 vdd.n8406 vss 0.00324f
C8855 vdd.n8407 vss 0.0424f
C8856 vdd.n8408 vss 0.00324f
C8857 vdd.n8409 vss 0.0128f
C8858 vdd.n8410 vss 0.02f
C8859 vdd.n8411 vss 0.0132f
C8860 vdd.n8412 vss 0.00925f
C8861 vdd.n8413 vss 0.00425f
C8862 vdd.n8415 vss 0.0471f
C8863 vdd.n8416 vss 0.00425f
C8864 vdd.n8417 vss 0.00413f
C8865 vdd.n8418 vss 0.00251f
C8866 vdd.n8419 vss 0.0471f
C8867 vdd.n8420 vss 0.00251f
C8868 vdd.n8421 vss 0.00517f
C8869 vdd.n8422 vss 0.00679f
C8870 vdd.n8423 vss 0.00324f
C8871 vdd.n8424 vss 0.00324f
C8872 vdd.n8425 vss 0.0132f
C8873 vdd.n8426 vss 0.0424f
C8874 vdd.n8427 vss 0.02f
C8875 vdd.n8428 vss 0.00425f
C8876 vdd.n8430 vss 0.0471f
C8877 vdd.n8431 vss 0.00425f
C8878 vdd.n8432 vss 0.00925f
C8879 vdd.n8433 vss 0.00679f
C8880 vdd.n8434 vss 0.00517f
C8881 vdd.n8435 vss 0.00251f
C8882 vdd.n8436 vss 0.0471f
C8883 vdd.n8437 vss 0.00251f
C8884 vdd.n8438 vss 0.0112f
C8885 vdd.n8439 vss 0.0128f
C8886 vdd.n8440 vss 0.00324f
C8887 vdd.n8441 vss 0.0112f
C8888 vdd.n8442 vss 0.0128f
C8889 vdd.n8443 vss 0.00413f
C8890 vdd.n8444 vss 0.00413f
C8891 vdd.n8445 vss 0.0471f
C8892 vdd.n8446 vss 0.0471f
C8893 vdd.n8447 vss 0.00324f
C8894 vdd.n8448 vss 0.00413f
C8895 vdd.n8449 vss 0.00413f
C8896 vdd.n8450 vss 0.00679f
C8897 vdd.n8451 vss 0.00413f
C8898 vdd.n8452 vss 0.0471f
C8899 vdd.n8453 vss 0.00324f
C8900 vdd.n8454 vss 0.0424f
C8901 vdd.n8455 vss 0.00324f
C8902 vdd.n8456 vss 0.0128f
C8903 vdd.n8457 vss 0.02f
C8904 vdd.n8458 vss 0.0132f
C8905 vdd.n8459 vss 0.00925f
C8906 vdd.n8460 vss 0.00425f
C8907 vdd.n8462 vss 0.0471f
C8908 vdd.n8463 vss 0.00425f
C8909 vdd.n8464 vss 0.00413f
C8910 vdd.n8465 vss 0.00251f
C8911 vdd.n8466 vss 0.0471f
C8912 vdd.n8467 vss 0.00251f
C8913 vdd.n8468 vss 0.00517f
C8914 vdd.n8469 vss 0.00679f
C8915 vdd.n8470 vss 0.00324f
C8916 vdd.n8471 vss 0.00324f
C8917 vdd.n8472 vss 0.0132f
C8918 vdd.n8473 vss 0.0424f
C8919 vdd.n8474 vss 0.02f
C8920 vdd.n8475 vss 0.00425f
C8921 vdd.n8477 vss 0.0471f
C8922 vdd.n8478 vss 0.00425f
C8923 vdd.n8479 vss 0.00925f
C8924 vdd.n8480 vss 0.00679f
C8925 vdd.n8481 vss 0.00517f
C8926 vdd.n8482 vss 0.00251f
C8927 vdd.n8483 vss 0.0471f
C8928 vdd.n8484 vss 0.00251f
C8929 vdd.n8485 vss 0.0112f
C8930 vdd.n8486 vss 0.0128f
C8931 vdd.n8487 vss 0.144f
C8932 vdd.n8488 vss 0.143f
C8933 vdd.n8489 vss 0.0608f
C8934 vdd.n8490 vss 0.00324f
C8935 vdd.n8491 vss 0.0112f
C8936 vdd.n8492 vss 0.0128f
C8937 vdd.n8493 vss 0.00413f
C8938 vdd.n8494 vss 0.00413f
C8939 vdd.n8495 vss 0.0471f
C8940 vdd.n8496 vss 0.0471f
C8941 vdd.n8497 vss 0.00324f
C8942 vdd.n8498 vss 0.00413f
C8943 vdd.n8499 vss 0.00413f
C8944 vdd.n8500 vss 0.00679f
C8945 vdd.n8501 vss 0.00413f
C8946 vdd.n8502 vss 0.0471f
C8947 vdd.n8503 vss 0.00324f
C8948 vdd.n8504 vss 0.0424f
C8949 vdd.n8505 vss 0.00324f
C8950 vdd.n8506 vss 0.0128f
C8951 vdd.n8507 vss 0.02f
C8952 vdd.n8508 vss 0.0132f
C8953 vdd.n8509 vss 0.00925f
C8954 vdd.n8510 vss 0.00425f
C8955 vdd.n8512 vss 0.0471f
C8956 vdd.n8513 vss 0.00425f
C8957 vdd.n8514 vss 0.00413f
C8958 vdd.n8515 vss 0.00251f
C8959 vdd.n8516 vss 0.0471f
C8960 vdd.n8517 vss 0.00251f
C8961 vdd.n8518 vss 0.00517f
C8962 vdd.n8519 vss 0.00679f
C8963 vdd.n8520 vss 0.00324f
C8964 vdd.n8521 vss 0.00324f
C8965 vdd.n8522 vss 0.0132f
C8966 vdd.n8523 vss 0.0424f
C8967 vdd.n8524 vss 0.02f
C8968 vdd.n8525 vss 0.00425f
C8969 vdd.n8527 vss 0.0471f
C8970 vdd.n8528 vss 0.00425f
C8971 vdd.n8529 vss 0.00925f
C8972 vdd.n8530 vss 0.00679f
C8973 vdd.n8531 vss 0.00517f
C8974 vdd.n8532 vss 0.00251f
C8975 vdd.n8533 vss 0.0471f
C8976 vdd.n8534 vss 0.00251f
C8977 vdd.n8535 vss 0.0112f
C8978 vdd.n8536 vss 0.0128f
C8979 vdd.n8537 vss 0.0666f
C8980 vdd.n8538 vss 0.118f
C8981 vdd.n8539 vss 0.121f
C8982 vdd.n8540 vss 0.00324f
C8983 vdd.n8541 vss 0.0112f
C8984 vdd.n8542 vss 0.0128f
C8985 vdd.n8543 vss 0.00413f
C8986 vdd.n8544 vss 0.00413f
C8987 vdd.n8545 vss 0.0471f
C8988 vdd.n8546 vss 0.0471f
C8989 vdd.n8547 vss 0.00324f
C8990 vdd.n8548 vss 0.00413f
C8991 vdd.n8549 vss 0.00413f
C8992 vdd.n8550 vss 0.00679f
C8993 vdd.n8551 vss 0.00413f
C8994 vdd.n8552 vss 0.0471f
C8995 vdd.n8553 vss 0.00324f
C8996 vdd.n8554 vss 0.0424f
C8997 vdd.n8555 vss 0.00324f
C8998 vdd.n8556 vss 0.0128f
C8999 vdd.n8557 vss 0.02f
C9000 vdd.n8558 vss 0.0132f
C9001 vdd.n8559 vss 0.00925f
C9002 vdd.n8560 vss 0.00425f
C9003 vdd.n8562 vss 0.0471f
C9004 vdd.n8563 vss 0.00425f
C9005 vdd.n8564 vss 0.00413f
C9006 vdd.n8565 vss 0.00251f
C9007 vdd.n8566 vss 0.0471f
C9008 vdd.n8567 vss 0.00251f
C9009 vdd.n8568 vss 0.00517f
C9010 vdd.n8569 vss 0.00679f
C9011 vdd.n8570 vss 0.00324f
C9012 vdd.n8571 vss 0.00324f
C9013 vdd.n8572 vss 0.0132f
C9014 vdd.n8573 vss 0.0424f
C9015 vdd.n8574 vss 0.02f
C9016 vdd.n8575 vss 0.00425f
C9017 vdd.n8577 vss 0.0471f
C9018 vdd.n8578 vss 0.00425f
C9019 vdd.n8579 vss 0.00925f
C9020 vdd.n8580 vss 0.00679f
C9021 vdd.n8581 vss 0.00517f
C9022 vdd.n8582 vss 0.00251f
C9023 vdd.n8583 vss 0.0471f
C9024 vdd.n8584 vss 0.00251f
C9025 vdd.n8585 vss 0.0112f
C9026 vdd.n8586 vss 0.0955f
C9027 vdd.n8587 vss 0.0608f
C9028 vdd.n8588 vss 0.00324f
C9029 vdd.n8589 vss 0.0112f
C9030 vdd.n8590 vss 0.0128f
C9031 vdd.n8591 vss 0.00413f
C9032 vdd.n8592 vss 0.00413f
C9033 vdd.n8593 vss 0.0471f
C9034 vdd.n8594 vss 0.0471f
C9035 vdd.n8595 vss 0.00324f
C9036 vdd.n8596 vss 0.00413f
C9037 vdd.n8597 vss 0.00413f
C9038 vdd.n8598 vss 0.00679f
C9039 vdd.n8599 vss 0.00413f
C9040 vdd.n8600 vss 0.0471f
C9041 vdd.n8601 vss 0.00324f
C9042 vdd.n8602 vss 0.0424f
C9043 vdd.n8603 vss 0.00324f
C9044 vdd.n8604 vss 0.0128f
C9045 vdd.n8605 vss 0.02f
C9046 vdd.n8606 vss 0.0132f
C9047 vdd.n8607 vss 0.00925f
C9048 vdd.n8608 vss 0.00425f
C9049 vdd.n8610 vss 0.0471f
C9050 vdd.n8611 vss 0.00425f
C9051 vdd.n8612 vss 0.00413f
C9052 vdd.n8613 vss 0.00251f
C9053 vdd.n8614 vss 0.0471f
C9054 vdd.n8615 vss 0.00251f
C9055 vdd.n8616 vss 0.00517f
C9056 vdd.n8617 vss 0.00679f
C9057 vdd.n8618 vss 0.00324f
C9058 vdd.n8619 vss 0.00324f
C9059 vdd.n8620 vss 0.0132f
C9060 vdd.n8621 vss 0.0424f
C9061 vdd.n8622 vss 0.02f
C9062 vdd.n8623 vss 0.00425f
C9063 vdd.n8625 vss 0.0471f
C9064 vdd.n8626 vss 0.00425f
C9065 vdd.n8627 vss 0.00925f
C9066 vdd.n8628 vss 0.00679f
C9067 vdd.n8629 vss 0.00517f
C9068 vdd.n8630 vss 0.00251f
C9069 vdd.n8631 vss 0.0471f
C9070 vdd.n8632 vss 0.00251f
C9071 vdd.n8633 vss 0.0112f
C9072 vdd.n8634 vss 0.0128f
C9073 vdd.n8635 vss 0.0666f
C9074 vdd.n8636 vss 0.0912f
C9075 vdd.n8637 vss 0.0824f
C9076 vdd.n8638 vss 0.0567f
C9077 vdd.n8639 vss 0.00324f
C9078 vdd.n8640 vss 0.0112f
C9079 vdd.n8641 vss 0.0128f
C9080 vdd.n8642 vss 0.00413f
C9081 vdd.n8643 vss 0.00413f
C9082 vdd.n8644 vss 0.0471f
C9083 vdd.n8645 vss 0.0471f
C9084 vdd.n8646 vss 0.00324f
C9085 vdd.n8647 vss 0.00413f
C9086 vdd.n8648 vss 0.00413f
C9087 vdd.n8649 vss 0.00679f
C9088 vdd.n8650 vss 0.00413f
C9089 vdd.n8651 vss 0.0471f
C9090 vdd.n8652 vss 0.00324f
C9091 vdd.n8653 vss 0.0424f
C9092 vdd.n8654 vss 0.00324f
C9093 vdd.n8655 vss 0.0128f
C9094 vdd.n8656 vss 0.02f
C9095 vdd.n8657 vss 0.0132f
C9096 vdd.n8658 vss 0.00925f
C9097 vdd.n8659 vss 0.00425f
C9098 vdd.n8661 vss 0.0471f
C9099 vdd.n8662 vss 0.00425f
C9100 vdd.n8663 vss 0.00413f
C9101 vdd.n8664 vss 0.00251f
C9102 vdd.n8665 vss 0.0471f
C9103 vdd.n8666 vss 0.00251f
C9104 vdd.n8667 vss 0.00517f
C9105 vdd.n8668 vss 0.00679f
C9106 vdd.n8669 vss 0.00324f
C9107 vdd.n8670 vss 0.00324f
C9108 vdd.n8671 vss 0.0132f
C9109 vdd.n8672 vss 0.0424f
C9110 vdd.n8673 vss 0.02f
C9111 vdd.n8674 vss 0.00425f
C9112 vdd.n8676 vss 0.0471f
C9113 vdd.n8677 vss 0.00425f
C9114 vdd.n8678 vss 0.00925f
C9115 vdd.n8679 vss 0.00679f
C9116 vdd.n8680 vss 0.00517f
C9117 vdd.n8681 vss 0.00251f
C9118 vdd.n8682 vss 0.0471f
C9119 vdd.n8683 vss 0.00251f
C9120 vdd.n8684 vss 0.0112f
C9121 vdd.n8685 vss 0.0128f
C9122 vdd.n8686 vss 0.00324f
C9123 vdd.n8687 vss 0.0112f
C9124 vdd.n8688 vss 0.0128f
C9125 vdd.n8689 vss 0.00413f
C9126 vdd.n8690 vss 0.00413f
C9127 vdd.n8691 vss 0.0471f
C9128 vdd.n8692 vss 0.0471f
C9129 vdd.n8693 vss 0.00324f
C9130 vdd.n8694 vss 0.00413f
C9131 vdd.n8695 vss 0.00413f
C9132 vdd.n8696 vss 0.00679f
C9133 vdd.n8697 vss 0.00413f
C9134 vdd.n8698 vss 0.0471f
C9135 vdd.n8699 vss 0.00324f
C9136 vdd.n8700 vss 0.0424f
C9137 vdd.n8701 vss 0.00324f
C9138 vdd.n8702 vss 0.0128f
C9139 vdd.n8703 vss 0.02f
C9140 vdd.n8704 vss 0.0132f
C9141 vdd.n8705 vss 0.00925f
C9142 vdd.n8706 vss 0.00425f
C9143 vdd.n8708 vss 0.0471f
C9144 vdd.n8709 vss 0.00425f
C9145 vdd.n8710 vss 0.00413f
C9146 vdd.n8711 vss 0.00251f
C9147 vdd.n8712 vss 0.0471f
C9148 vdd.n8713 vss 0.00251f
C9149 vdd.n8714 vss 0.00517f
C9150 vdd.n8715 vss 0.00679f
C9151 vdd.n8716 vss 0.00324f
C9152 vdd.n8717 vss 0.00324f
C9153 vdd.n8718 vss 0.0132f
C9154 vdd.n8719 vss 0.0424f
C9155 vdd.n8720 vss 0.02f
C9156 vdd.n8721 vss 0.00425f
C9157 vdd.n8723 vss 0.0471f
C9158 vdd.n8724 vss 0.00425f
C9159 vdd.n8725 vss 0.00925f
C9160 vdd.n8726 vss 0.00679f
C9161 vdd.n8727 vss 0.00517f
C9162 vdd.n8728 vss 0.00251f
C9163 vdd.n8729 vss 0.0471f
C9164 vdd.n8730 vss 0.00251f
C9165 vdd.n8731 vss 0.0112f
C9166 vdd.n8732 vss 0.0128f
C9167 vdd.n8733 vss 0.144f
C9168 vdd.n8734 vss 0.143f
C9169 vdd.n8735 vss 0.0608f
C9170 vdd.n8736 vss 0.00324f
C9171 vdd.n8737 vss 0.0112f
C9172 vdd.n8738 vss 0.0128f
C9173 vdd.n8739 vss 0.00413f
C9174 vdd.n8740 vss 0.00413f
C9175 vdd.n8741 vss 0.0471f
C9176 vdd.n8742 vss 0.0471f
C9177 vdd.n8743 vss 0.00324f
C9178 vdd.n8744 vss 0.00413f
C9179 vdd.n8745 vss 0.00413f
C9180 vdd.n8746 vss 0.00679f
C9181 vdd.n8747 vss 0.00413f
C9182 vdd.n8748 vss 0.0471f
C9183 vdd.n8749 vss 0.00324f
C9184 vdd.n8750 vss 0.0424f
C9185 vdd.n8751 vss 0.00324f
C9186 vdd.n8752 vss 0.0128f
C9187 vdd.n8753 vss 0.02f
C9188 vdd.n8754 vss 0.0132f
C9189 vdd.n8755 vss 0.00925f
C9190 vdd.n8756 vss 0.00425f
C9191 vdd.n8758 vss 0.0471f
C9192 vdd.n8759 vss 0.00425f
C9193 vdd.n8760 vss 0.00413f
C9194 vdd.n8761 vss 0.00251f
C9195 vdd.n8762 vss 0.0471f
C9196 vdd.n8763 vss 0.00251f
C9197 vdd.n8764 vss 0.00517f
C9198 vdd.n8765 vss 0.00679f
C9199 vdd.n8766 vss 0.00324f
C9200 vdd.n8767 vss 0.00324f
C9201 vdd.n8768 vss 0.0132f
C9202 vdd.n8769 vss 0.0424f
C9203 vdd.n8770 vss 0.02f
C9204 vdd.n8771 vss 0.00425f
C9205 vdd.n8773 vss 0.0471f
C9206 vdd.n8774 vss 0.00425f
C9207 vdd.n8775 vss 0.00925f
C9208 vdd.n8776 vss 0.00679f
C9209 vdd.n8777 vss 0.00517f
C9210 vdd.n8778 vss 0.00251f
C9211 vdd.n8779 vss 0.0471f
C9212 vdd.n8780 vss 0.00251f
C9213 vdd.n8781 vss 0.0112f
C9214 vdd.n8782 vss 0.0128f
C9215 vdd.n8783 vss 0.0666f
C9216 vdd.n8784 vss 0.118f
C9217 vdd.n8785 vss 0.121f
C9218 vdd.n8786 vss 0.00324f
C9219 vdd.n8787 vss 0.0112f
C9220 vdd.n8788 vss 0.0128f
C9221 vdd.n8789 vss 0.00413f
C9222 vdd.n8790 vss 0.00413f
C9223 vdd.n8791 vss 0.0471f
C9224 vdd.n8792 vss 0.0471f
C9225 vdd.n8793 vss 0.00324f
C9226 vdd.n8794 vss 0.00413f
C9227 vdd.n8795 vss 0.00413f
C9228 vdd.n8796 vss 0.00679f
C9229 vdd.n8797 vss 0.00413f
C9230 vdd.n8798 vss 0.0471f
C9231 vdd.n8799 vss 0.00324f
C9232 vdd.n8800 vss 0.0424f
C9233 vdd.n8801 vss 0.00324f
C9234 vdd.n8802 vss 0.0128f
C9235 vdd.n8803 vss 0.02f
C9236 vdd.n8804 vss 0.0132f
C9237 vdd.n8805 vss 0.00925f
C9238 vdd.n8806 vss 0.00425f
C9239 vdd.n8808 vss 0.0471f
C9240 vdd.n8809 vss 0.00425f
C9241 vdd.n8810 vss 0.00413f
C9242 vdd.n8811 vss 0.00251f
C9243 vdd.n8812 vss 0.0471f
C9244 vdd.n8813 vss 0.00251f
C9245 vdd.n8814 vss 0.00517f
C9246 vdd.n8815 vss 0.00679f
C9247 vdd.n8816 vss 0.00324f
C9248 vdd.n8817 vss 0.00324f
C9249 vdd.n8818 vss 0.0132f
C9250 vdd.n8819 vss 0.0424f
C9251 vdd.n8820 vss 0.02f
C9252 vdd.n8821 vss 0.00425f
C9253 vdd.n8823 vss 0.0471f
C9254 vdd.n8824 vss 0.00425f
C9255 vdd.n8825 vss 0.00925f
C9256 vdd.n8826 vss 0.00679f
C9257 vdd.n8827 vss 0.00517f
C9258 vdd.n8828 vss 0.00251f
C9259 vdd.n8829 vss 0.0471f
C9260 vdd.n8830 vss 0.00251f
C9261 vdd.n8831 vss 0.0112f
C9262 vdd.n8832 vss 0.0955f
C9263 vdd.n8833 vss 0.0608f
C9264 vdd.n8834 vss 0.00324f
C9265 vdd.n8835 vss 0.0112f
C9266 vdd.n8836 vss 0.0128f
C9267 vdd.n8837 vss 0.00413f
C9268 vdd.n8838 vss 0.00413f
C9269 vdd.n8839 vss 0.0471f
C9270 vdd.n8840 vss 0.0471f
C9271 vdd.n8841 vss 0.00324f
C9272 vdd.n8842 vss 0.00413f
C9273 vdd.n8843 vss 0.00413f
C9274 vdd.n8844 vss 0.00679f
C9275 vdd.n8845 vss 0.00413f
C9276 vdd.n8846 vss 0.0471f
C9277 vdd.n8847 vss 0.00324f
C9278 vdd.n8848 vss 0.0424f
C9279 vdd.n8849 vss 0.00324f
C9280 vdd.n8850 vss 0.0128f
C9281 vdd.n8851 vss 0.02f
C9282 vdd.n8852 vss 0.0132f
C9283 vdd.n8853 vss 0.00925f
C9284 vdd.n8854 vss 0.00425f
C9285 vdd.n8856 vss 0.0471f
C9286 vdd.n8857 vss 0.00425f
C9287 vdd.n8858 vss 0.00413f
C9288 vdd.n8859 vss 0.00251f
C9289 vdd.n8860 vss 0.0471f
C9290 vdd.n8861 vss 0.00251f
C9291 vdd.n8862 vss 0.00517f
C9292 vdd.n8863 vss 0.00679f
C9293 vdd.n8864 vss 0.00324f
C9294 vdd.n8865 vss 0.00324f
C9295 vdd.n8866 vss 0.0132f
C9296 vdd.n8867 vss 0.0424f
C9297 vdd.n8868 vss 0.02f
C9298 vdd.n8869 vss 0.00425f
C9299 vdd.n8871 vss 0.0471f
C9300 vdd.n8872 vss 0.00425f
C9301 vdd.n8873 vss 0.00925f
C9302 vdd.n8874 vss 0.00679f
C9303 vdd.n8875 vss 0.00517f
C9304 vdd.n8876 vss 0.00251f
C9305 vdd.n8877 vss 0.0471f
C9306 vdd.n8878 vss 0.00251f
C9307 vdd.n8879 vss 0.0112f
C9308 vdd.n8880 vss 0.0128f
C9309 vdd.n8881 vss 0.0666f
C9310 vdd.n8882 vss 0.299f
C9311 vdd.n8883 vss 0.00324f
C9312 vdd.n8884 vss 0.0112f
C9313 vdd.n8885 vss 0.0128f
C9314 vdd.n8886 vss 0.00413f
C9315 vdd.n8887 vss 0.00413f
C9316 vdd.n8888 vss 0.0471f
C9317 vdd.n8889 vss 0.0471f
C9318 vdd.n8890 vss 0.00324f
C9319 vdd.n8891 vss 0.00413f
C9320 vdd.n8892 vss 0.00413f
C9321 vdd.n8893 vss 0.00679f
C9322 vdd.n8894 vss 0.00413f
C9323 vdd.n8895 vss 0.0471f
C9324 vdd.n8896 vss 0.00324f
C9325 vdd.n8898 vss 0.00925f
C9326 vdd.n8899 vss 0.0471f
C9327 vdd.n8900 vss 0.00425f
C9328 vdd.n8901 vss 0.0424f
C9329 vdd.n8902 vss 0.0132f
C9330 vdd.n8903 vss 0.00324f
C9331 vdd.n8904 vss 0.0128f
C9332 vdd.n8905 vss 0.02f
C9333 vdd.n8906 vss 0.00425f
C9334 vdd.n8907 vss 0.00413f
C9335 vdd.n8908 vss 0.00251f
C9336 vdd.n8909 vss 0.0471f
C9337 vdd.n8910 vss 0.00251f
C9338 vdd.n8911 vss 0.00517f
C9339 vdd.n8912 vss 0.00679f
C9340 vdd.n8913 vss 0.00324f
C9341 vdd.n8914 vss 0.00324f
C9342 vdd.n8915 vss 0.0132f
C9343 vdd.n8916 vss 0.0424f
C9344 vdd.n8917 vss 0.02f
C9345 vdd.n8918 vss 0.00425f
C9346 vdd.n8919 vss 0.0471f
C9347 vdd.n8921 vss 0.00425f
C9348 vdd.n8922 vss 0.00925f
C9349 vdd.n8923 vss 0.00679f
C9350 vdd.n8924 vss 0.00517f
C9351 vdd.n8925 vss 0.00251f
C9352 vdd.n8926 vss 0.0471f
C9353 vdd.n8927 vss 0.00251f
C9354 vdd.n8928 vss 0.0112f
C9355 vdd.n8929 vss 0.0128f
C9356 vdd.n8930 vss 0.0619f
C9357 vdd.n8931 vss 0.262f
C9358 vdd.n8932 vss 0.00324f
C9359 vdd.n8933 vss 0.0112f
C9360 vdd.n8934 vss 0.0128f
C9361 vdd.n8935 vss 0.00413f
C9362 vdd.n8936 vss 0.00413f
C9363 vdd.n8937 vss 0.0471f
C9364 vdd.n8938 vss 0.0471f
C9365 vdd.n8939 vss 0.00324f
C9366 vdd.n8940 vss 0.00413f
C9367 vdd.n8941 vss 0.00413f
C9368 vdd.n8942 vss 0.00679f
C9369 vdd.n8943 vss 0.00413f
C9370 vdd.n8944 vss 0.0471f
C9371 vdd.n8945 vss 0.00324f
C9372 vdd.n8947 vss 0.00925f
C9373 vdd.n8948 vss 0.0471f
C9374 vdd.n8949 vss 0.00425f
C9375 vdd.n8950 vss 0.0424f
C9376 vdd.n8951 vss 0.0132f
C9377 vdd.n8952 vss 0.00324f
C9378 vdd.n8953 vss 0.0128f
C9379 vdd.n8954 vss 0.02f
C9380 vdd.n8955 vss 0.00425f
C9381 vdd.n8956 vss 0.00413f
C9382 vdd.n8957 vss 0.00251f
C9383 vdd.n8958 vss 0.0471f
C9384 vdd.n8959 vss 0.00251f
C9385 vdd.n8960 vss 0.00517f
C9386 vdd.n8961 vss 0.00679f
C9387 vdd.n8962 vss 0.00324f
C9388 vdd.n8963 vss 0.00324f
C9389 vdd.n8964 vss 0.0132f
C9390 vdd.n8965 vss 0.0424f
C9391 vdd.n8966 vss 0.02f
C9392 vdd.n8967 vss 0.00425f
C9393 vdd.n8968 vss 0.0471f
C9394 vdd.n8970 vss 0.00425f
C9395 vdd.n8971 vss 0.00925f
C9396 vdd.n8972 vss 0.00679f
C9397 vdd.n8973 vss 0.00517f
C9398 vdd.n8974 vss 0.00251f
C9399 vdd.n8975 vss 0.0471f
C9400 vdd.n8976 vss 0.00251f
C9401 vdd.n8977 vss 0.0112f
C9402 vdd.n8978 vss 0.0128f
C9403 vdd.n8979 vss 0.146f
C9404 vdd.n8980 vss 0.00324f
C9405 vdd.n8981 vss 0.0112f
C9406 vdd.n8982 vss 0.0128f
C9407 vdd.n8983 vss 0.00413f
C9408 vdd.n8984 vss 0.00413f
C9409 vdd.n8985 vss 0.0471f
C9410 vdd.n8986 vss 0.0471f
C9411 vdd.n8987 vss 0.00324f
C9412 vdd.n8988 vss 0.00413f
C9413 vdd.n8989 vss 0.00413f
C9414 vdd.n8990 vss 0.00679f
C9415 vdd.n8991 vss 0.00413f
C9416 vdd.n8992 vss 0.0471f
C9417 vdd.n8993 vss 0.00324f
C9418 vdd.n8995 vss 0.00925f
C9419 vdd.n8996 vss 0.0471f
C9420 vdd.n8997 vss 0.00425f
C9421 vdd.n8998 vss 0.0424f
C9422 vdd.n8999 vss 0.0132f
C9423 vdd.n9000 vss 0.00324f
C9424 vdd.n9001 vss 0.0128f
C9425 vdd.n9002 vss 0.02f
C9426 vdd.n9003 vss 0.00425f
C9427 vdd.n9004 vss 0.00413f
C9428 vdd.n9005 vss 0.00251f
C9429 vdd.n9006 vss 0.0471f
C9430 vdd.n9007 vss 0.00251f
C9431 vdd.n9008 vss 0.00517f
C9432 vdd.n9009 vss 0.00679f
C9433 vdd.n9010 vss 0.00324f
C9434 vdd.n9011 vss 0.00324f
C9435 vdd.n9012 vss 0.0132f
C9436 vdd.n9013 vss 0.0424f
C9437 vdd.n9014 vss 0.02f
C9438 vdd.n9015 vss 0.00425f
C9439 vdd.n9016 vss 0.0471f
C9440 vdd.n9018 vss 0.00425f
C9441 vdd.n9019 vss 0.00925f
C9442 vdd.n9020 vss 0.00679f
C9443 vdd.n9021 vss 0.00517f
C9444 vdd.n9022 vss 0.00251f
C9445 vdd.n9023 vss 0.0471f
C9446 vdd.n9024 vss 0.00251f
C9447 vdd.n9025 vss 0.0112f
C9448 vdd.n9026 vss 0.0128f
C9449 vdd.n9027 vss 0.146f
C9450 vdd.n9028 vss 0.0596f
C9451 vdd.n9029 vss 0.00324f
C9452 vdd.n9030 vss 0.0112f
C9453 vdd.n9031 vss 0.0128f
C9454 vdd.n9032 vss 0.00413f
C9455 vdd.n9033 vss 0.00413f
C9456 vdd.n9034 vss 0.0471f
C9457 vdd.n9035 vss 0.0471f
C9458 vdd.n9036 vss 0.00324f
C9459 vdd.n9037 vss 0.00413f
C9460 vdd.n9038 vss 0.00413f
C9461 vdd.n9039 vss 0.00679f
C9462 vdd.n9040 vss 0.00413f
C9463 vdd.n9041 vss 0.0471f
C9464 vdd.n9042 vss 0.00324f
C9465 vdd.n9044 vss 0.00925f
C9466 vdd.n9045 vss 0.0471f
C9467 vdd.n9046 vss 0.00425f
C9468 vdd.n9047 vss 0.0424f
C9469 vdd.n9048 vss 0.0132f
C9470 vdd.n9049 vss 0.00324f
C9471 vdd.n9050 vss 0.0128f
C9472 vdd.n9051 vss 0.02f
C9473 vdd.n9052 vss 0.00425f
C9474 vdd.n9053 vss 0.00413f
C9475 vdd.n9054 vss 0.00251f
C9476 vdd.n9055 vss 0.0471f
C9477 vdd.n9056 vss 0.00251f
C9478 vdd.n9057 vss 0.00517f
C9479 vdd.n9058 vss 0.00679f
C9480 vdd.n9059 vss 0.00324f
C9481 vdd.n9060 vss 0.00324f
C9482 vdd.n9061 vss 0.0132f
C9483 vdd.n9062 vss 0.0424f
C9484 vdd.n9063 vss 0.02f
C9485 vdd.n9064 vss 0.00425f
C9486 vdd.n9065 vss 0.0471f
C9487 vdd.n9067 vss 0.00425f
C9488 vdd.n9068 vss 0.00925f
C9489 vdd.n9069 vss 0.00679f
C9490 vdd.n9070 vss 0.00517f
C9491 vdd.n9071 vss 0.00251f
C9492 vdd.n9072 vss 0.0471f
C9493 vdd.n9073 vss 0.00251f
C9494 vdd.n9074 vss 0.0112f
C9495 vdd.n9075 vss 0.0128f
C9496 vdd.n9076 vss 0.0692f
C9497 vdd.n9077 vss 0.118f
C9498 vdd.n9078 vss 0.121f
C9499 vdd.n9079 vss 0.00324f
C9500 vdd.n9080 vss 0.0112f
C9501 vdd.n9081 vss 0.0128f
C9502 vdd.n9082 vss 0.00413f
C9503 vdd.n9083 vss 0.00413f
C9504 vdd.n9084 vss 0.0471f
C9505 vdd.n9085 vss 0.0471f
C9506 vdd.n9086 vss 0.00324f
C9507 vdd.n9087 vss 0.00413f
C9508 vdd.n9088 vss 0.00413f
C9509 vdd.n9089 vss 0.00679f
C9510 vdd.n9090 vss 0.00413f
C9511 vdd.n9091 vss 0.0471f
C9512 vdd.n9092 vss 0.00324f
C9513 vdd.n9094 vss 0.00925f
C9514 vdd.n9095 vss 0.0471f
C9515 vdd.n9096 vss 0.00425f
C9516 vdd.n9097 vss 0.0424f
C9517 vdd.n9098 vss 0.0132f
C9518 vdd.n9099 vss 0.00324f
C9519 vdd.n9100 vss 0.0128f
C9520 vdd.n9101 vss 0.02f
C9521 vdd.n9102 vss 0.00425f
C9522 vdd.n9103 vss 0.00413f
C9523 vdd.n9104 vss 0.00251f
C9524 vdd.n9105 vss 0.0471f
C9525 vdd.n9106 vss 0.00251f
C9526 vdd.n9107 vss 0.00517f
C9527 vdd.n9108 vss 0.00679f
C9528 vdd.n9109 vss 0.00324f
C9529 vdd.n9110 vss 0.00324f
C9530 vdd.n9111 vss 0.0132f
C9531 vdd.n9112 vss 0.0424f
C9532 vdd.n9113 vss 0.02f
C9533 vdd.n9114 vss 0.00425f
C9534 vdd.n9115 vss 0.0471f
C9535 vdd.n9117 vss 0.00425f
C9536 vdd.n9118 vss 0.00925f
C9537 vdd.n9119 vss 0.00679f
C9538 vdd.n9120 vss 0.00517f
C9539 vdd.n9121 vss 0.00251f
C9540 vdd.n9122 vss 0.0471f
C9541 vdd.n9123 vss 0.00251f
C9542 vdd.n9124 vss 0.0112f
C9543 vdd.n9125 vss 0.098f
C9544 vdd.n9126 vss 0.0596f
C9545 vdd.n9127 vss 0.00324f
C9546 vdd.n9128 vss 0.0112f
C9547 vdd.n9129 vss 0.0128f
C9548 vdd.n9130 vss 0.00413f
C9549 vdd.n9131 vss 0.00413f
C9550 vdd.n9132 vss 0.0471f
C9551 vdd.n9133 vss 0.0471f
C9552 vdd.n9134 vss 0.00324f
C9553 vdd.n9135 vss 0.00413f
C9554 vdd.n9136 vss 0.00413f
C9555 vdd.n9137 vss 0.00679f
C9556 vdd.n9138 vss 0.00413f
C9557 vdd.n9139 vss 0.0471f
C9558 vdd.n9140 vss 0.00324f
C9559 vdd.n9142 vss 0.00925f
C9560 vdd.n9143 vss 0.0471f
C9561 vdd.n9144 vss 0.00425f
C9562 vdd.n9145 vss 0.0424f
C9563 vdd.n9146 vss 0.0132f
C9564 vdd.n9147 vss 0.00324f
C9565 vdd.n9148 vss 0.0128f
C9566 vdd.n9149 vss 0.02f
C9567 vdd.n9150 vss 0.00425f
C9568 vdd.n9151 vss 0.00413f
C9569 vdd.n9152 vss 0.00251f
C9570 vdd.n9153 vss 0.0471f
C9571 vdd.n9154 vss 0.00251f
C9572 vdd.n9155 vss 0.00517f
C9573 vdd.n9156 vss 0.00679f
C9574 vdd.n9157 vss 0.00324f
C9575 vdd.n9158 vss 0.00324f
C9576 vdd.n9159 vss 0.0132f
C9577 vdd.n9160 vss 0.0424f
C9578 vdd.n9161 vss 0.02f
C9579 vdd.n9162 vss 0.00425f
C9580 vdd.n9163 vss 0.0471f
C9581 vdd.n9165 vss 0.00425f
C9582 vdd.n9166 vss 0.00925f
C9583 vdd.n9167 vss 0.00679f
C9584 vdd.n9168 vss 0.00517f
C9585 vdd.n9169 vss 0.00251f
C9586 vdd.n9170 vss 0.0471f
C9587 vdd.n9171 vss 0.00251f
C9588 vdd.n9172 vss 0.0112f
C9589 vdd.n9173 vss 0.0128f
C9590 vdd.n9174 vss 0.0692f
C9591 vdd.n9175 vss 0.0912f
C9592 vdd.n9176 vss 0.0824f
C9593 vdd.n9177 vss 0.059f
C9594 vdd.n9178 vss 0.00324f
C9595 vdd.n9179 vss 0.0112f
C9596 vdd.n9180 vss 0.0128f
C9597 vdd.n9181 vss 0.00413f
C9598 vdd.n9182 vss 0.00413f
C9599 vdd.n9183 vss 0.0471f
C9600 vdd.n9184 vss 0.0471f
C9601 vdd.n9185 vss 0.00324f
C9602 vdd.n9186 vss 0.00413f
C9603 vdd.n9187 vss 0.00413f
C9604 vdd.n9188 vss 0.00679f
C9605 vdd.n9189 vss 0.00413f
C9606 vdd.n9190 vss 0.0471f
C9607 vdd.n9191 vss 0.00324f
C9608 vdd.n9193 vss 0.00925f
C9609 vdd.n9194 vss 0.0471f
C9610 vdd.n9195 vss 0.00425f
C9611 vdd.n9196 vss 0.0424f
C9612 vdd.n9197 vss 0.0132f
C9613 vdd.n9198 vss 0.00324f
C9614 vdd.n9199 vss 0.0128f
C9615 vdd.n9200 vss 0.02f
C9616 vdd.n9201 vss 0.00425f
C9617 vdd.n9202 vss 0.00413f
C9618 vdd.n9203 vss 0.00251f
C9619 vdd.n9204 vss 0.0471f
C9620 vdd.n9205 vss 0.00251f
C9621 vdd.n9206 vss 0.00517f
C9622 vdd.n9207 vss 0.00679f
C9623 vdd.n9208 vss 0.00324f
C9624 vdd.n9209 vss 0.00324f
C9625 vdd.n9210 vss 0.0132f
C9626 vdd.n9211 vss 0.0424f
C9627 vdd.n9212 vss 0.02f
C9628 vdd.n9213 vss 0.00425f
C9629 vdd.n9214 vss 0.0471f
C9630 vdd.n9216 vss 0.00425f
C9631 vdd.n9217 vss 0.00925f
C9632 vdd.n9218 vss 0.00679f
C9633 vdd.n9219 vss 0.00517f
C9634 vdd.n9220 vss 0.00251f
C9635 vdd.n9221 vss 0.0471f
C9636 vdd.n9222 vss 0.00251f
C9637 vdd.n9223 vss 0.0112f
C9638 vdd.n9224 vss 0.0128f
C9639 vdd.n9225 vss 0.185f
C9640 vdd.n9226 vss 0.00324f
C9641 vdd.n9227 vss 0.0112f
C9642 vdd.n9228 vss 0.0128f
C9643 vdd.n9229 vss 0.00413f
C9644 vdd.n9230 vss 0.00413f
C9645 vdd.n9231 vss 0.0471f
C9646 vdd.n9232 vss 0.0471f
C9647 vdd.n9233 vss 0.00324f
C9648 vdd.n9234 vss 0.00413f
C9649 vdd.n9235 vss 0.00413f
C9650 vdd.n9236 vss 0.00679f
C9651 vdd.n9237 vss 0.00413f
C9652 vdd.n9238 vss 0.0471f
C9653 vdd.n9239 vss 0.00324f
C9654 vdd.n9241 vss 0.00925f
C9655 vdd.n9242 vss 0.0471f
C9656 vdd.n9243 vss 0.00425f
C9657 vdd.n9244 vss 0.0424f
C9658 vdd.n9245 vss 0.0132f
C9659 vdd.n9246 vss 0.00324f
C9660 vdd.n9247 vss 0.0128f
C9661 vdd.n9248 vss 0.02f
C9662 vdd.n9249 vss 0.00425f
C9663 vdd.n9250 vss 0.00413f
C9664 vdd.n9251 vss 0.00251f
C9665 vdd.n9252 vss 0.0471f
C9666 vdd.n9253 vss 0.00251f
C9667 vdd.n9254 vss 0.00517f
C9668 vdd.n9255 vss 0.00679f
C9669 vdd.n9256 vss 0.00324f
C9670 vdd.n9257 vss 0.00324f
C9671 vdd.n9258 vss 0.0132f
C9672 vdd.n9259 vss 0.0424f
C9673 vdd.n9260 vss 0.02f
C9674 vdd.n9261 vss 0.00425f
C9675 vdd.n9262 vss 0.0471f
C9676 vdd.n9264 vss 0.00425f
C9677 vdd.n9265 vss 0.00925f
C9678 vdd.n9266 vss 0.00679f
C9679 vdd.n9267 vss 0.00517f
C9680 vdd.n9268 vss 0.00251f
C9681 vdd.n9269 vss 0.0471f
C9682 vdd.n9270 vss 0.00251f
C9683 vdd.n9271 vss 0.0112f
C9684 vdd.n9272 vss 0.0128f
C9685 vdd.n9273 vss 0.059f
C9686 vdd.n9274 vss 0.256f
C9687 vdd.n9275 vss 0.00324f
C9688 vdd.n9276 vss 0.0112f
C9689 vdd.n9277 vss 0.0128f
C9690 vdd.n9278 vss 0.00413f
C9691 vdd.n9279 vss 0.00413f
C9692 vdd.n9280 vss 0.0471f
C9693 vdd.n9281 vss 0.0471f
C9694 vdd.n9282 vss 0.00324f
C9695 vdd.n9283 vss 0.00413f
C9696 vdd.n9284 vss 0.00413f
C9697 vdd.n9285 vss 0.00679f
C9698 vdd.n9286 vss 0.00413f
C9699 vdd.n9287 vss 0.0471f
C9700 vdd.n9288 vss 0.00324f
C9701 vdd.n9290 vss 0.00925f
C9702 vdd.n9291 vss 0.0471f
C9703 vdd.n9292 vss 0.00425f
C9704 vdd.n9293 vss 0.0424f
C9705 vdd.n9294 vss 0.0132f
C9706 vdd.n9295 vss 0.00324f
C9707 vdd.n9296 vss 0.0128f
C9708 vdd.n9297 vss 0.02f
C9709 vdd.n9298 vss 0.00425f
C9710 vdd.n9299 vss 0.00413f
C9711 vdd.n9300 vss 0.00251f
C9712 vdd.n9301 vss 0.0471f
C9713 vdd.n9302 vss 0.00251f
C9714 vdd.n9303 vss 0.00517f
C9715 vdd.n9304 vss 0.00679f
C9716 vdd.n9305 vss 0.00324f
C9717 vdd.n9306 vss 0.00324f
C9718 vdd.n9307 vss 0.0132f
C9719 vdd.n9308 vss 0.0424f
C9720 vdd.n9309 vss 0.02f
C9721 vdd.n9310 vss 0.00425f
C9722 vdd.n9311 vss 0.0471f
C9723 vdd.n9313 vss 0.00425f
C9724 vdd.n9314 vss 0.00925f
C9725 vdd.n9315 vss 0.00679f
C9726 vdd.n9316 vss 0.00517f
C9727 vdd.n9317 vss 0.00251f
C9728 vdd.n9318 vss 0.0471f
C9729 vdd.n9319 vss 0.00251f
C9730 vdd.n9320 vss 0.0112f
C9731 vdd.n9321 vss 0.0128f
C9732 vdd.n9322 vss 0.123f
C9733 vdd.n9323 vss 0.0596f
C9734 vdd.n9324 vss 0.00324f
C9735 vdd.n9325 vss 0.0112f
C9736 vdd.n9326 vss 0.0128f
C9737 vdd.n9327 vss 0.00413f
C9738 vdd.n9328 vss 0.00413f
C9739 vdd.n9329 vss 0.0471f
C9740 vdd.n9330 vss 0.0471f
C9741 vdd.n9331 vss 0.00324f
C9742 vdd.n9332 vss 0.00413f
C9743 vdd.n9333 vss 0.00413f
C9744 vdd.n9334 vss 0.00679f
C9745 vdd.n9335 vss 0.00413f
C9746 vdd.n9336 vss 0.0471f
C9747 vdd.n9337 vss 0.00324f
C9748 vdd.n9339 vss 0.00925f
C9749 vdd.n9340 vss 0.0471f
C9750 vdd.n9341 vss 0.00425f
C9751 vdd.n9342 vss 0.0424f
C9752 vdd.n9343 vss 0.0132f
C9753 vdd.n9344 vss 0.00324f
C9754 vdd.n9345 vss 0.0128f
C9755 vdd.n9346 vss 0.02f
C9756 vdd.n9347 vss 0.00425f
C9757 vdd.n9348 vss 0.00413f
C9758 vdd.n9349 vss 0.00251f
C9759 vdd.n9350 vss 0.0471f
C9760 vdd.n9351 vss 0.00251f
C9761 vdd.n9352 vss 0.00517f
C9762 vdd.n9353 vss 0.00679f
C9763 vdd.n9354 vss 0.00324f
C9764 vdd.n9355 vss 0.00324f
C9765 vdd.n9356 vss 0.0132f
C9766 vdd.n9357 vss 0.0424f
C9767 vdd.n9358 vss 0.02f
C9768 vdd.n9359 vss 0.00425f
C9769 vdd.n9360 vss 0.0471f
C9770 vdd.n9362 vss 0.00425f
C9771 vdd.n9363 vss 0.00925f
C9772 vdd.n9364 vss 0.00679f
C9773 vdd.n9365 vss 0.00517f
C9774 vdd.n9366 vss 0.00251f
C9775 vdd.n9367 vss 0.0471f
C9776 vdd.n9368 vss 0.00251f
C9777 vdd.n9369 vss 0.0112f
C9778 vdd.n9370 vss 0.0128f
C9779 vdd.n9371 vss 0.0692f
C9780 vdd.n9372 vss 0.118f
C9781 vdd.n9373 vss 0.121f
C9782 vdd.n9374 vss 0.00324f
C9783 vdd.n9375 vss 0.0112f
C9784 vdd.n9376 vss 0.0128f
C9785 vdd.n9377 vss 0.00413f
C9786 vdd.n9378 vss 0.00413f
C9787 vdd.n9379 vss 0.0471f
C9788 vdd.n9380 vss 0.0471f
C9789 vdd.n9381 vss 0.00324f
C9790 vdd.n9382 vss 0.00413f
C9791 vdd.n9383 vss 0.00413f
C9792 vdd.n9384 vss 0.00679f
C9793 vdd.n9385 vss 0.00413f
C9794 vdd.n9386 vss 0.0471f
C9795 vdd.n9387 vss 0.00324f
C9796 vdd.n9389 vss 0.00925f
C9797 vdd.n9390 vss 0.0471f
C9798 vdd.n9391 vss 0.00425f
C9799 vdd.n9392 vss 0.0424f
C9800 vdd.n9393 vss 0.0132f
C9801 vdd.n9394 vss 0.00324f
C9802 vdd.n9395 vss 0.0128f
C9803 vdd.n9396 vss 0.02f
C9804 vdd.n9397 vss 0.00425f
C9805 vdd.n9398 vss 0.00413f
C9806 vdd.n9399 vss 0.00251f
C9807 vdd.n9400 vss 0.0471f
C9808 vdd.n9401 vss 0.00251f
C9809 vdd.n9402 vss 0.00517f
C9810 vdd.n9403 vss 0.00679f
C9811 vdd.n9404 vss 0.00324f
C9812 vdd.n9405 vss 0.00324f
C9813 vdd.n9406 vss 0.0132f
C9814 vdd.n9407 vss 0.0424f
C9815 vdd.n9408 vss 0.02f
C9816 vdd.n9409 vss 0.00425f
C9817 vdd.n9410 vss 0.0471f
C9818 vdd.n9412 vss 0.00425f
C9819 vdd.n9413 vss 0.00925f
C9820 vdd.n9414 vss 0.00679f
C9821 vdd.n9415 vss 0.00517f
C9822 vdd.n9416 vss 0.00251f
C9823 vdd.n9417 vss 0.0471f
C9824 vdd.n9418 vss 0.00251f
C9825 vdd.n9419 vss 0.0112f
C9826 vdd.n9420 vss 0.098f
C9827 vdd.n9421 vss 0.0596f
C9828 vdd.n9422 vss 0.00324f
C9829 vdd.n9423 vss 0.0112f
C9830 vdd.n9424 vss 0.0128f
C9831 vdd.n9425 vss 0.00413f
C9832 vdd.n9426 vss 0.00413f
C9833 vdd.n9427 vss 0.0471f
C9834 vdd.n9428 vss 0.0471f
C9835 vdd.n9429 vss 0.00324f
C9836 vdd.n9430 vss 0.00413f
C9837 vdd.n9431 vss 0.00413f
C9838 vdd.n9432 vss 0.00679f
C9839 vdd.n9433 vss 0.00413f
C9840 vdd.n9434 vss 0.0471f
C9841 vdd.n9435 vss 0.00324f
C9842 vdd.n9437 vss 0.00925f
C9843 vdd.n9438 vss 0.0471f
C9844 vdd.n9439 vss 0.00425f
C9845 vdd.n9440 vss 0.0424f
C9846 vdd.n9441 vss 0.0132f
C9847 vdd.n9442 vss 0.00324f
C9848 vdd.n9443 vss 0.0128f
C9849 vdd.n9444 vss 0.02f
C9850 vdd.n9445 vss 0.00425f
C9851 vdd.n9446 vss 0.00413f
C9852 vdd.n9447 vss 0.00251f
C9853 vdd.n9448 vss 0.0471f
C9854 vdd.n9449 vss 0.00251f
C9855 vdd.n9450 vss 0.00517f
C9856 vdd.n9451 vss 0.00679f
C9857 vdd.n9452 vss 0.00324f
C9858 vdd.n9453 vss 0.00324f
C9859 vdd.n9454 vss 0.0132f
C9860 vdd.n9455 vss 0.0424f
C9861 vdd.n9456 vss 0.02f
C9862 vdd.n9457 vss 0.00425f
C9863 vdd.n9458 vss 0.0471f
C9864 vdd.n9460 vss 0.00425f
C9865 vdd.n9461 vss 0.00925f
C9866 vdd.n9462 vss 0.00679f
C9867 vdd.n9463 vss 0.00517f
C9868 vdd.n9464 vss 0.00251f
C9869 vdd.n9465 vss 0.0471f
C9870 vdd.n9466 vss 0.00251f
C9871 vdd.n9467 vss 0.0112f
C9872 vdd.n9468 vss 0.0128f
C9873 vdd.n9469 vss 0.0692f
C9874 vdd.n9470 vss 0.118f
C9875 vdd.n9471 vss 0.0951f
C9876 vdd.n9472 vss 0.00324f
C9877 vdd.n9473 vss 0.0112f
C9878 vdd.n9474 vss 0.0128f
C9879 vdd.n9475 vss 0.00413f
C9880 vdd.n9476 vss 0.00413f
C9881 vdd.n9477 vss 0.0471f
C9882 vdd.n9478 vss 0.0471f
C9883 vdd.n9479 vss 0.00324f
C9884 vdd.n9480 vss 0.00413f
C9885 vdd.n9481 vss 0.00413f
C9886 vdd.n9482 vss 0.00679f
C9887 vdd.n9483 vss 0.00413f
C9888 vdd.n9484 vss 0.0471f
C9889 vdd.n9485 vss 0.00324f
C9890 vdd.n9487 vss 0.00925f
C9891 vdd.n9488 vss 0.0471f
C9892 vdd.n9489 vss 0.00425f
C9893 vdd.n9490 vss 0.0424f
C9894 vdd.n9491 vss 0.0132f
C9895 vdd.n9492 vss 0.00324f
C9896 vdd.n9493 vss 0.0128f
C9897 vdd.n9494 vss 0.02f
C9898 vdd.n9495 vss 0.00425f
C9899 vdd.n9496 vss 0.00413f
C9900 vdd.n9497 vss 0.00251f
C9901 vdd.n9498 vss 0.0471f
C9902 vdd.n9499 vss 0.00251f
C9903 vdd.n9500 vss 0.00517f
C9904 vdd.n9501 vss 0.00679f
C9905 vdd.n9502 vss 0.00324f
C9906 vdd.n9503 vss 0.00324f
C9907 vdd.n9504 vss 0.0132f
C9908 vdd.n9505 vss 0.0424f
C9909 vdd.n9506 vss 0.02f
C9910 vdd.n9507 vss 0.00425f
C9911 vdd.n9508 vss 0.0471f
C9912 vdd.n9510 vss 0.00425f
C9913 vdd.n9511 vss 0.00925f
C9914 vdd.n9512 vss 0.00679f
C9915 vdd.n9513 vss 0.00517f
C9916 vdd.n9514 vss 0.00251f
C9917 vdd.n9515 vss 0.0471f
C9918 vdd.n9516 vss 0.00251f
C9919 vdd.n9517 vss 0.0112f
C9920 vdd.n9518 vss 0.0128f
C9921 vdd.n9519 vss 0.146f
C9922 vdd.n9520 vss 0.00324f
C9923 vdd.n9521 vss 0.0112f
C9924 vdd.n9522 vss 0.0128f
C9925 vdd.n9523 vss 0.00413f
C9926 vdd.n9524 vss 0.00413f
C9927 vdd.n9525 vss 0.0471f
C9928 vdd.n9526 vss 0.0471f
C9929 vdd.n9527 vss 0.00324f
C9930 vdd.n9528 vss 0.00413f
C9931 vdd.n9529 vss 0.00413f
C9932 vdd.n9530 vss 0.00679f
C9933 vdd.n9531 vss 0.00413f
C9934 vdd.n9532 vss 0.0471f
C9935 vdd.n9533 vss 0.00324f
C9936 vdd.n9535 vss 0.00925f
C9937 vdd.n9536 vss 0.0471f
C9938 vdd.n9537 vss 0.00425f
C9939 vdd.n9538 vss 0.0424f
C9940 vdd.n9539 vss 0.0132f
C9941 vdd.n9540 vss 0.00324f
C9942 vdd.n9541 vss 0.0128f
C9943 vdd.n9542 vss 0.02f
C9944 vdd.n9543 vss 0.00425f
C9945 vdd.n9544 vss 0.00413f
C9946 vdd.n9545 vss 0.00251f
C9947 vdd.n9546 vss 0.0471f
C9948 vdd.n9547 vss 0.00251f
C9949 vdd.n9548 vss 0.00517f
C9950 vdd.n9549 vss 0.00679f
C9951 vdd.n9550 vss 0.00324f
C9952 vdd.n9551 vss 0.00324f
C9953 vdd.n9552 vss 0.0132f
C9954 vdd.n9553 vss 0.0424f
C9955 vdd.n9554 vss 0.02f
C9956 vdd.n9555 vss 0.00425f
C9957 vdd.n9556 vss 0.0471f
C9958 vdd.n9558 vss 0.00425f
C9959 vdd.n9559 vss 0.00925f
C9960 vdd.n9560 vss 0.00679f
C9961 vdd.n9561 vss 0.00517f
C9962 vdd.n9562 vss 0.00251f
C9963 vdd.n9563 vss 0.0471f
C9964 vdd.n9564 vss 0.00251f
C9965 vdd.n9565 vss 0.0112f
C9966 vdd.n9566 vss 0.0128f
C9967 vdd.n9567 vss 0.146f
C9968 vdd.n9568 vss 0.0596f
C9969 vdd.n9569 vss 0.00324f
C9970 vdd.n9570 vss 0.0112f
C9971 vdd.n9571 vss 0.0128f
C9972 vdd.n9572 vss 0.00413f
C9973 vdd.n9573 vss 0.00413f
C9974 vdd.n9574 vss 0.0471f
C9975 vdd.n9575 vss 0.0471f
C9976 vdd.n9576 vss 0.00324f
C9977 vdd.n9577 vss 0.00413f
C9978 vdd.n9578 vss 0.00413f
C9979 vdd.n9579 vss 0.00679f
C9980 vdd.n9580 vss 0.00413f
C9981 vdd.n9581 vss 0.0471f
C9982 vdd.n9582 vss 0.00324f
C9983 vdd.n9584 vss 0.00925f
C9984 vdd.n9585 vss 0.0471f
C9985 vdd.n9586 vss 0.00425f
C9986 vdd.n9587 vss 0.0424f
C9987 vdd.n9588 vss 0.0132f
C9988 vdd.n9589 vss 0.00324f
C9989 vdd.n9590 vss 0.0128f
C9990 vdd.n9591 vss 0.02f
C9991 vdd.n9592 vss 0.00425f
C9992 vdd.n9593 vss 0.00413f
C9993 vdd.n9594 vss 0.00251f
C9994 vdd.n9595 vss 0.0471f
C9995 vdd.n9596 vss 0.00251f
C9996 vdd.n9597 vss 0.00517f
C9997 vdd.n9598 vss 0.00679f
C9998 vdd.n9599 vss 0.00324f
C9999 vdd.n9600 vss 0.00324f
C10000 vdd.n9601 vss 0.0132f
C10001 vdd.n9602 vss 0.0424f
C10002 vdd.n9603 vss 0.02f
C10003 vdd.n9604 vss 0.00425f
C10004 vdd.n9605 vss 0.0471f
C10005 vdd.n9607 vss 0.00425f
C10006 vdd.n9608 vss 0.00925f
C10007 vdd.n9609 vss 0.00679f
C10008 vdd.n9610 vss 0.00517f
C10009 vdd.n9611 vss 0.00251f
C10010 vdd.n9612 vss 0.0471f
C10011 vdd.n9613 vss 0.00251f
C10012 vdd.n9614 vss 0.0112f
C10013 vdd.n9615 vss 0.0128f
C10014 vdd.n9616 vss 0.0692f
C10015 vdd.n9617 vss 0.118f
C10016 vdd.n9618 vss 0.121f
C10017 vdd.n9619 vss 0.00324f
C10018 vdd.n9620 vss 0.0112f
C10019 vdd.n9621 vss 0.0128f
C10020 vdd.n9622 vss 0.00413f
C10021 vdd.n9623 vss 0.00413f
C10022 vdd.n9624 vss 0.0471f
C10023 vdd.n9625 vss 0.0471f
C10024 vdd.n9626 vss 0.00324f
C10025 vdd.n9627 vss 0.00413f
C10026 vdd.n9628 vss 0.00413f
C10027 vdd.n9629 vss 0.00679f
C10028 vdd.n9630 vss 0.00413f
C10029 vdd.n9631 vss 0.0471f
C10030 vdd.n9632 vss 0.00324f
C10031 vdd.n9634 vss 0.00925f
C10032 vdd.n9635 vss 0.0471f
C10033 vdd.n9636 vss 0.00425f
C10034 vdd.n9637 vss 0.0424f
C10035 vdd.n9638 vss 0.0132f
C10036 vdd.n9639 vss 0.00324f
C10037 vdd.n9640 vss 0.0128f
C10038 vdd.n9641 vss 0.02f
C10039 vdd.n9642 vss 0.00425f
C10040 vdd.n9643 vss 0.00413f
C10041 vdd.n9644 vss 0.00251f
C10042 vdd.n9645 vss 0.0471f
C10043 vdd.n9646 vss 0.00251f
C10044 vdd.n9647 vss 0.00517f
C10045 vdd.n9648 vss 0.00679f
C10046 vdd.n9649 vss 0.00324f
C10047 vdd.n9650 vss 0.00324f
C10048 vdd.n9651 vss 0.0132f
C10049 vdd.n9652 vss 0.0424f
C10050 vdd.n9653 vss 0.02f
C10051 vdd.n9654 vss 0.00425f
C10052 vdd.n9655 vss 0.0471f
C10053 vdd.n9657 vss 0.00425f
C10054 vdd.n9658 vss 0.00925f
C10055 vdd.n9659 vss 0.00679f
C10056 vdd.n9660 vss 0.00517f
C10057 vdd.n9661 vss 0.00251f
C10058 vdd.n9662 vss 0.0471f
C10059 vdd.n9663 vss 0.00251f
C10060 vdd.n9664 vss 0.0112f
C10061 vdd.n9665 vss 0.098f
C10062 vdd.n9666 vss 0.0596f
C10063 vdd.n9667 vss 0.00324f
C10064 vdd.n9668 vss 0.0112f
C10065 vdd.n9669 vss 0.0128f
C10066 vdd.n9670 vss 0.00413f
C10067 vdd.n9671 vss 0.00413f
C10068 vdd.n9672 vss 0.0471f
C10069 vdd.n9673 vss 0.0471f
C10070 vdd.n9674 vss 0.00324f
C10071 vdd.n9675 vss 0.00413f
C10072 vdd.n9676 vss 0.00413f
C10073 vdd.n9677 vss 0.00679f
C10074 vdd.n9678 vss 0.00413f
C10075 vdd.n9679 vss 0.0471f
C10076 vdd.n9680 vss 0.00324f
C10077 vdd.n9682 vss 0.00925f
C10078 vdd.n9683 vss 0.0471f
C10079 vdd.n9684 vss 0.00425f
C10080 vdd.n9685 vss 0.0424f
C10081 vdd.n9686 vss 0.0132f
C10082 vdd.n9687 vss 0.00324f
C10083 vdd.n9688 vss 0.0128f
C10084 vdd.n9689 vss 0.02f
C10085 vdd.n9690 vss 0.00425f
C10086 vdd.n9691 vss 0.00413f
C10087 vdd.n9692 vss 0.00251f
C10088 vdd.n9693 vss 0.0471f
C10089 vdd.n9694 vss 0.00251f
C10090 vdd.n9695 vss 0.00517f
C10091 vdd.n9696 vss 0.00679f
C10092 vdd.n9697 vss 0.00324f
C10093 vdd.n9698 vss 0.00324f
C10094 vdd.n9699 vss 0.0132f
C10095 vdd.n9700 vss 0.0424f
C10096 vdd.n9701 vss 0.02f
C10097 vdd.n9702 vss 0.00425f
C10098 vdd.n9703 vss 0.0471f
C10099 vdd.n9705 vss 0.00425f
C10100 vdd.n9706 vss 0.00925f
C10101 vdd.n9707 vss 0.00679f
C10102 vdd.n9708 vss 0.00517f
C10103 vdd.n9709 vss 0.00251f
C10104 vdd.n9710 vss 0.0471f
C10105 vdd.n9711 vss 0.00251f
C10106 vdd.n9712 vss 0.0112f
C10107 vdd.n9713 vss 0.0128f
C10108 vdd.n9714 vss 0.0692f
C10109 vdd.n9715 vss 0.0912f
C10110 vdd.n9716 vss 0.0824f
C10111 vdd.n9717 vss 0.059f
C10112 vdd.n9718 vss 0.00324f
C10113 vdd.n9719 vss 0.0112f
C10114 vdd.n9720 vss 0.0128f
C10115 vdd.n9721 vss 0.00413f
C10116 vdd.n9722 vss 0.00413f
C10117 vdd.n9723 vss 0.0471f
C10118 vdd.n9724 vss 0.0471f
C10119 vdd.n9725 vss 0.00324f
C10120 vdd.n9726 vss 0.00413f
C10121 vdd.n9727 vss 0.00413f
C10122 vdd.n9728 vss 0.00679f
C10123 vdd.n9729 vss 0.00413f
C10124 vdd.n9730 vss 0.0471f
C10125 vdd.n9731 vss 0.00324f
C10126 vdd.n9733 vss 0.00925f
C10127 vdd.n9734 vss 0.0471f
C10128 vdd.n9735 vss 0.00425f
C10129 vdd.n9736 vss 0.0424f
C10130 vdd.n9737 vss 0.0132f
C10131 vdd.n9738 vss 0.00324f
C10132 vdd.n9739 vss 0.0128f
C10133 vdd.n9740 vss 0.02f
C10134 vdd.n9741 vss 0.00425f
C10135 vdd.n9742 vss 0.00413f
C10136 vdd.n9743 vss 0.00251f
C10137 vdd.n9744 vss 0.0471f
C10138 vdd.n9745 vss 0.00251f
C10139 vdd.n9746 vss 0.00517f
C10140 vdd.n9747 vss 0.00679f
C10141 vdd.n9748 vss 0.00324f
C10142 vdd.n9749 vss 0.00324f
C10143 vdd.n9750 vss 0.0132f
C10144 vdd.n9751 vss 0.0424f
C10145 vdd.n9752 vss 0.02f
C10146 vdd.n9753 vss 0.00425f
C10147 vdd.n9754 vss 0.0471f
C10148 vdd.n9756 vss 0.00425f
C10149 vdd.n9757 vss 0.00925f
C10150 vdd.n9758 vss 0.00679f
C10151 vdd.n9759 vss 0.00517f
C10152 vdd.n9760 vss 0.00251f
C10153 vdd.n9761 vss 0.0471f
C10154 vdd.n9762 vss 0.00251f
C10155 vdd.n9763 vss 0.0112f
C10156 vdd.n9764 vss 0.0128f
C10157 vdd.n9765 vss 0.146f
C10158 vdd.n9766 vss 0.00324f
C10159 vdd.n9767 vss 0.0112f
C10160 vdd.n9768 vss 0.0128f
C10161 vdd.n9769 vss 0.00413f
C10162 vdd.n9770 vss 0.00413f
C10163 vdd.n9771 vss 0.0471f
C10164 vdd.n9772 vss 0.0471f
C10165 vdd.n9773 vss 0.00324f
C10166 vdd.n9774 vss 0.00413f
C10167 vdd.n9775 vss 0.00413f
C10168 vdd.n9776 vss 0.00679f
C10169 vdd.n9777 vss 0.00413f
C10170 vdd.n9778 vss 0.0471f
C10171 vdd.n9779 vss 0.00324f
C10172 vdd.n9781 vss 0.00925f
C10173 vdd.n9782 vss 0.0471f
C10174 vdd.n9783 vss 0.00425f
C10175 vdd.n9784 vss 0.0424f
C10176 vdd.n9785 vss 0.0132f
C10177 vdd.n9786 vss 0.00324f
C10178 vdd.n9787 vss 0.0128f
C10179 vdd.n9788 vss 0.02f
C10180 vdd.n9789 vss 0.00425f
C10181 vdd.n9790 vss 0.00413f
C10182 vdd.n9791 vss 0.00251f
C10183 vdd.n9792 vss 0.0471f
C10184 vdd.n9793 vss 0.00251f
C10185 vdd.n9794 vss 0.00517f
C10186 vdd.n9795 vss 0.00679f
C10187 vdd.n9796 vss 0.00324f
C10188 vdd.n9797 vss 0.00324f
C10189 vdd.n9798 vss 0.0132f
C10190 vdd.n9799 vss 0.0424f
C10191 vdd.n9800 vss 0.02f
C10192 vdd.n9801 vss 0.00425f
C10193 vdd.n9802 vss 0.0471f
C10194 vdd.n9804 vss 0.00425f
C10195 vdd.n9805 vss 0.00925f
C10196 vdd.n9806 vss 0.00679f
C10197 vdd.n9807 vss 0.00517f
C10198 vdd.n9808 vss 0.00251f
C10199 vdd.n9809 vss 0.0471f
C10200 vdd.n9810 vss 0.00251f
C10201 vdd.n9811 vss 0.0112f
C10202 vdd.n9812 vss 0.0128f
C10203 vdd.n9813 vss 0.146f
C10204 vdd.n9814 vss 0.0596f
C10205 vdd.n9815 vss 0.00324f
C10206 vdd.n9816 vss 0.0112f
C10207 vdd.n9817 vss 0.0128f
C10208 vdd.n9818 vss 0.00413f
C10209 vdd.n9819 vss 0.00413f
C10210 vdd.n9820 vss 0.0471f
C10211 vdd.n9821 vss 0.0471f
C10212 vdd.n9822 vss 0.00324f
C10213 vdd.n9823 vss 0.00413f
C10214 vdd.n9824 vss 0.00413f
C10215 vdd.n9825 vss 0.00679f
C10216 vdd.n9826 vss 0.00413f
C10217 vdd.n9827 vss 0.0471f
C10218 vdd.n9828 vss 0.00324f
C10219 vdd.n9830 vss 0.00925f
C10220 vdd.n9831 vss 0.0471f
C10221 vdd.n9832 vss 0.00425f
C10222 vdd.n9833 vss 0.0424f
C10223 vdd.n9834 vss 0.0132f
C10224 vdd.n9835 vss 0.00324f
C10225 vdd.n9836 vss 0.0128f
C10226 vdd.n9837 vss 0.02f
C10227 vdd.n9838 vss 0.00425f
C10228 vdd.n9839 vss 0.00413f
C10229 vdd.n9840 vss 0.00251f
C10230 vdd.n9841 vss 0.0471f
C10231 vdd.n9842 vss 0.00251f
C10232 vdd.n9843 vss 0.00517f
C10233 vdd.n9844 vss 0.00679f
C10234 vdd.n9845 vss 0.00324f
C10235 vdd.n9846 vss 0.00324f
C10236 vdd.n9847 vss 0.0132f
C10237 vdd.n9848 vss 0.0424f
C10238 vdd.n9849 vss 0.02f
C10239 vdd.n9850 vss 0.00425f
C10240 vdd.n9851 vss 0.0471f
C10241 vdd.n9853 vss 0.00425f
C10242 vdd.n9854 vss 0.00925f
C10243 vdd.n9855 vss 0.00679f
C10244 vdd.n9856 vss 0.00517f
C10245 vdd.n9857 vss 0.00251f
C10246 vdd.n9858 vss 0.0471f
C10247 vdd.n9859 vss 0.00251f
C10248 vdd.n9860 vss 0.0112f
C10249 vdd.n9861 vss 0.0128f
C10250 vdd.n9862 vss 0.0692f
C10251 vdd.n9863 vss 0.118f
C10252 vdd.n9864 vss 0.121f
C10253 vdd.n9865 vss 0.00324f
C10254 vdd.n9866 vss 0.0112f
C10255 vdd.n9867 vss 0.0128f
C10256 vdd.n9868 vss 0.00413f
C10257 vdd.n9869 vss 0.00413f
C10258 vdd.n9870 vss 0.0471f
C10259 vdd.n9871 vss 0.0471f
C10260 vdd.n9872 vss 0.00324f
C10261 vdd.n9873 vss 0.00413f
C10262 vdd.n9874 vss 0.00413f
C10263 vdd.n9875 vss 0.00679f
C10264 vdd.n9876 vss 0.00413f
C10265 vdd.n9877 vss 0.0471f
C10266 vdd.n9878 vss 0.00324f
C10267 vdd.n9880 vss 0.00925f
C10268 vdd.n9881 vss 0.0471f
C10269 vdd.n9882 vss 0.00425f
C10270 vdd.n9883 vss 0.0424f
C10271 vdd.n9884 vss 0.0132f
C10272 vdd.n9885 vss 0.00324f
C10273 vdd.n9886 vss 0.0128f
C10274 vdd.n9887 vss 0.02f
C10275 vdd.n9888 vss 0.00425f
C10276 vdd.n9889 vss 0.00413f
C10277 vdd.n9890 vss 0.00251f
C10278 vdd.n9891 vss 0.0471f
C10279 vdd.n9892 vss 0.00251f
C10280 vdd.n9893 vss 0.00517f
C10281 vdd.n9894 vss 0.00679f
C10282 vdd.n9895 vss 0.00324f
C10283 vdd.n9896 vss 0.00324f
C10284 vdd.n9897 vss 0.0132f
C10285 vdd.n9898 vss 0.0424f
C10286 vdd.n9899 vss 0.02f
C10287 vdd.n9900 vss 0.00425f
C10288 vdd.n9901 vss 0.0471f
C10289 vdd.n9903 vss 0.00425f
C10290 vdd.n9904 vss 0.00925f
C10291 vdd.n9905 vss 0.00679f
C10292 vdd.n9906 vss 0.00517f
C10293 vdd.n9907 vss 0.00251f
C10294 vdd.n9908 vss 0.0471f
C10295 vdd.n9909 vss 0.00251f
C10296 vdd.n9910 vss 0.0112f
C10297 vdd.n9911 vss 0.098f
C10298 vdd.n9912 vss 0.0596f
C10299 vdd.n9913 vss 0.00324f
C10300 vdd.n9914 vss 0.0112f
C10301 vdd.n9915 vss 0.0128f
C10302 vdd.n9916 vss 0.00413f
C10303 vdd.n9917 vss 0.00413f
C10304 vdd.n9918 vss 0.0471f
C10305 vdd.n9919 vss 0.0471f
C10306 vdd.n9920 vss 0.00324f
C10307 vdd.n9921 vss 0.00413f
C10308 vdd.n9922 vss 0.00413f
C10309 vdd.n9923 vss 0.00679f
C10310 vdd.n9924 vss 0.00413f
C10311 vdd.n9925 vss 0.0471f
C10312 vdd.n9926 vss 0.00324f
C10313 vdd.n9928 vss 0.00925f
C10314 vdd.n9929 vss 0.0471f
C10315 vdd.n9930 vss 0.00425f
C10316 vdd.n9931 vss 0.0424f
C10317 vdd.n9932 vss 0.0132f
C10318 vdd.n9933 vss 0.00324f
C10319 vdd.n9934 vss 0.0128f
C10320 vdd.n9935 vss 0.02f
C10321 vdd.n9936 vss 0.00425f
C10322 vdd.n9937 vss 0.00413f
C10323 vdd.n9938 vss 0.00251f
C10324 vdd.n9939 vss 0.0471f
C10325 vdd.n9940 vss 0.00251f
C10326 vdd.n9941 vss 0.00517f
C10327 vdd.n9942 vss 0.00679f
C10328 vdd.n9943 vss 0.00324f
C10329 vdd.n9944 vss 0.00324f
C10330 vdd.n9945 vss 0.0132f
C10331 vdd.n9946 vss 0.0424f
C10332 vdd.n9947 vss 0.02f
C10333 vdd.n9948 vss 0.00425f
C10334 vdd.n9949 vss 0.0471f
C10335 vdd.n9951 vss 0.00425f
C10336 vdd.n9952 vss 0.00925f
C10337 vdd.n9953 vss 0.00679f
C10338 vdd.n9954 vss 0.00517f
C10339 vdd.n9955 vss 0.00251f
C10340 vdd.n9956 vss 0.0471f
C10341 vdd.n9957 vss 0.00251f
C10342 vdd.n9958 vss 0.0112f
C10343 vdd.n9959 vss 0.0128f
C10344 vdd.n9960 vss 0.0692f
C10345 vdd.n9961 vss 0.121f
C10346 vdd.n9962 vss 0.291f
C10347 vdd.n9963 vss 0.227f
C10348 vdd.n9964 vss 0.00324f
C10349 vdd.n9965 vss 0.0112f
C10350 vdd.n9966 vss 0.0128f
C10351 vdd.n9967 vss 0.00413f
C10352 vdd.n9968 vss 0.00413f
C10353 vdd.n9969 vss 0.0471f
C10354 vdd.n9970 vss 0.0471f
C10355 vdd.n9971 vss 0.00324f
C10356 vdd.n9972 vss 0.00413f
C10357 vdd.n9973 vss 0.00413f
C10358 vdd.n9974 vss 0.00679f
C10359 vdd.n9975 vss 0.00413f
C10360 vdd.n9976 vss 0.0471f
C10361 vdd.n9977 vss 0.00324f
C10362 vdd.n9979 vss 0.00925f
C10363 vdd.n9980 vss 0.0471f
C10364 vdd.n9981 vss 0.00425f
C10365 vdd.n9982 vss 0.0424f
C10366 vdd.n9983 vss 0.0132f
C10367 vdd.n9984 vss 0.00324f
C10368 vdd.n9985 vss 0.0128f
C10369 vdd.n9986 vss 0.02f
C10370 vdd.n9987 vss 0.00425f
C10371 vdd.n9988 vss 0.00413f
C10372 vdd.n9989 vss 0.00251f
C10373 vdd.n9990 vss 0.0471f
C10374 vdd.n9991 vss 0.00251f
C10375 vdd.n9992 vss 0.00517f
C10376 vdd.n9993 vss 0.00679f
C10377 vdd.n9994 vss 0.00324f
C10378 vdd.n9995 vss 0.00324f
C10379 vdd.n9996 vss 0.0132f
C10380 vdd.n9997 vss 0.0424f
C10381 vdd.n9998 vss 0.02f
C10382 vdd.n9999 vss 0.00425f
C10383 vdd.n10000 vss 0.0471f
C10384 vdd.n10002 vss 0.00425f
C10385 vdd.n10003 vss 0.00925f
C10386 vdd.n10004 vss 0.00679f
C10387 vdd.n10005 vss 0.00517f
C10388 vdd.n10006 vss 0.00251f
C10389 vdd.n10007 vss 0.0471f
C10390 vdd.n10008 vss 0.00251f
C10391 vdd.n10009 vss 0.0112f
C10392 vdd.n10010 vss 0.0128f
C10393 vdd.n10011 vss 0.18f
C10394 vdd.n10012 vss 0.00324f
C10395 vdd.n10013 vss 0.0112f
C10396 vdd.n10014 vss 0.0128f
C10397 vdd.n10015 vss 0.00413f
C10398 vdd.n10016 vss 0.00413f
C10399 vdd.n10017 vss 0.0471f
C10400 vdd.n10018 vss 0.0471f
C10401 vdd.n10019 vss 0.00324f
C10402 vdd.n10020 vss 0.00413f
C10403 vdd.n10021 vss 0.00413f
C10404 vdd.n10022 vss 0.00679f
C10405 vdd.n10023 vss 0.00413f
C10406 vdd.n10024 vss 0.0471f
C10407 vdd.n10025 vss 0.00324f
C10408 vdd.n10027 vss 0.00925f
C10409 vdd.n10028 vss 0.0471f
C10410 vdd.n10029 vss 0.00425f
C10411 vdd.n10030 vss 0.0424f
C10412 vdd.n10031 vss 0.0132f
C10413 vdd.n10032 vss 0.00324f
C10414 vdd.n10033 vss 0.0128f
C10415 vdd.n10034 vss 0.02f
C10416 vdd.n10035 vss 0.00425f
C10417 vdd.n10036 vss 0.00413f
C10418 vdd.n10037 vss 0.00251f
C10419 vdd.n10038 vss 0.0471f
C10420 vdd.n10039 vss 0.00251f
C10421 vdd.n10040 vss 0.00517f
C10422 vdd.n10041 vss 0.00679f
C10423 vdd.n10042 vss 0.00324f
C10424 vdd.n10043 vss 0.00324f
C10425 vdd.n10044 vss 0.0132f
C10426 vdd.n10045 vss 0.0424f
C10427 vdd.n10046 vss 0.02f
C10428 vdd.n10047 vss 0.00425f
C10429 vdd.n10048 vss 0.0471f
C10430 vdd.n10050 vss 0.00425f
C10431 vdd.n10051 vss 0.00925f
C10432 vdd.n10052 vss 0.00679f
C10433 vdd.n10053 vss 0.00517f
C10434 vdd.n10054 vss 0.00251f
C10435 vdd.n10055 vss 0.0471f
C10436 vdd.n10056 vss 0.00251f
C10437 vdd.n10057 vss 0.0112f
C10438 vdd.n10058 vss 0.0128f
C10439 vdd.n10059 vss 0.248f
C10440 vdd.n10060 vss 0.00324f
C10441 vdd.n10061 vss 0.0112f
C10442 vdd.n10062 vss 0.0128f
C10443 vdd.n10063 vss 0.00413f
C10444 vdd.n10064 vss 0.00413f
C10445 vdd.n10065 vss 0.0471f
C10446 vdd.n10066 vss 0.0471f
C10447 vdd.n10067 vss 0.00324f
C10448 vdd.n10068 vss 0.00413f
C10449 vdd.n10069 vss 0.00413f
C10450 vdd.n10070 vss 0.00679f
C10451 vdd.n10071 vss 0.00413f
C10452 vdd.n10072 vss 0.0471f
C10453 vdd.n10073 vss 0.00324f
C10454 vdd.n10075 vss 0.00925f
C10455 vdd.n10076 vss 0.0471f
C10456 vdd.n10077 vss 0.00425f
C10457 vdd.n10078 vss 0.0424f
C10458 vdd.n10079 vss 0.0132f
C10459 vdd.n10080 vss 0.00324f
C10460 vdd.n10081 vss 0.0128f
C10461 vdd.n10082 vss 0.02f
C10462 vdd.n10083 vss 0.00425f
C10463 vdd.n10084 vss 0.00413f
C10464 vdd.n10085 vss 0.00251f
C10465 vdd.n10086 vss 0.0471f
C10466 vdd.n10087 vss 0.00251f
C10467 vdd.n10088 vss 0.00517f
C10468 vdd.n10089 vss 0.00679f
C10469 vdd.n10090 vss 0.00324f
C10470 vdd.n10091 vss 0.00324f
C10471 vdd.n10092 vss 0.0132f
C10472 vdd.n10093 vss 0.0424f
C10473 vdd.n10094 vss 0.02f
C10474 vdd.n10095 vss 0.00425f
C10475 vdd.n10096 vss 0.0471f
C10476 vdd.n10098 vss 0.00425f
C10477 vdd.n10099 vss 0.00925f
C10478 vdd.n10100 vss 0.00679f
C10479 vdd.n10101 vss 0.00517f
C10480 vdd.n10102 vss 0.00251f
C10481 vdd.n10103 vss 0.0471f
C10482 vdd.n10104 vss 0.00251f
C10483 vdd.n10105 vss 0.0112f
C10484 vdd.n10106 vss 0.0128f
C10485 vdd.n10107 vss 0.0692f
C10486 vdd.n10108 vss 0.00324f
C10487 vdd.n10109 vss 0.0112f
C10488 vdd.n10110 vss 0.0128f
C10489 vdd.n10111 vss 0.00413f
C10490 vdd.n10112 vss 0.00413f
C10491 vdd.n10113 vss 0.0471f
C10492 vdd.n10114 vss 0.0471f
C10493 vdd.n10115 vss 0.00324f
C10494 vdd.n10116 vss 0.00413f
C10495 vdd.n10117 vss 0.00413f
C10496 vdd.n10118 vss 0.00679f
C10497 vdd.n10119 vss 0.00413f
C10498 vdd.n10120 vss 0.0471f
C10499 vdd.n10121 vss 0.00324f
C10500 vdd.n10123 vss 0.00925f
C10501 vdd.n10124 vss 0.0471f
C10502 vdd.n10125 vss 0.00425f
C10503 vdd.n10126 vss 0.0424f
C10504 vdd.n10127 vss 0.0132f
C10505 vdd.n10128 vss 0.00324f
C10506 vdd.n10129 vss 0.0128f
C10507 vdd.n10130 vss 0.02f
C10508 vdd.n10131 vss 0.00425f
C10509 vdd.n10132 vss 0.00413f
C10510 vdd.n10133 vss 0.00251f
C10511 vdd.n10134 vss 0.0471f
C10512 vdd.n10135 vss 0.00251f
C10513 vdd.n10136 vss 0.00517f
C10514 vdd.n10137 vss 0.00679f
C10515 vdd.n10138 vss 0.00324f
C10516 vdd.n10139 vss 0.00324f
C10517 vdd.n10140 vss 0.0132f
C10518 vdd.n10141 vss 0.0424f
C10519 vdd.n10142 vss 0.02f
C10520 vdd.n10143 vss 0.00425f
C10521 vdd.n10144 vss 0.0471f
C10522 vdd.n10146 vss 0.00425f
C10523 vdd.n10147 vss 0.00925f
C10524 vdd.n10148 vss 0.00679f
C10525 vdd.n10149 vss 0.00517f
C10526 vdd.n10150 vss 0.00251f
C10527 vdd.n10151 vss 0.0471f
C10528 vdd.n10152 vss 0.00251f
C10529 vdd.n10153 vss 0.0112f
C10530 vdd.n10154 vss 0.0128f
C10531 vdd.n10155 vss 0.0619f
C10532 vdd.n10156 vss 0.00335f
C10533 vdd.n10157 vss 0.0855f
C10534 vdd.n10158 vss 0.00991f
C10535 vdd.n10159 vss 0.0424f
C10536 vdd.n10160 vss 0.00679f
C10537 vdd.n10161 vss 0.00413f
C10538 vdd.n10162 vss 0.0471f
C10539 vdd.n10163 vss 0.00251f
C10540 vdd.n10164 vss 0.00679f
C10541 vdd.n10165 vss 0.00413f
C10542 vdd.n10166 vss 0.00413f
C10543 vdd.n10167 vss 0.0471f
C10544 vdd.n10168 vss 0.00251f
C10545 vdd.n10169 vss 0.00413f
C10546 vdd.n10170 vss 0.00324f
C10547 vdd.n10171 vss 0.0132f
C10548 vdd.n10172 vss 0.0424f
C10549 vdd.n10173 vss 0.00324f
C10550 vdd.n10174 vss 0.00413f
C10551 vdd.n10175 vss 0.00517f
C10552 vdd.n10176 vss 0.00679f
C10553 vdd.n10177 vss 0.00925f
C10554 vdd.n10178 vss 0.00425f
C10555 vdd.n10179 vss 0.0471f
C10556 vdd.n10181 vss 0.00425f
C10557 vdd.n10182 vss 0.02f
C10558 vdd.n10183 vss 0.0128f
C10559 vdd.n10184 vss 0.0105f
C10560 vdd.n10185 vss 0.00251f
C10561 vdd.n10186 vss 0.0471f
C10562 vdd.n10187 vss 0.00517f
C10563 vdd.n10188 vss 0.00251f
C10564 vdd.n10189 vss 0.0471f
C10565 vdd.n10190 vss 0.0471f
C10566 vdd.n10191 vss 0.00324f
C10567 vdd.n10192 vss 0.00324f
C10568 vdd.n10193 vss 0.00805f
C10569 vdd.n10194 vss 0.0112f
C10570 vdd.n10195 vss 0.0128f
C10571 vdd.n10196 vss 0.00324f
C10572 vdd.n10197 vss 0.00324f
C10573 vdd.n10198 vss 0.00413f
C10574 vdd.n10199 vss 0.00425f
C10575 vdd.n10200 vss 0.0471f
C10576 vdd.n10202 vss 0.00425f
C10577 vdd.n10203 vss 0.00925f
C10578 vdd.n10204 vss 0.0107f
C10579 vdd.n10205 vss 0.0126f
C10580 vdd.n10206 vss 0.0516f
C10581 vdd.n10207 vss 0.00163f
C10582 vdd.n10208 vss 0.00145f
C10583 vdd.n10209 vss 0.0271f
C10584 vdd.n10210 vss 0.00324f
C10585 vdd.n10211 vss 0.0112f
C10586 vdd.n10212 vss 0.0128f
C10587 vdd.n10213 vss 0.00413f
C10588 vdd.n10214 vss 0.00413f
C10589 vdd.n10215 vss 0.0471f
C10590 vdd.n10216 vss 0.0471f
C10591 vdd.n10217 vss 0.00324f
C10592 vdd.n10218 vss 0.00413f
C10593 vdd.n10219 vss 0.00413f
C10594 vdd.n10220 vss 0.00679f
C10595 vdd.n10221 vss 0.00413f
C10596 vdd.n10222 vss 0.0471f
C10597 vdd.n10223 vss 0.00324f
C10598 vdd.n10225 vss 0.00925f
C10599 vdd.n10226 vss 0.0471f
C10600 vdd.n10227 vss 0.00425f
C10601 vdd.n10228 vss 0.0424f
C10602 vdd.n10229 vss 0.0132f
C10603 vdd.n10230 vss 0.00324f
C10604 vdd.n10231 vss 0.0128f
C10605 vdd.n10232 vss 0.02f
C10606 vdd.n10233 vss 0.00425f
C10607 vdd.n10234 vss 0.00413f
C10608 vdd.n10235 vss 0.00251f
C10609 vdd.n10236 vss 0.0471f
C10610 vdd.n10237 vss 0.00251f
C10611 vdd.n10238 vss 0.00517f
C10612 vdd.n10239 vss 0.00679f
C10613 vdd.n10240 vss 0.00324f
C10614 vdd.n10241 vss 0.00324f
C10615 vdd.n10242 vss 0.0132f
C10616 vdd.n10243 vss 0.0424f
C10617 vdd.n10244 vss 0.02f
C10618 vdd.n10245 vss 0.00425f
C10619 vdd.n10246 vss 0.0471f
C10620 vdd.n10248 vss 0.00425f
C10621 vdd.n10249 vss 0.00925f
C10622 vdd.n10250 vss 0.00679f
C10623 vdd.n10251 vss 0.00517f
C10624 vdd.n10252 vss 0.00251f
C10625 vdd.n10253 vss 0.0471f
C10626 vdd.n10254 vss 0.00251f
C10627 vdd.n10255 vss 0.0112f
C10628 vdd.n10256 vss 0.0128f
C10629 vdd.n10257 vss 0.0692f
C10630 vdd.n10258 vss 0.00324f
C10631 vdd.n10259 vss 0.0112f
C10632 vdd.n10260 vss 0.0128f
C10633 vdd.n10261 vss 0.00413f
C10634 vdd.n10262 vss 0.00413f
C10635 vdd.n10263 vss 0.0471f
C10636 vdd.n10264 vss 0.0471f
C10637 vdd.n10265 vss 0.00324f
C10638 vdd.n10266 vss 0.00413f
C10639 vdd.n10267 vss 0.00413f
C10640 vdd.n10268 vss 0.00679f
C10641 vdd.n10269 vss 0.00413f
C10642 vdd.n10270 vss 0.0471f
C10643 vdd.n10271 vss 0.00324f
C10644 vdd.n10273 vss 0.00925f
C10645 vdd.n10274 vss 0.0471f
C10646 vdd.n10275 vss 0.00425f
C10647 vdd.n10276 vss 0.0424f
C10648 vdd.n10277 vss 0.0132f
C10649 vdd.n10278 vss 0.00324f
C10650 vdd.n10279 vss 0.0128f
C10651 vdd.n10280 vss 0.02f
C10652 vdd.n10281 vss 0.00425f
C10653 vdd.n10282 vss 0.00413f
C10654 vdd.n10283 vss 0.00251f
C10655 vdd.n10284 vss 0.0471f
C10656 vdd.n10285 vss 0.00251f
C10657 vdd.n10286 vss 0.00517f
C10658 vdd.n10287 vss 0.00679f
C10659 vdd.n10288 vss 0.00324f
C10660 vdd.n10289 vss 0.00324f
C10661 vdd.n10290 vss 0.0132f
C10662 vdd.n10291 vss 0.0424f
C10663 vdd.n10292 vss 0.02f
C10664 vdd.n10293 vss 0.00425f
C10665 vdd.n10294 vss 0.0471f
C10666 vdd.n10296 vss 0.00425f
C10667 vdd.n10297 vss 0.00925f
C10668 vdd.n10298 vss 0.00679f
C10669 vdd.n10299 vss 0.00517f
C10670 vdd.n10300 vss 0.00251f
C10671 vdd.n10301 vss 0.0471f
C10672 vdd.n10302 vss 0.00251f
C10673 vdd.n10303 vss 0.0112f
C10674 vdd.n10304 vss 0.0128f
C10675 vdd.n10305 vss 0.0619f
C10676 vdd.n10306 vss 0.00324f
C10677 vdd.n10307 vss 0.0112f
C10678 vdd.n10308 vss 0.0128f
C10679 vdd.n10309 vss 0.00413f
C10680 vdd.n10310 vss 0.00413f
C10681 vdd.n10311 vss 0.0471f
C10682 vdd.n10312 vss 0.0471f
C10683 vdd.n10313 vss 0.00324f
C10684 vdd.n10314 vss 0.00413f
C10685 vdd.n10315 vss 0.00413f
C10686 vdd.n10316 vss 0.00679f
C10687 vdd.n10317 vss 0.00413f
C10688 vdd.n10318 vss 0.0471f
C10689 vdd.n10319 vss 0.00324f
C10690 vdd.n10321 vss 0.00925f
C10691 vdd.n10322 vss 0.0471f
C10692 vdd.n10323 vss 0.00425f
C10693 vdd.n10324 vss 0.0424f
C10694 vdd.n10325 vss 0.0132f
C10695 vdd.n10326 vss 0.00324f
C10696 vdd.n10327 vss 0.0128f
C10697 vdd.n10328 vss 0.02f
C10698 vdd.n10329 vss 0.00425f
C10699 vdd.n10330 vss 0.00413f
C10700 vdd.n10331 vss 0.00251f
C10701 vdd.n10332 vss 0.0471f
C10702 vdd.n10333 vss 0.00251f
C10703 vdd.n10334 vss 0.00517f
C10704 vdd.n10335 vss 0.00679f
C10705 vdd.n10336 vss 0.00324f
C10706 vdd.n10337 vss 0.00324f
C10707 vdd.n10338 vss 0.0132f
C10708 vdd.n10339 vss 0.0424f
C10709 vdd.n10340 vss 0.02f
C10710 vdd.n10341 vss 0.00425f
C10711 vdd.n10342 vss 0.0471f
C10712 vdd.n10344 vss 0.00425f
C10713 vdd.n10345 vss 0.00925f
C10714 vdd.n10346 vss 0.00679f
C10715 vdd.n10347 vss 0.00517f
C10716 vdd.n10348 vss 0.00251f
C10717 vdd.n10349 vss 0.0471f
C10718 vdd.n10350 vss 0.00251f
C10719 vdd.n10351 vss 0.0112f
C10720 vdd.n10352 vss 0.0128f
C10721 vdd.n10353 vss 0.0692f
C10722 vdd.n10354 vss 0.00324f
C10723 vdd.n10355 vss 0.0112f
C10724 vdd.n10356 vss 0.0128f
C10725 vdd.n10357 vss 0.00413f
C10726 vdd.n10358 vss 0.00413f
C10727 vdd.n10359 vss 0.0471f
C10728 vdd.n10360 vss 0.0471f
C10729 vdd.n10361 vss 0.00324f
C10730 vdd.n10362 vss 0.00413f
C10731 vdd.n10363 vss 0.00413f
C10732 vdd.n10364 vss 0.00679f
C10733 vdd.n10365 vss 0.00413f
C10734 vdd.n10366 vss 0.0471f
C10735 vdd.n10367 vss 0.00324f
C10736 vdd.n10369 vss 0.00925f
C10737 vdd.n10370 vss 0.0471f
C10738 vdd.n10371 vss 0.00425f
C10739 vdd.n10372 vss 0.0424f
C10740 vdd.n10373 vss 0.0132f
C10741 vdd.n10374 vss 0.00324f
C10742 vdd.n10375 vss 0.0128f
C10743 vdd.n10376 vss 0.02f
C10744 vdd.n10377 vss 0.00425f
C10745 vdd.n10378 vss 0.00413f
C10746 vdd.n10379 vss 0.00251f
C10747 vdd.n10380 vss 0.0471f
C10748 vdd.n10381 vss 0.00251f
C10749 vdd.n10382 vss 0.00517f
C10750 vdd.n10383 vss 0.00679f
C10751 vdd.n10384 vss 0.00324f
C10752 vdd.n10385 vss 0.00324f
C10753 vdd.n10386 vss 0.0132f
C10754 vdd.n10387 vss 0.0424f
C10755 vdd.n10388 vss 0.02f
C10756 vdd.n10389 vss 0.00425f
C10757 vdd.n10390 vss 0.0471f
C10758 vdd.n10392 vss 0.00425f
C10759 vdd.n10393 vss 0.00925f
C10760 vdd.n10394 vss 0.00679f
C10761 vdd.n10395 vss 0.00517f
C10762 vdd.n10396 vss 0.00251f
C10763 vdd.n10397 vss 0.0471f
C10764 vdd.n10398 vss 0.00251f
C10765 vdd.n10399 vss 0.0112f
C10766 vdd.n10400 vss 0.0128f
C10767 vdd.n10401 vss 0.0619f
C10768 vdd.n10402 vss 0.00335f
C10769 vdd.n10403 vss 0.0855f
C10770 vdd.n10404 vss 0.00991f
C10771 vdd.n10405 vss 0.0424f
C10772 vdd.n10406 vss 0.00679f
C10773 vdd.n10407 vss 0.00413f
C10774 vdd.n10408 vss 0.0471f
C10775 vdd.n10409 vss 0.00251f
C10776 vdd.n10410 vss 0.00679f
C10777 vdd.n10411 vss 0.00413f
C10778 vdd.n10412 vss 0.00413f
C10779 vdd.n10413 vss 0.0471f
C10780 vdd.n10414 vss 0.00251f
C10781 vdd.n10415 vss 0.00413f
C10782 vdd.n10416 vss 0.00324f
C10783 vdd.n10417 vss 0.0132f
C10784 vdd.n10418 vss 0.0424f
C10785 vdd.n10419 vss 0.00324f
C10786 vdd.n10420 vss 0.00413f
C10787 vdd.n10421 vss 0.00517f
C10788 vdd.n10422 vss 0.00679f
C10789 vdd.n10423 vss 0.00925f
C10790 vdd.n10424 vss 0.00425f
C10791 vdd.n10425 vss 0.0471f
C10792 vdd.n10427 vss 0.00425f
C10793 vdd.n10428 vss 0.02f
C10794 vdd.n10429 vss 0.0128f
C10795 vdd.n10430 vss 0.0105f
C10796 vdd.n10431 vss 0.00251f
C10797 vdd.n10432 vss 0.0471f
C10798 vdd.n10433 vss 0.00517f
C10799 vdd.n10434 vss 0.00251f
C10800 vdd.n10435 vss 0.0471f
C10801 vdd.n10436 vss 0.0471f
C10802 vdd.n10437 vss 0.00324f
C10803 vdd.n10438 vss 0.00324f
C10804 vdd.n10439 vss 0.00805f
C10805 vdd.n10440 vss 0.0112f
C10806 vdd.n10441 vss 0.0128f
C10807 vdd.n10442 vss 0.00324f
C10808 vdd.n10443 vss 0.00324f
C10809 vdd.n10444 vss 0.00413f
C10810 vdd.n10445 vss 0.00425f
C10811 vdd.n10446 vss 0.0471f
C10812 vdd.n10448 vss 0.00425f
C10813 vdd.n10449 vss 0.00925f
C10814 vdd.n10450 vss 0.0107f
C10815 vdd.n10451 vss 0.0126f
C10816 vdd.n10452 vss 0.0516f
C10817 vdd.n10453 vss 0.00163f
C10818 vdd.n10454 vss 0.00145f
C10819 vdd.n10455 vss 0.0271f
C10820 vdd.n10456 vss 0.00324f
C10821 vdd.n10457 vss 0.0112f
C10822 vdd.n10458 vss 0.0128f
C10823 vdd.n10459 vss 0.00413f
C10824 vdd.n10460 vss 0.00413f
C10825 vdd.n10461 vss 0.0471f
C10826 vdd.n10462 vss 0.0471f
C10827 vdd.n10463 vss 0.00324f
C10828 vdd.n10464 vss 0.00413f
C10829 vdd.n10465 vss 0.00413f
C10830 vdd.n10466 vss 0.00679f
C10831 vdd.n10467 vss 0.00413f
C10832 vdd.n10468 vss 0.0471f
C10833 vdd.n10469 vss 0.00324f
C10834 vdd.n10471 vss 0.00925f
C10835 vdd.n10472 vss 0.0471f
C10836 vdd.n10473 vss 0.00425f
C10837 vdd.n10474 vss 0.0424f
C10838 vdd.n10475 vss 0.0132f
C10839 vdd.n10476 vss 0.00324f
C10840 vdd.n10477 vss 0.0128f
C10841 vdd.n10478 vss 0.02f
C10842 vdd.n10479 vss 0.00425f
C10843 vdd.n10480 vss 0.00413f
C10844 vdd.n10481 vss 0.00251f
C10845 vdd.n10482 vss 0.0471f
C10846 vdd.n10483 vss 0.00251f
C10847 vdd.n10484 vss 0.00517f
C10848 vdd.n10485 vss 0.00679f
C10849 vdd.n10486 vss 0.00324f
C10850 vdd.n10487 vss 0.00324f
C10851 vdd.n10488 vss 0.0132f
C10852 vdd.n10489 vss 0.0424f
C10853 vdd.n10490 vss 0.02f
C10854 vdd.n10491 vss 0.00425f
C10855 vdd.n10492 vss 0.0471f
C10856 vdd.n10494 vss 0.00425f
C10857 vdd.n10495 vss 0.00925f
C10858 vdd.n10496 vss 0.00679f
C10859 vdd.n10497 vss 0.00517f
C10860 vdd.n10498 vss 0.00251f
C10861 vdd.n10499 vss 0.0471f
C10862 vdd.n10500 vss 0.00251f
C10863 vdd.n10501 vss 0.0112f
C10864 vdd.n10502 vss 0.0128f
C10865 vdd.n10503 vss 0.0692f
C10866 vdd.n10504 vss 0.00324f
C10867 vdd.n10505 vss 0.0112f
C10868 vdd.n10506 vss 0.0128f
C10869 vdd.n10507 vss 0.00413f
C10870 vdd.n10508 vss 0.00413f
C10871 vdd.n10509 vss 0.0471f
C10872 vdd.n10510 vss 0.0471f
C10873 vdd.n10511 vss 0.00324f
C10874 vdd.n10512 vss 0.00413f
C10875 vdd.n10513 vss 0.00413f
C10876 vdd.n10514 vss 0.00679f
C10877 vdd.n10515 vss 0.00413f
C10878 vdd.n10516 vss 0.0471f
C10879 vdd.n10517 vss 0.00324f
C10880 vdd.n10519 vss 0.00925f
C10881 vdd.n10520 vss 0.0471f
C10882 vdd.n10521 vss 0.00425f
C10883 vdd.n10522 vss 0.0424f
C10884 vdd.n10523 vss 0.0132f
C10885 vdd.n10524 vss 0.00324f
C10886 vdd.n10525 vss 0.0128f
C10887 vdd.n10526 vss 0.02f
C10888 vdd.n10527 vss 0.00425f
C10889 vdd.n10528 vss 0.00413f
C10890 vdd.n10529 vss 0.00251f
C10891 vdd.n10530 vss 0.0471f
C10892 vdd.n10531 vss 0.00251f
C10893 vdd.n10532 vss 0.00517f
C10894 vdd.n10533 vss 0.00679f
C10895 vdd.n10534 vss 0.00324f
C10896 vdd.n10535 vss 0.00324f
C10897 vdd.n10536 vss 0.0132f
C10898 vdd.n10537 vss 0.0424f
C10899 vdd.n10538 vss 0.02f
C10900 vdd.n10539 vss 0.00425f
C10901 vdd.n10540 vss 0.0471f
C10902 vdd.n10542 vss 0.00425f
C10903 vdd.n10543 vss 0.00925f
C10904 vdd.n10544 vss 0.00679f
C10905 vdd.n10545 vss 0.00517f
C10906 vdd.n10546 vss 0.00251f
C10907 vdd.n10547 vss 0.0471f
C10908 vdd.n10548 vss 0.00251f
C10909 vdd.n10549 vss 0.0112f
C10910 vdd.n10550 vss 0.0128f
C10911 vdd.n10551 vss 0.0692f
C10912 vdd.n10552 vss 0.118f
C10913 vdd.n10553 vss 0.121f
C10914 vdd.n10554 vss 0.00324f
C10915 vdd.n10555 vss 0.0112f
C10916 vdd.n10556 vss 0.0128f
C10917 vdd.n10557 vss 0.00413f
C10918 vdd.n10558 vss 0.00413f
C10919 vdd.n10559 vss 0.0471f
C10920 vdd.n10560 vss 0.0471f
C10921 vdd.n10561 vss 0.00324f
C10922 vdd.n10562 vss 0.00413f
C10923 vdd.n10563 vss 0.00413f
C10924 vdd.n10564 vss 0.00679f
C10925 vdd.n10565 vss 0.00413f
C10926 vdd.n10566 vss 0.0471f
C10927 vdd.n10567 vss 0.00324f
C10928 vdd.n10569 vss 0.00925f
C10929 vdd.n10570 vss 0.0471f
C10930 vdd.n10571 vss 0.00425f
C10931 vdd.n10572 vss 0.0424f
C10932 vdd.n10573 vss 0.0132f
C10933 vdd.n10574 vss 0.00324f
C10934 vdd.n10575 vss 0.0128f
C10935 vdd.n10576 vss 0.02f
C10936 vdd.n10577 vss 0.00425f
C10937 vdd.n10578 vss 0.00413f
C10938 vdd.n10579 vss 0.00251f
C10939 vdd.n10580 vss 0.0471f
C10940 vdd.n10581 vss 0.00251f
C10941 vdd.n10582 vss 0.00517f
C10942 vdd.n10583 vss 0.00679f
C10943 vdd.n10584 vss 0.00324f
C10944 vdd.n10585 vss 0.00324f
C10945 vdd.n10586 vss 0.0132f
C10946 vdd.n10587 vss 0.0424f
C10947 vdd.n10588 vss 0.02f
C10948 vdd.n10589 vss 0.00425f
C10949 vdd.n10590 vss 0.0471f
C10950 vdd.n10592 vss 0.00425f
C10951 vdd.n10593 vss 0.00925f
C10952 vdd.n10594 vss 0.00679f
C10953 vdd.n10595 vss 0.00517f
C10954 vdd.n10596 vss 0.00251f
C10955 vdd.n10597 vss 0.0471f
C10956 vdd.n10598 vss 0.00251f
C10957 vdd.n10599 vss 0.0112f
C10958 vdd.n10600 vss 0.098f
C10959 vdd.n10601 vss 0.0596f
C10960 vdd.n10602 vss 0.00324f
C10961 vdd.n10603 vss 0.0112f
C10962 vdd.n10604 vss 0.0128f
C10963 vdd.n10605 vss 0.00413f
C10964 vdd.n10606 vss 0.00413f
C10965 vdd.n10607 vss 0.0471f
C10966 vdd.n10608 vss 0.0471f
C10967 vdd.n10609 vss 0.00324f
C10968 vdd.n10610 vss 0.00413f
C10969 vdd.n10611 vss 0.00413f
C10970 vdd.n10612 vss 0.00679f
C10971 vdd.n10613 vss 0.00413f
C10972 vdd.n10614 vss 0.0471f
C10973 vdd.n10615 vss 0.00324f
C10974 vdd.n10617 vss 0.00925f
C10975 vdd.n10618 vss 0.0471f
C10976 vdd.n10619 vss 0.00425f
C10977 vdd.n10620 vss 0.0424f
C10978 vdd.n10621 vss 0.0132f
C10979 vdd.n10622 vss 0.00324f
C10980 vdd.n10623 vss 0.0128f
C10981 vdd.n10624 vss 0.02f
C10982 vdd.n10625 vss 0.00425f
C10983 vdd.n10626 vss 0.00413f
C10984 vdd.n10627 vss 0.00251f
C10985 vdd.n10628 vss 0.0471f
C10986 vdd.n10629 vss 0.00251f
C10987 vdd.n10630 vss 0.00517f
C10988 vdd.n10631 vss 0.00679f
C10989 vdd.n10632 vss 0.00324f
C10990 vdd.n10633 vss 0.00324f
C10991 vdd.n10634 vss 0.0132f
C10992 vdd.n10635 vss 0.0424f
C10993 vdd.n10636 vss 0.02f
C10994 vdd.n10637 vss 0.00425f
C10995 vdd.n10638 vss 0.0471f
C10996 vdd.n10640 vss 0.00425f
C10997 vdd.n10641 vss 0.00925f
C10998 vdd.n10642 vss 0.00679f
C10999 vdd.n10643 vss 0.00517f
C11000 vdd.n10644 vss 0.00251f
C11001 vdd.n10645 vss 0.0471f
C11002 vdd.n10646 vss 0.00251f
C11003 vdd.n10647 vss 0.0112f
C11004 vdd.n10648 vss 0.0128f
C11005 vdd.n10649 vss 0.0692f
C11006 vdd.n10650 vss 0.0912f
C11007 vdd.n10651 vss 0.0824f
C11008 vdd.n10652 vss 0.059f
C11009 vdd.n10653 vss 0.00324f
C11010 vdd.n10654 vss 0.0112f
C11011 vdd.n10655 vss 0.0128f
C11012 vdd.n10656 vss 0.00413f
C11013 vdd.n10657 vss 0.00413f
C11014 vdd.n10658 vss 0.0471f
C11015 vdd.n10659 vss 0.0471f
C11016 vdd.n10660 vss 0.00324f
C11017 vdd.n10661 vss 0.00413f
C11018 vdd.n10662 vss 0.00413f
C11019 vdd.n10663 vss 0.00679f
C11020 vdd.n10664 vss 0.00413f
C11021 vdd.n10665 vss 0.0471f
C11022 vdd.n10666 vss 0.00324f
C11023 vdd.n10668 vss 0.00925f
C11024 vdd.n10669 vss 0.0471f
C11025 vdd.n10670 vss 0.00425f
C11026 vdd.n10671 vss 0.0424f
C11027 vdd.n10672 vss 0.0132f
C11028 vdd.n10673 vss 0.00324f
C11029 vdd.n10674 vss 0.0128f
C11030 vdd.n10675 vss 0.02f
C11031 vdd.n10676 vss 0.00425f
C11032 vdd.n10677 vss 0.00413f
C11033 vdd.n10678 vss 0.00251f
C11034 vdd.n10679 vss 0.0471f
C11035 vdd.n10680 vss 0.00251f
C11036 vdd.n10681 vss 0.00517f
C11037 vdd.n10682 vss 0.00679f
C11038 vdd.n10683 vss 0.00324f
C11039 vdd.n10684 vss 0.00324f
C11040 vdd.n10685 vss 0.0132f
C11041 vdd.n10686 vss 0.0424f
C11042 vdd.n10687 vss 0.02f
C11043 vdd.n10688 vss 0.00425f
C11044 vdd.n10689 vss 0.0471f
C11045 vdd.n10691 vss 0.00425f
C11046 vdd.n10692 vss 0.00925f
C11047 vdd.n10693 vss 0.00679f
C11048 vdd.n10694 vss 0.00517f
C11049 vdd.n10695 vss 0.00251f
C11050 vdd.n10696 vss 0.0471f
C11051 vdd.n10697 vss 0.00251f
C11052 vdd.n10698 vss 0.0112f
C11053 vdd.n10699 vss 0.0128f
C11054 vdd.n10700 vss 0.185f
C11055 vdd.n10701 vss 0.00324f
C11056 vdd.n10702 vss 0.0112f
C11057 vdd.n10703 vss 0.0128f
C11058 vdd.n10704 vss 0.00413f
C11059 vdd.n10705 vss 0.00413f
C11060 vdd.n10706 vss 0.0471f
C11061 vdd.n10707 vss 0.0471f
C11062 vdd.n10708 vss 0.00324f
C11063 vdd.n10709 vss 0.00413f
C11064 vdd.n10710 vss 0.00413f
C11065 vdd.n10711 vss 0.00679f
C11066 vdd.n10712 vss 0.00413f
C11067 vdd.n10713 vss 0.0471f
C11068 vdd.n10714 vss 0.00324f
C11069 vdd.n10716 vss 0.00925f
C11070 vdd.n10717 vss 0.0471f
C11071 vdd.n10718 vss 0.00425f
C11072 vdd.n10719 vss 0.0424f
C11073 vdd.n10720 vss 0.0132f
C11074 vdd.n10721 vss 0.00324f
C11075 vdd.n10722 vss 0.0128f
C11076 vdd.n10723 vss 0.02f
C11077 vdd.n10724 vss 0.00425f
C11078 vdd.n10725 vss 0.00413f
C11079 vdd.n10726 vss 0.00251f
C11080 vdd.n10727 vss 0.0471f
C11081 vdd.n10728 vss 0.00251f
C11082 vdd.n10729 vss 0.00517f
C11083 vdd.n10730 vss 0.00679f
C11084 vdd.n10731 vss 0.00324f
C11085 vdd.n10732 vss 0.00324f
C11086 vdd.n10733 vss 0.0132f
C11087 vdd.n10734 vss 0.0424f
C11088 vdd.n10735 vss 0.02f
C11089 vdd.n10736 vss 0.00425f
C11090 vdd.n10737 vss 0.0471f
C11091 vdd.n10739 vss 0.00425f
C11092 vdd.n10740 vss 0.00925f
C11093 vdd.n10741 vss 0.00679f
C11094 vdd.n10742 vss 0.00517f
C11095 vdd.n10743 vss 0.00251f
C11096 vdd.n10744 vss 0.0471f
C11097 vdd.n10745 vss 0.00251f
C11098 vdd.n10746 vss 0.0112f
C11099 vdd.n10747 vss 0.0128f
C11100 vdd.n10748 vss 0.059f
C11101 vdd.n10749 vss 0.256f
C11102 vdd.n10750 vss 0.00324f
C11103 vdd.n10751 vss 0.0112f
C11104 vdd.n10752 vss 0.0128f
C11105 vdd.n10753 vss 0.00413f
C11106 vdd.n10754 vss 0.00413f
C11107 vdd.n10755 vss 0.0471f
C11108 vdd.n10756 vss 0.0471f
C11109 vdd.n10757 vss 0.00324f
C11110 vdd.n10758 vss 0.00413f
C11111 vdd.n10759 vss 0.00413f
C11112 vdd.n10760 vss 0.00679f
C11113 vdd.n10761 vss 0.00413f
C11114 vdd.n10762 vss 0.0471f
C11115 vdd.n10763 vss 0.00324f
C11116 vdd.n10765 vss 0.00925f
C11117 vdd.n10766 vss 0.0471f
C11118 vdd.n10767 vss 0.00425f
C11119 vdd.n10768 vss 0.0424f
C11120 vdd.n10769 vss 0.0132f
C11121 vdd.n10770 vss 0.00324f
C11122 vdd.n10771 vss 0.0128f
C11123 vdd.n10772 vss 0.02f
C11124 vdd.n10773 vss 0.00425f
C11125 vdd.n10774 vss 0.00413f
C11126 vdd.n10775 vss 0.00251f
C11127 vdd.n10776 vss 0.0471f
C11128 vdd.n10777 vss 0.00251f
C11129 vdd.n10778 vss 0.00517f
C11130 vdd.n10779 vss 0.00679f
C11131 vdd.n10780 vss 0.00324f
C11132 vdd.n10781 vss 0.00324f
C11133 vdd.n10782 vss 0.0132f
C11134 vdd.n10783 vss 0.0424f
C11135 vdd.n10784 vss 0.02f
C11136 vdd.n10785 vss 0.00425f
C11137 vdd.n10786 vss 0.0471f
C11138 vdd.n10788 vss 0.00425f
C11139 vdd.n10789 vss 0.00925f
C11140 vdd.n10790 vss 0.00679f
C11141 vdd.n10791 vss 0.00517f
C11142 vdd.n10792 vss 0.00251f
C11143 vdd.n10793 vss 0.0471f
C11144 vdd.n10794 vss 0.00251f
C11145 vdd.n10795 vss 0.0112f
C11146 vdd.n10796 vss 0.0128f
C11147 vdd.n10797 vss 0.123f
C11148 vdd.n10798 vss 0.0596f
C11149 vdd.n10799 vss 0.00324f
C11150 vdd.n10800 vss 0.0112f
C11151 vdd.n10801 vss 0.0128f
C11152 vdd.n10802 vss 0.00413f
C11153 vdd.n10803 vss 0.00413f
C11154 vdd.n10804 vss 0.0471f
C11155 vdd.n10805 vss 0.0471f
C11156 vdd.n10806 vss 0.00324f
C11157 vdd.n10807 vss 0.00413f
C11158 vdd.n10808 vss 0.00413f
C11159 vdd.n10809 vss 0.00679f
C11160 vdd.n10810 vss 0.00413f
C11161 vdd.n10811 vss 0.0471f
C11162 vdd.n10812 vss 0.00324f
C11163 vdd.n10814 vss 0.00925f
C11164 vdd.n10815 vss 0.0471f
C11165 vdd.n10816 vss 0.00425f
C11166 vdd.n10817 vss 0.0424f
C11167 vdd.n10818 vss 0.0132f
C11168 vdd.n10819 vss 0.00324f
C11169 vdd.n10820 vss 0.0128f
C11170 vdd.n10821 vss 0.02f
C11171 vdd.n10822 vss 0.00425f
C11172 vdd.n10823 vss 0.00413f
C11173 vdd.n10824 vss 0.00251f
C11174 vdd.n10825 vss 0.0471f
C11175 vdd.n10826 vss 0.00251f
C11176 vdd.n10827 vss 0.00517f
C11177 vdd.n10828 vss 0.00679f
C11178 vdd.n10829 vss 0.00324f
C11179 vdd.n10830 vss 0.00324f
C11180 vdd.n10831 vss 0.0132f
C11181 vdd.n10832 vss 0.0424f
C11182 vdd.n10833 vss 0.02f
C11183 vdd.n10834 vss 0.00425f
C11184 vdd.n10835 vss 0.0471f
C11185 vdd.n10837 vss 0.00425f
C11186 vdd.n10838 vss 0.00925f
C11187 vdd.n10839 vss 0.00679f
C11188 vdd.n10840 vss 0.00517f
C11189 vdd.n10841 vss 0.00251f
C11190 vdd.n10842 vss 0.0471f
C11191 vdd.n10843 vss 0.00251f
C11192 vdd.n10844 vss 0.0112f
C11193 vdd.n10845 vss 0.0128f
C11194 vdd.n10846 vss 0.0692f
C11195 vdd.n10847 vss 0.118f
C11196 vdd.n10848 vss 0.121f
C11197 vdd.n10849 vss 0.00324f
C11198 vdd.n10850 vss 0.0112f
C11199 vdd.n10851 vss 0.0128f
C11200 vdd.n10852 vss 0.00413f
C11201 vdd.n10853 vss 0.00413f
C11202 vdd.n10854 vss 0.0471f
C11203 vdd.n10855 vss 0.0471f
C11204 vdd.n10856 vss 0.00324f
C11205 vdd.n10857 vss 0.00413f
C11206 vdd.n10858 vss 0.00413f
C11207 vdd.n10859 vss 0.00679f
C11208 vdd.n10860 vss 0.00413f
C11209 vdd.n10861 vss 0.0471f
C11210 vdd.n10862 vss 0.00324f
C11211 vdd.n10864 vss 0.00925f
C11212 vdd.n10865 vss 0.0471f
C11213 vdd.n10866 vss 0.00425f
C11214 vdd.n10867 vss 0.0424f
C11215 vdd.n10868 vss 0.0132f
C11216 vdd.n10869 vss 0.00324f
C11217 vdd.n10870 vss 0.0128f
C11218 vdd.n10871 vss 0.02f
C11219 vdd.n10872 vss 0.00425f
C11220 vdd.n10873 vss 0.00413f
C11221 vdd.n10874 vss 0.00251f
C11222 vdd.n10875 vss 0.0471f
C11223 vdd.n10876 vss 0.00251f
C11224 vdd.n10877 vss 0.00517f
C11225 vdd.n10878 vss 0.00679f
C11226 vdd.n10879 vss 0.00324f
C11227 vdd.n10880 vss 0.00324f
C11228 vdd.n10881 vss 0.0132f
C11229 vdd.n10882 vss 0.0424f
C11230 vdd.n10883 vss 0.02f
C11231 vdd.n10884 vss 0.00425f
C11232 vdd.n10885 vss 0.0471f
C11233 vdd.n10887 vss 0.00425f
C11234 vdd.n10888 vss 0.00925f
C11235 vdd.n10889 vss 0.00679f
C11236 vdd.n10890 vss 0.00517f
C11237 vdd.n10891 vss 0.00251f
C11238 vdd.n10892 vss 0.0471f
C11239 vdd.n10893 vss 0.00251f
C11240 vdd.n10894 vss 0.0112f
C11241 vdd.n10895 vss 0.098f
C11242 vdd.n10896 vss 0.0596f
C11243 vdd.n10897 vss 0.00324f
C11244 vdd.n10898 vss 0.0112f
C11245 vdd.n10899 vss 0.0128f
C11246 vdd.n10900 vss 0.00413f
C11247 vdd.n10901 vss 0.00413f
C11248 vdd.n10902 vss 0.0471f
C11249 vdd.n10903 vss 0.0471f
C11250 vdd.n10904 vss 0.00324f
C11251 vdd.n10905 vss 0.00413f
C11252 vdd.n10906 vss 0.00413f
C11253 vdd.n10907 vss 0.00679f
C11254 vdd.n10908 vss 0.00413f
C11255 vdd.n10909 vss 0.0471f
C11256 vdd.n10910 vss 0.00324f
C11257 vdd.n10912 vss 0.00925f
C11258 vdd.n10913 vss 0.0471f
C11259 vdd.n10914 vss 0.00425f
C11260 vdd.n10915 vss 0.0424f
C11261 vdd.n10916 vss 0.0132f
C11262 vdd.n10917 vss 0.00324f
C11263 vdd.n10918 vss 0.0128f
C11264 vdd.n10919 vss 0.02f
C11265 vdd.n10920 vss 0.00425f
C11266 vdd.n10921 vss 0.00413f
C11267 vdd.n10922 vss 0.00251f
C11268 vdd.n10923 vss 0.0471f
C11269 vdd.n10924 vss 0.00251f
C11270 vdd.n10925 vss 0.00517f
C11271 vdd.n10926 vss 0.00679f
C11272 vdd.n10927 vss 0.00324f
C11273 vdd.n10928 vss 0.00324f
C11274 vdd.n10929 vss 0.0132f
C11275 vdd.n10930 vss 0.0424f
C11276 vdd.n10931 vss 0.02f
C11277 vdd.n10932 vss 0.00425f
C11278 vdd.n10933 vss 0.0471f
C11279 vdd.n10935 vss 0.00425f
C11280 vdd.n10936 vss 0.00925f
C11281 vdd.n10937 vss 0.00679f
C11282 vdd.n10938 vss 0.00517f
C11283 vdd.n10939 vss 0.00251f
C11284 vdd.n10940 vss 0.0471f
C11285 vdd.n10941 vss 0.00251f
C11286 vdd.n10942 vss 0.0112f
C11287 vdd.n10943 vss 0.0128f
C11288 vdd.n10944 vss 0.0692f
C11289 vdd.n10945 vss 0.118f
C11290 vdd.n10946 vss 0.0951f
C11291 vdd.n10947 vss 0.00324f
C11292 vdd.n10948 vss 0.0112f
C11293 vdd.n10949 vss 0.0128f
C11294 vdd.n10950 vss 0.00413f
C11295 vdd.n10951 vss 0.00413f
C11296 vdd.n10952 vss 0.0471f
C11297 vdd.n10953 vss 0.0471f
C11298 vdd.n10954 vss 0.00324f
C11299 vdd.n10955 vss 0.00413f
C11300 vdd.n10956 vss 0.00413f
C11301 vdd.n10957 vss 0.00679f
C11302 vdd.n10958 vss 0.00413f
C11303 vdd.n10959 vss 0.0471f
C11304 vdd.n10960 vss 0.00324f
C11305 vdd.n10962 vss 0.00925f
C11306 vdd.n10963 vss 0.0471f
C11307 vdd.n10964 vss 0.00425f
C11308 vdd.n10965 vss 0.0424f
C11309 vdd.n10966 vss 0.0132f
C11310 vdd.n10967 vss 0.00324f
C11311 vdd.n10968 vss 0.0128f
C11312 vdd.n10969 vss 0.02f
C11313 vdd.n10970 vss 0.00425f
C11314 vdd.n10971 vss 0.00413f
C11315 vdd.n10972 vss 0.00251f
C11316 vdd.n10973 vss 0.0471f
C11317 vdd.n10974 vss 0.00251f
C11318 vdd.n10975 vss 0.00517f
C11319 vdd.n10976 vss 0.00679f
C11320 vdd.n10977 vss 0.00324f
C11321 vdd.n10978 vss 0.00324f
C11322 vdd.n10979 vss 0.0132f
C11323 vdd.n10980 vss 0.0424f
C11324 vdd.n10981 vss 0.02f
C11325 vdd.n10982 vss 0.00425f
C11326 vdd.n10983 vss 0.0471f
C11327 vdd.n10985 vss 0.00425f
C11328 vdd.n10986 vss 0.00925f
C11329 vdd.n10987 vss 0.00679f
C11330 vdd.n10988 vss 0.00517f
C11331 vdd.n10989 vss 0.00251f
C11332 vdd.n10990 vss 0.0471f
C11333 vdd.n10991 vss 0.00251f
C11334 vdd.n10992 vss 0.0112f
C11335 vdd.n10993 vss 0.0128f
C11336 vdd.n10994 vss 0.146f
C11337 vdd.n10995 vss 0.00324f
C11338 vdd.n10996 vss 0.0112f
C11339 vdd.n10997 vss 0.0128f
C11340 vdd.n10998 vss 0.00413f
C11341 vdd.n10999 vss 0.00413f
C11342 vdd.n11000 vss 0.0471f
C11343 vdd.n11001 vss 0.0471f
C11344 vdd.n11002 vss 0.00324f
C11345 vdd.n11003 vss 0.00413f
C11346 vdd.n11004 vss 0.00413f
C11347 vdd.n11005 vss 0.00679f
C11348 vdd.n11006 vss 0.00413f
C11349 vdd.n11007 vss 0.0471f
C11350 vdd.n11008 vss 0.00324f
C11351 vdd.n11010 vss 0.00925f
C11352 vdd.n11011 vss 0.0471f
C11353 vdd.n11012 vss 0.00425f
C11354 vdd.n11013 vss 0.0424f
C11355 vdd.n11014 vss 0.0132f
C11356 vdd.n11015 vss 0.00324f
C11357 vdd.n11016 vss 0.0128f
C11358 vdd.n11017 vss 0.02f
C11359 vdd.n11018 vss 0.00425f
C11360 vdd.n11019 vss 0.00413f
C11361 vdd.n11020 vss 0.00251f
C11362 vdd.n11021 vss 0.0471f
C11363 vdd.n11022 vss 0.00251f
C11364 vdd.n11023 vss 0.00517f
C11365 vdd.n11024 vss 0.00679f
C11366 vdd.n11025 vss 0.00324f
C11367 vdd.n11026 vss 0.00324f
C11368 vdd.n11027 vss 0.0132f
C11369 vdd.n11028 vss 0.0424f
C11370 vdd.n11029 vss 0.02f
C11371 vdd.n11030 vss 0.00425f
C11372 vdd.n11031 vss 0.0471f
C11373 vdd.n11033 vss 0.00425f
C11374 vdd.n11034 vss 0.00925f
C11375 vdd.n11035 vss 0.00679f
C11376 vdd.n11036 vss 0.00517f
C11377 vdd.n11037 vss 0.00251f
C11378 vdd.n11038 vss 0.0471f
C11379 vdd.n11039 vss 0.00251f
C11380 vdd.n11040 vss 0.0112f
C11381 vdd.n11041 vss 0.0128f
C11382 vdd.n11042 vss 0.146f
C11383 vdd.n11043 vss 0.0596f
C11384 vdd.n11044 vss 0.00324f
C11385 vdd.n11045 vss 0.0112f
C11386 vdd.n11046 vss 0.0128f
C11387 vdd.n11047 vss 0.00413f
C11388 vdd.n11048 vss 0.00413f
C11389 vdd.n11049 vss 0.0471f
C11390 vdd.n11050 vss 0.0471f
C11391 vdd.n11051 vss 0.00324f
C11392 vdd.n11052 vss 0.00413f
C11393 vdd.n11053 vss 0.00413f
C11394 vdd.n11054 vss 0.00679f
C11395 vdd.n11055 vss 0.00413f
C11396 vdd.n11056 vss 0.0471f
C11397 vdd.n11057 vss 0.00324f
C11398 vdd.n11059 vss 0.00925f
C11399 vdd.n11060 vss 0.0471f
C11400 vdd.n11061 vss 0.00425f
C11401 vdd.n11062 vss 0.0424f
C11402 vdd.n11063 vss 0.0132f
C11403 vdd.n11064 vss 0.00324f
C11404 vdd.n11065 vss 0.0128f
C11405 vdd.n11066 vss 0.02f
C11406 vdd.n11067 vss 0.00425f
C11407 vdd.n11068 vss 0.00413f
C11408 vdd.n11069 vss 0.00251f
C11409 vdd.n11070 vss 0.0471f
C11410 vdd.n11071 vss 0.00251f
C11411 vdd.n11072 vss 0.00517f
C11412 vdd.n11073 vss 0.00679f
C11413 vdd.n11074 vss 0.00324f
C11414 vdd.n11075 vss 0.00324f
C11415 vdd.n11076 vss 0.0132f
C11416 vdd.n11077 vss 0.0424f
C11417 vdd.n11078 vss 0.02f
C11418 vdd.n11079 vss 0.00425f
C11419 vdd.n11080 vss 0.0471f
C11420 vdd.n11082 vss 0.00425f
C11421 vdd.n11083 vss 0.00925f
C11422 vdd.n11084 vss 0.00679f
C11423 vdd.n11085 vss 0.00517f
C11424 vdd.n11086 vss 0.00251f
C11425 vdd.n11087 vss 0.0471f
C11426 vdd.n11088 vss 0.00251f
C11427 vdd.n11089 vss 0.0112f
C11428 vdd.n11090 vss 0.0128f
C11429 vdd.n11091 vss 0.0692f
C11430 vdd.n11092 vss 0.118f
C11431 vdd.n11093 vss 0.121f
C11432 vdd.n11094 vss 0.00324f
C11433 vdd.n11095 vss 0.0112f
C11434 vdd.n11096 vss 0.0128f
C11435 vdd.n11097 vss 0.00413f
C11436 vdd.n11098 vss 0.00413f
C11437 vdd.n11099 vss 0.0471f
C11438 vdd.n11100 vss 0.0471f
C11439 vdd.n11101 vss 0.00324f
C11440 vdd.n11102 vss 0.00413f
C11441 vdd.n11103 vss 0.00413f
C11442 vdd.n11104 vss 0.00679f
C11443 vdd.n11105 vss 0.00413f
C11444 vdd.n11106 vss 0.0471f
C11445 vdd.n11107 vss 0.00324f
C11446 vdd.n11109 vss 0.00925f
C11447 vdd.n11110 vss 0.0471f
C11448 vdd.n11111 vss 0.00425f
C11449 vdd.n11112 vss 0.0424f
C11450 vdd.n11113 vss 0.0132f
C11451 vdd.n11114 vss 0.00324f
C11452 vdd.n11115 vss 0.0128f
C11453 vdd.n11116 vss 0.02f
C11454 vdd.n11117 vss 0.00425f
C11455 vdd.n11118 vss 0.00413f
C11456 vdd.n11119 vss 0.00251f
C11457 vdd.n11120 vss 0.0471f
C11458 vdd.n11121 vss 0.00251f
C11459 vdd.n11122 vss 0.00517f
C11460 vdd.n11123 vss 0.00679f
C11461 vdd.n11124 vss 0.00324f
C11462 vdd.n11125 vss 0.00324f
C11463 vdd.n11126 vss 0.0132f
C11464 vdd.n11127 vss 0.0424f
C11465 vdd.n11128 vss 0.02f
C11466 vdd.n11129 vss 0.00425f
C11467 vdd.n11130 vss 0.0471f
C11468 vdd.n11132 vss 0.00425f
C11469 vdd.n11133 vss 0.00925f
C11470 vdd.n11134 vss 0.00679f
C11471 vdd.n11135 vss 0.00517f
C11472 vdd.n11136 vss 0.00251f
C11473 vdd.n11137 vss 0.0471f
C11474 vdd.n11138 vss 0.00251f
C11475 vdd.n11139 vss 0.0112f
C11476 vdd.n11140 vss 0.098f
C11477 vdd.n11141 vss 0.0596f
C11478 vdd.n11142 vss 0.00324f
C11479 vdd.n11143 vss 0.0112f
C11480 vdd.n11144 vss 0.0128f
C11481 vdd.n11145 vss 0.00413f
C11482 vdd.n11146 vss 0.00413f
C11483 vdd.n11147 vss 0.0471f
C11484 vdd.n11148 vss 0.0471f
C11485 vdd.n11149 vss 0.00324f
C11486 vdd.n11150 vss 0.00413f
C11487 vdd.n11151 vss 0.00413f
C11488 vdd.n11152 vss 0.00679f
C11489 vdd.n11153 vss 0.00413f
C11490 vdd.n11154 vss 0.0471f
C11491 vdd.n11155 vss 0.00324f
C11492 vdd.n11157 vss 0.00925f
C11493 vdd.n11158 vss 0.0471f
C11494 vdd.n11159 vss 0.00425f
C11495 vdd.n11160 vss 0.0424f
C11496 vdd.n11161 vss 0.0132f
C11497 vdd.n11162 vss 0.00324f
C11498 vdd.n11163 vss 0.0128f
C11499 vdd.n11164 vss 0.02f
C11500 vdd.n11165 vss 0.00425f
C11501 vdd.n11166 vss 0.00413f
C11502 vdd.n11167 vss 0.00251f
C11503 vdd.n11168 vss 0.0471f
C11504 vdd.n11169 vss 0.00251f
C11505 vdd.n11170 vss 0.00517f
C11506 vdd.n11171 vss 0.00679f
C11507 vdd.n11172 vss 0.00324f
C11508 vdd.n11173 vss 0.00324f
C11509 vdd.n11174 vss 0.0132f
C11510 vdd.n11175 vss 0.0424f
C11511 vdd.n11176 vss 0.02f
C11512 vdd.n11177 vss 0.00425f
C11513 vdd.n11178 vss 0.0471f
C11514 vdd.n11180 vss 0.00425f
C11515 vdd.n11181 vss 0.00925f
C11516 vdd.n11182 vss 0.00679f
C11517 vdd.n11183 vss 0.00517f
C11518 vdd.n11184 vss 0.00251f
C11519 vdd.n11185 vss 0.0471f
C11520 vdd.n11186 vss 0.00251f
C11521 vdd.n11187 vss 0.0112f
C11522 vdd.n11188 vss 0.0128f
C11523 vdd.n11189 vss 0.0692f
C11524 vdd.n11190 vss 0.0912f
C11525 vdd.n11191 vss 0.0824f
C11526 vdd.n11192 vss 0.059f
C11527 vdd.n11193 vss 0.00324f
C11528 vdd.n11194 vss 0.0112f
C11529 vdd.n11195 vss 0.0128f
C11530 vdd.n11196 vss 0.00413f
C11531 vdd.n11197 vss 0.00413f
C11532 vdd.n11198 vss 0.0471f
C11533 vdd.n11199 vss 0.0471f
C11534 vdd.n11200 vss 0.00324f
C11535 vdd.n11201 vss 0.00413f
C11536 vdd.n11202 vss 0.00413f
C11537 vdd.n11203 vss 0.00679f
C11538 vdd.n11204 vss 0.00413f
C11539 vdd.n11205 vss 0.0471f
C11540 vdd.n11206 vss 0.00324f
C11541 vdd.n11208 vss 0.00925f
C11542 vdd.n11209 vss 0.0471f
C11543 vdd.n11210 vss 0.00425f
C11544 vdd.n11211 vss 0.0424f
C11545 vdd.n11212 vss 0.0132f
C11546 vdd.n11213 vss 0.00324f
C11547 vdd.n11214 vss 0.0128f
C11548 vdd.n11215 vss 0.02f
C11549 vdd.n11216 vss 0.00425f
C11550 vdd.n11217 vss 0.00413f
C11551 vdd.n11218 vss 0.00251f
C11552 vdd.n11219 vss 0.0471f
C11553 vdd.n11220 vss 0.00251f
C11554 vdd.n11221 vss 0.00517f
C11555 vdd.n11222 vss 0.00679f
C11556 vdd.n11223 vss 0.00324f
C11557 vdd.n11224 vss 0.00324f
C11558 vdd.n11225 vss 0.0132f
C11559 vdd.n11226 vss 0.0424f
C11560 vdd.n11227 vss 0.02f
C11561 vdd.n11228 vss 0.00425f
C11562 vdd.n11229 vss 0.0471f
C11563 vdd.n11231 vss 0.00425f
C11564 vdd.n11232 vss 0.00925f
C11565 vdd.n11233 vss 0.00679f
C11566 vdd.n11234 vss 0.00517f
C11567 vdd.n11235 vss 0.00251f
C11568 vdd.n11236 vss 0.0471f
C11569 vdd.n11237 vss 0.00251f
C11570 vdd.n11238 vss 0.0112f
C11571 vdd.n11239 vss 0.0128f
C11572 vdd.n11240 vss 0.146f
C11573 vdd.n11241 vss 0.00324f
C11574 vdd.n11242 vss 0.0112f
C11575 vdd.n11243 vss 0.0128f
C11576 vdd.n11244 vss 0.00413f
C11577 vdd.n11245 vss 0.00413f
C11578 vdd.n11246 vss 0.0471f
C11579 vdd.n11247 vss 0.0471f
C11580 vdd.n11248 vss 0.00324f
C11581 vdd.n11249 vss 0.00413f
C11582 vdd.n11250 vss 0.00413f
C11583 vdd.n11251 vss 0.00679f
C11584 vdd.n11252 vss 0.00413f
C11585 vdd.n11253 vss 0.0471f
C11586 vdd.n11254 vss 0.00324f
C11587 vdd.n11256 vss 0.00925f
C11588 vdd.n11257 vss 0.0471f
C11589 vdd.n11258 vss 0.00425f
C11590 vdd.n11259 vss 0.0424f
C11591 vdd.n11260 vss 0.0132f
C11592 vdd.n11261 vss 0.00324f
C11593 vdd.n11262 vss 0.0128f
C11594 vdd.n11263 vss 0.02f
C11595 vdd.n11264 vss 0.00425f
C11596 vdd.n11265 vss 0.00413f
C11597 vdd.n11266 vss 0.00251f
C11598 vdd.n11267 vss 0.0471f
C11599 vdd.n11268 vss 0.00251f
C11600 vdd.n11269 vss 0.00517f
C11601 vdd.n11270 vss 0.00679f
C11602 vdd.n11271 vss 0.00324f
C11603 vdd.n11272 vss 0.00324f
C11604 vdd.n11273 vss 0.0132f
C11605 vdd.n11274 vss 0.0424f
C11606 vdd.n11275 vss 0.02f
C11607 vdd.n11276 vss 0.00425f
C11608 vdd.n11277 vss 0.0471f
C11609 vdd.n11279 vss 0.00425f
C11610 vdd.n11280 vss 0.00925f
C11611 vdd.n11281 vss 0.00679f
C11612 vdd.n11282 vss 0.00517f
C11613 vdd.n11283 vss 0.00251f
C11614 vdd.n11284 vss 0.0471f
C11615 vdd.n11285 vss 0.00251f
C11616 vdd.n11286 vss 0.0112f
C11617 vdd.n11287 vss 0.0128f
C11618 vdd.n11288 vss 0.146f
C11619 vdd.n11289 vss 0.0596f
C11620 vdd.n11290 vss 0.00324f
C11621 vdd.n11291 vss 0.0112f
C11622 vdd.n11292 vss 0.0128f
C11623 vdd.n11293 vss 0.00413f
C11624 vdd.n11294 vss 0.00413f
C11625 vdd.n11295 vss 0.0471f
C11626 vdd.n11296 vss 0.0471f
C11627 vdd.n11297 vss 0.00324f
C11628 vdd.n11298 vss 0.00413f
C11629 vdd.n11299 vss 0.00413f
C11630 vdd.n11300 vss 0.00679f
C11631 vdd.n11301 vss 0.00413f
C11632 vdd.n11302 vss 0.0471f
C11633 vdd.n11303 vss 0.00324f
C11634 vdd.n11305 vss 0.00925f
C11635 vdd.n11306 vss 0.0471f
C11636 vdd.n11307 vss 0.00425f
C11637 vdd.n11308 vss 0.0424f
C11638 vdd.n11309 vss 0.0132f
C11639 vdd.n11310 vss 0.00324f
C11640 vdd.n11311 vss 0.0128f
C11641 vdd.n11312 vss 0.02f
C11642 vdd.n11313 vss 0.00425f
C11643 vdd.n11314 vss 0.00413f
C11644 vdd.n11315 vss 0.00251f
C11645 vdd.n11316 vss 0.0471f
C11646 vdd.n11317 vss 0.00251f
C11647 vdd.n11318 vss 0.00517f
C11648 vdd.n11319 vss 0.00679f
C11649 vdd.n11320 vss 0.00324f
C11650 vdd.n11321 vss 0.00324f
C11651 vdd.n11322 vss 0.0132f
C11652 vdd.n11323 vss 0.0424f
C11653 vdd.n11324 vss 0.02f
C11654 vdd.n11325 vss 0.00425f
C11655 vdd.n11326 vss 0.0471f
C11656 vdd.n11328 vss 0.00425f
C11657 vdd.n11329 vss 0.00925f
C11658 vdd.n11330 vss 0.00679f
C11659 vdd.n11331 vss 0.00517f
C11660 vdd.n11332 vss 0.00251f
C11661 vdd.n11333 vss 0.0471f
C11662 vdd.n11334 vss 0.00251f
C11663 vdd.n11335 vss 0.0112f
C11664 vdd.n11336 vss 0.0128f
C11665 vdd.n11337 vss 0.0692f
C11666 vdd.n11338 vss 0.118f
C11667 vdd.n11339 vss 0.121f
C11668 vdd.n11340 vss 0.00324f
C11669 vdd.n11341 vss 0.0112f
C11670 vdd.n11342 vss 0.0128f
C11671 vdd.n11343 vss 0.00413f
C11672 vdd.n11344 vss 0.00413f
C11673 vdd.n11345 vss 0.0471f
C11674 vdd.n11346 vss 0.0471f
C11675 vdd.n11347 vss 0.00324f
C11676 vdd.n11348 vss 0.00413f
C11677 vdd.n11349 vss 0.00413f
C11678 vdd.n11350 vss 0.00679f
C11679 vdd.n11351 vss 0.00413f
C11680 vdd.n11352 vss 0.0471f
C11681 vdd.n11353 vss 0.00324f
C11682 vdd.n11355 vss 0.00925f
C11683 vdd.n11356 vss 0.0471f
C11684 vdd.n11357 vss 0.00425f
C11685 vdd.n11358 vss 0.0424f
C11686 vdd.n11359 vss 0.0132f
C11687 vdd.n11360 vss 0.00324f
C11688 vdd.n11361 vss 0.0128f
C11689 vdd.n11362 vss 0.02f
C11690 vdd.n11363 vss 0.00425f
C11691 vdd.n11364 vss 0.00413f
C11692 vdd.n11365 vss 0.00251f
C11693 vdd.n11366 vss 0.0471f
C11694 vdd.n11367 vss 0.00251f
C11695 vdd.n11368 vss 0.00517f
C11696 vdd.n11369 vss 0.00679f
C11697 vdd.n11370 vss 0.00324f
C11698 vdd.n11371 vss 0.00324f
C11699 vdd.n11372 vss 0.0132f
C11700 vdd.n11373 vss 0.0424f
C11701 vdd.n11374 vss 0.02f
C11702 vdd.n11375 vss 0.00425f
C11703 vdd.n11376 vss 0.0471f
C11704 vdd.n11378 vss 0.00425f
C11705 vdd.n11379 vss 0.00925f
C11706 vdd.n11380 vss 0.00679f
C11707 vdd.n11381 vss 0.00517f
C11708 vdd.n11382 vss 0.00251f
C11709 vdd.n11383 vss 0.0471f
C11710 vdd.n11384 vss 0.00251f
C11711 vdd.n11385 vss 0.0112f
C11712 vdd.n11386 vss 0.098f
C11713 vdd.n11387 vss 0.0596f
C11714 vdd.n11388 vss 0.00324f
C11715 vdd.n11389 vss 0.0112f
C11716 vdd.n11390 vss 0.0128f
C11717 vdd.n11391 vss 0.00413f
C11718 vdd.n11392 vss 0.00413f
C11719 vdd.n11393 vss 0.0471f
C11720 vdd.n11394 vss 0.0471f
C11721 vdd.n11395 vss 0.00324f
C11722 vdd.n11396 vss 0.00413f
C11723 vdd.n11397 vss 0.00413f
C11724 vdd.n11398 vss 0.00679f
C11725 vdd.n11399 vss 0.00413f
C11726 vdd.n11400 vss 0.0471f
C11727 vdd.n11401 vss 0.00324f
C11728 vdd.n11403 vss 0.00925f
C11729 vdd.n11404 vss 0.0471f
C11730 vdd.n11405 vss 0.00425f
C11731 vdd.n11406 vss 0.0424f
C11732 vdd.n11407 vss 0.0132f
C11733 vdd.n11408 vss 0.00324f
C11734 vdd.n11409 vss 0.0128f
C11735 vdd.n11410 vss 0.02f
C11736 vdd.n11411 vss 0.00425f
C11737 vdd.n11412 vss 0.00413f
C11738 vdd.n11413 vss 0.00251f
C11739 vdd.n11414 vss 0.0471f
C11740 vdd.n11415 vss 0.00251f
C11741 vdd.n11416 vss 0.00517f
C11742 vdd.n11417 vss 0.00679f
C11743 vdd.n11418 vss 0.00324f
C11744 vdd.n11419 vss 0.00324f
C11745 vdd.n11420 vss 0.0132f
C11746 vdd.n11421 vss 0.0424f
C11747 vdd.n11422 vss 0.02f
C11748 vdd.n11423 vss 0.00425f
C11749 vdd.n11424 vss 0.0471f
C11750 vdd.n11426 vss 0.00425f
C11751 vdd.n11427 vss 0.00925f
C11752 vdd.n11428 vss 0.00679f
C11753 vdd.n11429 vss 0.00517f
C11754 vdd.n11430 vss 0.00251f
C11755 vdd.n11431 vss 0.0471f
C11756 vdd.n11432 vss 0.00251f
C11757 vdd.n11433 vss 0.0112f
C11758 vdd.n11434 vss 0.0128f
C11759 vdd.n11435 vss 0.0692f
C11760 vdd.n11436 vss 0.121f
C11761 vdd.n11437 vss 0.32f
C11762 vdd.n11438 vss 0.202f
C11763 vdd.n11439 vss 0.00324f
C11764 vdd.n11440 vss 0.0112f
C11765 vdd.n11441 vss 0.0128f
C11766 vdd.n11442 vss 0.00413f
C11767 vdd.n11443 vss 0.00413f
C11768 vdd.n11444 vss 0.0471f
C11769 vdd.n11445 vss 0.0471f
C11770 vdd.n11446 vss 0.00324f
C11771 vdd.n11447 vss 0.00413f
C11772 vdd.n11448 vss 0.00413f
C11773 vdd.n11449 vss 0.00679f
C11774 vdd.n11450 vss 0.00413f
C11775 vdd.n11451 vss 0.0471f
C11776 vdd.n11452 vss 0.00324f
C11777 vdd.n11453 vss 0.0424f
C11778 vdd.n11454 vss 0.00324f
C11779 vdd.n11455 vss 0.0128f
C11780 vdd.n11456 vss 0.02f
C11781 vdd.n11457 vss 0.0132f
C11782 vdd.n11458 vss 0.00925f
C11783 vdd.n11459 vss 0.00425f
C11784 vdd.n11461 vss 0.0471f
C11785 vdd.n11462 vss 0.00425f
C11786 vdd.n11463 vss 0.00413f
C11787 vdd.n11464 vss 0.00251f
C11788 vdd.n11465 vss 0.0471f
C11789 vdd.n11466 vss 0.00251f
C11790 vdd.n11467 vss 0.00517f
C11791 vdd.n11468 vss 0.00679f
C11792 vdd.n11469 vss 0.00324f
C11793 vdd.n11470 vss 0.00324f
C11794 vdd.n11471 vss 0.0132f
C11795 vdd.n11472 vss 0.0424f
C11796 vdd.n11473 vss 0.02f
C11797 vdd.n11474 vss 0.00425f
C11798 vdd.n11476 vss 0.0471f
C11799 vdd.n11477 vss 0.00425f
C11800 vdd.n11478 vss 0.00925f
C11801 vdd.n11479 vss 0.00679f
C11802 vdd.n11480 vss 0.00517f
C11803 vdd.n11481 vss 0.00251f
C11804 vdd.n11482 vss 0.0471f
C11805 vdd.n11483 vss 0.00251f
C11806 vdd.n11484 vss 0.0112f
C11807 vdd.n11485 vss 0.0128f
C11808 vdd.n11486 vss 0.00324f
C11809 vdd.n11487 vss 0.0112f
C11810 vdd.n11488 vss 0.0128f
C11811 vdd.n11489 vss 0.00413f
C11812 vdd.n11490 vss 0.00413f
C11813 vdd.n11491 vss 0.0471f
C11814 vdd.n11492 vss 0.0471f
C11815 vdd.n11493 vss 0.00324f
C11816 vdd.n11494 vss 0.00413f
C11817 vdd.n11495 vss 0.00413f
C11818 vdd.n11496 vss 0.00679f
C11819 vdd.n11497 vss 0.00413f
C11820 vdd.n11498 vss 0.0471f
C11821 vdd.n11499 vss 0.00324f
C11822 vdd.n11500 vss 0.0424f
C11823 vdd.n11501 vss 0.00324f
C11824 vdd.n11502 vss 0.0128f
C11825 vdd.n11503 vss 0.02f
C11826 vdd.n11504 vss 0.0132f
C11827 vdd.n11505 vss 0.00925f
C11828 vdd.n11506 vss 0.00425f
C11829 vdd.n11508 vss 0.0471f
C11830 vdd.n11509 vss 0.00425f
C11831 vdd.n11510 vss 0.00413f
C11832 vdd.n11511 vss 0.00251f
C11833 vdd.n11512 vss 0.0471f
C11834 vdd.n11513 vss 0.00251f
C11835 vdd.n11514 vss 0.00517f
C11836 vdd.n11515 vss 0.00679f
C11837 vdd.n11516 vss 0.00324f
C11838 vdd.n11517 vss 0.00324f
C11839 vdd.n11518 vss 0.0132f
C11840 vdd.n11519 vss 0.0424f
C11841 vdd.n11520 vss 0.02f
C11842 vdd.n11521 vss 0.00425f
C11843 vdd.n11523 vss 0.0471f
C11844 vdd.n11524 vss 0.00425f
C11845 vdd.n11525 vss 0.00925f
C11846 vdd.n11526 vss 0.00679f
C11847 vdd.n11527 vss 0.00517f
C11848 vdd.n11528 vss 0.00251f
C11849 vdd.n11529 vss 0.0471f
C11850 vdd.n11530 vss 0.00251f
C11851 vdd.n11531 vss 0.0112f
C11852 vdd.n11532 vss 0.0128f
C11853 vdd.n11533 vss 0.144f
C11854 vdd.n11534 vss 0.143f
C11855 vdd.n11535 vss 0.0608f
C11856 vdd.n11536 vss 0.00324f
C11857 vdd.n11537 vss 0.0112f
C11858 vdd.n11538 vss 0.0128f
C11859 vdd.n11539 vss 0.00413f
C11860 vdd.n11540 vss 0.00413f
C11861 vdd.n11541 vss 0.0471f
C11862 vdd.n11542 vss 0.0471f
C11863 vdd.n11543 vss 0.00324f
C11864 vdd.n11544 vss 0.00413f
C11865 vdd.n11545 vss 0.00413f
C11866 vdd.n11546 vss 0.00679f
C11867 vdd.n11547 vss 0.00413f
C11868 vdd.n11548 vss 0.0471f
C11869 vdd.n11549 vss 0.00324f
C11870 vdd.n11550 vss 0.0424f
C11871 vdd.n11551 vss 0.00324f
C11872 vdd.n11552 vss 0.0128f
C11873 vdd.n11553 vss 0.02f
C11874 vdd.n11554 vss 0.0132f
C11875 vdd.n11555 vss 0.00925f
C11876 vdd.n11556 vss 0.00425f
C11877 vdd.n11558 vss 0.0471f
C11878 vdd.n11559 vss 0.00425f
C11879 vdd.n11560 vss 0.00413f
C11880 vdd.n11561 vss 0.00251f
C11881 vdd.n11562 vss 0.0471f
C11882 vdd.n11563 vss 0.00251f
C11883 vdd.n11564 vss 0.00517f
C11884 vdd.n11565 vss 0.00679f
C11885 vdd.n11566 vss 0.00324f
C11886 vdd.n11567 vss 0.00324f
C11887 vdd.n11568 vss 0.0132f
C11888 vdd.n11569 vss 0.0424f
C11889 vdd.n11570 vss 0.02f
C11890 vdd.n11571 vss 0.00425f
C11891 vdd.n11573 vss 0.0471f
C11892 vdd.n11574 vss 0.00425f
C11893 vdd.n11575 vss 0.00925f
C11894 vdd.n11576 vss 0.00679f
C11895 vdd.n11577 vss 0.00517f
C11896 vdd.n11578 vss 0.00251f
C11897 vdd.n11579 vss 0.0471f
C11898 vdd.n11580 vss 0.00251f
C11899 vdd.n11581 vss 0.0112f
C11900 vdd.n11582 vss 0.0128f
C11901 vdd.n11583 vss 0.0666f
C11902 vdd.n11584 vss 0.118f
C11903 vdd.n11585 vss 0.121f
C11904 vdd.n11586 vss 0.00324f
C11905 vdd.n11587 vss 0.0112f
C11906 vdd.n11588 vss 0.0128f
C11907 vdd.n11589 vss 0.00413f
C11908 vdd.n11590 vss 0.00413f
C11909 vdd.n11591 vss 0.0471f
C11910 vdd.n11592 vss 0.0471f
C11911 vdd.n11593 vss 0.00324f
C11912 vdd.n11594 vss 0.00413f
C11913 vdd.n11595 vss 0.00413f
C11914 vdd.n11596 vss 0.00679f
C11915 vdd.n11597 vss 0.00413f
C11916 vdd.n11598 vss 0.0471f
C11917 vdd.n11599 vss 0.00324f
C11918 vdd.n11600 vss 0.0424f
C11919 vdd.n11601 vss 0.00324f
C11920 vdd.n11602 vss 0.0128f
C11921 vdd.n11603 vss 0.02f
C11922 vdd.n11604 vss 0.0132f
C11923 vdd.n11605 vss 0.00925f
C11924 vdd.n11606 vss 0.00425f
C11925 vdd.n11608 vss 0.0471f
C11926 vdd.n11609 vss 0.00425f
C11927 vdd.n11610 vss 0.00413f
C11928 vdd.n11611 vss 0.00251f
C11929 vdd.n11612 vss 0.0471f
C11930 vdd.n11613 vss 0.00251f
C11931 vdd.n11614 vss 0.00517f
C11932 vdd.n11615 vss 0.00679f
C11933 vdd.n11616 vss 0.00324f
C11934 vdd.n11617 vss 0.00324f
C11935 vdd.n11618 vss 0.0132f
C11936 vdd.n11619 vss 0.0424f
C11937 vdd.n11620 vss 0.02f
C11938 vdd.n11621 vss 0.00425f
C11939 vdd.n11623 vss 0.0471f
C11940 vdd.n11624 vss 0.00425f
C11941 vdd.n11625 vss 0.00925f
C11942 vdd.n11626 vss 0.00679f
C11943 vdd.n11627 vss 0.00517f
C11944 vdd.n11628 vss 0.00251f
C11945 vdd.n11629 vss 0.0471f
C11946 vdd.n11630 vss 0.00251f
C11947 vdd.n11631 vss 0.0112f
C11948 vdd.n11632 vss 0.0955f
C11949 vdd.n11633 vss 0.0608f
C11950 vdd.n11634 vss 0.00324f
C11951 vdd.n11635 vss 0.0112f
C11952 vdd.n11636 vss 0.0128f
C11953 vdd.n11637 vss 0.00413f
C11954 vdd.n11638 vss 0.00413f
C11955 vdd.n11639 vss 0.0471f
C11956 vdd.n11640 vss 0.0471f
C11957 vdd.n11641 vss 0.00324f
C11958 vdd.n11642 vss 0.00413f
C11959 vdd.n11643 vss 0.00413f
C11960 vdd.n11644 vss 0.00679f
C11961 vdd.n11645 vss 0.00413f
C11962 vdd.n11646 vss 0.0471f
C11963 vdd.n11647 vss 0.00324f
C11964 vdd.n11648 vss 0.0424f
C11965 vdd.n11649 vss 0.00324f
C11966 vdd.n11650 vss 0.0128f
C11967 vdd.n11651 vss 0.02f
C11968 vdd.n11652 vss 0.0132f
C11969 vdd.n11653 vss 0.00925f
C11970 vdd.n11654 vss 0.00425f
C11971 vdd.n11656 vss 0.0471f
C11972 vdd.n11657 vss 0.00425f
C11973 vdd.n11658 vss 0.00413f
C11974 vdd.n11659 vss 0.00251f
C11975 vdd.n11660 vss 0.0471f
C11976 vdd.n11661 vss 0.00251f
C11977 vdd.n11662 vss 0.00517f
C11978 vdd.n11663 vss 0.00679f
C11979 vdd.n11664 vss 0.00324f
C11980 vdd.n11665 vss 0.00324f
C11981 vdd.n11666 vss 0.0132f
C11982 vdd.n11667 vss 0.0424f
C11983 vdd.n11668 vss 0.02f
C11984 vdd.n11669 vss 0.00425f
C11985 vdd.n11671 vss 0.0471f
C11986 vdd.n11672 vss 0.00425f
C11987 vdd.n11673 vss 0.00925f
C11988 vdd.n11674 vss 0.00679f
C11989 vdd.n11675 vss 0.00517f
C11990 vdd.n11676 vss 0.00251f
C11991 vdd.n11677 vss 0.0471f
C11992 vdd.n11678 vss 0.00251f
C11993 vdd.n11679 vss 0.0112f
C11994 vdd.n11680 vss 0.0128f
C11995 vdd.n11681 vss 0.0666f
C11996 vdd.n11682 vss 0.0912f
C11997 vdd.n11683 vss 0.0824f
C11998 vdd.n11684 vss 0.0567f
C11999 vdd.n11685 vss 0.00324f
C12000 vdd.n11686 vss 0.0112f
C12001 vdd.n11687 vss 0.0128f
C12002 vdd.n11688 vss 0.00413f
C12003 vdd.n11689 vss 0.00413f
C12004 vdd.n11690 vss 0.0471f
C12005 vdd.n11691 vss 0.0471f
C12006 vdd.n11692 vss 0.00324f
C12007 vdd.n11693 vss 0.00413f
C12008 vdd.n11694 vss 0.00413f
C12009 vdd.n11695 vss 0.00679f
C12010 vdd.n11696 vss 0.00413f
C12011 vdd.n11697 vss 0.0471f
C12012 vdd.n11698 vss 0.00324f
C12013 vdd.n11699 vss 0.0424f
C12014 vdd.n11700 vss 0.00324f
C12015 vdd.n11701 vss 0.0128f
C12016 vdd.n11702 vss 0.02f
C12017 vdd.n11703 vss 0.0132f
C12018 vdd.n11704 vss 0.00925f
C12019 vdd.n11705 vss 0.00425f
C12020 vdd.n11707 vss 0.0471f
C12021 vdd.n11708 vss 0.00425f
C12022 vdd.n11709 vss 0.00413f
C12023 vdd.n11710 vss 0.00251f
C12024 vdd.n11711 vss 0.0471f
C12025 vdd.n11712 vss 0.00251f
C12026 vdd.n11713 vss 0.00517f
C12027 vdd.n11714 vss 0.00679f
C12028 vdd.n11715 vss 0.00324f
C12029 vdd.n11716 vss 0.00324f
C12030 vdd.n11717 vss 0.0132f
C12031 vdd.n11718 vss 0.0424f
C12032 vdd.n11719 vss 0.02f
C12033 vdd.n11720 vss 0.00425f
C12034 vdd.n11722 vss 0.0471f
C12035 vdd.n11723 vss 0.00425f
C12036 vdd.n11724 vss 0.00925f
C12037 vdd.n11725 vss 0.00679f
C12038 vdd.n11726 vss 0.00517f
C12039 vdd.n11727 vss 0.00251f
C12040 vdd.n11728 vss 0.0471f
C12041 vdd.n11729 vss 0.00251f
C12042 vdd.n11730 vss 0.0112f
C12043 vdd.n11731 vss 0.0128f
C12044 vdd.n11732 vss 0.00324f
C12045 vdd.n11733 vss 0.0112f
C12046 vdd.n11734 vss 0.0128f
C12047 vdd.n11735 vss 0.00413f
C12048 vdd.n11736 vss 0.00413f
C12049 vdd.n11737 vss 0.0471f
C12050 vdd.n11738 vss 0.0471f
C12051 vdd.n11739 vss 0.00324f
C12052 vdd.n11740 vss 0.00413f
C12053 vdd.n11741 vss 0.00413f
C12054 vdd.n11742 vss 0.00679f
C12055 vdd.n11743 vss 0.00413f
C12056 vdd.n11744 vss 0.0471f
C12057 vdd.n11745 vss 0.00324f
C12058 vdd.n11746 vss 0.0424f
C12059 vdd.n11747 vss 0.00324f
C12060 vdd.n11748 vss 0.0128f
C12061 vdd.n11749 vss 0.02f
C12062 vdd.n11750 vss 0.0132f
C12063 vdd.n11751 vss 0.00925f
C12064 vdd.n11752 vss 0.00425f
C12065 vdd.n11754 vss 0.0471f
C12066 vdd.n11755 vss 0.00425f
C12067 vdd.n11756 vss 0.00413f
C12068 vdd.n11757 vss 0.00251f
C12069 vdd.n11758 vss 0.0471f
C12070 vdd.n11759 vss 0.00251f
C12071 vdd.n11760 vss 0.00517f
C12072 vdd.n11761 vss 0.00679f
C12073 vdd.n11762 vss 0.00324f
C12074 vdd.n11763 vss 0.00324f
C12075 vdd.n11764 vss 0.0132f
C12076 vdd.n11765 vss 0.0424f
C12077 vdd.n11766 vss 0.02f
C12078 vdd.n11767 vss 0.00425f
C12079 vdd.n11769 vss 0.0471f
C12080 vdd.n11770 vss 0.00425f
C12081 vdd.n11771 vss 0.00925f
C12082 vdd.n11772 vss 0.00679f
C12083 vdd.n11773 vss 0.00517f
C12084 vdd.n11774 vss 0.00251f
C12085 vdd.n11775 vss 0.0471f
C12086 vdd.n11776 vss 0.00251f
C12087 vdd.n11777 vss 0.0112f
C12088 vdd.n11778 vss 0.0128f
C12089 vdd.n11779 vss 0.0564f
C12090 vdd.n11780 vss 0.00324f
C12091 vdd.n11781 vss 0.0112f
C12092 vdd.n11782 vss 0.0128f
C12093 vdd.n11783 vss 0.00413f
C12094 vdd.n11784 vss 0.00413f
C12095 vdd.n11785 vss 0.0471f
C12096 vdd.n11786 vss 0.0471f
C12097 vdd.n11787 vss 0.00324f
C12098 vdd.n11788 vss 0.00413f
C12099 vdd.n11789 vss 0.00413f
C12100 vdd.n11790 vss 0.00679f
C12101 vdd.n11791 vss 0.00413f
C12102 vdd.n11792 vss 0.0471f
C12103 vdd.n11793 vss 0.00324f
C12104 vdd.n11794 vss 0.0424f
C12105 vdd.n11795 vss 0.00324f
C12106 vdd.n11796 vss 0.0128f
C12107 vdd.n11797 vss 0.02f
C12108 vdd.n11798 vss 0.0132f
C12109 vdd.n11799 vss 0.00925f
C12110 vdd.n11800 vss 0.00425f
C12111 vdd.n11802 vss 0.0471f
C12112 vdd.n11803 vss 0.00425f
C12113 vdd.n11804 vss 0.00413f
C12114 vdd.n11805 vss 0.00251f
C12115 vdd.n11806 vss 0.0471f
C12116 vdd.n11807 vss 0.00251f
C12117 vdd.n11808 vss 0.00517f
C12118 vdd.n11809 vss 0.00679f
C12119 vdd.n11810 vss 0.00324f
C12120 vdd.n11811 vss 0.00324f
C12121 vdd.n11812 vss 0.0132f
C12122 vdd.n11813 vss 0.0424f
C12123 vdd.n11814 vss 0.02f
C12124 vdd.n11815 vss 0.00425f
C12125 vdd.n11817 vss 0.0471f
C12126 vdd.n11818 vss 0.00425f
C12127 vdd.n11819 vss 0.00925f
C12128 vdd.n11820 vss 0.00679f
C12129 vdd.n11821 vss 0.00517f
C12130 vdd.n11822 vss 0.00251f
C12131 vdd.n11823 vss 0.0471f
C12132 vdd.n11824 vss 0.00251f
C12133 vdd.n11825 vss 0.0112f
C12134 vdd.n11826 vss 0.0128f
C12135 vdd.n11827 vss 0.183f
C12136 vdd.n11828 vss 0.256f
C12137 vdd.n11829 vss 0.12f
C12138 vdd.n11830 vss 0.0608f
C12139 vdd.n11831 vss 0.00324f
C12140 vdd.n11832 vss 0.0112f
C12141 vdd.n11833 vss 0.0128f
C12142 vdd.n11834 vss 0.00413f
C12143 vdd.n11835 vss 0.00413f
C12144 vdd.n11836 vss 0.0471f
C12145 vdd.n11837 vss 0.0471f
C12146 vdd.n11838 vss 0.00324f
C12147 vdd.n11839 vss 0.00413f
C12148 vdd.n11840 vss 0.00413f
C12149 vdd.n11841 vss 0.00679f
C12150 vdd.n11842 vss 0.00413f
C12151 vdd.n11843 vss 0.0471f
C12152 vdd.n11844 vss 0.00324f
C12153 vdd.n11845 vss 0.0424f
C12154 vdd.n11846 vss 0.00324f
C12155 vdd.n11847 vss 0.0128f
C12156 vdd.n11848 vss 0.02f
C12157 vdd.n11849 vss 0.0132f
C12158 vdd.n11850 vss 0.00925f
C12159 vdd.n11851 vss 0.00425f
C12160 vdd.n11853 vss 0.0471f
C12161 vdd.n11854 vss 0.00425f
C12162 vdd.n11855 vss 0.00413f
C12163 vdd.n11856 vss 0.00251f
C12164 vdd.n11857 vss 0.0471f
C12165 vdd.n11858 vss 0.00251f
C12166 vdd.n11859 vss 0.00517f
C12167 vdd.n11860 vss 0.00679f
C12168 vdd.n11861 vss 0.00324f
C12169 vdd.n11862 vss 0.00324f
C12170 vdd.n11863 vss 0.0132f
C12171 vdd.n11864 vss 0.0424f
C12172 vdd.n11865 vss 0.02f
C12173 vdd.n11866 vss 0.00425f
C12174 vdd.n11868 vss 0.0471f
C12175 vdd.n11869 vss 0.00425f
C12176 vdd.n11870 vss 0.00925f
C12177 vdd.n11871 vss 0.00679f
C12178 vdd.n11872 vss 0.00517f
C12179 vdd.n11873 vss 0.00251f
C12180 vdd.n11874 vss 0.0471f
C12181 vdd.n11875 vss 0.00251f
C12182 vdd.n11876 vss 0.0112f
C12183 vdd.n11877 vss 0.0128f
C12184 vdd.n11878 vss 0.0666f
C12185 vdd.n11879 vss 0.118f
C12186 vdd.n11880 vss 0.121f
C12187 vdd.n11881 vss 0.00324f
C12188 vdd.n11882 vss 0.0112f
C12189 vdd.n11883 vss 0.0128f
C12190 vdd.n11884 vss 0.00413f
C12191 vdd.n11885 vss 0.00413f
C12192 vdd.n11886 vss 0.0471f
C12193 vdd.n11887 vss 0.0471f
C12194 vdd.n11888 vss 0.00324f
C12195 vdd.n11889 vss 0.00413f
C12196 vdd.n11890 vss 0.00413f
C12197 vdd.n11891 vss 0.00679f
C12198 vdd.n11892 vss 0.00413f
C12199 vdd.n11893 vss 0.0471f
C12200 vdd.n11894 vss 0.00324f
C12201 vdd.n11895 vss 0.0424f
C12202 vdd.n11896 vss 0.00324f
C12203 vdd.n11897 vss 0.0128f
C12204 vdd.n11898 vss 0.02f
C12205 vdd.n11899 vss 0.0132f
C12206 vdd.n11900 vss 0.00925f
C12207 vdd.n11901 vss 0.00425f
C12208 vdd.n11903 vss 0.0471f
C12209 vdd.n11904 vss 0.00425f
C12210 vdd.n11905 vss 0.00413f
C12211 vdd.n11906 vss 0.00251f
C12212 vdd.n11907 vss 0.0471f
C12213 vdd.n11908 vss 0.00251f
C12214 vdd.n11909 vss 0.00517f
C12215 vdd.n11910 vss 0.00679f
C12216 vdd.n11911 vss 0.00324f
C12217 vdd.n11912 vss 0.00324f
C12218 vdd.n11913 vss 0.0132f
C12219 vdd.n11914 vss 0.0424f
C12220 vdd.n11915 vss 0.02f
C12221 vdd.n11916 vss 0.00425f
C12222 vdd.n11918 vss 0.0471f
C12223 vdd.n11919 vss 0.00425f
C12224 vdd.n11920 vss 0.00925f
C12225 vdd.n11921 vss 0.00679f
C12226 vdd.n11922 vss 0.00517f
C12227 vdd.n11923 vss 0.00251f
C12228 vdd.n11924 vss 0.0471f
C12229 vdd.n11925 vss 0.00251f
C12230 vdd.n11926 vss 0.0112f
C12231 vdd.n11927 vss 0.0955f
C12232 vdd.n11928 vss 0.0608f
C12233 vdd.n11929 vss 0.00324f
C12234 vdd.n11930 vss 0.0112f
C12235 vdd.n11931 vss 0.0128f
C12236 vdd.n11932 vss 0.00413f
C12237 vdd.n11933 vss 0.00413f
C12238 vdd.n11934 vss 0.0471f
C12239 vdd.n11935 vss 0.0471f
C12240 vdd.n11936 vss 0.00324f
C12241 vdd.n11937 vss 0.00413f
C12242 vdd.n11938 vss 0.00413f
C12243 vdd.n11939 vss 0.00679f
C12244 vdd.n11940 vss 0.00413f
C12245 vdd.n11941 vss 0.0471f
C12246 vdd.n11942 vss 0.00324f
C12247 vdd.n11943 vss 0.0424f
C12248 vdd.n11944 vss 0.00324f
C12249 vdd.n11945 vss 0.0128f
C12250 vdd.n11946 vss 0.02f
C12251 vdd.n11947 vss 0.0132f
C12252 vdd.n11948 vss 0.00925f
C12253 vdd.n11949 vss 0.00425f
C12254 vdd.n11951 vss 0.0471f
C12255 vdd.n11952 vss 0.00425f
C12256 vdd.n11953 vss 0.00413f
C12257 vdd.n11954 vss 0.00251f
C12258 vdd.n11955 vss 0.0471f
C12259 vdd.n11956 vss 0.00251f
C12260 vdd.n11957 vss 0.00517f
C12261 vdd.n11958 vss 0.00679f
C12262 vdd.n11959 vss 0.00324f
C12263 vdd.n11960 vss 0.00324f
C12264 vdd.n11961 vss 0.0132f
C12265 vdd.n11962 vss 0.0424f
C12266 vdd.n11963 vss 0.02f
C12267 vdd.n11964 vss 0.00425f
C12268 vdd.n11966 vss 0.0471f
C12269 vdd.n11967 vss 0.00425f
C12270 vdd.n11968 vss 0.00925f
C12271 vdd.n11969 vss 0.00679f
C12272 vdd.n11970 vss 0.00517f
C12273 vdd.n11971 vss 0.00251f
C12274 vdd.n11972 vss 0.0471f
C12275 vdd.n11973 vss 0.00251f
C12276 vdd.n11974 vss 0.0112f
C12277 vdd.n11975 vss 0.0128f
C12278 vdd.n11976 vss 0.0666f
C12279 vdd.n11977 vss 0.118f
C12280 vdd.n11978 vss 0.0935f
C12281 vdd.n11979 vss 0.00324f
C12282 vdd.n11980 vss 0.0112f
C12283 vdd.n11981 vss 0.0128f
C12284 vdd.n11982 vss 0.00413f
C12285 vdd.n11983 vss 0.00413f
C12286 vdd.n11984 vss 0.0471f
C12287 vdd.n11985 vss 0.0471f
C12288 vdd.n11986 vss 0.00324f
C12289 vdd.n11987 vss 0.00413f
C12290 vdd.n11988 vss 0.00413f
C12291 vdd.n11989 vss 0.00679f
C12292 vdd.n11990 vss 0.00413f
C12293 vdd.n11991 vss 0.0471f
C12294 vdd.n11992 vss 0.00324f
C12295 vdd.n11993 vss 0.0424f
C12296 vdd.n11994 vss 0.00324f
C12297 vdd.n11995 vss 0.0128f
C12298 vdd.n11996 vss 0.02f
C12299 vdd.n11997 vss 0.0132f
C12300 vdd.n11998 vss 0.00925f
C12301 vdd.n11999 vss 0.00425f
C12302 vdd.n12001 vss 0.0471f
C12303 vdd.n12002 vss 0.00425f
C12304 vdd.n12003 vss 0.00413f
C12305 vdd.n12004 vss 0.00251f
C12306 vdd.n12005 vss 0.0471f
C12307 vdd.n12006 vss 0.00251f
C12308 vdd.n12007 vss 0.00517f
C12309 vdd.n12008 vss 0.00679f
C12310 vdd.n12009 vss 0.00324f
C12311 vdd.n12010 vss 0.00324f
C12312 vdd.n12011 vss 0.0132f
C12313 vdd.n12012 vss 0.0424f
C12314 vdd.n12013 vss 0.02f
C12315 vdd.n12014 vss 0.00425f
C12316 vdd.n12016 vss 0.0471f
C12317 vdd.n12017 vss 0.00425f
C12318 vdd.n12018 vss 0.00925f
C12319 vdd.n12019 vss 0.00679f
C12320 vdd.n12020 vss 0.00517f
C12321 vdd.n12021 vss 0.00251f
C12322 vdd.n12022 vss 0.0471f
C12323 vdd.n12023 vss 0.00251f
C12324 vdd.n12024 vss 0.0112f
C12325 vdd.n12025 vss 0.0128f
C12326 vdd.n12026 vss 0.00324f
C12327 vdd.n12027 vss 0.0112f
C12328 vdd.n12028 vss 0.0128f
C12329 vdd.n12029 vss 0.00413f
C12330 vdd.n12030 vss 0.00413f
C12331 vdd.n12031 vss 0.0471f
C12332 vdd.n12032 vss 0.0471f
C12333 vdd.n12033 vss 0.00324f
C12334 vdd.n12034 vss 0.00413f
C12335 vdd.n12035 vss 0.00413f
C12336 vdd.n12036 vss 0.00679f
C12337 vdd.n12037 vss 0.00413f
C12338 vdd.n12038 vss 0.0471f
C12339 vdd.n12039 vss 0.00324f
C12340 vdd.n12040 vss 0.0424f
C12341 vdd.n12041 vss 0.00324f
C12342 vdd.n12042 vss 0.0128f
C12343 vdd.n12043 vss 0.02f
C12344 vdd.n12044 vss 0.0132f
C12345 vdd.n12045 vss 0.00925f
C12346 vdd.n12046 vss 0.00425f
C12347 vdd.n12048 vss 0.0471f
C12348 vdd.n12049 vss 0.00425f
C12349 vdd.n12050 vss 0.00413f
C12350 vdd.n12051 vss 0.00251f
C12351 vdd.n12052 vss 0.0471f
C12352 vdd.n12053 vss 0.00251f
C12353 vdd.n12054 vss 0.00517f
C12354 vdd.n12055 vss 0.00679f
C12355 vdd.n12056 vss 0.00324f
C12356 vdd.n12057 vss 0.00324f
C12357 vdd.n12058 vss 0.0132f
C12358 vdd.n12059 vss 0.0424f
C12359 vdd.n12060 vss 0.02f
C12360 vdd.n12061 vss 0.00425f
C12361 vdd.n12063 vss 0.0471f
C12362 vdd.n12064 vss 0.00425f
C12363 vdd.n12065 vss 0.00925f
C12364 vdd.n12066 vss 0.00679f
C12365 vdd.n12067 vss 0.00517f
C12366 vdd.n12068 vss 0.00251f
C12367 vdd.n12069 vss 0.0471f
C12368 vdd.n12070 vss 0.00251f
C12369 vdd.n12071 vss 0.0112f
C12370 vdd.n12072 vss 0.0128f
C12371 vdd.n12073 vss 0.144f
C12372 vdd.n12074 vss 0.143f
C12373 vdd.n12075 vss 0.0608f
C12374 vdd.n12076 vss 0.00324f
C12375 vdd.n12077 vss 0.0112f
C12376 vdd.n12078 vss 0.0128f
C12377 vdd.n12079 vss 0.00413f
C12378 vdd.n12080 vss 0.00413f
C12379 vdd.n12081 vss 0.0471f
C12380 vdd.n12082 vss 0.0471f
C12381 vdd.n12083 vss 0.00324f
C12382 vdd.n12084 vss 0.00413f
C12383 vdd.n12085 vss 0.00413f
C12384 vdd.n12086 vss 0.00679f
C12385 vdd.n12087 vss 0.00413f
C12386 vdd.n12088 vss 0.0471f
C12387 vdd.n12089 vss 0.00324f
C12388 vdd.n12090 vss 0.0424f
C12389 vdd.n12091 vss 0.00324f
C12390 vdd.n12092 vss 0.0128f
C12391 vdd.n12093 vss 0.02f
C12392 vdd.n12094 vss 0.0132f
C12393 vdd.n12095 vss 0.00925f
C12394 vdd.n12096 vss 0.00425f
C12395 vdd.n12098 vss 0.0471f
C12396 vdd.n12099 vss 0.00425f
C12397 vdd.n12100 vss 0.00413f
C12398 vdd.n12101 vss 0.00251f
C12399 vdd.n12102 vss 0.0471f
C12400 vdd.n12103 vss 0.00251f
C12401 vdd.n12104 vss 0.00517f
C12402 vdd.n12105 vss 0.00679f
C12403 vdd.n12106 vss 0.00324f
C12404 vdd.n12107 vss 0.00324f
C12405 vdd.n12108 vss 0.0132f
C12406 vdd.n12109 vss 0.0424f
C12407 vdd.n12110 vss 0.02f
C12408 vdd.n12111 vss 0.00425f
C12409 vdd.n12113 vss 0.0471f
C12410 vdd.n12114 vss 0.00425f
C12411 vdd.n12115 vss 0.00925f
C12412 vdd.n12116 vss 0.00679f
C12413 vdd.n12117 vss 0.00517f
C12414 vdd.n12118 vss 0.00251f
C12415 vdd.n12119 vss 0.0471f
C12416 vdd.n12120 vss 0.00251f
C12417 vdd.n12121 vss 0.0112f
C12418 vdd.n12122 vss 0.0128f
C12419 vdd.n12123 vss 0.0666f
C12420 vdd.n12124 vss 0.118f
C12421 vdd.n12125 vss 0.121f
C12422 vdd.n12126 vss 0.00324f
C12423 vdd.n12127 vss 0.0112f
C12424 vdd.n12128 vss 0.0128f
C12425 vdd.n12129 vss 0.00413f
C12426 vdd.n12130 vss 0.00413f
C12427 vdd.n12131 vss 0.0471f
C12428 vdd.n12132 vss 0.0471f
C12429 vdd.n12133 vss 0.00324f
C12430 vdd.n12134 vss 0.00413f
C12431 vdd.n12135 vss 0.00413f
C12432 vdd.n12136 vss 0.00679f
C12433 vdd.n12137 vss 0.00413f
C12434 vdd.n12138 vss 0.0471f
C12435 vdd.n12139 vss 0.00324f
C12436 vdd.n12140 vss 0.0424f
C12437 vdd.n12141 vss 0.00324f
C12438 vdd.n12142 vss 0.0128f
C12439 vdd.n12143 vss 0.02f
C12440 vdd.n12144 vss 0.0132f
C12441 vdd.n12145 vss 0.00925f
C12442 vdd.n12146 vss 0.00425f
C12443 vdd.n12148 vss 0.0471f
C12444 vdd.n12149 vss 0.00425f
C12445 vdd.n12150 vss 0.00413f
C12446 vdd.n12151 vss 0.00251f
C12447 vdd.n12152 vss 0.0471f
C12448 vdd.n12153 vss 0.00251f
C12449 vdd.n12154 vss 0.00517f
C12450 vdd.n12155 vss 0.00679f
C12451 vdd.n12156 vss 0.00324f
C12452 vdd.n12157 vss 0.00324f
C12453 vdd.n12158 vss 0.0132f
C12454 vdd.n12159 vss 0.0424f
C12455 vdd.n12160 vss 0.02f
C12456 vdd.n12161 vss 0.00425f
C12457 vdd.n12163 vss 0.0471f
C12458 vdd.n12164 vss 0.00425f
C12459 vdd.n12165 vss 0.00925f
C12460 vdd.n12166 vss 0.00679f
C12461 vdd.n12167 vss 0.00517f
C12462 vdd.n12168 vss 0.00251f
C12463 vdd.n12169 vss 0.0471f
C12464 vdd.n12170 vss 0.00251f
C12465 vdd.n12171 vss 0.0112f
C12466 vdd.n12172 vss 0.0955f
C12467 vdd.n12173 vss 0.0608f
C12468 vdd.n12174 vss 0.00324f
C12469 vdd.n12175 vss 0.0112f
C12470 vdd.n12176 vss 0.0128f
C12471 vdd.n12177 vss 0.00413f
C12472 vdd.n12178 vss 0.00413f
C12473 vdd.n12179 vss 0.0471f
C12474 vdd.n12180 vss 0.0471f
C12475 vdd.n12181 vss 0.00324f
C12476 vdd.n12182 vss 0.00413f
C12477 vdd.n12183 vss 0.00413f
C12478 vdd.n12184 vss 0.00679f
C12479 vdd.n12185 vss 0.00413f
C12480 vdd.n12186 vss 0.0471f
C12481 vdd.n12187 vss 0.00324f
C12482 vdd.n12188 vss 0.0424f
C12483 vdd.n12189 vss 0.00324f
C12484 vdd.n12190 vss 0.0128f
C12485 vdd.n12191 vss 0.02f
C12486 vdd.n12192 vss 0.0132f
C12487 vdd.n12193 vss 0.00925f
C12488 vdd.n12194 vss 0.00425f
C12489 vdd.n12196 vss 0.0471f
C12490 vdd.n12197 vss 0.00425f
C12491 vdd.n12198 vss 0.00413f
C12492 vdd.n12199 vss 0.00251f
C12493 vdd.n12200 vss 0.0471f
C12494 vdd.n12201 vss 0.00251f
C12495 vdd.n12202 vss 0.00517f
C12496 vdd.n12203 vss 0.00679f
C12497 vdd.n12204 vss 0.00324f
C12498 vdd.n12205 vss 0.00324f
C12499 vdd.n12206 vss 0.0132f
C12500 vdd.n12207 vss 0.0424f
C12501 vdd.n12208 vss 0.02f
C12502 vdd.n12209 vss 0.00425f
C12503 vdd.n12211 vss 0.0471f
C12504 vdd.n12212 vss 0.00425f
C12505 vdd.n12213 vss 0.00925f
C12506 vdd.n12214 vss 0.00679f
C12507 vdd.n12215 vss 0.00517f
C12508 vdd.n12216 vss 0.00251f
C12509 vdd.n12217 vss 0.0471f
C12510 vdd.n12218 vss 0.00251f
C12511 vdd.n12219 vss 0.0112f
C12512 vdd.n12220 vss 0.0128f
C12513 vdd.n12221 vss 0.0666f
C12514 vdd.n12222 vss 0.0912f
C12515 vdd.n12223 vss 0.0824f
C12516 vdd.n12224 vss 0.0567f
C12517 vdd.n12225 vss 0.00324f
C12518 vdd.n12226 vss 0.0112f
C12519 vdd.n12227 vss 0.0128f
C12520 vdd.n12228 vss 0.00413f
C12521 vdd.n12229 vss 0.00413f
C12522 vdd.n12230 vss 0.0471f
C12523 vdd.n12231 vss 0.0471f
C12524 vdd.n12232 vss 0.00324f
C12525 vdd.n12233 vss 0.00413f
C12526 vdd.n12234 vss 0.00413f
C12527 vdd.n12235 vss 0.00679f
C12528 vdd.n12236 vss 0.00413f
C12529 vdd.n12237 vss 0.0471f
C12530 vdd.n12238 vss 0.00324f
C12531 vdd.n12239 vss 0.0424f
C12532 vdd.n12240 vss 0.00324f
C12533 vdd.n12241 vss 0.0128f
C12534 vdd.n12242 vss 0.02f
C12535 vdd.n12243 vss 0.0132f
C12536 vdd.n12244 vss 0.00925f
C12537 vdd.n12245 vss 0.00425f
C12538 vdd.n12247 vss 0.0471f
C12539 vdd.n12248 vss 0.00425f
C12540 vdd.n12249 vss 0.00413f
C12541 vdd.n12250 vss 0.00251f
C12542 vdd.n12251 vss 0.0471f
C12543 vdd.n12252 vss 0.00251f
C12544 vdd.n12253 vss 0.00517f
C12545 vdd.n12254 vss 0.00679f
C12546 vdd.n12255 vss 0.00324f
C12547 vdd.n12256 vss 0.00324f
C12548 vdd.n12257 vss 0.0132f
C12549 vdd.n12258 vss 0.0424f
C12550 vdd.n12259 vss 0.02f
C12551 vdd.n12260 vss 0.00425f
C12552 vdd.n12262 vss 0.0471f
C12553 vdd.n12263 vss 0.00425f
C12554 vdd.n12264 vss 0.00925f
C12555 vdd.n12265 vss 0.00679f
C12556 vdd.n12266 vss 0.00517f
C12557 vdd.n12267 vss 0.00251f
C12558 vdd.n12268 vss 0.0471f
C12559 vdd.n12269 vss 0.00251f
C12560 vdd.n12270 vss 0.0112f
C12561 vdd.n12271 vss 0.0128f
C12562 vdd.n12272 vss 0.00324f
C12563 vdd.n12273 vss 0.0112f
C12564 vdd.n12274 vss 0.0128f
C12565 vdd.n12275 vss 0.00413f
C12566 vdd.n12276 vss 0.00413f
C12567 vdd.n12277 vss 0.0471f
C12568 vdd.n12278 vss 0.0471f
C12569 vdd.n12279 vss 0.00324f
C12570 vdd.n12280 vss 0.00413f
C12571 vdd.n12281 vss 0.00413f
C12572 vdd.n12282 vss 0.00679f
C12573 vdd.n12283 vss 0.00413f
C12574 vdd.n12284 vss 0.0471f
C12575 vdd.n12285 vss 0.00324f
C12576 vdd.n12286 vss 0.0424f
C12577 vdd.n12287 vss 0.00324f
C12578 vdd.n12288 vss 0.0128f
C12579 vdd.n12289 vss 0.02f
C12580 vdd.n12290 vss 0.0132f
C12581 vdd.n12291 vss 0.00925f
C12582 vdd.n12292 vss 0.00425f
C12583 vdd.n12294 vss 0.0471f
C12584 vdd.n12295 vss 0.00425f
C12585 vdd.n12296 vss 0.00413f
C12586 vdd.n12297 vss 0.00251f
C12587 vdd.n12298 vss 0.0471f
C12588 vdd.n12299 vss 0.00251f
C12589 vdd.n12300 vss 0.00517f
C12590 vdd.n12301 vss 0.00679f
C12591 vdd.n12302 vss 0.00324f
C12592 vdd.n12303 vss 0.00324f
C12593 vdd.n12304 vss 0.0132f
C12594 vdd.n12305 vss 0.0424f
C12595 vdd.n12306 vss 0.02f
C12596 vdd.n12307 vss 0.00425f
C12597 vdd.n12309 vss 0.0471f
C12598 vdd.n12310 vss 0.00425f
C12599 vdd.n12311 vss 0.00925f
C12600 vdd.n12312 vss 0.00679f
C12601 vdd.n12313 vss 0.00517f
C12602 vdd.n12314 vss 0.00251f
C12603 vdd.n12315 vss 0.0471f
C12604 vdd.n12316 vss 0.00251f
C12605 vdd.n12317 vss 0.0112f
C12606 vdd.n12318 vss 0.0128f
C12607 vdd.n12319 vss 0.144f
C12608 vdd.n12320 vss 0.143f
C12609 vdd.n12321 vss 0.0608f
C12610 vdd.n12322 vss 0.00324f
C12611 vdd.n12323 vss 0.0112f
C12612 vdd.n12324 vss 0.0128f
C12613 vdd.n12325 vss 0.00413f
C12614 vdd.n12326 vss 0.00413f
C12615 vdd.n12327 vss 0.0471f
C12616 vdd.n12328 vss 0.0471f
C12617 vdd.n12329 vss 0.00324f
C12618 vdd.n12330 vss 0.00413f
C12619 vdd.n12331 vss 0.00413f
C12620 vdd.n12332 vss 0.00679f
C12621 vdd.n12333 vss 0.00413f
C12622 vdd.n12334 vss 0.0471f
C12623 vdd.n12335 vss 0.00324f
C12624 vdd.n12336 vss 0.0424f
C12625 vdd.n12337 vss 0.00324f
C12626 vdd.n12338 vss 0.0128f
C12627 vdd.n12339 vss 0.02f
C12628 vdd.n12340 vss 0.0132f
C12629 vdd.n12341 vss 0.00925f
C12630 vdd.n12342 vss 0.00425f
C12631 vdd.n12344 vss 0.0471f
C12632 vdd.n12345 vss 0.00425f
C12633 vdd.n12346 vss 0.00413f
C12634 vdd.n12347 vss 0.00251f
C12635 vdd.n12348 vss 0.0471f
C12636 vdd.n12349 vss 0.00251f
C12637 vdd.n12350 vss 0.00517f
C12638 vdd.n12351 vss 0.00679f
C12639 vdd.n12352 vss 0.00324f
C12640 vdd.n12353 vss 0.00324f
C12641 vdd.n12354 vss 0.0132f
C12642 vdd.n12355 vss 0.0424f
C12643 vdd.n12356 vss 0.02f
C12644 vdd.n12357 vss 0.00425f
C12645 vdd.n12359 vss 0.0471f
C12646 vdd.n12360 vss 0.00425f
C12647 vdd.n12361 vss 0.00925f
C12648 vdd.n12362 vss 0.00679f
C12649 vdd.n12363 vss 0.00517f
C12650 vdd.n12364 vss 0.00251f
C12651 vdd.n12365 vss 0.0471f
C12652 vdd.n12366 vss 0.00251f
C12653 vdd.n12367 vss 0.0112f
C12654 vdd.n12368 vss 0.0128f
C12655 vdd.n12369 vss 0.0666f
C12656 vdd.n12370 vss 0.118f
C12657 vdd.n12371 vss 0.121f
C12658 vdd.n12372 vss 0.00324f
C12659 vdd.n12373 vss 0.0112f
C12660 vdd.n12374 vss 0.0128f
C12661 vdd.n12375 vss 0.00413f
C12662 vdd.n12376 vss 0.00413f
C12663 vdd.n12377 vss 0.0471f
C12664 vdd.n12378 vss 0.0471f
C12665 vdd.n12379 vss 0.00324f
C12666 vdd.n12380 vss 0.00413f
C12667 vdd.n12381 vss 0.00413f
C12668 vdd.n12382 vss 0.00679f
C12669 vdd.n12383 vss 0.00413f
C12670 vdd.n12384 vss 0.0471f
C12671 vdd.n12385 vss 0.00324f
C12672 vdd.n12386 vss 0.0424f
C12673 vdd.n12387 vss 0.00324f
C12674 vdd.n12388 vss 0.0128f
C12675 vdd.n12389 vss 0.02f
C12676 vdd.n12390 vss 0.0132f
C12677 vdd.n12391 vss 0.00925f
C12678 vdd.n12392 vss 0.00425f
C12679 vdd.n12394 vss 0.0471f
C12680 vdd.n12395 vss 0.00425f
C12681 vdd.n12396 vss 0.00413f
C12682 vdd.n12397 vss 0.00251f
C12683 vdd.n12398 vss 0.0471f
C12684 vdd.n12399 vss 0.00251f
C12685 vdd.n12400 vss 0.00517f
C12686 vdd.n12401 vss 0.00679f
C12687 vdd.n12402 vss 0.00324f
C12688 vdd.n12403 vss 0.00324f
C12689 vdd.n12404 vss 0.0132f
C12690 vdd.n12405 vss 0.0424f
C12691 vdd.n12406 vss 0.02f
C12692 vdd.n12407 vss 0.00425f
C12693 vdd.n12409 vss 0.0471f
C12694 vdd.n12410 vss 0.00425f
C12695 vdd.n12411 vss 0.00925f
C12696 vdd.n12412 vss 0.00679f
C12697 vdd.n12413 vss 0.00517f
C12698 vdd.n12414 vss 0.00251f
C12699 vdd.n12415 vss 0.0471f
C12700 vdd.n12416 vss 0.00251f
C12701 vdd.n12417 vss 0.0112f
C12702 vdd.n12418 vss 0.0955f
C12703 vdd.n12419 vss 0.0608f
C12704 vdd.n12420 vss 0.00324f
C12705 vdd.n12421 vss 0.0112f
C12706 vdd.n12422 vss 0.0128f
C12707 vdd.n12423 vss 0.00413f
C12708 vdd.n12424 vss 0.00413f
C12709 vdd.n12425 vss 0.0471f
C12710 vdd.n12426 vss 0.0471f
C12711 vdd.n12427 vss 0.00324f
C12712 vdd.n12428 vss 0.00413f
C12713 vdd.n12429 vss 0.00413f
C12714 vdd.n12430 vss 0.00679f
C12715 vdd.n12431 vss 0.00413f
C12716 vdd.n12432 vss 0.0471f
C12717 vdd.n12433 vss 0.00324f
C12718 vdd.n12434 vss 0.0424f
C12719 vdd.n12435 vss 0.00324f
C12720 vdd.n12436 vss 0.0128f
C12721 vdd.n12437 vss 0.02f
C12722 vdd.n12438 vss 0.0132f
C12723 vdd.n12439 vss 0.00925f
C12724 vdd.n12440 vss 0.00425f
C12725 vdd.n12442 vss 0.0471f
C12726 vdd.n12443 vss 0.00425f
C12727 vdd.n12444 vss 0.00413f
C12728 vdd.n12445 vss 0.00251f
C12729 vdd.n12446 vss 0.0471f
C12730 vdd.n12447 vss 0.00251f
C12731 vdd.n12448 vss 0.00517f
C12732 vdd.n12449 vss 0.00679f
C12733 vdd.n12450 vss 0.00324f
C12734 vdd.n12451 vss 0.00324f
C12735 vdd.n12452 vss 0.0132f
C12736 vdd.n12453 vss 0.0424f
C12737 vdd.n12454 vss 0.02f
C12738 vdd.n12455 vss 0.00425f
C12739 vdd.n12457 vss 0.0471f
C12740 vdd.n12458 vss 0.00425f
C12741 vdd.n12459 vss 0.00925f
C12742 vdd.n12460 vss 0.00679f
C12743 vdd.n12461 vss 0.00517f
C12744 vdd.n12462 vss 0.00251f
C12745 vdd.n12463 vss 0.0471f
C12746 vdd.n12464 vss 0.00251f
C12747 vdd.n12465 vss 0.0112f
C12748 vdd.n12466 vss 0.0128f
C12749 vdd.n12467 vss 0.0666f
C12750 vdd.n12468 vss 0.299f
C12751 vdd.n12469 vss 0.262f
C12752 vdd.n12470 vss 0.0471f
C12753 vdd.n12471 vss 0.00324f
C12754 vdd.n12472 vss 0.00324f
C12755 vdd.n12473 vss 0.0471f
C12756 vdd.n12474 vss 0.00324f
C12757 vdd.n12475 vss 0.00324f
C12758 vdd.n12476 vss 0.0424f
C12759 vdd.n12477 vss 0.0132f
C12760 vdd.n12478 vss 0.00925f
C12761 vdd.n12479 vss 0.00425f
C12762 vdd.n12480 vss 0.0471f
C12763 vdd.n12482 vss 0.00425f
C12764 vdd.n12483 vss 0.02f
C12765 vdd.n12484 vss 0.0128f
C12766 vdd.n12485 vss 0.00413f
C12767 vdd.n12486 vss 0.00413f
C12768 vdd.n12487 vss 0.00413f
C12769 vdd.n12488 vss 0.00413f
C12770 vdd.n12489 vss 0.00679f
C12771 vdd.n12490 vss 0.00679f
C12772 vdd.n12491 vss 0.00517f
C12773 vdd.n12492 vss 0.00251f
C12774 vdd.n12493 vss 0.0471f
C12775 vdd.n12494 vss 0.00251f
C12776 vdd.n12495 vss 0.0112f
C12777 vdd.n12496 vss 0.0471f
C12778 vdd.n12497 vss 0.00324f
C12779 vdd.n12498 vss 0.00324f
C12780 vdd.n12499 vss 0.0424f
C12781 vdd.n12500 vss 0.0132f
C12782 vdd.n12501 vss 0.00925f
C12783 vdd.n12502 vss 0.00425f
C12784 vdd.n12504 vss 0.0471f
C12785 vdd.n12505 vss 0.00425f
C12786 vdd.n12506 vss 0.02f
C12787 vdd.n12507 vss 0.0128f
C12788 vdd.n12508 vss 0.00413f
C12789 vdd.n12509 vss 0.00413f
C12790 vdd.n12510 vss 0.00679f
C12791 vdd.n12511 vss 0.00517f
C12792 vdd.n12512 vss 0.00251f
C12793 vdd.n12513 vss 0.0471f
C12794 vdd.n12514 vss 0.00251f
C12795 vdd.n12515 vss 0.0112f
C12796 vdd.n12516 vss 0.0128f
C12797 vdd.n12517 vss 0.0624f
C12798 d0.t0 vss 0.0286f
C12799 d0.t1 vss 0.0175f
C12800 d0.n0 vss 0.217f
C12801 d0.t4 vss 0.0286f
C12802 d0.t5 vss 0.0175f
C12803 d0.n1 vss 0.217f
C12804 d0.n2 vss 0.0134f
C12805 d0.t8 vss 0.0286f
C12806 d0.t9 vss 0.0175f
C12807 d0.n3 vss 0.217f
C12808 d0.n4 vss 0.0134f
C12809 d0.t12 vss 0.0286f
C12810 d0.t13 vss 0.0175f
C12811 d0.n5 vss 0.217f
C12812 d0.n6 vss 0.0134f
C12813 d0.t16 vss 0.0286f
C12814 d0.t17 vss 0.0175f
C12815 d0.n7 vss 0.217f
C12816 d0.n8 vss 0.0134f
C12817 d0.t20 vss 0.0286f
C12818 d0.t21 vss 0.0175f
C12819 d0.n9 vss 0.217f
C12820 d0.n10 vss 0.0134f
C12821 d0.t24 vss 0.0286f
C12822 d0.t25 vss 0.0175f
C12823 d0.n11 vss 0.217f
C12824 d0.n12 vss 0.0134f
C12825 d0.t28 vss 0.0286f
C12826 d0.t29 vss 0.0175f
C12827 d0.n13 vss 0.217f
C12828 d0.n14 vss 0.0134f
C12829 d0.t255 vss 0.0175f
C12830 d0.t254 vss 0.0286f
C12831 d0.n15 vss 0.217f
C12832 d0.t253 vss 0.0175f
C12833 d0.t252 vss 0.0286f
C12834 d0.n16 vss 0.217f
C12835 d0.n17 vss 0.46f
C12836 d0.t251 vss 0.0175f
C12837 d0.t250 vss 0.0286f
C12838 d0.n18 vss 0.214f
C12839 d0.n19 vss 0.459f
C12840 d0.t249 vss 0.0175f
C12841 d0.t248 vss 0.0286f
C12842 d0.n20 vss 0.217f
C12843 d0.n21 vss 0.457f
C12844 d0.t247 vss 0.0175f
C12845 d0.t246 vss 0.0286f
C12846 d0.n22 vss 0.217f
C12847 d0.n23 vss 0.459f
C12848 d0.t245 vss 0.0175f
C12849 d0.t244 vss 0.0286f
C12850 d0.n24 vss 0.217f
C12851 d0.n25 vss 0.457f
C12852 d0.t243 vss 0.0175f
C12853 d0.t242 vss 0.0286f
C12854 d0.n26 vss 0.214f
C12855 d0.n27 vss 0.459f
C12856 d0.t241 vss 0.0175f
C12857 d0.t240 vss 0.0286f
C12858 d0.n28 vss 0.217f
C12859 d0.n29 vss 0.457f
C12860 d0.t239 vss 0.0175f
C12861 d0.t238 vss 0.0286f
C12862 d0.n30 vss 0.217f
C12863 d0.n31 vss 0.459f
C12864 d0.t237 vss 0.0175f
C12865 d0.t236 vss 0.0286f
C12866 d0.n32 vss 0.217f
C12867 d0.n33 vss 0.457f
C12868 d0.t235 vss 0.0175f
C12869 d0.t234 vss 0.0286f
C12870 d0.n34 vss 0.214f
C12871 d0.n35 vss 0.459f
C12872 d0.t233 vss 0.0175f
C12873 d0.t232 vss 0.0286f
C12874 d0.n36 vss 0.217f
C12875 d0.n37 vss 0.457f
C12876 d0.t231 vss 0.0175f
C12877 d0.t230 vss 0.0286f
C12878 d0.n38 vss 0.217f
C12879 d0.n39 vss 0.459f
C12880 d0.t229 vss 0.0175f
C12881 d0.t228 vss 0.0286f
C12882 d0.n40 vss 0.217f
C12883 d0.n41 vss 0.457f
C12884 d0.t227 vss 0.0175f
C12885 d0.t226 vss 0.0286f
C12886 d0.n42 vss 0.214f
C12887 d0.n43 vss 0.459f
C12888 d0.t225 vss 0.0175f
C12889 d0.t224 vss 0.0286f
C12890 d0.n44 vss 0.214f
C12891 d0.n45 vss 1.26f
C12892 d0.t192 vss 0.0286f
C12893 d0.t193 vss 0.0175f
C12894 d0.n46 vss 0.217f
C12895 d0.n47 vss 0.143f
C12896 d0.t194 vss 0.0286f
C12897 d0.t195 vss 0.0175f
C12898 d0.n48 vss 0.217f
C12899 d0.n49 vss 0.0134f
C12900 d0.n50 vss 0.459f
C12901 d0.t196 vss 0.0286f
C12902 d0.t197 vss 0.0175f
C12903 d0.n51 vss 0.217f
C12904 d0.n52 vss 0.0134f
C12905 d0.n53 vss 0.457f
C12906 d0.t198 vss 0.0286f
C12907 d0.t199 vss 0.0175f
C12908 d0.n54 vss 0.217f
C12909 d0.n55 vss 0.0134f
C12910 d0.n56 vss 0.459f
C12911 d0.t200 vss 0.0286f
C12912 d0.t201 vss 0.0175f
C12913 d0.n57 vss 0.217f
C12914 d0.n58 vss 0.0134f
C12915 d0.n59 vss 0.457f
C12916 d0.t202 vss 0.0286f
C12917 d0.t203 vss 0.0175f
C12918 d0.n60 vss 0.217f
C12919 d0.n61 vss 0.0134f
C12920 d0.n62 vss 0.459f
C12921 d0.t204 vss 0.0286f
C12922 d0.t205 vss 0.0175f
C12923 d0.n63 vss 0.217f
C12924 d0.n64 vss 0.0134f
C12925 d0.n65 vss 0.457f
C12926 d0.t206 vss 0.0286f
C12927 d0.t207 vss 0.0175f
C12928 d0.n66 vss 0.217f
C12929 d0.n67 vss 0.0134f
C12930 d0.n68 vss 0.459f
C12931 d0.t208 vss 0.0286f
C12932 d0.t209 vss 0.0175f
C12933 d0.n69 vss 0.217f
C12934 d0.n70 vss 0.0134f
C12935 d0.n71 vss 0.457f
C12936 d0.t210 vss 0.0286f
C12937 d0.t211 vss 0.0175f
C12938 d0.n72 vss 0.217f
C12939 d0.n73 vss 0.0134f
C12940 d0.n74 vss 0.459f
C12941 d0.t212 vss 0.0286f
C12942 d0.t213 vss 0.0175f
C12943 d0.n75 vss 0.217f
C12944 d0.n76 vss 0.0134f
C12945 d0.n77 vss 0.457f
C12946 d0.t214 vss 0.0286f
C12947 d0.t215 vss 0.0175f
C12948 d0.n78 vss 0.217f
C12949 d0.n79 vss 0.0134f
C12950 d0.n80 vss 0.459f
C12951 d0.t216 vss 0.0286f
C12952 d0.t217 vss 0.0175f
C12953 d0.n81 vss 0.217f
C12954 d0.n82 vss 0.0134f
C12955 d0.n83 vss 0.457f
C12956 d0.t218 vss 0.0286f
C12957 d0.t219 vss 0.0175f
C12958 d0.n84 vss 0.217f
C12959 d0.n85 vss 0.0134f
C12960 d0.n86 vss 0.459f
C12961 d0.t220 vss 0.0286f
C12962 d0.t221 vss 0.0175f
C12963 d0.n87 vss 0.217f
C12964 d0.n88 vss 0.0134f
C12965 d0.n89 vss 0.457f
C12966 d0.t222 vss 0.0286f
C12967 d0.t223 vss 0.0175f
C12968 d0.n90 vss 0.217f
C12969 d0.n91 vss 0.0134f
C12970 d0.n92 vss 0.358f
C12971 d0.n93 vss 1.44f
C12972 d0.t191 vss 0.0175f
C12973 d0.t190 vss 0.0286f
C12974 d0.n94 vss 0.217f
C12975 d0.t189 vss 0.0175f
C12976 d0.t188 vss 0.0286f
C12977 d0.n95 vss 0.217f
C12978 d0.n96 vss 0.46f
C12979 d0.t187 vss 0.0175f
C12980 d0.t186 vss 0.0286f
C12981 d0.n97 vss 0.214f
C12982 d0.n98 vss 0.459f
C12983 d0.t185 vss 0.0175f
C12984 d0.t184 vss 0.0286f
C12985 d0.n99 vss 0.217f
C12986 d0.n100 vss 0.457f
C12987 d0.t183 vss 0.0175f
C12988 d0.t182 vss 0.0286f
C12989 d0.n101 vss 0.217f
C12990 d0.n102 vss 0.459f
C12991 d0.t181 vss 0.0175f
C12992 d0.t180 vss 0.0286f
C12993 d0.n103 vss 0.217f
C12994 d0.n104 vss 0.457f
C12995 d0.t179 vss 0.0175f
C12996 d0.t178 vss 0.0286f
C12997 d0.n105 vss 0.214f
C12998 d0.n106 vss 0.459f
C12999 d0.t177 vss 0.0175f
C13000 d0.t176 vss 0.0286f
C13001 d0.n107 vss 0.217f
C13002 d0.n108 vss 0.457f
C13003 d0.t175 vss 0.0175f
C13004 d0.t174 vss 0.0286f
C13005 d0.n109 vss 0.217f
C13006 d0.n110 vss 0.459f
C13007 d0.t173 vss 0.0175f
C13008 d0.t172 vss 0.0286f
C13009 d0.n111 vss 0.217f
C13010 d0.n112 vss 0.457f
C13011 d0.t171 vss 0.0175f
C13012 d0.t170 vss 0.0286f
C13013 d0.n113 vss 0.214f
C13014 d0.n114 vss 0.459f
C13015 d0.t169 vss 0.0175f
C13016 d0.t168 vss 0.0286f
C13017 d0.n115 vss 0.217f
C13018 d0.n116 vss 0.457f
C13019 d0.t167 vss 0.0175f
C13020 d0.t166 vss 0.0286f
C13021 d0.n117 vss 0.217f
C13022 d0.n118 vss 0.459f
C13023 d0.t165 vss 0.0175f
C13024 d0.t164 vss 0.0286f
C13025 d0.n119 vss 0.217f
C13026 d0.n120 vss 0.457f
C13027 d0.t163 vss 0.0175f
C13028 d0.t162 vss 0.0286f
C13029 d0.n121 vss 0.214f
C13030 d0.n122 vss 0.459f
C13031 d0.t161 vss 0.0175f
C13032 d0.t160 vss 0.0286f
C13033 d0.n123 vss 0.214f
C13034 d0.n124 vss 0.363f
C13035 d0.n125 vss 1.22f
C13036 d0.t128 vss 0.0286f
C13037 d0.t129 vss 0.0175f
C13038 d0.n126 vss 0.217f
C13039 d0.n127 vss 0.142f
C13040 d0.t130 vss 0.0286f
C13041 d0.t131 vss 0.0175f
C13042 d0.n128 vss 0.217f
C13043 d0.n129 vss 0.0134f
C13044 d0.n130 vss 0.459f
C13045 d0.t132 vss 0.0286f
C13046 d0.t133 vss 0.0175f
C13047 d0.n131 vss 0.217f
C13048 d0.n132 vss 0.0134f
C13049 d0.n133 vss 0.457f
C13050 d0.t134 vss 0.0286f
C13051 d0.t135 vss 0.0175f
C13052 d0.n134 vss 0.217f
C13053 d0.n135 vss 0.0134f
C13054 d0.n136 vss 0.459f
C13055 d0.t136 vss 0.0286f
C13056 d0.t137 vss 0.0175f
C13057 d0.n137 vss 0.217f
C13058 d0.n138 vss 0.0134f
C13059 d0.n139 vss 0.457f
C13060 d0.t138 vss 0.0286f
C13061 d0.t139 vss 0.0175f
C13062 d0.n140 vss 0.217f
C13063 d0.n141 vss 0.0134f
C13064 d0.n142 vss 0.459f
C13065 d0.t140 vss 0.0286f
C13066 d0.t141 vss 0.0175f
C13067 d0.n143 vss 0.217f
C13068 d0.n144 vss 0.0134f
C13069 d0.n145 vss 0.457f
C13070 d0.t142 vss 0.0286f
C13071 d0.t143 vss 0.0175f
C13072 d0.n146 vss 0.217f
C13073 d0.n147 vss 0.0134f
C13074 d0.n148 vss 0.459f
C13075 d0.t144 vss 0.0286f
C13076 d0.t145 vss 0.0175f
C13077 d0.n149 vss 0.217f
C13078 d0.n150 vss 0.0134f
C13079 d0.n151 vss 0.457f
C13080 d0.t146 vss 0.0286f
C13081 d0.t147 vss 0.0175f
C13082 d0.n152 vss 0.217f
C13083 d0.n153 vss 0.0134f
C13084 d0.n154 vss 0.459f
C13085 d0.t148 vss 0.0286f
C13086 d0.t149 vss 0.0175f
C13087 d0.n155 vss 0.217f
C13088 d0.n156 vss 0.0134f
C13089 d0.n157 vss 0.457f
C13090 d0.t150 vss 0.0286f
C13091 d0.t151 vss 0.0175f
C13092 d0.n158 vss 0.217f
C13093 d0.n159 vss 0.0134f
C13094 d0.n160 vss 0.459f
C13095 d0.t152 vss 0.0286f
C13096 d0.t153 vss 0.0175f
C13097 d0.n161 vss 0.217f
C13098 d0.n162 vss 0.0134f
C13099 d0.n163 vss 0.457f
C13100 d0.t154 vss 0.0286f
C13101 d0.t155 vss 0.0175f
C13102 d0.n164 vss 0.217f
C13103 d0.n165 vss 0.0134f
C13104 d0.n166 vss 0.459f
C13105 d0.t156 vss 0.0286f
C13106 d0.t157 vss 0.0175f
C13107 d0.n167 vss 0.217f
C13108 d0.n168 vss 0.0134f
C13109 d0.n169 vss 0.457f
C13110 d0.t158 vss 0.0286f
C13111 d0.t159 vss 0.0175f
C13112 d0.n170 vss 0.217f
C13113 d0.n171 vss 0.0134f
C13114 d0.n172 vss 0.358f
C13115 d0.n173 vss 1.21f
C13116 d0.t127 vss 0.0175f
C13117 d0.t126 vss 0.0286f
C13118 d0.n174 vss 0.217f
C13119 d0.t125 vss 0.0175f
C13120 d0.t124 vss 0.0286f
C13121 d0.n175 vss 0.217f
C13122 d0.n176 vss 0.46f
C13123 d0.t123 vss 0.0175f
C13124 d0.t122 vss 0.0286f
C13125 d0.n177 vss 0.214f
C13126 d0.n178 vss 0.459f
C13127 d0.t121 vss 0.0175f
C13128 d0.t120 vss 0.0286f
C13129 d0.n179 vss 0.217f
C13130 d0.n180 vss 0.457f
C13131 d0.t119 vss 0.0175f
C13132 d0.t118 vss 0.0286f
C13133 d0.n181 vss 0.217f
C13134 d0.n182 vss 0.459f
C13135 d0.t117 vss 0.0175f
C13136 d0.t116 vss 0.0286f
C13137 d0.n183 vss 0.217f
C13138 d0.n184 vss 0.457f
C13139 d0.t115 vss 0.0175f
C13140 d0.t114 vss 0.0286f
C13141 d0.n185 vss 0.214f
C13142 d0.n186 vss 0.459f
C13143 d0.t113 vss 0.0175f
C13144 d0.t112 vss 0.0286f
C13145 d0.n187 vss 0.217f
C13146 d0.n188 vss 0.457f
C13147 d0.t111 vss 0.0175f
C13148 d0.t110 vss 0.0286f
C13149 d0.n189 vss 0.217f
C13150 d0.n190 vss 0.459f
C13151 d0.t109 vss 0.0175f
C13152 d0.t108 vss 0.0286f
C13153 d0.n191 vss 0.217f
C13154 d0.n192 vss 0.457f
C13155 d0.t107 vss 0.0175f
C13156 d0.t106 vss 0.0286f
C13157 d0.n193 vss 0.214f
C13158 d0.n194 vss 0.459f
C13159 d0.t105 vss 0.0175f
C13160 d0.t104 vss 0.0286f
C13161 d0.n195 vss 0.217f
C13162 d0.n196 vss 0.457f
C13163 d0.t103 vss 0.0175f
C13164 d0.t102 vss 0.0286f
C13165 d0.n197 vss 0.217f
C13166 d0.n198 vss 0.459f
C13167 d0.t101 vss 0.0175f
C13168 d0.t100 vss 0.0286f
C13169 d0.n199 vss 0.217f
C13170 d0.n200 vss 0.457f
C13171 d0.t99 vss 0.0175f
C13172 d0.t98 vss 0.0286f
C13173 d0.n201 vss 0.214f
C13174 d0.n202 vss 0.459f
C13175 d0.t97 vss 0.0175f
C13176 d0.t96 vss 0.0286f
C13177 d0.n203 vss 0.214f
C13178 d0.n204 vss 0.363f
C13179 d0.n205 vss 1.22f
C13180 d0.t64 vss 0.0286f
C13181 d0.t65 vss 0.0175f
C13182 d0.n206 vss 0.217f
C13183 d0.n207 vss 0.143f
C13184 d0.t66 vss 0.0286f
C13185 d0.t67 vss 0.0175f
C13186 d0.n208 vss 0.217f
C13187 d0.n209 vss 0.0134f
C13188 d0.n210 vss 0.459f
C13189 d0.t68 vss 0.0286f
C13190 d0.t69 vss 0.0175f
C13191 d0.n211 vss 0.217f
C13192 d0.n212 vss 0.0134f
C13193 d0.n213 vss 0.457f
C13194 d0.t70 vss 0.0286f
C13195 d0.t71 vss 0.0175f
C13196 d0.n214 vss 0.217f
C13197 d0.n215 vss 0.0134f
C13198 d0.n216 vss 0.459f
C13199 d0.t72 vss 0.0286f
C13200 d0.t73 vss 0.0175f
C13201 d0.n217 vss 0.217f
C13202 d0.n218 vss 0.0134f
C13203 d0.n219 vss 0.457f
C13204 d0.t74 vss 0.0286f
C13205 d0.t75 vss 0.0175f
C13206 d0.n220 vss 0.217f
C13207 d0.n221 vss 0.0134f
C13208 d0.n222 vss 0.459f
C13209 d0.t76 vss 0.0286f
C13210 d0.t77 vss 0.0175f
C13211 d0.n223 vss 0.217f
C13212 d0.n224 vss 0.0134f
C13213 d0.n225 vss 0.457f
C13214 d0.t78 vss 0.0286f
C13215 d0.t79 vss 0.0175f
C13216 d0.n226 vss 0.217f
C13217 d0.n227 vss 0.0134f
C13218 d0.n228 vss 0.459f
C13219 d0.t80 vss 0.0286f
C13220 d0.t81 vss 0.0175f
C13221 d0.n229 vss 0.217f
C13222 d0.n230 vss 0.0134f
C13223 d0.n231 vss 0.457f
C13224 d0.t82 vss 0.0286f
C13225 d0.t83 vss 0.0175f
C13226 d0.n232 vss 0.217f
C13227 d0.n233 vss 0.0134f
C13228 d0.n234 vss 0.459f
C13229 d0.t84 vss 0.0286f
C13230 d0.t85 vss 0.0175f
C13231 d0.n235 vss 0.217f
C13232 d0.n236 vss 0.0134f
C13233 d0.n237 vss 0.457f
C13234 d0.t86 vss 0.0286f
C13235 d0.t87 vss 0.0175f
C13236 d0.n238 vss 0.217f
C13237 d0.n239 vss 0.0134f
C13238 d0.n240 vss 0.459f
C13239 d0.t88 vss 0.0286f
C13240 d0.t89 vss 0.0175f
C13241 d0.n241 vss 0.217f
C13242 d0.n242 vss 0.0134f
C13243 d0.n243 vss 0.457f
C13244 d0.t90 vss 0.0286f
C13245 d0.t91 vss 0.0175f
C13246 d0.n244 vss 0.217f
C13247 d0.n245 vss 0.0134f
C13248 d0.n246 vss 0.459f
C13249 d0.t92 vss 0.0286f
C13250 d0.t93 vss 0.0175f
C13251 d0.n247 vss 0.217f
C13252 d0.n248 vss 0.0134f
C13253 d0.n249 vss 0.457f
C13254 d0.t94 vss 0.0286f
C13255 d0.t95 vss 0.0175f
C13256 d0.n250 vss 0.217f
C13257 d0.n251 vss 0.0134f
C13258 d0.n252 vss 0.358f
C13259 d0.n253 vss 1.21f
C13260 d0.t63 vss 0.0175f
C13261 d0.t62 vss 0.0286f
C13262 d0.n254 vss 0.217f
C13263 d0.t61 vss 0.0175f
C13264 d0.t60 vss 0.0286f
C13265 d0.n255 vss 0.217f
C13266 d0.n256 vss 0.46f
C13267 d0.t59 vss 0.0175f
C13268 d0.t58 vss 0.0286f
C13269 d0.n257 vss 0.214f
C13270 d0.n258 vss 0.459f
C13271 d0.t57 vss 0.0175f
C13272 d0.t56 vss 0.0286f
C13273 d0.n259 vss 0.217f
C13274 d0.n260 vss 0.457f
C13275 d0.t55 vss 0.0175f
C13276 d0.t54 vss 0.0286f
C13277 d0.n261 vss 0.217f
C13278 d0.n262 vss 0.459f
C13279 d0.t53 vss 0.0175f
C13280 d0.t52 vss 0.0286f
C13281 d0.n263 vss 0.217f
C13282 d0.n264 vss 0.457f
C13283 d0.t51 vss 0.0175f
C13284 d0.t50 vss 0.0286f
C13285 d0.n265 vss 0.214f
C13286 d0.n266 vss 0.459f
C13287 d0.t49 vss 0.0175f
C13288 d0.t48 vss 0.0286f
C13289 d0.n267 vss 0.217f
C13290 d0.n268 vss 0.457f
C13291 d0.t47 vss 0.0175f
C13292 d0.t46 vss 0.0286f
C13293 d0.n269 vss 0.217f
C13294 d0.n270 vss 0.459f
C13295 d0.t45 vss 0.0175f
C13296 d0.t44 vss 0.0286f
C13297 d0.n271 vss 0.217f
C13298 d0.n272 vss 0.457f
C13299 d0.t43 vss 0.0175f
C13300 d0.t42 vss 0.0286f
C13301 d0.n273 vss 0.214f
C13302 d0.n274 vss 0.459f
C13303 d0.t41 vss 0.0175f
C13304 d0.t40 vss 0.0286f
C13305 d0.n275 vss 0.217f
C13306 d0.n276 vss 0.457f
C13307 d0.t39 vss 0.0175f
C13308 d0.t38 vss 0.0286f
C13309 d0.n277 vss 0.217f
C13310 d0.n278 vss 0.459f
C13311 d0.t37 vss 0.0175f
C13312 d0.t36 vss 0.0286f
C13313 d0.n279 vss 0.217f
C13314 d0.n280 vss 0.457f
C13315 d0.t35 vss 0.0175f
C13316 d0.t34 vss 0.0286f
C13317 d0.n281 vss 0.214f
C13318 d0.n282 vss 0.459f
C13319 d0.t33 vss 0.0175f
C13320 d0.t32 vss 0.0286f
C13321 d0.n283 vss 0.214f
C13322 d0.n284 vss 0.363f
C13323 d0.n285 vss 1.45f
C13324 d0.t30 vss 0.0286f
C13325 d0.t31 vss 0.0175f
C13326 d0.n286 vss 0.217f
C13327 d0.n287 vss 0.0134f
C13328 d0.n288 vss 1.25f
C13329 d0.n289 vss 0.457f
C13330 d0.t26 vss 0.0286f
C13331 d0.t27 vss 0.0175f
C13332 d0.n290 vss 0.217f
C13333 d0.n291 vss 0.0134f
C13334 d0.n292 vss 0.459f
C13335 d0.n293 vss 0.457f
C13336 d0.t22 vss 0.0286f
C13337 d0.t23 vss 0.0175f
C13338 d0.n294 vss 0.217f
C13339 d0.n295 vss 0.0134f
C13340 d0.n296 vss 0.459f
C13341 d0.n297 vss 0.457f
C13342 d0.t18 vss 0.0286f
C13343 d0.t19 vss 0.0175f
C13344 d0.n298 vss 0.217f
C13345 d0.n299 vss 0.0134f
C13346 d0.n300 vss 0.459f
C13347 d0.n301 vss 0.457f
C13348 d0.t14 vss 0.0286f
C13349 d0.t15 vss 0.0175f
C13350 d0.n302 vss 0.217f
C13351 d0.n303 vss 0.0134f
C13352 d0.n304 vss 0.459f
C13353 d0.n305 vss 0.457f
C13354 d0.t10 vss 0.0286f
C13355 d0.t11 vss 0.0175f
C13356 d0.n306 vss 0.217f
C13357 d0.n307 vss 0.0134f
C13358 d0.n308 vss 0.459f
C13359 d0.n309 vss 0.457f
C13360 d0.t6 vss 0.0286f
C13361 d0.t7 vss 0.0175f
C13362 d0.n310 vss 0.217f
C13363 d0.n311 vss 0.0134f
C13364 d0.n312 vss 0.459f
C13365 d0.n313 vss 0.457f
C13366 d0.t2 vss 0.0286f
C13367 d0.t3 vss 0.0175f
C13368 d0.n314 vss 0.217f
C13369 d0.n315 vss 0.0134f
C13370 d0.n316 vss 0.459f
C13371 d0.n317 vss 0.142f
C13372 d7 vss 0.613f
C13373 vout vss 0.2f
C13374 X3/m1_688_n494# vss 0.858f
C13375 X3/m1_994_178# vss 1.15f
C13376 d6 vss 15.5f
C13377 X3/vin2 vss 2.58f
C13378 X2/X3/m1_688_n494# vss 0.856f
C13379 X2/X3/m1_994_178# vss 1.15f
C13380 X2/X3/vin2 vss 2.16f
C13381 X2/X2/X3/m1_688_n494# vss 0.858f
C13382 X2/X2/X3/m1_994_178# vss 1.15f
C13383 X2/X2/X3/vin2 vss 1.27f
C13384 X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13385 X2/X2/X2/X3/m1_994_178# vss 1.15f
C13386 X2/X2/X2/X3/vin2 vss 1.85f
C13387 X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13388 X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C13389 X2/X2/X2/X2/X3/vin2 vss 1.75f
C13390 X2/X2/X2/X2/X2/sw_0/m1_688_n494# vss 0.858f
C13391 X2/X2/X2/X2/X2/sw_0/m1_994_178# vss 1.15f
C13392 X2/X2/X2/X2/X2/X2/vout vss 0.868f
C13393 X2/X2/X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13394 X2/X2/X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C13395 X2/X2/X2/X2/X2/X2/X2/vin1 vss 1.46f
C13396 X2/X2/X2/X2/X2/X2/X3/vin2 vss 1.23f
C13397 X2/X2/X2/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C13398 X2/X2/X2/X2/X2/X2/X2/m1_994_178# vss 1.15f
C13399 vrefl vss 2.39f
C13400 X2/X2/X2/X2/X2/X2/X1/vin1 vss 1.91f
C13401 X2/X2/X2/X2/X2/X2/X3/vin1 vss 0.816f
C13402 X2/X2/X2/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C13403 X2/X2/X2/X2/X2/X2/X1/m1_994_178# vss 1.15f
C13404 X2/X2/X2/X2/X2/X2/X1/vin2 vss 1.73f
C13405 X2/X2/X2/X2/X2/X1/vout vss 0.607f
C13406 X2/X2/X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13407 X2/X2/X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C13408 X2/X2/X2/X2/X2/X1/X2/vin1 vss 1.46f
C13409 X2/X2/X2/X2/X2/X1/X3/vin2 vss 1.23f
C13410 X2/X2/X2/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C13411 X2/X2/X2/X2/X2/X1/X2/m1_994_178# vss 1.15f
C13412 X2/X2/X2/X2/X2/X2/vrefh vss 3.27f
C13413 X2/X2/X2/X2/X2/X1/X1/vin1 vss 1.91f
C13414 X2/X2/X2/X2/X2/X1/X3/vin1 vss 0.816f
C13415 X2/X2/X2/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C13416 X2/X2/X2/X2/X2/X1/X1/m1_994_178# vss 1.15f
C13417 X2/X2/X2/X2/X2/X1/X1/vin2 vss 1.73f
C13418 X2/X2/X2/X2/X3/vin1 vss 1.49f
C13419 X2/X2/X2/X2/X1/sw_0/m1_688_n494# vss 0.858f
C13420 X2/X2/X2/X2/X1/sw_0/m1_994_178# vss 1.15f
C13421 X2/X2/X2/X2/X1/X2/vout vss 0.868f
C13422 X2/X2/X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C13423 X2/X2/X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C13424 X2/X2/X2/X2/X1/X2/X2/vin1 vss 1.46f
C13425 X2/X2/X2/X2/X1/X2/X3/vin2 vss 1.23f
C13426 X2/X2/X2/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C13427 X2/X2/X2/X2/X1/X2/X2/m1_994_178# vss 1.15f
C13428 X2/X2/X2/X2/X2/vrefh vss 3.27f
C13429 X2/X2/X2/X2/X1/X2/X1/vin1 vss 1.91f
C13430 X2/X2/X2/X2/X1/X2/X3/vin1 vss 0.816f
C13431 X2/X2/X2/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C13432 X2/X2/X2/X2/X1/X2/X1/m1_994_178# vss 1.15f
C13433 X2/X2/X2/X2/X1/X2/X1/vin2 vss 1.73f
C13434 X2/X2/X2/X2/X1/X1/vout vss 0.607f
C13435 X2/X2/X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C13436 X2/X2/X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C13437 X2/X2/X2/X2/X1/X1/X2/vin1 vss 1.46f
C13438 X2/X2/X2/X2/X1/X1/X3/vin2 vss 1.23f
C13439 X2/X2/X2/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C13440 X2/X2/X2/X2/X1/X1/X2/m1_994_178# vss 1.15f
C13441 X2/X2/X2/X2/X1/X2/vrefh vss 3.27f
C13442 X2/X2/X2/X2/X1/X1/X1/vin1 vss 1.91f
C13443 X2/X2/X2/X2/X1/X1/X3/vin1 vss 0.816f
C13444 X2/X2/X2/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C13445 X2/X2/X2/X2/X1/X1/X1/m1_994_178# vss 1.15f
C13446 X2/X2/X2/X2/X1/X1/X1/vin2 vss 1.73f
C13447 X2/X2/X2/X3/vin1 vss 1.6f
C13448 X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13449 X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C13450 X2/X2/X2/X1/X3/vin2 vss 1.75f
C13451 X2/X2/X2/X1/X2/sw_0/m1_688_n494# vss 0.858f
C13452 X2/X2/X2/X1/X2/sw_0/m1_994_178# vss 1.15f
C13453 X2/X2/X2/X1/X2/X2/vout vss 0.868f
C13454 X2/X2/X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C13455 X2/X2/X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C13456 X2/X2/X2/X1/X2/X2/X2/vin1 vss 1.46f
C13457 X2/X2/X2/X1/X2/X2/X3/vin2 vss 1.23f
C13458 X2/X2/X2/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C13459 X2/X2/X2/X1/X2/X2/X2/m1_994_178# vss 1.15f
C13460 X2/X2/X2/X2/vrefh vss 3.27f
C13461 X2/X2/X2/X1/X2/X2/X1/vin1 vss 1.91f
C13462 X2/X2/X2/X1/X2/X2/X3/vin1 vss 0.816f
C13463 X2/X2/X2/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C13464 X2/X2/X2/X1/X2/X2/X1/m1_994_178# vss 1.15f
C13465 X2/X2/X2/X1/X2/X2/X1/vin2 vss 1.73f
C13466 X2/X2/X2/X1/X2/X1/vout vss 0.607f
C13467 X2/X2/X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C13468 X2/X2/X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C13469 X2/X2/X2/X1/X2/X1/X2/vin1 vss 1.46f
C13470 X2/X2/X2/X1/X2/X1/X3/vin2 vss 1.23f
C13471 X2/X2/X2/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C13472 X2/X2/X2/X1/X2/X1/X2/m1_994_178# vss 1.15f
C13473 X2/X2/X2/X1/X2/X2/vrefh vss 3.27f
C13474 X2/X2/X2/X1/X2/X1/X1/vin1 vss 1.91f
C13475 X2/X2/X2/X1/X2/X1/X3/vin1 vss 0.816f
C13476 X2/X2/X2/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C13477 X2/X2/X2/X1/X2/X1/X1/m1_994_178# vss 1.15f
C13478 X2/X2/X2/X1/X2/X1/X1/vin2 vss 1.73f
C13479 X2/X2/X2/X1/X3/vin1 vss 1.49f
C13480 X2/X2/X2/X1/X1/sw_0/m1_688_n494# vss 0.858f
C13481 X2/X2/X2/X1/X1/sw_0/m1_994_178# vss 1.15f
C13482 X2/X2/X2/X1/X1/X2/vout vss 0.868f
C13483 X2/X2/X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C13484 X2/X2/X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C13485 X2/X2/X2/X1/X1/X2/X2/vin1 vss 1.46f
C13486 X2/X2/X2/X1/X1/X2/X3/vin2 vss 1.23f
C13487 X2/X2/X2/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C13488 X2/X2/X2/X1/X1/X2/X2/m1_994_178# vss 1.15f
C13489 X2/X2/X2/X1/X2/vrefh vss 3.27f
C13490 X2/X2/X2/X1/X1/X2/X1/vin1 vss 1.91f
C13491 X2/X2/X2/X1/X1/X2/X3/vin1 vss 0.816f
C13492 X2/X2/X2/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C13493 X2/X2/X2/X1/X1/X2/X1/m1_994_178# vss 1.15f
C13494 X2/X2/X2/X1/X1/X2/X1/vin2 vss 1.73f
C13495 X2/X2/X2/X1/X1/X1/vout vss 0.607f
C13496 X2/X2/X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C13497 X2/X2/X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C13498 X2/X2/X2/X1/X1/X1/X2/vin1 vss 1.46f
C13499 X2/X2/X2/X1/X1/X1/X3/vin2 vss 1.23f
C13500 X2/X2/X2/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C13501 X2/X2/X2/X1/X1/X1/X2/m1_994_178# vss 1.15f
C13502 X2/X2/X2/X1/X1/X2/vrefh vss 3.27f
C13503 X2/X2/X2/X1/X1/X1/X1/vin1 vss 1.91f
C13504 X2/X2/X2/X1/X1/X1/X3/vin1 vss 0.816f
C13505 X2/X2/X2/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C13506 X2/X2/X2/X1/X1/X1/X1/m1_994_178# vss 1.15f
C13507 X2/X2/X2/X1/X1/X1/X1/vin2 vss 1.73f
C13508 X2/X2/X3/vin1 vss 1.12f
C13509 X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13510 X2/X2/X1/X3/m1_994_178# vss 1.15f
C13511 X2/X2/X1/X3/vin2 vss 1.85f
C13512 X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C13513 X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C13514 X2/X2/X1/X2/X3/vin2 vss 1.75f
C13515 X2/X2/X1/X2/X2/sw_0/m1_688_n494# vss 0.858f
C13516 X2/X2/X1/X2/X2/sw_0/m1_994_178# vss 1.15f
C13517 X2/X2/X1/X2/X2/X2/vout vss 0.868f
C13518 X2/X2/X1/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13519 X2/X2/X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C13520 X2/X2/X1/X2/X2/X2/X2/vin1 vss 1.46f
C13521 X2/X2/X1/X2/X2/X2/X3/vin2 vss 1.23f
C13522 X2/X2/X1/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C13523 X2/X2/X1/X2/X2/X2/X2/m1_994_178# vss 1.15f
C13524 X2/X2/X2/vrefh vss 6.35f
C13525 X2/X2/X1/X2/X2/X2/X1/vin1 vss 1.91f
C13526 X2/X2/X1/X2/X2/X2/X3/vin1 vss 0.816f
C13527 X2/X2/X1/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C13528 X2/X2/X1/X2/X2/X2/X1/m1_994_178# vss 1.15f
C13529 X2/X2/X1/X2/X2/X2/X1/vin2 vss 1.73f
C13530 X2/X2/X1/X2/X2/X1/vout vss 0.607f
C13531 X2/X2/X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13532 X2/X2/X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C13533 X2/X2/X1/X2/X2/X1/X2/vin1 vss 1.46f
C13534 X2/X2/X1/X2/X2/X1/X3/vin2 vss 1.23f
C13535 X2/X2/X1/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C13536 X2/X2/X1/X2/X2/X1/X2/m1_994_178# vss 1.15f
C13537 X2/X2/X1/X2/X2/X2/vrefh vss 3.27f
C13538 X2/X2/X1/X2/X2/X1/X1/vin1 vss 1.91f
C13539 X2/X2/X1/X2/X2/X1/X3/vin1 vss 0.816f
C13540 X2/X2/X1/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C13541 X2/X2/X1/X2/X2/X1/X1/m1_994_178# vss 1.15f
C13542 X2/X2/X1/X2/X2/X1/X1/vin2 vss 1.73f
C13543 X2/X2/X1/X2/X3/vin1 vss 1.49f
C13544 X2/X2/X1/X2/X1/sw_0/m1_688_n494# vss 0.858f
C13545 X2/X2/X1/X2/X1/sw_0/m1_994_178# vss 1.15f
C13546 X2/X2/X1/X2/X1/X2/vout vss 0.868f
C13547 X2/X2/X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C13548 X2/X2/X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C13549 X2/X2/X1/X2/X1/X2/X2/vin1 vss 1.46f
C13550 X2/X2/X1/X2/X1/X2/X3/vin2 vss 1.23f
C13551 X2/X2/X1/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C13552 X2/X2/X1/X2/X1/X2/X2/m1_994_178# vss 1.15f
C13553 X2/X2/X1/X2/X2/vrefh vss 3.27f
C13554 X2/X2/X1/X2/X1/X2/X1/vin1 vss 1.91f
C13555 X2/X2/X1/X2/X1/X2/X3/vin1 vss 0.816f
C13556 X2/X2/X1/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C13557 X2/X2/X1/X2/X1/X2/X1/m1_994_178# vss 1.15f
C13558 X2/X2/X1/X2/X1/X2/X1/vin2 vss 1.73f
C13559 X2/X2/X1/X2/X1/X1/vout vss 0.607f
C13560 X2/X2/X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C13561 X2/X2/X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C13562 X2/X2/X1/X2/X1/X1/X2/vin1 vss 1.46f
C13563 X2/X2/X1/X2/X1/X1/X3/vin2 vss 1.23f
C13564 X2/X2/X1/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C13565 X2/X2/X1/X2/X1/X1/X2/m1_994_178# vss 1.15f
C13566 X2/X2/X1/X2/X1/X2/vrefh vss 3.27f
C13567 X2/X2/X1/X2/X1/X1/X1/vin1 vss 1.91f
C13568 X2/X2/X1/X2/X1/X1/X3/vin1 vss 0.816f
C13569 X2/X2/X1/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C13570 X2/X2/X1/X2/X1/X1/X1/m1_994_178# vss 1.15f
C13571 X2/X2/X1/X2/X1/X1/X1/vin2 vss 1.73f
C13572 X2/X2/X1/X3/vin1 vss 1.6f
C13573 X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C13574 X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C13575 X2/X2/X1/X1/X3/vin2 vss 1.75f
C13576 X2/X2/X1/X1/X2/sw_0/m1_688_n494# vss 0.858f
C13577 X2/X2/X1/X1/X2/sw_0/m1_994_178# vss 1.15f
C13578 X2/X2/X1/X1/X2/X2/vout vss 0.868f
C13579 X2/X2/X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C13580 X2/X2/X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C13581 X2/X2/X1/X1/X2/X2/X2/vin1 vss 1.46f
C13582 X2/X2/X1/X1/X2/X2/X3/vin2 vss 1.23f
C13583 X2/X2/X1/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C13584 X2/X2/X1/X1/X2/X2/X2/m1_994_178# vss 1.15f
C13585 X2/X2/X1/X2/vrefh vss 3.27f
C13586 X2/X2/X1/X1/X2/X2/X1/vin1 vss 1.91f
C13587 X2/X2/X1/X1/X2/X2/X3/vin1 vss 0.816f
C13588 X2/X2/X1/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C13589 X2/X2/X1/X1/X2/X2/X1/m1_994_178# vss 1.15f
C13590 X2/X2/X1/X1/X2/X2/X1/vin2 vss 1.73f
C13591 X2/X2/X1/X1/X2/X1/vout vss 0.607f
C13592 X2/X2/X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C13593 X2/X2/X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C13594 X2/X2/X1/X1/X2/X1/X2/vin1 vss 1.46f
C13595 X2/X2/X1/X1/X2/X1/X3/vin2 vss 1.23f
C13596 X2/X2/X1/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C13597 X2/X2/X1/X1/X2/X1/X2/m1_994_178# vss 1.15f
C13598 X2/X2/X1/X1/X2/X2/vrefh vss 3.27f
C13599 X2/X2/X1/X1/X2/X1/X1/vin1 vss 1.91f
C13600 X2/X2/X1/X1/X2/X1/X3/vin1 vss 0.816f
C13601 X2/X2/X1/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C13602 X2/X2/X1/X1/X2/X1/X1/m1_994_178# vss 1.15f
C13603 X2/X2/X1/X1/X2/X1/X1/vin2 vss 1.73f
C13604 X2/X2/X1/X1/X3/vin1 vss 1.49f
C13605 X2/X2/X1/X1/X1/sw_0/m1_688_n494# vss 0.858f
C13606 X2/X2/X1/X1/X1/sw_0/m1_994_178# vss 1.15f
C13607 X2/X2/X1/X1/X1/X2/vout vss 0.868f
C13608 X2/X2/X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C13609 X2/X2/X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C13610 X2/X2/X1/X1/X1/X2/X2/vin1 vss 1.46f
C13611 X2/X2/X1/X1/X1/X2/X3/vin2 vss 1.23f
C13612 X2/X2/X1/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C13613 X2/X2/X1/X1/X1/X2/X2/m1_994_178# vss 1.15f
C13614 X2/X2/X1/X1/X2/vrefh vss 3.27f
C13615 X2/X2/X1/X1/X1/X2/X1/vin1 vss 1.91f
C13616 X2/X2/X1/X1/X1/X2/X3/vin1 vss 0.816f
C13617 X2/X2/X1/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C13618 X2/X2/X1/X1/X1/X2/X1/m1_994_178# vss 1.15f
C13619 X2/X2/X1/X1/X1/X2/X1/vin2 vss 1.73f
C13620 X2/X2/X1/X1/X1/X1/vout vss 0.607f
C13621 X2/X2/X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C13622 X2/X2/X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C13623 X2/X2/X1/X1/X1/X1/X2/vin1 vss 1.46f
C13624 X2/X2/X1/X1/X1/X1/X3/vin2 vss 1.23f
C13625 X2/X2/X1/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C13626 X2/X2/X1/X1/X1/X1/X2/m1_994_178# vss 1.15f
C13627 X2/X2/X1/X1/X1/X2/vrefh vss 3.27f
C13628 X2/X2/X1/X1/X1/X1/X1/vin1 vss 1.96f
C13629 X2/X2/X1/X1/X1/X1/X3/vin1 vss 0.816f
C13630 X2/X2/X1/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C13631 X2/X2/X1/X1/X1/X1/X1/m1_994_178# vss 1.15f
C13632 X2/X2/X1/X1/X1/X1/X1/vin2 vss 1.74f
C13633 X2/X3/vin1 vss 1.34f
C13634 X2/X1/X3/m1_688_n494# vss 0.858f
C13635 X2/X1/X3/m1_994_178# vss 1.15f
C13636 X2/X1/X3/vin2 vss 1.27f
C13637 X2/X1/X2/X3/m1_688_n494# vss 0.858f
C13638 X2/X1/X2/X3/m1_994_178# vss 1.15f
C13639 X2/X1/X2/X3/vin2 vss 1.85f
C13640 X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C13641 X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C13642 X2/X1/X2/X2/X3/vin2 vss 1.75f
C13643 X2/X1/X2/X2/X2/sw_0/m1_688_n494# vss 0.858f
C13644 X2/X1/X2/X2/X2/sw_0/m1_994_178# vss 1.15f
C13645 X2/X1/X2/X2/X2/X2/vout vss 0.868f
C13646 X2/X1/X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13647 X2/X1/X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C13648 X2/X1/X2/X2/X2/X2/X2/vin1 vss 1.46f
C13649 X2/X1/X2/X2/X2/X2/X3/vin2 vss 1.24f
C13650 X2/X1/X2/X2/X2/X2/X2/m1_688_n494# vss 0.859f
C13651 X2/X1/X2/X2/X2/X2/X2/m1_994_178# vss 1.15f
C13652 X2/X2/vrefh vss 4.1f
C13653 X2/X1/X2/X2/X2/X2/X1/vin1 vss 1.91f
C13654 X2/X1/X2/X2/X2/X2/X3/vin1 vss 0.816f
C13655 X2/X1/X2/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C13656 X2/X1/X2/X2/X2/X2/X1/m1_994_178# vss 1.15f
C13657 X2/X1/X2/X2/X2/X2/X1/vin2 vss 1.73f
C13658 X2/X1/X2/X2/X2/X1/vout vss 0.607f
C13659 X2/X1/X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13660 X2/X1/X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C13661 X2/X1/X2/X2/X2/X1/X2/vin1 vss 1.46f
C13662 X2/X1/X2/X2/X2/X1/X3/vin2 vss 1.23f
C13663 X2/X1/X2/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C13664 X2/X1/X2/X2/X2/X1/X2/m1_994_178# vss 1.15f
C13665 X2/X1/X2/X2/X2/X2/vrefh vss 3.27f
C13666 X2/X1/X2/X2/X2/X1/X1/vin1 vss 1.91f
C13667 X2/X1/X2/X2/X2/X1/X3/vin1 vss 0.816f
C13668 X2/X1/X2/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C13669 X2/X1/X2/X2/X2/X1/X1/m1_994_178# vss 1.15f
C13670 X2/X1/X2/X2/X2/X1/X1/vin2 vss 1.73f
C13671 X2/X1/X2/X2/X3/vin1 vss 1.49f
C13672 X2/X1/X2/X2/X1/sw_0/m1_688_n494# vss 0.858f
C13673 X2/X1/X2/X2/X1/sw_0/m1_994_178# vss 1.15f
C13674 X2/X1/X2/X2/X1/X2/vout vss 0.868f
C13675 X2/X1/X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C13676 X2/X1/X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C13677 X2/X1/X2/X2/X1/X2/X2/vin1 vss 1.46f
C13678 X2/X1/X2/X2/X1/X2/X3/vin2 vss 1.23f
C13679 X2/X1/X2/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C13680 X2/X1/X2/X2/X1/X2/X2/m1_994_178# vss 1.15f
C13681 X2/X1/X2/X2/X2/vrefh vss 3.27f
C13682 X2/X1/X2/X2/X1/X2/X1/vin1 vss 1.91f
C13683 X2/X1/X2/X2/X1/X2/X3/vin1 vss 0.816f
C13684 X2/X1/X2/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C13685 X2/X1/X2/X2/X1/X2/X1/m1_994_178# vss 1.15f
C13686 X2/X1/X2/X2/X1/X2/X1/vin2 vss 1.73f
C13687 X2/X1/X2/X2/X1/X1/vout vss 0.607f
C13688 X2/X1/X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C13689 X2/X1/X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C13690 X2/X1/X2/X2/X1/X1/X2/vin1 vss 1.46f
C13691 X2/X1/X2/X2/X1/X1/X3/vin2 vss 1.23f
C13692 X2/X1/X2/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C13693 X2/X1/X2/X2/X1/X1/X2/m1_994_178# vss 1.15f
C13694 X2/X1/X2/X2/X1/X2/vrefh vss 3.27f
C13695 X2/X1/X2/X2/X1/X1/X1/vin1 vss 1.91f
C13696 X2/X1/X2/X2/X1/X1/X3/vin1 vss 0.816f
C13697 X2/X1/X2/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C13698 X2/X1/X2/X2/X1/X1/X1/m1_994_178# vss 1.15f
C13699 X2/X1/X2/X2/X1/X1/X1/vin2 vss 1.73f
C13700 X2/X1/X2/X3/vin1 vss 1.6f
C13701 X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C13702 X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C13703 X2/X1/X2/X1/X3/vin2 vss 1.75f
C13704 X2/X1/X2/X1/X2/sw_0/m1_688_n494# vss 0.858f
C13705 X2/X1/X2/X1/X2/sw_0/m1_994_178# vss 1.15f
C13706 X2/X1/X2/X1/X2/X2/vout vss 0.868f
C13707 X2/X1/X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C13708 X2/X1/X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C13709 X2/X1/X2/X1/X2/X2/X2/vin1 vss 1.46f
C13710 X2/X1/X2/X1/X2/X2/X3/vin2 vss 1.23f
C13711 X2/X1/X2/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C13712 X2/X1/X2/X1/X2/X2/X2/m1_994_178# vss 1.15f
C13713 X2/X1/X2/X2/vrefh vss 3.27f
C13714 X2/X1/X2/X1/X2/X2/X1/vin1 vss 1.91f
C13715 X2/X1/X2/X1/X2/X2/X3/vin1 vss 0.816f
C13716 X2/X1/X2/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C13717 X2/X1/X2/X1/X2/X2/X1/m1_994_178# vss 1.15f
C13718 X2/X1/X2/X1/X2/X2/X1/vin2 vss 1.73f
C13719 X2/X1/X2/X1/X2/X1/vout vss 0.607f
C13720 X2/X1/X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C13721 X2/X1/X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C13722 X2/X1/X2/X1/X2/X1/X2/vin1 vss 1.46f
C13723 X2/X1/X2/X1/X2/X1/X3/vin2 vss 1.23f
C13724 X2/X1/X2/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C13725 X2/X1/X2/X1/X2/X1/X2/m1_994_178# vss 1.15f
C13726 X2/X1/X2/X1/X2/X2/vrefh vss 3.27f
C13727 X2/X1/X2/X1/X2/X1/X1/vin1 vss 1.91f
C13728 X2/X1/X2/X1/X2/X1/X3/vin1 vss 0.816f
C13729 X2/X1/X2/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C13730 X2/X1/X2/X1/X2/X1/X1/m1_994_178# vss 1.15f
C13731 X2/X1/X2/X1/X2/X1/X1/vin2 vss 1.73f
C13732 X2/X1/X2/X1/X3/vin1 vss 1.49f
C13733 X2/X1/X2/X1/X1/sw_0/m1_688_n494# vss 0.858f
C13734 X2/X1/X2/X1/X1/sw_0/m1_994_178# vss 1.15f
C13735 X2/X1/X2/X1/X1/X2/vout vss 0.868f
C13736 X2/X1/X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C13737 X2/X1/X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C13738 X2/X1/X2/X1/X1/X2/X2/vin1 vss 1.46f
C13739 X2/X1/X2/X1/X1/X2/X3/vin2 vss 1.23f
C13740 X2/X1/X2/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C13741 X2/X1/X2/X1/X1/X2/X2/m1_994_178# vss 1.15f
C13742 X2/X1/X2/X1/X2/vrefh vss 3.27f
C13743 X2/X1/X2/X1/X1/X2/X1/vin1 vss 1.91f
C13744 X2/X1/X2/X1/X1/X2/X3/vin1 vss 0.816f
C13745 X2/X1/X2/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C13746 X2/X1/X2/X1/X1/X2/X1/m1_994_178# vss 1.15f
C13747 X2/X1/X2/X1/X1/X2/X1/vin2 vss 1.73f
C13748 X2/X1/X2/X1/X1/X1/vout vss 0.607f
C13749 X2/X1/X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C13750 X2/X1/X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C13751 X2/X1/X2/X1/X1/X1/X2/vin1 vss 1.46f
C13752 X2/X1/X2/X1/X1/X1/X3/vin2 vss 1.23f
C13753 X2/X1/X2/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C13754 X2/X1/X2/X1/X1/X1/X2/m1_994_178# vss 1.15f
C13755 X2/X1/X2/X1/X1/X2/vrefh vss 3.27f
C13756 X2/X1/X2/X1/X1/X1/X1/vin1 vss 1.91f
C13757 X2/X1/X2/X1/X1/X1/X3/vin1 vss 0.816f
C13758 X2/X1/X2/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C13759 X2/X1/X2/X1/X1/X1/X1/m1_994_178# vss 1.15f
C13760 X2/X1/X2/X1/X1/X1/X1/vin2 vss 1.73f
C13761 X2/X1/X3/vin1 vss 1.12f
C13762 X2/X1/X1/X3/m1_688_n494# vss 0.858f
C13763 X2/X1/X1/X3/m1_994_178# vss 1.15f
C13764 X2/X1/X1/X3/vin2 vss 1.85f
C13765 X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C13766 X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C13767 X2/X1/X1/X2/X3/vin2 vss 1.75f
C13768 X2/X1/X1/X2/X2/sw_0/m1_688_n494# vss 0.858f
C13769 X2/X1/X1/X2/X2/sw_0/m1_994_178# vss 1.15f
C13770 X2/X1/X1/X2/X2/X2/vout vss 0.868f
C13771 X2/X1/X1/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13772 X2/X1/X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C13773 X2/X1/X1/X2/X2/X2/X2/vin1 vss 1.46f
C13774 X2/X1/X1/X2/X2/X2/X3/vin2 vss 1.23f
C13775 X2/X1/X1/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C13776 X2/X1/X1/X2/X2/X2/X2/m1_994_178# vss 1.15f
C13777 X2/X1/X2/vrefh vss 6.36f
C13778 X2/X1/X1/X2/X2/X2/X1/vin1 vss 1.91f
C13779 X2/X1/X1/X2/X2/X2/X3/vin1 vss 0.816f
C13780 X2/X1/X1/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C13781 X2/X1/X1/X2/X2/X2/X1/m1_994_178# vss 1.15f
C13782 X2/X1/X1/X2/X2/X2/X1/vin2 vss 1.74f
C13783 X2/X1/X1/X2/X2/X1/vout vss 0.607f
C13784 X2/X1/X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13785 X2/X1/X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C13786 X2/X1/X1/X2/X2/X1/X2/vin1 vss 1.46f
C13787 X2/X1/X1/X2/X2/X1/X3/vin2 vss 1.23f
C13788 X2/X1/X1/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C13789 X2/X1/X1/X2/X2/X1/X2/m1_994_178# vss 1.15f
C13790 X2/X1/X1/X2/X2/X2/vrefh vss 3.27f
C13791 X2/X1/X1/X2/X2/X1/X1/vin1 vss 1.91f
C13792 X2/X1/X1/X2/X2/X1/X3/vin1 vss 0.816f
C13793 X2/X1/X1/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C13794 X2/X1/X1/X2/X2/X1/X1/m1_994_178# vss 1.15f
C13795 X2/X1/X1/X2/X2/X1/X1/vin2 vss 1.74f
C13796 X2/X1/X1/X2/X3/vin1 vss 1.49f
C13797 X2/X1/X1/X2/X1/sw_0/m1_688_n494# vss 0.858f
C13798 X2/X1/X1/X2/X1/sw_0/m1_994_178# vss 1.15f
C13799 X2/X1/X1/X2/X1/X2/vout vss 0.868f
C13800 X2/X1/X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C13801 X2/X1/X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C13802 X2/X1/X1/X2/X1/X2/X2/vin1 vss 1.46f
C13803 X2/X1/X1/X2/X1/X2/X3/vin2 vss 1.23f
C13804 X2/X1/X1/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C13805 X2/X1/X1/X2/X1/X2/X2/m1_994_178# vss 1.15f
C13806 X2/X1/X1/X2/X2/vrefh vss 3.27f
C13807 X2/X1/X1/X2/X1/X2/X1/vin1 vss 1.91f
C13808 X2/X1/X1/X2/X1/X2/X3/vin1 vss 0.816f
C13809 X2/X1/X1/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C13810 X2/X1/X1/X2/X1/X2/X1/m1_994_178# vss 1.15f
C13811 X2/X1/X1/X2/X1/X2/X1/vin2 vss 1.74f
C13812 X2/X1/X1/X2/X1/X1/vout vss 0.607f
C13813 X2/X1/X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C13814 X2/X1/X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C13815 X2/X1/X1/X2/X1/X1/X2/vin1 vss 1.46f
C13816 X2/X1/X1/X2/X1/X1/X3/vin2 vss 1.23f
C13817 X2/X1/X1/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C13818 X2/X1/X1/X2/X1/X1/X2/m1_994_178# vss 1.15f
C13819 X2/X1/X1/X2/X1/X2/vrefh vss 3.27f
C13820 X2/X1/X1/X2/X1/X1/X1/vin1 vss 1.91f
C13821 X2/X1/X1/X2/X1/X1/X3/vin1 vss 0.816f
C13822 X2/X1/X1/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C13823 X2/X1/X1/X2/X1/X1/X1/m1_994_178# vss 1.15f
C13824 X2/X1/X1/X2/X1/X1/X1/vin2 vss 1.74f
C13825 X2/X1/X1/X3/vin1 vss 1.6f
C13826 X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C13827 X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C13828 X2/X1/X1/X1/X3/vin2 vss 1.75f
C13829 X2/X1/X1/X1/X2/sw_0/m1_688_n494# vss 0.858f
C13830 X2/X1/X1/X1/X2/sw_0/m1_994_178# vss 1.15f
C13831 X2/X1/X1/X1/X2/X2/vout vss 0.868f
C13832 X2/X1/X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C13833 X2/X1/X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C13834 X2/X1/X1/X1/X2/X2/X2/vin1 vss 1.46f
C13835 X2/X1/X1/X1/X2/X2/X3/vin2 vss 1.23f
C13836 X2/X1/X1/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C13837 X2/X1/X1/X1/X2/X2/X2/m1_994_178# vss 1.15f
C13838 X2/X1/X1/X2/vrefh vss 3.27f
C13839 X2/X1/X1/X1/X2/X2/X1/vin1 vss 1.91f
C13840 X2/X1/X1/X1/X2/X2/X3/vin1 vss 0.816f
C13841 X2/X1/X1/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C13842 X2/X1/X1/X1/X2/X2/X1/m1_994_178# vss 1.15f
C13843 X2/X1/X1/X1/X2/X2/X1/vin2 vss 1.74f
C13844 X2/X1/X1/X1/X2/X1/vout vss 0.607f
C13845 X2/X1/X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C13846 X2/X1/X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C13847 X2/X1/X1/X1/X2/X1/X2/vin1 vss 1.46f
C13848 X2/X1/X1/X1/X2/X1/X3/vin2 vss 1.23f
C13849 X2/X1/X1/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C13850 X2/X1/X1/X1/X2/X1/X2/m1_994_178# vss 1.15f
C13851 X2/X1/X1/X1/X2/X2/vrefh vss 3.27f
C13852 X2/X1/X1/X1/X2/X1/X1/vin1 vss 1.91f
C13853 X2/X1/X1/X1/X2/X1/X3/vin1 vss 0.816f
C13854 X2/X1/X1/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C13855 X2/X1/X1/X1/X2/X1/X1/m1_994_178# vss 1.15f
C13856 X2/X1/X1/X1/X2/X1/X1/vin2 vss 1.74f
C13857 X2/X1/X1/X1/X3/vin1 vss 1.49f
C13858 X2/X1/X1/X1/X1/sw_0/m1_688_n494# vss 0.858f
C13859 X2/X1/X1/X1/X1/sw_0/m1_994_178# vss 1.15f
C13860 X2/X1/X1/X1/X1/X2/vout vss 0.868f
C13861 X2/X1/X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C13862 X2/X1/X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C13863 X2/X1/X1/X1/X1/X2/X2/vin1 vss 1.46f
C13864 X2/X1/X1/X1/X1/X2/X3/vin2 vss 1.23f
C13865 X2/X1/X1/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C13866 X2/X1/X1/X1/X1/X2/X2/m1_994_178# vss 1.15f
C13867 X2/X1/X1/X1/X2/vrefh vss 3.27f
C13868 X2/X1/X1/X1/X1/X2/X1/vin1 vss 1.91f
C13869 X2/X1/X1/X1/X1/X2/X3/vin1 vss 0.816f
C13870 X2/X1/X1/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C13871 X2/X1/X1/X1/X1/X2/X1/m1_994_178# vss 1.15f
C13872 X2/X1/X1/X1/X1/X2/X1/vin2 vss 1.74f
C13873 X2/X1/X1/X1/X1/X1/vout vss 0.607f
C13874 X2/X1/X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C13875 X2/X1/X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C13876 X2/X1/X1/X1/X1/X1/X2/vin1 vss 1.46f
C13877 X2/X1/X1/X1/X1/X1/X3/vin2 vss 1.23f
C13878 X2/X1/X1/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C13879 X2/X1/X1/X1/X1/X1/X2/m1_994_178# vss 1.15f
C13880 X2/X1/X1/X1/X1/X2/vrefh vss 3.27f
C13881 X2/X1/X1/X1/X1/X1/X1/vin1 vss 1.96f
C13882 X2/X1/X1/X1/X1/X1/X3/vin1 vss 0.816f
C13883 X2/X1/X1/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C13884 X2/X1/X1/X1/X1/X1/X1/m1_994_178# vss 1.15f
C13885 X2/X1/X1/X1/X1/X1/X1/vin2 vss 1.74f
C13886 X3/vin1 vss 1.77f
C13887 X1/X3/m1_688_n494# vss 0.856f
C13888 X1/X3/m1_994_178# vss 1.15f
C13889 d5 vss 12.5f
C13890 X1/X3/vin2 vss 2.16f
C13891 X1/X2/X3/m1_688_n494# vss 0.858f
C13892 X1/X2/X3/m1_994_178# vss 1.15f
C13893 X1/X2/X3/vin2 vss 1.27f
C13894 X1/X2/X2/X3/m1_688_n494# vss 0.858f
C13895 X1/X2/X2/X3/m1_994_178# vss 1.15f
C13896 X1/X2/X2/X3/vin2 vss 1.85f
C13897 X1/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13898 X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C13899 X1/X2/X2/X2/X3/vin2 vss 1.75f
C13900 X1/X2/X2/X2/X2/sw_0/m1_688_n494# vss 0.858f
C13901 X1/X2/X2/X2/X2/sw_0/m1_994_178# vss 1.15f
C13902 X1/X2/X2/X2/X2/X2/vout vss 0.868f
C13903 X1/X2/X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C13904 X1/X2/X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C13905 X1/X2/X2/X2/X2/X2/X2/vin1 vss 1.46f
C13906 X1/X2/X2/X2/X2/X2/X3/vin2 vss 1.24f
C13907 X1/X2/X2/X2/X2/X2/X2/m1_688_n494# vss 0.859f
C13908 X1/X2/X2/X2/X2/X2/X2/m1_994_178# vss 1.15f
C13909 X2/vrefh vss 3.92f
C13910 X1/X2/X2/X2/X2/X2/X1/vin1 vss 1.91f
C13911 X1/X2/X2/X2/X2/X2/X3/vin1 vss 0.816f
C13912 X1/X2/X2/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C13913 X1/X2/X2/X2/X2/X2/X1/m1_994_178# vss 1.15f
C13914 X1/X2/X2/X2/X2/X2/X1/vin2 vss 1.74f
C13915 X1/X2/X2/X2/X2/X1/vout vss 0.607f
C13916 X1/X2/X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13917 X1/X2/X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C13918 X1/X2/X2/X2/X2/X1/X2/vin1 vss 1.46f
C13919 X1/X2/X2/X2/X2/X1/X3/vin2 vss 1.23f
C13920 X1/X2/X2/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C13921 X1/X2/X2/X2/X2/X1/X2/m1_994_178# vss 1.15f
C13922 X1/X2/X2/X2/X2/X2/vrefh vss 3.27f
C13923 X1/X2/X2/X2/X2/X1/X1/vin1 vss 1.91f
C13924 X1/X2/X2/X2/X2/X1/X3/vin1 vss 0.816f
C13925 X1/X2/X2/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C13926 X1/X2/X2/X2/X2/X1/X1/m1_994_178# vss 1.15f
C13927 X1/X2/X2/X2/X2/X1/X1/vin2 vss 1.74f
C13928 X1/X2/X2/X2/X3/vin1 vss 1.49f
C13929 X1/X2/X2/X2/X1/sw_0/m1_688_n494# vss 0.858f
C13930 X1/X2/X2/X2/X1/sw_0/m1_994_178# vss 1.15f
C13931 X1/X2/X2/X2/X1/X2/vout vss 0.868f
C13932 X1/X2/X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C13933 X1/X2/X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C13934 X1/X2/X2/X2/X1/X2/X2/vin1 vss 1.46f
C13935 X1/X2/X2/X2/X1/X2/X3/vin2 vss 1.23f
C13936 X1/X2/X2/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C13937 X1/X2/X2/X2/X1/X2/X2/m1_994_178# vss 1.15f
C13938 X1/X2/X2/X2/X2/vrefh vss 3.27f
C13939 X1/X2/X2/X2/X1/X2/X1/vin1 vss 1.91f
C13940 X1/X2/X2/X2/X1/X2/X3/vin1 vss 0.816f
C13941 X1/X2/X2/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C13942 X1/X2/X2/X2/X1/X2/X1/m1_994_178# vss 1.15f
C13943 X1/X2/X2/X2/X1/X2/X1/vin2 vss 1.74f
C13944 X1/X2/X2/X2/X1/X1/vout vss 0.607f
C13945 X1/X2/X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C13946 X1/X2/X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C13947 X1/X2/X2/X2/X1/X1/X2/vin1 vss 1.46f
C13948 X1/X2/X2/X2/X1/X1/X3/vin2 vss 1.23f
C13949 X1/X2/X2/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C13950 X1/X2/X2/X2/X1/X1/X2/m1_994_178# vss 1.15f
C13951 X1/X2/X2/X2/X1/X2/vrefh vss 3.27f
C13952 X1/X2/X2/X2/X1/X1/X1/vin1 vss 1.91f
C13953 X1/X2/X2/X2/X1/X1/X3/vin1 vss 0.816f
C13954 X1/X2/X2/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C13955 X1/X2/X2/X2/X1/X1/X1/m1_994_178# vss 1.15f
C13956 X1/X2/X2/X2/X1/X1/X1/vin2 vss 1.74f
C13957 X1/X2/X2/X3/vin1 vss 1.6f
C13958 X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C13959 X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C13960 X1/X2/X2/X1/X3/vin2 vss 1.75f
C13961 X1/X2/X2/X1/X2/sw_0/m1_688_n494# vss 0.858f
C13962 X1/X2/X2/X1/X2/sw_0/m1_994_178# vss 1.15f
C13963 X1/X2/X2/X1/X2/X2/vout vss 0.868f
C13964 X1/X2/X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C13965 X1/X2/X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C13966 X1/X2/X2/X1/X2/X2/X2/vin1 vss 1.46f
C13967 X1/X2/X2/X1/X2/X2/X3/vin2 vss 1.23f
C13968 X1/X2/X2/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C13969 X1/X2/X2/X1/X2/X2/X2/m1_994_178# vss 1.15f
C13970 X1/X2/X2/X2/vrefh vss 3.27f
C13971 X1/X2/X2/X1/X2/X2/X1/vin1 vss 1.91f
C13972 X1/X2/X2/X1/X2/X2/X3/vin1 vss 0.816f
C13973 X1/X2/X2/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C13974 X1/X2/X2/X1/X2/X2/X1/m1_994_178# vss 1.15f
C13975 X1/X2/X2/X1/X2/X2/X1/vin2 vss 1.74f
C13976 X1/X2/X2/X1/X2/X1/vout vss 0.607f
C13977 X1/X2/X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C13978 X1/X2/X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C13979 X1/X2/X2/X1/X2/X1/X2/vin1 vss 1.46f
C13980 X1/X2/X2/X1/X2/X1/X3/vin2 vss 1.23f
C13981 X1/X2/X2/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C13982 X1/X2/X2/X1/X2/X1/X2/m1_994_178# vss 1.15f
C13983 X1/X2/X2/X1/X2/X2/vrefh vss 3.27f
C13984 X1/X2/X2/X1/X2/X1/X1/vin1 vss 1.91f
C13985 X1/X2/X2/X1/X2/X1/X3/vin1 vss 0.816f
C13986 X1/X2/X2/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C13987 X1/X2/X2/X1/X2/X1/X1/m1_994_178# vss 1.15f
C13988 X1/X2/X2/X1/X2/X1/X1/vin2 vss 1.74f
C13989 X1/X2/X2/X1/X3/vin1 vss 1.49f
C13990 X1/X2/X2/X1/X1/sw_0/m1_688_n494# vss 0.858f
C13991 X1/X2/X2/X1/X1/sw_0/m1_994_178# vss 1.15f
C13992 X1/X2/X2/X1/X1/X2/vout vss 0.868f
C13993 X1/X2/X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C13994 X1/X2/X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C13995 X1/X2/X2/X1/X1/X2/X2/vin1 vss 1.46f
C13996 X1/X2/X2/X1/X1/X2/X3/vin2 vss 1.23f
C13997 X1/X2/X2/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C13998 X1/X2/X2/X1/X1/X2/X2/m1_994_178# vss 1.15f
C13999 X1/X2/X2/X1/X2/vrefh vss 3.27f
C14000 X1/X2/X2/X1/X1/X2/X1/vin1 vss 1.91f
C14001 X1/X2/X2/X1/X1/X2/X3/vin1 vss 0.816f
C14002 X1/X2/X2/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C14003 X1/X2/X2/X1/X1/X2/X1/m1_994_178# vss 1.15f
C14004 X1/X2/X2/X1/X1/X2/X1/vin2 vss 1.74f
C14005 X1/X2/X2/X1/X1/X1/vout vss 0.607f
C14006 X1/X2/X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C14007 X1/X2/X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C14008 X1/X2/X2/X1/X1/X1/X2/vin1 vss 1.46f
C14009 X1/X2/X2/X1/X1/X1/X3/vin2 vss 1.23f
C14010 X1/X2/X2/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C14011 X1/X2/X2/X1/X1/X1/X2/m1_994_178# vss 1.15f
C14012 X1/X2/X2/X1/X1/X2/vrefh vss 3.27f
C14013 X1/X2/X2/X1/X1/X1/X1/vin1 vss 1.91f
C14014 X1/X2/X2/X1/X1/X1/X3/vin1 vss 0.816f
C14015 X1/X2/X2/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C14016 X1/X2/X2/X1/X1/X1/X1/m1_994_178# vss 1.15f
C14017 X1/X2/X2/X1/X1/X1/X1/vin2 vss 1.74f
C14018 X1/X2/X3/vin1 vss 1.12f
C14019 X1/X2/X1/X3/m1_688_n494# vss 0.858f
C14020 X1/X2/X1/X3/m1_994_178# vss 1.15f
C14021 X1/X2/X1/X3/vin2 vss 1.85f
C14022 X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C14023 X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C14024 X1/X2/X1/X2/X3/vin2 vss 1.75f
C14025 X1/X2/X1/X2/X2/sw_0/m1_688_n494# vss 0.858f
C14026 X1/X2/X1/X2/X2/sw_0/m1_994_178# vss 1.15f
C14027 X1/X2/X1/X2/X2/X2/vout vss 0.868f
C14028 X1/X2/X1/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C14029 X1/X2/X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C14030 X1/X2/X1/X2/X2/X2/X2/vin1 vss 1.46f
C14031 X1/X2/X1/X2/X2/X2/X3/vin2 vss 1.23f
C14032 X1/X2/X1/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C14033 X1/X2/X1/X2/X2/X2/X2/m1_994_178# vss 1.15f
C14034 X1/X2/X2/vrefh vss 6.35f
C14035 X1/X2/X1/X2/X2/X2/X1/vin1 vss 1.91f
C14036 X1/X2/X1/X2/X2/X2/X3/vin1 vss 0.816f
C14037 X1/X2/X1/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C14038 X1/X2/X1/X2/X2/X2/X1/m1_994_178# vss 1.15f
C14039 X1/X2/X1/X2/X2/X2/X1/vin2 vss 1.73f
C14040 X1/X2/X1/X2/X2/X1/vout vss 0.607f
C14041 X1/X2/X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C14042 X1/X2/X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C14043 X1/X2/X1/X2/X2/X1/X2/vin1 vss 1.46f
C14044 X1/X2/X1/X2/X2/X1/X3/vin2 vss 1.23f
C14045 X1/X2/X1/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C14046 X1/X2/X1/X2/X2/X1/X2/m1_994_178# vss 1.15f
C14047 X1/X2/X1/X2/X2/X2/vrefh vss 3.27f
C14048 X1/X2/X1/X2/X2/X1/X1/vin1 vss 1.91f
C14049 X1/X2/X1/X2/X2/X1/X3/vin1 vss 0.816f
C14050 X1/X2/X1/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C14051 X1/X2/X1/X2/X2/X1/X1/m1_994_178# vss 1.15f
C14052 X1/X2/X1/X2/X2/X1/X1/vin2 vss 1.73f
C14053 X1/X2/X1/X2/X3/vin1 vss 1.49f
C14054 X1/X2/X1/X2/X1/sw_0/m1_688_n494# vss 0.858f
C14055 X1/X2/X1/X2/X1/sw_0/m1_994_178# vss 1.15f
C14056 X1/X2/X1/X2/X1/X2/vout vss 0.868f
C14057 X1/X2/X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C14058 X1/X2/X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C14059 X1/X2/X1/X2/X1/X2/X2/vin1 vss 1.46f
C14060 X1/X2/X1/X2/X1/X2/X3/vin2 vss 1.23f
C14061 X1/X2/X1/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C14062 X1/X2/X1/X2/X1/X2/X2/m1_994_178# vss 1.15f
C14063 X1/X2/X1/X2/X2/vrefh vss 3.27f
C14064 X1/X2/X1/X2/X1/X2/X1/vin1 vss 1.91f
C14065 X1/X2/X1/X2/X1/X2/X3/vin1 vss 0.816f
C14066 X1/X2/X1/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C14067 X1/X2/X1/X2/X1/X2/X1/m1_994_178# vss 1.15f
C14068 X1/X2/X1/X2/X1/X2/X1/vin2 vss 1.73f
C14069 X1/X2/X1/X2/X1/X1/vout vss 0.607f
C14070 X1/X2/X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C14071 X1/X2/X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C14072 X1/X2/X1/X2/X1/X1/X2/vin1 vss 1.46f
C14073 X1/X2/X1/X2/X1/X1/X3/vin2 vss 1.23f
C14074 X1/X2/X1/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C14075 X1/X2/X1/X2/X1/X1/X2/m1_994_178# vss 1.15f
C14076 X1/X2/X1/X2/X1/X2/vrefh vss 3.27f
C14077 X1/X2/X1/X2/X1/X1/X1/vin1 vss 1.91f
C14078 X1/X2/X1/X2/X1/X1/X3/vin1 vss 0.816f
C14079 X1/X2/X1/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C14080 X1/X2/X1/X2/X1/X1/X1/m1_994_178# vss 1.15f
C14081 X1/X2/X1/X2/X1/X1/X1/vin2 vss 1.73f
C14082 X1/X2/X1/X3/vin1 vss 1.6f
C14083 X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C14084 X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C14085 X1/X2/X1/X1/X3/vin2 vss 1.75f
C14086 X1/X2/X1/X1/X2/sw_0/m1_688_n494# vss 0.858f
C14087 X1/X2/X1/X1/X2/sw_0/m1_994_178# vss 1.15f
C14088 X1/X2/X1/X1/X2/X2/vout vss 0.868f
C14089 X1/X2/X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C14090 X1/X2/X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C14091 X1/X2/X1/X1/X2/X2/X2/vin1 vss 1.46f
C14092 X1/X2/X1/X1/X2/X2/X3/vin2 vss 1.23f
C14093 X1/X2/X1/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C14094 X1/X2/X1/X1/X2/X2/X2/m1_994_178# vss 1.15f
C14095 X1/X2/X1/X2/vrefh vss 3.27f
C14096 X1/X2/X1/X1/X2/X2/X1/vin1 vss 1.91f
C14097 X1/X2/X1/X1/X2/X2/X3/vin1 vss 0.816f
C14098 X1/X2/X1/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C14099 X1/X2/X1/X1/X2/X2/X1/m1_994_178# vss 1.15f
C14100 X1/X2/X1/X1/X2/X2/X1/vin2 vss 1.73f
C14101 X1/X2/X1/X1/X2/X1/vout vss 0.607f
C14102 X1/X2/X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C14103 X1/X2/X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C14104 X1/X2/X1/X1/X2/X1/X2/vin1 vss 1.46f
C14105 X1/X2/X1/X1/X2/X1/X3/vin2 vss 1.23f
C14106 X1/X2/X1/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C14107 X1/X2/X1/X1/X2/X1/X2/m1_994_178# vss 1.15f
C14108 X1/X2/X1/X1/X2/X2/vrefh vss 3.27f
C14109 X1/X2/X1/X1/X2/X1/X1/vin1 vss 1.91f
C14110 X1/X2/X1/X1/X2/X1/X3/vin1 vss 0.816f
C14111 X1/X2/X1/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C14112 X1/X2/X1/X1/X2/X1/X1/m1_994_178# vss 1.15f
C14113 X1/X2/X1/X1/X2/X1/X1/vin2 vss 1.73f
C14114 X1/X2/X1/X1/X3/vin1 vss 1.49f
C14115 X1/X2/X1/X1/X1/sw_0/m1_688_n494# vss 0.858f
C14116 X1/X2/X1/X1/X1/sw_0/m1_994_178# vss 1.15f
C14117 X1/X2/X1/X1/X1/X2/vout vss 0.868f
C14118 X1/X2/X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C14119 X1/X2/X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C14120 X1/X2/X1/X1/X1/X2/X2/vin1 vss 1.46f
C14121 X1/X2/X1/X1/X1/X2/X3/vin2 vss 1.23f
C14122 X1/X2/X1/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C14123 X1/X2/X1/X1/X1/X2/X2/m1_994_178# vss 1.15f
C14124 X1/X2/X1/X1/X2/vrefh vss 3.27f
C14125 X1/X2/X1/X1/X1/X2/X1/vin1 vss 1.91f
C14126 X1/X2/X1/X1/X1/X2/X3/vin1 vss 0.816f
C14127 X1/X2/X1/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C14128 X1/X2/X1/X1/X1/X2/X1/m1_994_178# vss 1.15f
C14129 X1/X2/X1/X1/X1/X2/X1/vin2 vss 1.73f
C14130 X1/X2/X1/X1/X1/X1/vout vss 0.607f
C14131 X1/X2/X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C14132 X1/X2/X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C14133 X1/X2/X1/X1/X1/X1/X2/vin1 vss 1.46f
C14134 X1/X2/X1/X1/X1/X1/X3/vin2 vss 1.23f
C14135 X1/X2/X1/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C14136 X1/X2/X1/X1/X1/X1/X2/m1_994_178# vss 1.15f
C14137 X1/X2/X1/X1/X1/X2/vrefh vss 3.27f
C14138 X1/X2/X1/X1/X1/X1/X1/vin1 vss 1.96f
C14139 X1/X2/X1/X1/X1/X1/X3/vin1 vss 0.816f
C14140 X1/X2/X1/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C14141 X1/X2/X1/X1/X1/X1/X1/m1_994_178# vss 1.15f
C14142 X1/X2/X1/X1/X1/X1/X1/vin2 vss 1.74f
C14143 X1/X3/vin1 vss 1.34f
C14144 X1/X1/X3/m1_688_n494# vss 0.858f
C14145 X1/X1/X3/m1_994_178# vss 1.15f
C14146 X1/X1/X3/vin2 vss 1.27f
C14147 X1/X1/X2/X3/m1_688_n494# vss 0.858f
C14148 X1/X1/X2/X3/m1_994_178# vss 1.15f
C14149 X1/X1/X2/X3/vin2 vss 1.85f
C14150 X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C14151 X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C14152 X1/X1/X2/X2/X3/vin2 vss 1.75f
C14153 X1/X1/X2/X2/X2/sw_0/m1_688_n494# vss 0.858f
C14154 X1/X1/X2/X2/X2/sw_0/m1_994_178# vss 1.15f
C14155 X1/X1/X2/X2/X2/X2/vout vss 0.868f
C14156 X1/X1/X2/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C14157 X1/X1/X2/X2/X2/X2/X3/m1_994_178# vss 1.15f
C14158 X1/X1/X2/X2/X2/X2/X2/vin1 vss 1.46f
C14159 X1/X1/X2/X2/X2/X2/X3/vin2 vss 1.24f
C14160 X1/X1/X2/X2/X2/X2/X2/m1_688_n494# vss 0.859f
C14161 X1/X1/X2/X2/X2/X2/X2/m1_994_178# vss 1.15f
C14162 X1/X2/vrefh vss 4.1f
C14163 X1/X1/X2/X2/X2/X2/X1/vin1 vss 1.91f
C14164 X1/X1/X2/X2/X2/X2/X3/vin1 vss 0.816f
C14165 X1/X1/X2/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C14166 X1/X1/X2/X2/X2/X2/X1/m1_994_178# vss 1.15f
C14167 X1/X1/X2/X2/X2/X2/X1/vin2 vss 1.73f
C14168 X1/X1/X2/X2/X2/X1/vout vss 0.607f
C14169 X1/X1/X2/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C14170 X1/X1/X2/X2/X2/X1/X3/m1_994_178# vss 1.15f
C14171 X1/X1/X2/X2/X2/X1/X2/vin1 vss 1.46f
C14172 X1/X1/X2/X2/X2/X1/X3/vin2 vss 1.23f
C14173 X1/X1/X2/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C14174 X1/X1/X2/X2/X2/X1/X2/m1_994_178# vss 1.15f
C14175 X1/X1/X2/X2/X2/X2/vrefh vss 3.27f
C14176 X1/X1/X2/X2/X2/X1/X1/vin1 vss 1.91f
C14177 X1/X1/X2/X2/X2/X1/X3/vin1 vss 0.816f
C14178 X1/X1/X2/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C14179 X1/X1/X2/X2/X2/X1/X1/m1_994_178# vss 1.15f
C14180 X1/X1/X2/X2/X2/X1/X1/vin2 vss 1.73f
C14181 X1/X1/X2/X2/X3/vin1 vss 1.49f
C14182 X1/X1/X2/X2/X1/sw_0/m1_688_n494# vss 0.858f
C14183 X1/X1/X2/X2/X1/sw_0/m1_994_178# vss 1.15f
C14184 X1/X1/X2/X2/X1/X2/vout vss 0.868f
C14185 X1/X1/X2/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C14186 X1/X1/X2/X2/X1/X2/X3/m1_994_178# vss 1.15f
C14187 X1/X1/X2/X2/X1/X2/X2/vin1 vss 1.46f
C14188 X1/X1/X2/X2/X1/X2/X3/vin2 vss 1.23f
C14189 X1/X1/X2/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C14190 X1/X1/X2/X2/X1/X2/X2/m1_994_178# vss 1.15f
C14191 X1/X1/X2/X2/X2/vrefh vss 3.27f
C14192 X1/X1/X2/X2/X1/X2/X1/vin1 vss 1.91f
C14193 X1/X1/X2/X2/X1/X2/X3/vin1 vss 0.816f
C14194 X1/X1/X2/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C14195 X1/X1/X2/X2/X1/X2/X1/m1_994_178# vss 1.15f
C14196 X1/X1/X2/X2/X1/X2/X1/vin2 vss 1.73f
C14197 X1/X1/X2/X2/X1/X1/vout vss 0.607f
C14198 X1/X1/X2/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C14199 X1/X1/X2/X2/X1/X1/X3/m1_994_178# vss 1.15f
C14200 X1/X1/X2/X2/X1/X1/X2/vin1 vss 1.46f
C14201 X1/X1/X2/X2/X1/X1/X3/vin2 vss 1.23f
C14202 X1/X1/X2/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C14203 X1/X1/X2/X2/X1/X1/X2/m1_994_178# vss 1.15f
C14204 X1/X1/X2/X2/X1/X2/vrefh vss 3.27f
C14205 X1/X1/X2/X2/X1/X1/X1/vin1 vss 1.91f
C14206 X1/X1/X2/X2/X1/X1/X3/vin1 vss 0.816f
C14207 X1/X1/X2/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C14208 X1/X1/X2/X2/X1/X1/X1/m1_994_178# vss 1.15f
C14209 X1/X1/X2/X2/X1/X1/X1/vin2 vss 1.73f
C14210 X1/X1/X2/X3/vin1 vss 1.6f
C14211 X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C14212 X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C14213 X1/X1/X2/X1/X3/vin2 vss 1.75f
C14214 X1/X1/X2/X1/X2/sw_0/m1_688_n494# vss 0.858f
C14215 X1/X1/X2/X1/X2/sw_0/m1_994_178# vss 1.15f
C14216 X1/X1/X2/X1/X2/X2/vout vss 0.868f
C14217 X1/X1/X2/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C14218 X1/X1/X2/X1/X2/X2/X3/m1_994_178# vss 1.15f
C14219 X1/X1/X2/X1/X2/X2/X2/vin1 vss 1.46f
C14220 X1/X1/X2/X1/X2/X2/X3/vin2 vss 1.23f
C14221 X1/X1/X2/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C14222 X1/X1/X2/X1/X2/X2/X2/m1_994_178# vss 1.15f
C14223 X1/X1/X2/X2/vrefh vss 3.27f
C14224 X1/X1/X2/X1/X2/X2/X1/vin1 vss 1.91f
C14225 X1/X1/X2/X1/X2/X2/X3/vin1 vss 0.816f
C14226 X1/X1/X2/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C14227 X1/X1/X2/X1/X2/X2/X1/m1_994_178# vss 1.15f
C14228 X1/X1/X2/X1/X2/X2/X1/vin2 vss 1.73f
C14229 X1/X1/X2/X1/X2/X1/vout vss 0.607f
C14230 X1/X1/X2/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C14231 X1/X1/X2/X1/X2/X1/X3/m1_994_178# vss 1.15f
C14232 X1/X1/X2/X1/X2/X1/X2/vin1 vss 1.46f
C14233 X1/X1/X2/X1/X2/X1/X3/vin2 vss 1.23f
C14234 X1/X1/X2/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C14235 X1/X1/X2/X1/X2/X1/X2/m1_994_178# vss 1.15f
C14236 X1/X1/X2/X1/X2/X2/vrefh vss 3.27f
C14237 X1/X1/X2/X1/X2/X1/X1/vin1 vss 1.91f
C14238 X1/X1/X2/X1/X2/X1/X3/vin1 vss 0.816f
C14239 X1/X1/X2/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C14240 X1/X1/X2/X1/X2/X1/X1/m1_994_178# vss 1.15f
C14241 X1/X1/X2/X1/X2/X1/X1/vin2 vss 1.73f
C14242 X1/X1/X2/X1/X3/vin1 vss 1.49f
C14243 X1/X1/X2/X1/X1/sw_0/m1_688_n494# vss 0.858f
C14244 X1/X1/X2/X1/X1/sw_0/m1_994_178# vss 1.15f
C14245 X1/X1/X2/X1/X1/X2/vout vss 0.868f
C14246 X1/X1/X2/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C14247 X1/X1/X2/X1/X1/X2/X3/m1_994_178# vss 1.15f
C14248 X1/X1/X2/X1/X1/X2/X2/vin1 vss 1.46f
C14249 X1/X1/X2/X1/X1/X2/X3/vin2 vss 1.23f
C14250 X1/X1/X2/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C14251 X1/X1/X2/X1/X1/X2/X2/m1_994_178# vss 1.15f
C14252 X1/X1/X2/X1/X2/vrefh vss 3.27f
C14253 X1/X1/X2/X1/X1/X2/X1/vin1 vss 1.91f
C14254 X1/X1/X2/X1/X1/X2/X3/vin1 vss 0.816f
C14255 X1/X1/X2/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C14256 X1/X1/X2/X1/X1/X2/X1/m1_994_178# vss 1.15f
C14257 X1/X1/X2/X1/X1/X2/X1/vin2 vss 1.73f
C14258 X1/X1/X2/X1/X1/X1/vout vss 0.607f
C14259 X1/X1/X2/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C14260 X1/X1/X2/X1/X1/X1/X3/m1_994_178# vss 1.15f
C14261 X1/X1/X2/X1/X1/X1/X2/vin1 vss 1.46f
C14262 X1/X1/X2/X1/X1/X1/X3/vin2 vss 1.23f
C14263 X1/X1/X2/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C14264 X1/X1/X2/X1/X1/X1/X2/m1_994_178# vss 1.15f
C14265 X1/X1/X2/X1/X1/X2/vrefh vss 3.27f
C14266 X1/X1/X2/X1/X1/X1/X1/vin1 vss 1.91f
C14267 X1/X1/X2/X1/X1/X1/X3/vin1 vss 0.816f
C14268 X1/X1/X2/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C14269 X1/X1/X2/X1/X1/X1/X1/m1_994_178# vss 1.15f
C14270 X1/X1/X2/X1/X1/X1/X1/vin2 vss 1.73f
C14271 d4 vss 8.18f
C14272 X1/X1/X3/vin1 vss 1.12f
C14273 X1/X1/X1/X3/m1_688_n494# vss 0.858f
C14274 X1/X1/X1/X3/m1_994_178# vss 1.15f
C14275 d3 vss 32.9f
C14276 X1/X1/X1/X3/vin2 vss 1.85f
C14277 X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C14278 X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C14279 d2 vss 51.4f
C14280 X1/X1/X1/X2/X3/vin2 vss 1.75f
C14281 X1/X1/X1/X2/X2/sw_0/m1_688_n494# vss 0.858f
C14282 X1/X1/X1/X2/X2/sw_0/m1_994_178# vss 1.15f
C14283 X1/X1/X1/X2/X2/X2/vout vss 0.868f
C14284 X1/X1/X1/X2/X2/X2/X3/m1_688_n494# vss 0.858f
C14285 X1/X1/X1/X2/X2/X2/X3/m1_994_178# vss 1.15f
C14286 d0 vss 0.147p
C14287 X1/X1/X1/X2/X2/X2/X2/vin1 vss 1.46f
C14288 X1/X1/X1/X2/X2/X2/X3/vin2 vss 1.23f
C14289 X1/X1/X1/X2/X2/X2/X2/m1_688_n494# vss 0.858f
C14290 X1/X1/X1/X2/X2/X2/X2/m1_994_178# vss 1.15f
C14291 X1/X1/X2/vrefh vss 6.35f
C14292 X1/X1/X1/X2/X2/X2/X1/vin1 vss 1.91f
C14293 X1/X1/X1/X2/X2/X2/X3/vin1 vss 0.816f
C14294 X1/X1/X1/X2/X2/X2/X1/m1_688_n494# vss 0.858f
C14295 X1/X1/X1/X2/X2/X2/X1/m1_994_178# vss 1.15f
C14296 X1/X1/X1/X2/X2/X2/X1/vin2 vss 1.73f
C14297 X1/X1/X1/X2/X2/X1/vout vss 0.607f
C14298 X1/X1/X1/X2/X2/X1/X3/m1_688_n494# vss 0.858f
C14299 X1/X1/X1/X2/X2/X1/X3/m1_994_178# vss 1.15f
C14300 X1/X1/X1/X2/X2/X1/X2/vin1 vss 1.46f
C14301 X1/X1/X1/X2/X2/X1/X3/vin2 vss 1.23f
C14302 X1/X1/X1/X2/X2/X1/X2/m1_688_n494# vss 0.858f
C14303 X1/X1/X1/X2/X2/X1/X2/m1_994_178# vss 1.15f
C14304 X1/X1/X1/X2/X2/X2/vrefh vss 3.27f
C14305 X1/X1/X1/X2/X2/X1/X1/vin1 vss 1.91f
C14306 X1/X1/X1/X2/X2/X1/X3/vin1 vss 0.816f
C14307 X1/X1/X1/X2/X2/X1/X1/m1_688_n494# vss 0.858f
C14308 X1/X1/X1/X2/X2/X1/X1/m1_994_178# vss 1.15f
C14309 X1/X1/X1/X2/X2/X1/X1/vin2 vss 1.73f
C14310 X1/X1/X1/X2/X3/vin1 vss 1.49f
C14311 X1/X1/X1/X2/X1/sw_0/m1_688_n494# vss 0.858f
C14312 X1/X1/X1/X2/X1/sw_0/m1_994_178# vss 1.15f
C14313 X1/X1/X1/X2/X1/X2/vout vss 0.868f
C14314 X1/X1/X1/X2/X1/X2/X3/m1_688_n494# vss 0.858f
C14315 X1/X1/X1/X2/X1/X2/X3/m1_994_178# vss 1.15f
C14316 X1/X1/X1/X2/X1/X2/X2/vin1 vss 1.46f
C14317 X1/X1/X1/X2/X1/X2/X3/vin2 vss 1.23f
C14318 X1/X1/X1/X2/X1/X2/X2/m1_688_n494# vss 0.858f
C14319 X1/X1/X1/X2/X1/X2/X2/m1_994_178# vss 1.15f
C14320 X1/X1/X1/X2/X2/vrefh vss 3.27f
C14321 X1/X1/X1/X2/X1/X2/X1/vin1 vss 1.91f
C14322 X1/X1/X1/X2/X1/X2/X3/vin1 vss 0.816f
C14323 X1/X1/X1/X2/X1/X2/X1/m1_688_n494# vss 0.858f
C14324 X1/X1/X1/X2/X1/X2/X1/m1_994_178# vss 1.15f
C14325 X1/X1/X1/X2/X1/X2/X1/vin2 vss 1.73f
C14326 X1/X1/X1/X2/X1/X1/vout vss 0.607f
C14327 X1/X1/X1/X2/X1/X1/X3/m1_688_n494# vss 0.858f
C14328 X1/X1/X1/X2/X1/X1/X3/m1_994_178# vss 1.15f
C14329 X1/X1/X1/X2/X1/X1/X2/vin1 vss 1.46f
C14330 X1/X1/X1/X2/X1/X1/X3/vin2 vss 1.23f
C14331 X1/X1/X1/X2/X1/X1/X2/m1_688_n494# vss 0.858f
C14332 X1/X1/X1/X2/X1/X1/X2/m1_994_178# vss 1.15f
C14333 X1/X1/X1/X2/X1/X2/vrefh vss 3.27f
C14334 X1/X1/X1/X2/X1/X1/X1/vin1 vss 1.91f
C14335 X1/X1/X1/X2/X1/X1/X3/vin1 vss 0.816f
C14336 X1/X1/X1/X2/X1/X1/X1/m1_688_n494# vss 0.858f
C14337 X1/X1/X1/X2/X1/X1/X1/m1_994_178# vss 1.15f
C14338 X1/X1/X1/X2/X1/X1/X1/vin2 vss 1.73f
C14339 X1/X1/X1/X3/vin1 vss 1.6f
C14340 X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C14341 X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C14342 X1/X1/X1/X1/X3/vin2 vss 1.75f
C14343 X1/X1/X1/X1/X2/sw_0/m1_688_n494# vss 0.858f
C14344 X1/X1/X1/X1/X2/sw_0/m1_994_178# vss 1.15f
C14345 X1/X1/X1/X1/X2/X2/vout vss 0.868f
C14346 X1/X1/X1/X1/X2/X2/X3/m1_688_n494# vss 0.858f
C14347 X1/X1/X1/X1/X2/X2/X3/m1_994_178# vss 1.15f
C14348 X1/X1/X1/X1/X2/X2/X2/vin1 vss 1.46f
C14349 X1/X1/X1/X1/X2/X2/X3/vin2 vss 1.23f
C14350 X1/X1/X1/X1/X2/X2/X2/m1_688_n494# vss 0.858f
C14351 X1/X1/X1/X1/X2/X2/X2/m1_994_178# vss 1.15f
C14352 X1/X1/X1/X2/vrefh vss 3.27f
C14353 X1/X1/X1/X1/X2/X2/X1/vin1 vss 1.91f
C14354 X1/X1/X1/X1/X2/X2/X3/vin1 vss 0.816f
C14355 X1/X1/X1/X1/X2/X2/X1/m1_688_n494# vss 0.858f
C14356 X1/X1/X1/X1/X2/X2/X1/m1_994_178# vss 1.15f
C14357 X1/X1/X1/X1/X2/X2/X1/vin2 vss 1.73f
C14358 X1/X1/X1/X1/X2/X1/vout vss 0.607f
C14359 X1/X1/X1/X1/X2/X1/X3/m1_688_n494# vss 0.858f
C14360 X1/X1/X1/X1/X2/X1/X3/m1_994_178# vss 1.15f
C14361 X1/X1/X1/X1/X2/X1/X2/vin1 vss 1.46f
C14362 X1/X1/X1/X1/X2/X1/X3/vin2 vss 1.23f
C14363 X1/X1/X1/X1/X2/X1/X2/m1_688_n494# vss 0.858f
C14364 X1/X1/X1/X1/X2/X1/X2/m1_994_178# vss 1.15f
C14365 X1/X1/X1/X1/X2/X2/vrefh vss 3.27f
C14366 X1/X1/X1/X1/X2/X1/X1/vin1 vss 1.91f
C14367 X1/X1/X1/X1/X2/X1/X3/vin1 vss 0.816f
C14368 X1/X1/X1/X1/X2/X1/X1/m1_688_n494# vss 0.858f
C14369 X1/X1/X1/X1/X2/X1/X1/m1_994_178# vss 1.15f
C14370 X1/X1/X1/X1/X2/X1/X1/vin2 vss 1.73f
C14371 X1/X1/X1/X1/X3/vin1 vss 1.49f
C14372 X1/X1/X1/X1/X1/sw_0/m1_688_n494# vss 0.858f
C14373 X1/X1/X1/X1/X1/sw_0/m1_994_178# vss 1.15f
C14374 d1 vss 65.4f
C14375 X1/X1/X1/X1/X1/X2/vout vss 0.868f
C14376 X1/X1/X1/X1/X1/X2/X3/m1_688_n494# vss 0.858f
C14377 X1/X1/X1/X1/X1/X2/X3/m1_994_178# vss 1.15f
C14378 X1/X1/X1/X1/X1/X2/X2/vin1 vss 1.46f
C14379 X1/X1/X1/X1/X1/X2/X3/vin2 vss 1.23f
C14380 X1/X1/X1/X1/X1/X2/X2/m1_688_n494# vss 0.858f
C14381 X1/X1/X1/X1/X1/X2/X2/m1_994_178# vss 1.15f
C14382 X1/X1/X1/X1/X2/vrefh vss 3.27f
C14383 X1/X1/X1/X1/X1/X2/X1/vin1 vss 1.91f
C14384 X1/X1/X1/X1/X1/X2/X3/vin1 vss 0.816f
C14385 X1/X1/X1/X1/X1/X2/X1/m1_688_n494# vss 0.858f
C14386 X1/X1/X1/X1/X1/X2/X1/m1_994_178# vss 1.15f
C14387 X1/X1/X1/X1/X1/X2/X1/vin2 vss 1.73f
C14388 X1/X1/X1/X1/X1/X1/vout vss 0.607f
C14389 X1/X1/X1/X1/X1/X1/X3/m1_688_n494# vss 0.858f
C14390 X1/X1/X1/X1/X1/X1/X3/m1_994_178# vss 1.15f
C14391 X1/X1/X1/X1/X1/X1/X2/vin1 vss 1.46f
C14392 X1/X1/X1/X1/X1/X1/X3/vin2 vss 1.23f
C14393 X1/X1/X1/X1/X1/X1/X2/m1_688_n494# vss 0.858f
C14394 X1/X1/X1/X1/X1/X1/X2/m1_994_178# vss 1.15f
C14395 X1/X1/X1/X1/X1/X2/vrefh vss 3.27f
C14396 X1/X1/X1/X1/X1/X1/X1/vin1 vss 1.91f
C14397 X1/X1/X1/X1/X1/X1/X3/vin1 vss 0.816f
C14398 X1/X1/X1/X1/X1/X1/X1/m1_688_n494# vss 0.858f
C14399 X1/X1/X1/X1/X1/X1/X1/m1_994_178# vss 1.15f
C14400 X1/X1/X1/X1/X1/X1/X1/vin2 vss 1.73f
C14401 vrefh vss 1.11f
.ends

