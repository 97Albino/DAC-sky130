** sch_path: /home/97ms/uci/ip/dac5v/1.schematics/sw.sch

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/corners/tt.spice
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /mnt/tools4/open_pdks/sky130/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice

.subckt sw vdd vss din vin1 vin2 vout
XM1 net1 din vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1
XM2 net2 net1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1
XM3 vout net1 vin1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1
XM4 vin2 net2 vout vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1
XM5 net1 din vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42
XM6 net2 net1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42
XM7 vout net1 vin2 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42
XM8 vin1 net2 vout vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.42
.ends
