** sch_path: /home/97ms/uci/ip/dac5v/1.schematics/7bit_dac.sch

.include 6bit_dac.spice

.subckt 7bit_dac vdd vss vrefh vrefl d0 d1 d2 d3 d4 d5 d6 vout
X1 vdd vss vrefh net3 d0 d1 d2 d3 d4 d5 net1 6bit_dac
X2 vdd vss net3 vrefl d0 d1 d2 d3 d4 d5 net2 6bit_dac
X3 vdd vss d6 net1 net2 vout sw
.ends
