magic
tech sky130B
magscale 1 2
timestamp 1687214045
<< checkpaint >>
rect -874 2311 2138 2392
rect -1313 -713 2138 2311
rect -1260 -766 2138 -713
rect -1260 -3260 1460 -766
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__nfet_01v8_ZFH27D  XM1
timestamp 0
transform 1 0 193 0 1 799
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_XPYSY6  XM2
timestamp 0
transform 1 0 632 0 1 813
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 out
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 p_body
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 n_body
port 5 nsew
<< end >>
